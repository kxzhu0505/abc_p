// Benchmark "merged" written by ABC on Fri Sep  8 10:27:45 2023

module merged ( 
    ys__n14, ys__n16, ys__n22, ys__n24, ys__n26, ys__n28, ys__n30, ys__n32,
    ys__n34, ys__n36, ys__n38, ys__n40, ys__n42, ys__n44, ys__n46, ys__n48,
    ys__n50, ys__n52, ys__n54, ys__n56, ys__n58, ys__n60, ys__n62, ys__n66,
    ys__n70, ys__n72, ys__n74, ys__n76, ys__n78, ys__n80, ys__n82, ys__n84,
    ys__n86, ys__n88, ys__n90, ys__n96, ys__n98, ys__n100, ys__n108,
    ys__n110, ys__n112, ys__n114, ys__n116, ys__n118, ys__n120, ys__n122,
    ys__n124, ys__n126, ys__n128, ys__n130, ys__n132, ys__n134, ys__n136,
    ys__n138, ys__n140, ys__n142, ys__n148, ys__n150, ys__n152, ys__n156,
    ys__n158, ys__n160, ys__n162, ys__n164, ys__n166, ys__n168, ys__n170,
    ys__n172, ys__n174, ys__n176, ys__n178, ys__n182, ys__n184, ys__n186,
    ys__n190, ys__n192, ys__n194, ys__n196, ys__n198, ys__n202, ys__n204,
    ys__n206, ys__n208, ys__n210, ys__n212, ys__n214, ys__n216, ys__n218,
    ys__n220, ys__n222, ys__n226, ys__n232, ys__n238, ys__n240, ys__n242,
    ys__n244, ys__n248, ys__n256, ys__n258, ys__n262, ys__n290, ys__n294,
    ys__n296, ys__n298, ys__n300, ys__n302, ys__n304, ys__n306, ys__n308,
    ys__n310, ys__n312, ys__n314, ys__n316, ys__n318, ys__n326, ys__n328,
    ys__n330, ys__n332, ys__n336, ys__n338, ys__n340, ys__n342, ys__n344,
    ys__n346, ys__n348, ys__n350, ys__n352, ys__n354, ys__n356, ys__n358,
    ys__n360, ys__n362, ys__n364, ys__n366, ys__n368, ys__n370, ys__n372,
    ys__n374, ys__n376, ys__n378, ys__n380, ys__n382, ys__n384, ys__n386,
    ys__n392, ys__n394, ys__n396, ys__n398, ys__n402, ys__n408, ys__n414,
    ys__n416, ys__n418, ys__n420, ys__n422, ys__n424, ys__n426, ys__n428,
    ys__n430, ys__n432, ys__n434, ys__n436, ys__n438, ys__n440, ys__n442,
    ys__n444, ys__n446, ys__n448, ys__n450, ys__n452, ys__n454, ys__n456,
    ys__n464, ys__n488, ys__n490, ys__n500, ys__n504, ys__n512, ys__n514,
    ys__n516, ys__n518, ys__n520, ys__n522, ys__n524, ys__n526, ys__n528,
    ys__n530, ys__n532, ys__n536, ys__n538, ys__n544, ys__n546, ys__n548,
    ys__n550, ys__n556, ys__n558, ys__n562, ys__n564, ys__n566, ys__n568,
    ys__n570, ys__n572, ys__n580, ys__n582, ys__n584, ys__n586, ys__n588,
    ys__n598, ys__n600, ys__n602, ys__n604, ys__n606, ys__n608, ys__n610,
    ys__n612, ys__n614, ys__n616, ys__n618, ys__n620, ys__n622, ys__n624,
    ys__n626, ys__n632, ys__n634, ys__n636, ys__n638, ys__n640, ys__n642,
    ys__n644, ys__n646, ys__n648, ys__n650, ys__n652, ys__n654, ys__n656,
    ys__n658, ys__n660, ys__n662, ys__n664, ys__n666, ys__n668, ys__n670,
    ys__n672, ys__n674, ys__n676, ys__n678, ys__n680, ys__n682, ys__n684,
    ys__n686, ys__n688, ys__n690, ys__n692, ys__n694, ys__n696, ys__n698,
    ys__n700, ys__n702, ys__n704, ys__n706, ys__n708, ys__n710, ys__n712,
    ys__n718, ys__n720, ys__n722, ys__n724, ys__n726, ys__n728, ys__n736,
    ys__n742, ys__n744, ys__n746, ys__n748, ys__n750, ys__n752, ys__n758,
    ys__n760, ys__n762, ys__n764, ys__n766, ys__n768, ys__n770, ys__n772,
    ys__n774, ys__n776, ys__n778, ys__n780, ys__n782, ys__n784, ys__n816,
    ys__n818, ys__n820, ys__n822, ys__n824, ys__n826, ys__n828, ys__n830,
    ys__n832, ys__n834, ys__n836, ys__n838, ys__n840, ys__n842, ys__n844,
    ys__n846, ys__n848, ys__n850, ys__n852, ys__n854, ys__n856, ys__n858,
    ys__n860, ys__n874, ys__n889, ys__n935, ys__n1029, ys__n1036,
    ys__n1038, ys__n1048, ys__n1072, ys__n1076, ys__n1078, ys__n1084,
    ys__n1094, ys__n1098, ys__n1099, ys__n1106, ys__n1107, ys__n1109,
    ys__n1110, ys__n1116, ys__n1117, ys__n1119, ys__n1120, ys__n1129,
    ys__n1147, ys__n1151, ys__n1153, ys__n1154, ys__n1156, ys__n1157,
    ys__n1301, ys__n1309, ys__n1489, ys__n1490, ys__n1492, ys__n1493,
    ys__n1495, ys__n1496, ys__n1498, ys__n1499, ys__n1502, ys__n1503,
    ys__n1505, ys__n1506, ys__n1508, ys__n1509, ys__n1511, ys__n1535,
    ys__n2024, ys__n2233, ys__n2239, ys__n2245, ys__n2247, ys__n2251,
    ys__n2276, ys__n2282, ys__n2306, ys__n2308, ys__n2312, ys__n2427,
    ys__n2429, ys__n2433, ys__n2644, ys__n2652, ys__n2693, ys__n2716,
    ys__n2779, ys__n2830, ys__n2924, ys__n3214, ys__n4168, ys__n4176,
    ys__n4177, ys__n4184, ys__n4185, ys__n4190, ys__n4291, ys__n4292,
    ys__n4294, ys__n4296, ys__n4297, ys__n4299, ys__n4300, ys__n4305,
    ys__n4340, ys__n4448, ys__n4449, ys__n4451, ys__n4452, ys__n4454,
    ys__n4455, ys__n4457, ys__n4458, ys__n4460, ys__n4461, ys__n4465,
    ys__n4478, ys__n4480, ys__n4488, ys__n4494, ys__n4496, ys__n4613,
    ys__n4625, ys__n4627, ys__n4688, ys__n4698, ys__n4736, ys__n4744,
    ys__n4746, ys__n4750, ys__n4751, ys__n4753, ys__n4754, ys__n4756,
    ys__n4757, ys__n4759, ys__n4761, ys__n4783, ys__n4784, ys__n4810,
    ys__n4826, ys__n4832, ys__n4833, ys__n4836, ys__n4837, ys__n6112,
    ys__n6113, ys__n6115, ys__n6118, ys__n6119, ys__n6120, ys__n6121,
    ys__n6123, ys__n6124, ys__n6126, ys__n6127, ys__n6129, ys__n6130,
    ys__n6133, ys__n6134, ys__n17803, ys__n17804, ys__n17806, ys__n17807,
    ys__n17809, ys__n17810, ys__n17812, ys__n17813, ys__n17815, ys__n17816,
    ys__n17818, ys__n17819, ys__n17821, ys__n17822, ys__n17824, ys__n17825,
    ys__n17827, ys__n17828, ys__n17830, ys__n17831, ys__n17833, ys__n17834,
    ys__n17836, ys__n17837, ys__n17839, ys__n17840, ys__n17842, ys__n17843,
    ys__n17845, ys__n17846, ys__n17848, ys__n17849, ys__n17866, ys__n17867,
    ys__n17869, ys__n17870, ys__n17872, ys__n17873, ys__n17875, ys__n17876,
    ys__n17878, ys__n17879, ys__n17881, ys__n17882, ys__n17884, ys__n17885,
    ys__n17887, ys__n17888, ys__n17890, ys__n17891, ys__n17893, ys__n17894,
    ys__n17896, ys__n17897, ys__n17899, ys__n17900, ys__n17902, ys__n17903,
    ys__n17905, ys__n17906, ys__n17908, ys__n17909, ys__n17911, ys__n17912,
    ys__n17941, ys__n17943, ys__n18041, ys__n18043, ys__n18045, ys__n18047,
    ys__n18049, ys__n18051, ys__n18053, ys__n18055, ys__n18057, ys__n18059,
    ys__n18061, ys__n18063, ys__n18065, ys__n18067, ys__n18070, ys__n18071,
    ys__n18090, ys__n18101, ys__n18105, ys__n18106, ys__n18109, ys__n18111,
    ys__n18112, ys__n18114, ys__n18116, ys__n18118, ys__n18121, ys__n18122,
    ys__n18124, ys__n18143, ys__n18149, ys__n18150, ys__n18156, ys__n18173,
    ys__n18208, ys__n18226, ys__n18229, ys__n18231, ys__n18240, ys__n18242,
    ys__n18243, ys__n18270, ys__n18271, ys__n18277, ys__n18280, ys__n18283,
    ys__n18286, ys__n18317, ys__n18378, ys__n18381, ys__n18384, ys__n18389,
    ys__n18393, ys__n18448, ys__n18451, ys__n18454, ys__n18457, ys__n18460,
    ys__n18463, ys__n18466, ys__n18469, ys__n18472, ys__n18475, ys__n18478,
    ys__n18481, ys__n18484, ys__n18487, ys__n18490, ys__n18493, ys__n18496,
    ys__n18499, ys__n18502, ys__n18505, ys__n18508, ys__n18511, ys__n18514,
    ys__n18517, ys__n18520, ys__n18523, ys__n18526, ys__n18529, ys__n18532,
    ys__n18535, ys__n18538, ys__n18541, ys__n18544, ys__n18546, ys__n18556,
    ys__n18558, ys__n18560, ys__n18562, ys__n18565, ys__n18568, ys__n18569,
    ys__n18571, ys__n18572, ys__n18574, ys__n18575, ys__n18577, ys__n18578,
    ys__n18580, ys__n18581, ys__n18583, ys__n18584, ys__n18586, ys__n18587,
    ys__n18589, ys__n18590, ys__n18592, ys__n18593, ys__n18595, ys__n18596,
    ys__n18598, ys__n18599, ys__n18601, ys__n18602, ys__n18604, ys__n18605,
    ys__n18607, ys__n18608, ys__n18610, ys__n18611, ys__n18613, ys__n18614,
    ys__n18616, ys__n18617, ys__n18619, ys__n18620, ys__n18622, ys__n18623,
    ys__n18625, ys__n18626, ys__n18628, ys__n18630, ys__n18632, ys__n18634,
    ys__n18636, ys__n18638, ys__n18639, ys__n18641, ys__n18642, ys__n18644,
    ys__n18645, ys__n18647, ys__n18650, ys__n18651, ys__n18749, ys__n18752,
    ys__n18755, ys__n18758, ys__n18761, ys__n18762, ys__n18765, ys__n18767,
    ys__n18769, ys__n18771, ys__n18773, ys__n18775, ys__n18777, ys__n18779,
    ys__n18781, ys__n18783, ys__n18785, ys__n18787, ys__n18789, ys__n18791,
    ys__n18793, ys__n18795, ys__n18797, ys__n18799, ys__n18801, ys__n18803,
    ys__n18805, ys__n18807, ys__n18809, ys__n18811, ys__n18813, ys__n18815,
    ys__n18817, ys__n18819, ys__n18821, ys__n18823, ys__n18825, ys__n18827,
    ys__n18829, ys__n18831, ys__n18833, ys__n18835, ys__n18837, ys__n18839,
    ys__n18841, ys__n18843, ys__n18845, ys__n18847, ys__n18849, ys__n18851,
    ys__n18853, ys__n18855, ys__n18857, ys__n18859, ys__n18861, ys__n18863,
    ys__n18865, ys__n18867, ys__n18869, ys__n18871, ys__n18873, ys__n18875,
    ys__n18877, ys__n18879, ys__n18881, ys__n18883, ys__n18885, ys__n18887,
    ys__n18889, ys__n18891, ys__n18956, ys__n18957, ys__n18958, ys__n18959,
    ys__n18960, ys__n18961, ys__n18962, ys__n18963, ys__n18964, ys__n18965,
    ys__n18966, ys__n18967, ys__n18968, ys__n18969, ys__n18970, ys__n18971,
    ys__n18972, ys__n18973, ys__n18974, ys__n18975, ys__n18976, ys__n18977,
    ys__n18978, ys__n18979, ys__n18980, ys__n18981, ys__n18982, ys__n18983,
    ys__n18984, ys__n18985, ys__n18986, ys__n18987, ys__n18989, ys__n18991,
    ys__n18993, ys__n18995, ys__n18997, ys__n18999, ys__n19001, ys__n19003,
    ys__n19005, ys__n19007, ys__n19009, ys__n19011, ys__n19013, ys__n19015,
    ys__n19017, ys__n19019, ys__n19021, ys__n19023, ys__n19025, ys__n19027,
    ys__n19029, ys__n19031, ys__n19033, ys__n19035, ys__n19037, ys__n19039,
    ys__n19041, ys__n19043, ys__n19045, ys__n19047, ys__n19049, ys__n19051,
    ys__n19116, ys__n19117, ys__n19118, ys__n19119, ys__n19120, ys__n19121,
    ys__n19122, ys__n19123, ys__n19124, ys__n19125, ys__n19126, ys__n19127,
    ys__n19128, ys__n19129, ys__n19130, ys__n19131, ys__n19132, ys__n19133,
    ys__n19134, ys__n19135, ys__n19136, ys__n19137, ys__n19138, ys__n19139,
    ys__n19140, ys__n19141, ys__n19142, ys__n19143, ys__n19144, ys__n19145,
    ys__n19146, ys__n19147, ys__n19156, ys__n19157, ys__n19166, ys__n19171,
    ys__n19203, ys__n19215, ys__n19245, ys__n19251, ys__n19253, ys__n19259,
    ys__n19261, ys__n19263, ys__n19843, ys__n19844, ys__n19845, ys__n19846,
    ys__n19847, ys__n19848, ys__n19849, ys__n19850, ys__n19851, ys__n19852,
    ys__n19853, ys__n19854, ys__n19855, ys__n19856, ys__n19857, ys__n19858,
    ys__n19859, ys__n19860, ys__n19861, ys__n19862, ys__n19863, ys__n19864,
    ys__n19865, ys__n19866, ys__n19867, ys__n19868, ys__n19869, ys__n19870,
    ys__n19871, ys__n19872, ys__n19873, ys__n19874, ys__n19875, ys__n19972,
    ys__n19973, ys__n19974, ys__n19975, ys__n19976, ys__n19977, ys__n19978,
    ys__n19979, ys__n19980, ys__n19981, ys__n19982, ys__n19983, ys__n19984,
    ys__n19985, ys__n19986, ys__n19987, ys__n19988, ys__n19989, ys__n19990,
    ys__n19991, ys__n19992, ys__n19993, ys__n19994, ys__n19995, ys__n19996,
    ys__n19997, ys__n19998, ys__n19999, ys__n20000, ys__n20001, ys__n20002,
    ys__n20003, ys__n20004, ys__n20035, ys__n20058, ys__n20061, ys__n20064,
    ys__n20067, ys__n20070, ys__n20073, ys__n20076, ys__n20079, ys__n20138,
    ys__n20140, ys__n20142, ys__n20144, ys__n20146, ys__n20148, ys__n20150,
    ys__n20152, ys__n20186, ys__n20188, ys__n20190, ys__n20192, ys__n20194,
    ys__n20196, ys__n20198, ys__n20200, ys__n20202, ys__n20204, ys__n20206,
    ys__n20208, ys__n20210, ys__n20212, ys__n20214, ys__n20216, ys__n20273,
    ys__n20279, ys__n20280, ys__n20540, ys__n20542, ys__n20544, ys__n20546,
    ys__n20548, ys__n20550, ys__n20552, ys__n20554, ys__n20556, ys__n20558,
    ys__n20560, ys__n20562, ys__n20564, ys__n20566, ys__n20568, ys__n20570,
    ys__n20572, ys__n20574, ys__n20576, ys__n20578, ys__n20580, ys__n20582,
    ys__n20584, ys__n20586, ys__n20588, ys__n20590, ys__n20592, ys__n20594,
    ys__n20596, ys__n20598, ys__n20600, ys__n20602, ys__n20604, ys__n20606,
    ys__n20608, ys__n20610, ys__n20612, ys__n20614, ys__n20616, ys__n20618,
    ys__n20620, ys__n20622, ys__n20624, ys__n20626, ys__n20628, ys__n20630,
    ys__n20632, ys__n20634, ys__n20636, ys__n20638, ys__n20640, ys__n20642,
    ys__n20644, ys__n20646, ys__n20648, ys__n20650, ys__n20652, ys__n20654,
    ys__n20656, ys__n20658, ys__n20660, ys__n20662, ys__n20664, ys__n20666,
    ys__n20668, ys__n20670, ys__n20672, ys__n20674, ys__n20676, ys__n20678,
    ys__n20680, ys__n20682, ys__n20684, ys__n20686, ys__n20688, ys__n20690,
    ys__n20692, ys__n20694, ys__n20696, ys__n20698, ys__n20700, ys__n20702,
    ys__n20704, ys__n20706, ys__n20708, ys__n20710, ys__n20712, ys__n20714,
    ys__n20716, ys__n20718, ys__n20720, ys__n20722, ys__n20724, ys__n20726,
    ys__n20728, ys__n20730, ys__n20732, ys__n20734, ys__n20736, ys__n20738,
    ys__n20740, ys__n20742, ys__n20744, ys__n20746, ys__n20748, ys__n20750,
    ys__n20752, ys__n20754, ys__n20756, ys__n20758, ys__n20760, ys__n20762,
    ys__n20764, ys__n20766, ys__n20768, ys__n20770, ys__n20772, ys__n20774,
    ys__n20776, ys__n20778, ys__n20780, ys__n20782, ys__n20784, ys__n20786,
    ys__n20788, ys__n20790, ys__n20792, ys__n20794, ys__n20796, ys__n20798,
    ys__n20800, ys__n20802, ys__n20804, ys__n20806, ys__n20808, ys__n20810,
    ys__n20812, ys__n20814, ys__n20816, ys__n20818, ys__n20820, ys__n20822,
    ys__n20824, ys__n20826, ys__n20828, ys__n20830, ys__n20832, ys__n20834,
    ys__n20836, ys__n20838, ys__n20840, ys__n20842, ys__n20844, ys__n20846,
    ys__n20848, ys__n20850, ys__n20852, ys__n20854, ys__n20856, ys__n20858,
    ys__n20860, ys__n20862, ys__n20864, ys__n20866, ys__n20868, ys__n20870,
    ys__n20872, ys__n20874, ys__n20876, ys__n20878, ys__n20880, ys__n20882,
    ys__n20884, ys__n20886, ys__n20888, ys__n20890, ys__n20892, ys__n20894,
    ys__n20896, ys__n20898, ys__n20900, ys__n20902, ys__n20904, ys__n20906,
    ys__n20908, ys__n20910, ys__n20912, ys__n20914, ys__n20916, ys__n20918,
    ys__n20920, ys__n20922, ys__n20924, ys__n20925, ys__n20926, ys__n20927,
    ys__n20928, ys__n20929, ys__n20930, ys__n20931, ys__n20932, ys__n20933,
    ys__n20934, ys__n20935, ys__n20936, ys__n20937, ys__n20938, ys__n20939,
    ys__n20940, ys__n20941, ys__n20942, ys__n20943, ys__n20944, ys__n20945,
    ys__n20946, ys__n20947, ys__n20948, ys__n20949, ys__n20950, ys__n20951,
    ys__n20952, ys__n20953, ys__n20954, ys__n20955, ys__n20956, ys__n20958,
    ys__n20960, ys__n20962, ys__n20964, ys__n20966, ys__n20968, ys__n20970,
    ys__n20972, ys__n20974, ys__n20976, ys__n20978, ys__n20980, ys__n20982,
    ys__n20984, ys__n20986, ys__n20988, ys__n20990, ys__n20992, ys__n20994,
    ys__n20996, ys__n20998, ys__n21000, ys__n21002, ys__n21004, ys__n21006,
    ys__n21008, ys__n21010, ys__n21012, ys__n21014, ys__n21016, ys__n21018,
    ys__n21020, ys__n21022, ys__n21024, ys__n21026, ys__n21028, ys__n21030,
    ys__n21032, ys__n21034, ys__n21036, ys__n21038, ys__n21040, ys__n21042,
    ys__n21044, ys__n21046, ys__n21048, ys__n21050, ys__n21052, ys__n21054,
    ys__n21056, ys__n21058, ys__n21060, ys__n21062, ys__n21064, ys__n21066,
    ys__n21068, ys__n21070, ys__n21072, ys__n21074, ys__n21076, ys__n21078,
    ys__n21080, ys__n21082, ys__n21084, ys__n21086, ys__n21088, ys__n21090,
    ys__n21092, ys__n21094, ys__n21096, ys__n21098, ys__n21100, ys__n21102,
    ys__n21104, ys__n21106, ys__n21108, ys__n21110, ys__n21112, ys__n21114,
    ys__n21116, ys__n21118, ys__n21120, ys__n21122, ys__n21124, ys__n21126,
    ys__n21128, ys__n21130, ys__n21132, ys__n21134, ys__n21136, ys__n21138,
    ys__n21140, ys__n21142, ys__n21144, ys__n21146, ys__n21148, ys__n21150,
    ys__n21152, ys__n21154, ys__n21156, ys__n21158, ys__n21160, ys__n21162,
    ys__n21164, ys__n21166, ys__n21168, ys__n21170, ys__n21172, ys__n21174,
    ys__n21176, ys__n21178, ys__n21180, ys__n21182, ys__n21184, ys__n21186,
    ys__n21188, ys__n21190, ys__n21192, ys__n21194, ys__n21196, ys__n21198,
    ys__n21200, ys__n21202, ys__n21204, ys__n21206, ys__n21208, ys__n21210,
    ys__n21212, ys__n21214, ys__n21216, ys__n21218, ys__n21220, ys__n21222,
    ys__n21224, ys__n21226, ys__n21228, ys__n21230, ys__n21232, ys__n21234,
    ys__n21236, ys__n21238, ys__n21240, ys__n21242, ys__n21244, ys__n21246,
    ys__n21248, ys__n21250, ys__n21252, ys__n21254, ys__n21256, ys__n21258,
    ys__n21260, ys__n21262, ys__n21264, ys__n21266, ys__n21268, ys__n21270,
    ys__n21272, ys__n21274, ys__n21276, ys__n21278, ys__n21280, ys__n21282,
    ys__n21284, ys__n21286, ys__n21288, ys__n21290, ys__n21292, ys__n21294,
    ys__n21296, ys__n21298, ys__n21300, ys__n21302, ys__n21304, ys__n21306,
    ys__n21308, ys__n21310, ys__n21312, ys__n21314, ys__n21316, ys__n21318,
    ys__n21320, ys__n21322, ys__n21324, ys__n21326, ys__n21328, ys__n21330,
    ys__n21332, ys__n21334, ys__n21336, ys__n21338, ys__n21340, ys__n21342,
    ys__n21344, ys__n21346, ys__n21348, ys__n21350, ys__n21352, ys__n21354,
    ys__n21356, ys__n21358, ys__n21360, ys__n21362, ys__n21364, ys__n21366,
    ys__n21368, ys__n21370, ys__n21372, ys__n21374, ys__n21376, ys__n21378,
    ys__n21380, ys__n21382, ys__n21384, ys__n21386, ys__n21388, ys__n21390,
    ys__n21392, ys__n21394, ys__n21396, ys__n21398, ys__n21400, ys__n21402,
    ys__n21404, ys__n21405, ys__n21406, ys__n21407, ys__n21408, ys__n21409,
    ys__n21410, ys__n21411, ys__n21412, ys__n21413, ys__n21414, ys__n21415,
    ys__n21416, ys__n21417, ys__n21418, ys__n21419, ys__n21420, ys__n21421,
    ys__n21422, ys__n21423, ys__n21424, ys__n21425, ys__n21426, ys__n21427,
    ys__n21428, ys__n21429, ys__n21430, ys__n21431, ys__n21432, ys__n21433,
    ys__n21434, ys__n21435, ys__n21500, ys__n21502, ys__n21504, ys__n21506,
    ys__n21508, ys__n21510, ys__n21512, ys__n21514, ys__n21516, ys__n21518,
    ys__n21520, ys__n21522, ys__n21524, ys__n21526, ys__n21528, ys__n21530,
    ys__n21532, ys__n21534, ys__n21536, ys__n21538, ys__n21540, ys__n21542,
    ys__n21544, ys__n21546, ys__n21548, ys__n21550, ys__n21552, ys__n21554,
    ys__n21556, ys__n21558, ys__n21560, ys__n21562, ys__n21564, ys__n21566,
    ys__n21568, ys__n21570, ys__n21572, ys__n21574, ys__n21576, ys__n21578,
    ys__n21580, ys__n21582, ys__n21584, ys__n21586, ys__n21588, ys__n21590,
    ys__n21592, ys__n21594, ys__n21596, ys__n21598, ys__n21600, ys__n21602,
    ys__n21604, ys__n21606, ys__n21608, ys__n21610, ys__n21612, ys__n21614,
    ys__n21616, ys__n21618, ys__n21620, ys__n21622, ys__n21624, ys__n21626,
    ys__n21628, ys__n21630, ys__n21632, ys__n21634, ys__n21636, ys__n21638,
    ys__n21640, ys__n21642, ys__n21644, ys__n21646, ys__n21648, ys__n21650,
    ys__n21652, ys__n21654, ys__n21656, ys__n21658, ys__n21660, ys__n21662,
    ys__n21664, ys__n21666, ys__n21668, ys__n21670, ys__n21672, ys__n21674,
    ys__n21676, ys__n21678, ys__n21680, ys__n21682, ys__n21684, ys__n21686,
    ys__n21688, ys__n21690, ys__n21692, ys__n21694, ys__n21696, ys__n21698,
    ys__n21700, ys__n21702, ys__n21704, ys__n21706, ys__n21708, ys__n21710,
    ys__n21712, ys__n21714, ys__n21716, ys__n21718, ys__n21720, ys__n21722,
    ys__n21724, ys__n21726, ys__n21728, ys__n21730, ys__n21732, ys__n21734,
    ys__n21736, ys__n21738, ys__n21740, ys__n21742, ys__n21744, ys__n21746,
    ys__n21748, ys__n21750, ys__n21752, ys__n21754, ys__n21756, ys__n21758,
    ys__n21760, ys__n21762, ys__n21764, ys__n21766, ys__n21768, ys__n21770,
    ys__n21772, ys__n21774, ys__n21776, ys__n21778, ys__n21780, ys__n21782,
    ys__n21784, ys__n21786, ys__n21788, ys__n21790, ys__n21792, ys__n21794,
    ys__n21796, ys__n21798, ys__n21800, ys__n21802, ys__n21804, ys__n21806,
    ys__n21808, ys__n21810, ys__n21812, ys__n21814, ys__n21816, ys__n21818,
    ys__n21820, ys__n21822, ys__n21824, ys__n21826, ys__n21828, ys__n21830,
    ys__n21832, ys__n21834, ys__n21836, ys__n21838, ys__n21840, ys__n21842,
    ys__n21844, ys__n21846, ys__n21848, ys__n21850, ys__n21852, ys__n21854,
    ys__n21856, ys__n21858, ys__n21860, ys__n21862, ys__n21864, ys__n21866,
    ys__n21868, ys__n21870, ys__n21872, ys__n21874, ys__n21876, ys__n21878,
    ys__n21880, ys__n21882, ys__n21884, ys__n21886, ys__n21888, ys__n21890,
    ys__n21892, ys__n21894, ys__n21896, ys__n21898, ys__n21900, ys__n21902,
    ys__n21904, ys__n21906, ys__n21908, ys__n21910, ys__n21912, ys__n21914,
    ys__n21916, ys__n21918, ys__n21920, ys__n21922, ys__n21924, ys__n21926,
    ys__n21928, ys__n21930, ys__n21932, ys__n21934, ys__n21936, ys__n21938,
    ys__n21940, ys__n21942, ys__n21944, ys__n21946, ys__n21948, ys__n21949,
    ys__n21950, ys__n21951, ys__n21952, ys__n21953, ys__n21954, ys__n21955,
    ys__n21956, ys__n21957, ys__n21958, ys__n21959, ys__n21960, ys__n21961,
    ys__n21962, ys__n21963, ys__n21964, ys__n21965, ys__n21966, ys__n21967,
    ys__n21968, ys__n21969, ys__n21970, ys__n21971, ys__n21972, ys__n21973,
    ys__n21974, ys__n21975, ys__n21976, ys__n21977, ys__n21978, ys__n21979,
    ys__n21980, ys__n21982, ys__n21984, ys__n21986, ys__n21988, ys__n21990,
    ys__n21992, ys__n21994, ys__n21996, ys__n21998, ys__n22000, ys__n22002,
    ys__n22004, ys__n22006, ys__n22008, ys__n22010, ys__n22012, ys__n22014,
    ys__n22016, ys__n22018, ys__n22020, ys__n22022, ys__n22024, ys__n22026,
    ys__n22028, ys__n22030, ys__n22032, ys__n22034, ys__n22036, ys__n22038,
    ys__n22040, ys__n22042, ys__n22044, ys__n22046, ys__n22048, ys__n22050,
    ys__n22052, ys__n22054, ys__n22056, ys__n22058, ys__n22060, ys__n22062,
    ys__n22064, ys__n22066, ys__n22068, ys__n22070, ys__n22072, ys__n22074,
    ys__n22076, ys__n22078, ys__n22080, ys__n22082, ys__n22084, ys__n22086,
    ys__n22088, ys__n22090, ys__n22092, ys__n22094, ys__n22096, ys__n22098,
    ys__n22100, ys__n22102, ys__n22104, ys__n22106, ys__n22108, ys__n22110,
    ys__n22112, ys__n22114, ys__n22116, ys__n22118, ys__n22120, ys__n22122,
    ys__n22124, ys__n22126, ys__n22128, ys__n22130, ys__n22132, ys__n22134,
    ys__n22136, ys__n22138, ys__n22140, ys__n22142, ys__n22144, ys__n22146,
    ys__n22148, ys__n22150, ys__n22152, ys__n22154, ys__n22156, ys__n22158,
    ys__n22160, ys__n22162, ys__n22164, ys__n22166, ys__n22168, ys__n22170,
    ys__n22172, ys__n22174, ys__n22176, ys__n22178, ys__n22180, ys__n22182,
    ys__n22184, ys__n22186, ys__n22188, ys__n22190, ys__n22192, ys__n22194,
    ys__n22196, ys__n22198, ys__n22200, ys__n22202, ys__n22204, ys__n22206,
    ys__n22208, ys__n22210, ys__n22212, ys__n22214, ys__n22216, ys__n22218,
    ys__n22220, ys__n22222, ys__n22224, ys__n22226, ys__n22228, ys__n22230,
    ys__n22232, ys__n22234, ys__n22236, ys__n22238, ys__n22240, ys__n22242,
    ys__n22244, ys__n22246, ys__n22248, ys__n22250, ys__n22252, ys__n22254,
    ys__n22256, ys__n22258, ys__n22260, ys__n22262, ys__n22264, ys__n22266,
    ys__n22268, ys__n22270, ys__n22272, ys__n22274, ys__n22276, ys__n22278,
    ys__n22280, ys__n22282, ys__n22284, ys__n22286, ys__n22288, ys__n22290,
    ys__n22292, ys__n22294, ys__n22296, ys__n22298, ys__n22300, ys__n22302,
    ys__n22304, ys__n22306, ys__n22308, ys__n22310, ys__n22312, ys__n22314,
    ys__n22316, ys__n22318, ys__n22320, ys__n22322, ys__n22324, ys__n22326,
    ys__n22328, ys__n22330, ys__n22332, ys__n22334, ys__n22336, ys__n22338,
    ys__n22340, ys__n22342, ys__n22344, ys__n22346, ys__n22348, ys__n22350,
    ys__n22352, ys__n22354, ys__n22356, ys__n22358, ys__n22360, ys__n22362,
    ys__n22364, ys__n22366, ys__n22368, ys__n22370, ys__n22372, ys__n22374,
    ys__n22376, ys__n22378, ys__n22380, ys__n22382, ys__n22384, ys__n22386,
    ys__n22388, ys__n22390, ys__n22392, ys__n22394, ys__n22396, ys__n22398,
    ys__n22400, ys__n22402, ys__n22404, ys__n22406, ys__n22408, ys__n22410,
    ys__n22412, ys__n22414, ys__n22416, ys__n22418, ys__n22420, ys__n22422,
    ys__n22424, ys__n22426, ys__n22428, ys__n22429, ys__n22430, ys__n22431,
    ys__n22432, ys__n22433, ys__n22434, ys__n22435, ys__n22436, ys__n22437,
    ys__n22438, ys__n22439, ys__n22440, ys__n22441, ys__n22442, ys__n22443,
    ys__n22444, ys__n22445, ys__n22446, ys__n22447, ys__n22448, ys__n22449,
    ys__n22450, ys__n22451, ys__n22452, ys__n22453, ys__n22454, ys__n22455,
    ys__n22456, ys__n22457, ys__n22458, ys__n22459, ys__n22464, ys__n22465,
    ys__n22564, ys__n22566, ys__n22568, ys__n22570, ys__n22572, ys__n22574,
    ys__n22576, ys__n22578, ys__n22580, ys__n22582, ys__n22584, ys__n22586,
    ys__n22588, ys__n22590, ys__n22592, ys__n22594, ys__n22596, ys__n22598,
    ys__n22600, ys__n22602, ys__n22604, ys__n22606, ys__n22608, ys__n22610,
    ys__n22612, ys__n22614, ys__n22616, ys__n22618, ys__n22620, ys__n22622,
    ys__n22624, ys__n22626, ys__n22630, ys__n22632, ys__n22634, ys__n22636,
    ys__n22640, ys__n22642, ys__n22644, ys__n22646, ys__n22648, ys__n22650,
    ys__n22652, ys__n22654, ys__n22668, ys__n22670, ys__n22673, ys__n22675,
    ys__n22677, ys__n22679, ys__n22681, ys__n22683, ys__n22685, ys__n22687,
    ys__n22689, ys__n22715, ys__n22717, ys__n22719, ys__n22721, ys__n22723,
    ys__n22725, ys__n22727, ys__n22729, ys__n22731, ys__n22733, ys__n22735,
    ys__n22737, ys__n22739, ys__n22741, ys__n22743, ys__n22745, ys__n22747,
    ys__n22749, ys__n22751, ys__n22753, ys__n22755, ys__n22757, ys__n22759,
    ys__n22761, ys__n22763, ys__n22765, ys__n22767, ys__n22769, ys__n22771,
    ys__n22773, ys__n22775, ys__n22777, ys__n22779, ys__n22781, ys__n22783,
    ys__n22785, ys__n22787, ys__n22789, ys__n22792, ys__n22794, ys__n22799,
    ys__n22818, ys__n22820, ys__n22822, ys__n22824, ys__n22826, ys__n22828,
    ys__n22830, ys__n22832, ys__n22834, ys__n22836, ys__n22838, ys__n22840,
    ys__n22842, ys__n22844, ys__n22846, ys__n22848, ys__n22850, ys__n22852,
    ys__n22854, ys__n22856, ys__n22858, ys__n22860, ys__n22862, ys__n22864,
    ys__n22866, ys__n22868, ys__n22870, ys__n22872, ys__n22874, ys__n22876,
    ys__n22878, ys__n22880, ys__n22882, ys__n22884, ys__n22885, ys__n22886,
    ys__n22887, ys__n22888, ys__n22889, ys__n22890, ys__n22891, ys__n22892,
    ys__n22893, ys__n22894, ys__n22895, ys__n22896, ys__n22897, ys__n22898,
    ys__n22899, ys__n22900, ys__n22901, ys__n22902, ys__n22903, ys__n22904,
    ys__n22905, ys__n22906, ys__n22907, ys__n22908, ys__n22909, ys__n22910,
    ys__n22911, ys__n22912, ys__n22913, ys__n22914, ys__n22915, ys__n22916,
    ys__n22918, ys__n22921, ys__n22924, ys__n22927, ys__n22930, ys__n22933,
    ys__n22936, ys__n22939, ys__n22942, ys__n22945, ys__n22948, ys__n22951,
    ys__n22954, ys__n22957, ys__n22960, ys__n22963, ys__n22966, ys__n22969,
    ys__n22972, ys__n22975, ys__n22978, ys__n22981, ys__n22984, ys__n22987,
    ys__n22990, ys__n22993, ys__n22996, ys__n22999, ys__n23002, ys__n23005,
    ys__n23008, ys__n23011, ys__n23014, ys__n23016, ys__n23018, ys__n23020,
    ys__n23022, ys__n23024, ys__n23026, ys__n23028, ys__n23030, ys__n23032,
    ys__n23034, ys__n23036, ys__n23038, ys__n23040, ys__n23042, ys__n23044,
    ys__n23046, ys__n23048, ys__n23050, ys__n23052, ys__n23054, ys__n23056,
    ys__n23058, ys__n23060, ys__n23062, ys__n23064, ys__n23066, ys__n23068,
    ys__n23070, ys__n23072, ys__n23074, ys__n23076, ys__n23077, ys__n23078,
    ys__n23079, ys__n23080, ys__n23081, ys__n23082, ys__n23083, ys__n23084,
    ys__n23085, ys__n23086, ys__n23087, ys__n23088, ys__n23089, ys__n23090,
    ys__n23091, ys__n23092, ys__n23093, ys__n23094, ys__n23095, ys__n23096,
    ys__n23097, ys__n23098, ys__n23099, ys__n23100, ys__n23101, ys__n23102,
    ys__n23103, ys__n23104, ys__n23105, ys__n23106, ys__n23107, ys__n23108,
    ys__n23111, ys__n23114, ys__n23117, ys__n23120, ys__n23123, ys__n23126,
    ys__n23129, ys__n23132, ys__n23135, ys__n23138, ys__n23141, ys__n23144,
    ys__n23147, ys__n23150, ys__n23153, ys__n23156, ys__n23159, ys__n23162,
    ys__n23165, ys__n23168, ys__n23171, ys__n23174, ys__n23177, ys__n23180,
    ys__n23183, ys__n23186, ys__n23189, ys__n23192, ys__n23195, ys__n23198,
    ys__n23203, ys__n23205, ys__n23207, ys__n23209, ys__n23211, ys__n23213,
    ys__n23215, ys__n23217, ys__n23219, ys__n23221, ys__n23223, ys__n23225,
    ys__n23227, ys__n23229, ys__n23231, ys__n23233, ys__n23235, ys__n23237,
    ys__n23239, ys__n23241, ys__n23243, ys__n23245, ys__n23247, ys__n23249,
    ys__n23251, ys__n23253, ys__n23255, ys__n23257, ys__n23259, ys__n23261,
    ys__n23269, ys__n23271, ys__n23272, ys__n23274, ys__n23276, ys__n23278,
    ys__n23280, ys__n23282, ys__n23284, ys__n23286, ys__n23288, ys__n23290,
    ys__n23292, ys__n23294, ys__n23296, ys__n23298, ys__n23300, ys__n23302,
    ys__n23304, ys__n23306, ys__n23308, ys__n23310, ys__n23312, ys__n23314,
    ys__n23316, ys__n23318, ys__n23320, ys__n23322, ys__n23324, ys__n23326,
    ys__n23328, ys__n23330, ys__n23332, ys__n23335, ys__n23339, ys__n23480,
    ys__n23548, ys__n23550, ys__n23552, ys__n23554, ys__n23556, ys__n23558,
    ys__n23560, ys__n23562, ys__n23564, ys__n23566, ys__n23568, ys__n23570,
    ys__n23572, ys__n23574, ys__n23627, ys__n23629, ys__n23641, ys__n23644,
    ys__n23645, ys__n23647, ys__n23650, ys__n23652, ys__n23655, ys__n23658,
    ys__n23661, ys__n23663, ys__n23705, ys__n23706, ys__n23707, ys__n23708,
    ys__n23709, ys__n23710, ys__n23711, ys__n23712, ys__n23713, ys__n23714,
    ys__n23715, ys__n23717, ys__n23729, ys__n23730, ys__n23763, ys__n23818,
    ys__n23819, ys__n23820, ys__n23821, ys__n23822, ys__n23834, ys__n23836,
    ys__n23838, ys__n23840, ys__n23842, ys__n23850, ys__n23888, ys__n23889,
    ys__n23890, ys__n23891, ys__n23892, ys__n23904, ys__n23906, ys__n23908,
    ys__n23910, ys__n23912, ys__n23956, ys__n23957, ys__n23958, ys__n23959,
    ys__n23960, ys__n23977, ys__n23979, ys__n23981, ys__n23983, ys__n23985,
    ys__n24106, ys__n24107, ys__n24108, ys__n24112, ys__n24123, ys__n24124,
    ys__n24131, ys__n24143, ys__n24158, ys__n24167, ys__n24168, ys__n24177,
    ys__n24197, ys__n24199, ys__n24201, ys__n24203, ys__n24205, ys__n24207,
    ys__n24209, ys__n24211, ys__n24213, ys__n24215, ys__n24217, ys__n24219,
    ys__n24228, ys__n24233, ys__n24235, ys__n24243, ys__n24248, ys__n24279,
    ys__n24280, ys__n24303, ys__n24306, ys__n24308, ys__n24310, ys__n24312,
    ys__n24314, ys__n24316, ys__n24318, ys__n24337, ys__n24340, ys__n24342,
    ys__n24344, ys__n24346, ys__n24348, ys__n24350, ys__n24352, ys__n24371,
    ys__n24374, ys__n24376, ys__n24378, ys__n24380, ys__n24382, ys__n24384,
    ys__n24386, ys__n24389, ys__n24406, ys__n24409, ys__n24411, ys__n24413,
    ys__n24415, ys__n24417, ys__n24419, ys__n24421, ys__n24427, ys__n24433,
    ys__n24434, ys__n24461, ys__n24463, ys__n24464, ys__n24483, ys__n24485,
    ys__n24506, ys__n24519, ys__n24567, ys__n24575, ys__n24578, ys__n24590,
    ys__n24591, ys__n24615, ys__n24616, ys__n24617, ys__n24618, ys__n24619,
    ys__n24620, ys__n24621, ys__n24622, ys__n24623, ys__n24624, ys__n24625,
    ys__n24626, ys__n24627, ys__n24628, ys__n24629, ys__n24630, ys__n24631,
    ys__n24632, ys__n24633, ys__n24634, ys__n24635, ys__n24636, ys__n24637,
    ys__n24638, ys__n24639, ys__n24640, ys__n24641, ys__n24642, ys__n24643,
    ys__n24644, ys__n24645, ys__n24646, ys__n24647, ys__n24648, ys__n24649,
    ys__n24650, ys__n24651, ys__n24652, ys__n24653, ys__n24654, ys__n24655,
    ys__n24656, ys__n24657, ys__n24658, ys__n24659, ys__n24660, ys__n24661,
    ys__n24662, ys__n24663, ys__n24664, ys__n24665, ys__n24666, ys__n24667,
    ys__n24668, ys__n24669, ys__n24670, ys__n24671, ys__n24672, ys__n24673,
    ys__n24674, ys__n24675, ys__n24677, ys__n24679, ys__n24681, ys__n24683,
    ys__n24684, ys__n24685, ys__n24686, ys__n24687, ys__n24688, ys__n24689,
    ys__n24690, ys__n24691, ys__n24692, ys__n24693, ys__n24694, ys__n24695,
    ys__n24696, ys__n24697, ys__n24698, ys__n24699, ys__n24700, ys__n24701,
    ys__n24702, ys__n24703, ys__n24704, ys__n24705, ys__n24706, ys__n24707,
    ys__n24708, ys__n24709, ys__n24710, ys__n24711, ys__n24712, ys__n24741,
    ys__n24744, ys__n24747, ys__n24750, ys__n24753, ys__n24756, ys__n24759,
    ys__n24762, ys__n24765, ys__n24768, ys__n24771, ys__n24774, ys__n24777,
    ys__n24780, ys__n24783, ys__n24786, ys__n24789, ys__n24792, ys__n24795,
    ys__n24798, ys__n24801, ys__n24804, ys__n24807, ys__n24810, ys__n24813,
    ys__n24816, ys__n24819, ys__n24822, ys__n24825, ys__n24828, ys__n24831,
    ys__n24834, ys__n25292, ys__n25300, ys__n25381, ys__n25382, ys__n25383,
    ys__n25384, ys__n25470, ys__n25564, ys__n25567, ys__n25570, ys__n25573,
    ys__n25576, ys__n25579, ys__n25582, ys__n25585, ys__n25588, ys__n25591,
    ys__n25594, ys__n25597, ys__n25600, ys__n25603, ys__n25606, ys__n25609,
    ys__n25612, ys__n25615, ys__n25618, ys__n25621, ys__n25624, ys__n25627,
    ys__n25630, ys__n25633, ys__n25636, ys__n25639, ys__n25642, ys__n25645,
    ys__n25648, ys__n25651, ys__n25654, ys__n25657, ys__n25727, ys__n25730,
    ys__n25733, ys__n25736, ys__n25853, ys__n25856, ys__n25859, ys__n25862,
    ys__n25980, ys__n25984, ys__n25987, ys__n25990, ys__n25993, ys__n25996,
    ys__n25999, ys__n26002, ys__n26005, ys__n26008, ys__n26011, ys__n26014,
    ys__n26017, ys__n26020, ys__n26023, ys__n26026, ys__n26029, ys__n26032,
    ys__n26035, ys__n26038, ys__n26041, ys__n26044, ys__n26047, ys__n26050,
    ys__n26053, ys__n26056, ys__n26059, ys__n26062, ys__n26065, ys__n26068,
    ys__n26071, ys__n26074, ys__n26143, ys__n26145, ys__n26147, ys__n26149,
    ys__n26151, ys__n26153, ys__n26155, ys__n26157, ys__n26159, ys__n26161,
    ys__n26162, ys__n26164, ys__n26166, ys__n26168, ys__n26170, ys__n26172,
    ys__n26174, ys__n26176, ys__n26178, ys__n26180, ys__n26182, ys__n26184,
    ys__n26186, ys__n26188, ys__n26190, ys__n26192, ys__n26194, ys__n26196,
    ys__n26198, ys__n26200, ys__n26202, ys__n26204, ys__n26206, ys__n26208,
    ys__n26210, ys__n26212, ys__n26214, ys__n26216, ys__n26218, ys__n26279,
    ys__n26285, ys__n26359, ys__n26362, ys__n26425, ys__n26428, ys__n26431,
    ys__n26434, ys__n26437, ys__n26440, ys__n26443, ys__n26446, ys__n26449,
    ys__n26452, ys__n26455, ys__n26460, ys__n26463, ys__n26466, ys__n26469,
    ys__n26472, ys__n26475, ys__n26478, ys__n26481, ys__n26484, ys__n26487,
    ys__n26490, ys__n26493, ys__n26496, ys__n26499, ys__n26502, ys__n26505,
    ys__n26508, ys__n26511, ys__n26514, ys__n26517, ys__n26552, ys__n26553,
    ys__n26554, ys__n26556, ys__n26557, ys__n26558, ys__n26559, ys__n26560,
    ys__n26561, ys__n26562, ys__n26563, ys__n26564, ys__n26565, ys__n26567,
    ys__n26568, ys__n26569, ys__n26570, ys__n26571, ys__n26572, ys__n26766,
    ys__n26768, ys__n26770, ys__n26772, ys__n27479, ys__n27481, ys__n27485,
    ys__n27488, ys__n27496, ys__n27498, ys__n27499, ys__n27507, ys__n27509,
    ys__n27510, ys__n27518, ys__n27520, ys__n27607, ys__n27608, ys__n27611,
    ys__n27612, ys__n27614, ys__n27615, ys__n27617, ys__n27618, ys__n27620,
    ys__n27621, ys__n27623, ys__n27624, ys__n27626, ys__n27627, ys__n27629,
    ys__n27630, ys__n27632, ys__n27633, ys__n27635, ys__n27636, ys__n27638,
    ys__n27639, ys__n27641, ys__n27642, ys__n27644, ys__n27645, ys__n27647,
    ys__n27648, ys__n27650, ys__n27651, ys__n27653, ys__n27654, ys__n27656,
    ys__n27657, ys__n27659, ys__n27660, ys__n27662, ys__n27663, ys__n27665,
    ys__n27666, ys__n27668, ys__n27669, ys__n27671, ys__n27672, ys__n27674,
    ys__n27675, ys__n27677, ys__n27678, ys__n27680, ys__n27681, ys__n27683,
    ys__n27684, ys__n27686, ys__n27687, ys__n27689, ys__n27690, ys__n27692,
    ys__n27693, ys__n27695, ys__n27696, ys__n27698, ys__n27699, ys__n27701,
    ys__n27702, ys__n27737, ys__n27738, ys__n27740, ys__n27743, ys__n27747,
    ys__n27750, ys__n27753, ys__n27756, ys__n27759, ys__n27762, ys__n27765,
    ys__n27768, ys__n27771, ys__n27774, ys__n27777, ys__n27780, ys__n27783,
    ys__n27786, ys__n27789, ys__n27792, ys__n27795, ys__n27798, ys__n27801,
    ys__n27804, ys__n27807, ys__n27810, ys__n27813, ys__n27816, ys__n27819,
    ys__n27822, ys__n27825, ys__n27828, ys__n27831, ys__n27834, ys__n27837,
    ys__n27855, ys__n27857, ys__n27859, ys__n27861, ys__n27863, ys__n27865,
    ys__n27867, ys__n27869, ys__n27871, ys__n27873, ys__n27875, ys__n27877,
    ys__n27879, ys__n27881, ys__n27883, ys__n27885, ys__n28015, ys__n28016,
    ys__n28017, ys__n28018, ys__n28019, ys__n28020, ys__n28021, ys__n28022,
    ys__n28023, ys__n28024, ys__n28025, ys__n28026, ys__n28027, ys__n28028,
    ys__n28029, ys__n28030, ys__n28243, ys__n28287, ys__n28288, ys__n28290,
    ys__n28292, ys__n28294, ys__n28296, ys__n28424, ys__n28426, ys__n28428,
    ys__n28430, ys__n28432, ys__n28434, ys__n28436, ys__n28438, ys__n28446,
    ys__n28453, ys__n28455, ys__n28457, ys__n28459, ys__n28462, ys__n28464,
    ys__n28466, ys__n28468, ys__n28470, ys__n28472, ys__n28632, ys__n28633,
    ys__n28634, ys__n28635, ys__n28636, ys__n28637, ys__n28638, ys__n28639,
    ys__n28640, ys__n28641, ys__n28718, ys__n28719, ys__n28720, ys__n28859,
    ys__n28863, ys__n28866, ys__n28869, ys__n28872, ys__n28875, ys__n28878,
    ys__n28881, ys__n28884, ys__n28887, ys__n28890, ys__n28893, ys__n28896,
    ys__n28899, ys__n28902, ys__n28905, ys__n28908, ys__n28911, ys__n28914,
    ys__n28917, ys__n28920, ys__n28923, ys__n28926, ys__n28929, ys__n28932,
    ys__n28935, ys__n28938, ys__n28941, ys__n28944, ys__n28947, ys__n28950,
    ys__n28953, ys__n29117, ys__n29119, ys__n29120, ys__n29121, ys__n29123,
    ys__n29124, ys__n29126, ys__n29127, ys__n29129, ys__n29130, ys__n29132,
    ys__n29133, ys__n29135, ys__n29136, ys__n29138, ys__n29139, ys__n29141,
    ys__n29142, ys__n29144, ys__n29145, ys__n29147, ys__n29148, ys__n29150,
    ys__n29151, ys__n29153, ys__n29154, ys__n29156, ys__n29157, ys__n29159,
    ys__n29160, ys__n29162, ys__n29163, ys__n29165, ys__n29166, ys__n29168,
    ys__n29169, ys__n29171, ys__n29172, ys__n29174, ys__n29175, ys__n29177,
    ys__n29178, ys__n29180, ys__n29181, ys__n29183, ys__n29184, ys__n29186,
    ys__n29187, ys__n29189, ys__n29190, ys__n29192, ys__n29193, ys__n29195,
    ys__n29196, ys__n29198, ys__n29199, ys__n29201, ys__n29202, ys__n29204,
    ys__n29205, ys__n29207, ys__n29208, ys__n29210, ys__n29211, ys__n29213,
    ys__n29214, ys__n29218, ys__n29220, ys__n29224, ys__n29237, ys__n29240,
    ys__n29242, ys__n29244, ys__n29246, ys__n29248, ys__n29250, ys__n29252,
    ys__n29254, ys__n29256, ys__n29258, ys__n29260, ys__n29262, ys__n29264,
    ys__n29266, ys__n29268, ys__n29270, ys__n29272, ys__n29274, ys__n29276,
    ys__n29278, ys__n29280, ys__n29282, ys__n29284, ys__n29286, ys__n29288,
    ys__n29290, ys__n29292, ys__n29294, ys__n29296, ys__n29298, ys__n29300,
    ys__n29432, ys__n29433, ys__n29434, ys__n29436, ys__n29437, ys__n29439,
    ys__n29440, ys__n29442, ys__n29443, ys__n29445, ys__n29446, ys__n29448,
    ys__n29449, ys__n29451, ys__n29452, ys__n29454, ys__n29455, ys__n29457,
    ys__n29458, ys__n29460, ys__n29461, ys__n29463, ys__n29464, ys__n29466,
    ys__n29467, ys__n29469, ys__n29470, ys__n29472, ys__n29473, ys__n29475,
    ys__n29476, ys__n29478, ys__n29479, ys__n29481, ys__n29482, ys__n29484,
    ys__n29485, ys__n29487, ys__n29488, ys__n29490, ys__n29491, ys__n29493,
    ys__n29494, ys__n29496, ys__n29497, ys__n29499, ys__n29500, ys__n29502,
    ys__n29503, ys__n29505, ys__n29506, ys__n29508, ys__n29509, ys__n29511,
    ys__n29512, ys__n29514, ys__n29515, ys__n29517, ys__n29518, ys__n29520,
    ys__n29521, ys__n29523, ys__n29524, ys__n29526, ys__n29527, ys__n29531,
    ys__n29533, ys__n29537, ys__n29550, ys__n29552, ys__n29553, ys__n29554,
    ys__n29555, ys__n29556, ys__n29557, ys__n29558, ys__n29559, ys__n29560,
    ys__n29561, ys__n29562, ys__n29563, ys__n29564, ys__n29565, ys__n29566,
    ys__n29567, ys__n29568, ys__n29569, ys__n29570, ys__n29571, ys__n29572,
    ys__n29573, ys__n29574, ys__n29575, ys__n29576, ys__n29577, ys__n29578,
    ys__n29579, ys__n29580, ys__n29581, ys__n29582, ys__n29583, ys__n29584,
    ys__n29585, ys__n29586, ys__n29587, ys__n29588, ys__n29589, ys__n29590,
    ys__n29591, ys__n29592, ys__n29593, ys__n29594, ys__n29595, ys__n29596,
    ys__n29597, ys__n29598, ys__n29599, ys__n29600, ys__n29601, ys__n29602,
    ys__n29603, ys__n29604, ys__n29605, ys__n29606, ys__n29607, ys__n29608,
    ys__n29707, ys__n29708, ys__n29709, ys__n29711, ys__n29712, ys__n29714,
    ys__n29715, ys__n29717, ys__n29718, ys__n29720, ys__n29721, ys__n29723,
    ys__n29724, ys__n29726, ys__n29727, ys__n29729, ys__n29730, ys__n29732,
    ys__n29733, ys__n29735, ys__n29736, ys__n29738, ys__n29739, ys__n29741,
    ys__n29742, ys__n29744, ys__n29745, ys__n29747, ys__n29748, ys__n29750,
    ys__n29751, ys__n29753, ys__n29754, ys__n29756, ys__n29757, ys__n29759,
    ys__n29760, ys__n29762, ys__n29763, ys__n29765, ys__n29766, ys__n29768,
    ys__n29769, ys__n29771, ys__n29772, ys__n29774, ys__n29775, ys__n29777,
    ys__n29778, ys__n29780, ys__n29781, ys__n29783, ys__n29784, ys__n29786,
    ys__n29787, ys__n29789, ys__n29790, ys__n29792, ys__n29793, ys__n29795,
    ys__n29796, ys__n29798, ys__n29799, ys__n29801, ys__n29802, ys__n29806,
    ys__n29808, ys__n29812, ys__n29846, ys__n29880, ys__n29881, ys__n29883,
    ys__n29884, ys__n29885, ys__n29886, ys__n29887, ys__n29888, ys__n29889,
    ys__n29890, ys__n29891, ys__n29892, ys__n29893, ys__n29894, ys__n29895,
    ys__n29896, ys__n29897, ys__n29898, ys__n29899, ys__n29900, ys__n29901,
    ys__n29902, ys__n29903, ys__n29904, ys__n29905, ys__n29906, ys__n29907,
    ys__n29908, ys__n29909, ys__n29910, ys__n29911, ys__n29912, ys__n29913,
    ys__n30011, ys__n30014, ys__n30016, ys__n30018, ys__n30020, ys__n30022,
    ys__n30024, ys__n30026, ys__n30028, ys__n30030, ys__n30032, ys__n30034,
    ys__n30036, ys__n30038, ys__n30040, ys__n30042, ys__n30044, ys__n30046,
    ys__n30048, ys__n30050, ys__n30052, ys__n30054, ys__n30056, ys__n30058,
    ys__n30060, ys__n30062, ys__n30064, ys__n30066, ys__n30068, ys__n30070,
    ys__n30072, ys__n30074, ys__n30214, ys__n30216, ys__n30217, ys__n30219,
    ys__n30220, ys__n30225, ys__n30230, ys__n30232, ys__n30333, ys__n30334,
    ys__n30553, ys__n30815, ys__n30816, ys__n30818, ys__n30819, ys__n30820,
    ys__n30837, ys__n30861, ys__n30862, ys__n30863, ys__n30865, ys__n30867,
    ys__n30869, ys__n30871, ys__n30877, ys__n30879, ys__n30881, ys__n30883,
    ys__n30885, ys__n30887, ys__n30889, ys__n30891, ys__n30893, ys__n30895,
    ys__n30897, ys__n30899, ys__n30901, ys__n30903, ys__n30905, ys__n30907,
    ys__n30909, ys__n30911, ys__n30913, ys__n30915, ys__n30917, ys__n30919,
    ys__n30921, ys__n30923, ys__n30925, ys__n30927, ys__n30929, ys__n30931,
    ys__n30933, ys__n30935, ys__n30937, ys__n30939, ys__n30941, ys__n30957,
    ys__n30960, ys__n30961, ys__n30962, ys__n30974, ys__n31031, ys__n33212,
    ys__n33214, ys__n33216, ys__n33218, ys__n33220, ys__n33222, ys__n33259,
    ys__n33261, ys__n33263, ys__n33265, ys__n33267, ys__n33269, ys__n33272,
    ys__n33274, ys__n33276, ys__n33278, ys__n33300, ys__n33309, ys__n33311,
    ys__n33313, ys__n33318, ys__n33320, ys__n33328, ys__n33330, ys__n33332,
    ys__n33334, ys__n33336, ys__n33338, ys__n33340, ys__n33342, ys__n33350,
    ys__n33352, ys__n33359, ys__n33364, ys__n33370, ys__n33375, ys__n33380,
    ys__n33384, ys__n33386, ys__n33389, ys__n33394, ys__n33396, ys__n33398,
    ys__n33403, ys__n33407, ys__n33409, ys__n33411, ys__n33423, ys__n33431,
    ys__n33442, ys__n33451, ys__n33464, ys__n33469, ys__n33471, ys__n33473,
    ys__n33475, ys__n33479, ys__n33481, ys__n33488, ys__n33491, ys__n33493,
    ys__n33495, ys__n33497, ys__n33499, ys__n33509, ys__n33511, ys__n33522,
    ys__n33532, ys__n33541, ys__n33545, ys__n33548, ys__n33552, ys__n33558,
    ys__n33563, ys__n33564, ys__n33566, ys__n33568, ys__n33570, ys__n33572,
    ys__n33574, ys__n33576, ys__n33579, ys__n33581, ys__n33614, ys__n33632,
    ys__n33634, ys__n33636, ys__n33638, ys__n33640, ys__n33642, ys__n33644,
    ys__n33646, ys__n33648, ys__n33650, ys__n33652, ys__n33654, ys__n33656,
    ys__n33658, ys__n33660, ys__n33662, ys__n33664, ys__n33666, ys__n33668,
    ys__n33670, ys__n33672, ys__n33674, ys__n33676, ys__n33678, ys__n33681,
    ys__n33683, ys__n33685, ys__n33687, ys__n33689, ys__n33691, ys__n33693,
    ys__n33695, ys__n33697, ys__n33699, ys__n33701, ys__n33703, ys__n33705,
    ys__n33707, ys__n33709, ys__n33711, ys__n33713, ys__n33715, ys__n33717,
    ys__n33719, ys__n33721, ys__n33723, ys__n33725, ys__n33727, ys__n33729,
    ys__n33731, ys__n33733, ys__n33735, ys__n33737, ys__n33739, ys__n33741,
    ys__n33743, ys__n33745, ys__n33747, ys__n33749, ys__n34666, ys__n34668,
    ys__n34670, ys__n34672, ys__n34674, ys__n34676, ys__n34678, ys__n34680,
    ys__n34682, ys__n34684, ys__n34686, ys__n34688, ys__n34690, ys__n34692,
    ys__n34694, ys__n34696, ys__n34698, ys__n34700, ys__n34702, ys__n34704,
    ys__n34706, ys__n34708, ys__n34710, ys__n34712, ys__n34714, ys__n34716,
    ys__n34718, ys__n34720, ys__n34722, ys__n34724, ys__n34726, ys__n34728,
    ys__n34730, ys__n34732, ys__n34734, ys__n34736, ys__n34738, ys__n34740,
    ys__n34742, ys__n34744, ys__n34746, ys__n34748, ys__n34750, ys__n34752,
    ys__n34754, ys__n34756, ys__n34758, ys__n34760, ys__n34762, ys__n34764,
    ys__n34766, ys__n34768, ys__n34770, ys__n34772, ys__n34774, ys__n34776,
    ys__n34778, ys__n34780, ys__n34782, ys__n34784, ys__n34786, ys__n34788,
    ys__n34790, ys__n34792, ys__n34794, ys__n34796, ys__n34798, ys__n34800,
    ys__n34802, ys__n34804, ys__n34806, ys__n34808, ys__n34810, ys__n34812,
    ys__n34814, ys__n34816, ys__n34818, ys__n34820, ys__n34822, ys__n34824,
    ys__n34826, ys__n34828, ys__n34830, ys__n34832, ys__n34834, ys__n34836,
    ys__n34838, ys__n34840, ys__n34842, ys__n34844, ys__n34846, ys__n34848,
    ys__n34850, ys__n34852, ys__n34854, ys__n34856, ys__n34858, ys__n34860,
    ys__n34862, ys__n34864, ys__n34866, ys__n34868, ys__n34870, ys__n34872,
    ys__n34874, ys__n34876, ys__n34878, ys__n34880, ys__n34882, ys__n34884,
    ys__n34886, ys__n34888, ys__n34890, ys__n34892, ys__n34894, ys__n34896,
    ys__n34898, ys__n34900, ys__n34902, ys__n34904, ys__n34906, ys__n34908,
    ys__n34910, ys__n34912, ys__n34914, ys__n34916, ys__n34918, ys__n34920,
    ys__n34922, ys__n34924, ys__n34926, ys__n34928, ys__n34930, ys__n34932,
    ys__n34934, ys__n34936, ys__n34938, ys__n34940, ys__n34942, ys__n34944,
    ys__n34946, ys__n34948, ys__n34950, ys__n34959, ys__n34966, ys__n34972,
    ys__n34976, ys__n34978, ys__n34984, ys__n34988, ys__n34990, ys__n34996,
    ys__n35000, ys__n35002, ys__n35008, ys__n35012, ys__n35014, ys__n35020,
    ys__n35024, ys__n35026, ys__n35028, ys__n35031, ys__n35033, ys__n35035,
    ys__n35037, ys__n35039, ys__n35041, ys__n35047, ys__n35049, ys__n35057,
    ys__n35059, ys__n35065, ys__n35076, ys__n35078, ys__n35080, ys__n35082,
    ys__n35084, ys__n35086, ys__n35088, ys__n35090, ys__n35092, ys__n35094,
    ys__n35096, ys__n35098, ys__n35102, ys__n35104, ys__n35106, ys__n35108,
    ys__n35110, ys__n35112, ys__n35114, ys__n35116, ys__n35118, ys__n35120,
    ys__n35122, ys__n35124, ys__n35413, ys__n35415, ys__n35417, ys__n35419,
    ys__n35421, ys__n35423, ys__n35426, ys__n35704, ys__n35717, ys__n35719,
    ys__n35721, ys__n35723, ys__n35725, ys__n35727, ys__n37668, ys__n37669,
    ys__n37670, ys__n37671, ys__n37672, ys__n37673, ys__n37674, ys__n37675,
    ys__n37678, ys__n37679, ys__n37682, ys__n37692, ys__n37694, ys__n37696,
    ys__n37710, ys__n37712, ys__n37713, ys__n37743, ys__n37744, ys__n37745,
    ys__n37746, ys__n37747, ys__n37748, ys__n37749, ys__n37750, ys__n37751,
    ys__n37752, ys__n37753, ys__n37754, ys__n37755, ys__n37756, ys__n37757,
    ys__n37758, ys__n37759, ys__n37760, ys__n37761, ys__n37762, ys__n37763,
    ys__n37764, ys__n37765, ys__n37766, ys__n37767, ys__n37768, ys__n37769,
    ys__n37770, ys__n37771, ys__n37772, ys__n37773, ys__n37774, ys__n37775,
    ys__n37776, ys__n37777, ys__n37778, ys__n37779, ys__n37780, ys__n37781,
    ys__n37782, ys__n37783, ys__n37784, ys__n37785, ys__n37786, ys__n37787,
    ys__n37788, ys__n37789, ys__n37790, ys__n37791, ys__n37792, ys__n37793,
    ys__n37794, ys__n37795, ys__n37796, ys__n37797, ys__n37798, ys__n37799,
    ys__n37800, ys__n37801, ys__n37802, ys__n37803, ys__n37804, ys__n37805,
    ys__n37806, ys__n37807, ys__n37808, ys__n37809, ys__n37810, ys__n37811,
    ys__n37812, ys__n37813, ys__n37814, ys__n37815, ys__n37816, ys__n37817,
    ys__n37818, ys__n37819, ys__n37820, ys__n37821, ys__n37822, ys__n37823,
    ys__n37824, ys__n37825, ys__n37826, ys__n37827, ys__n37828, ys__n37829,
    ys__n37830, ys__n37831, ys__n37832, ys__n37833, ys__n37834, ys__n37835,
    ys__n37836, ys__n37837, ys__n37838, ys__n37839, ys__n37840, ys__n37841,
    ys__n37842, ys__n37843, ys__n37844, ys__n37845, ys__n37846, ys__n37847,
    ys__n37848, ys__n37849, ys__n37850, ys__n37851, ys__n37852, ys__n37853,
    ys__n37854, ys__n37855, ys__n37856, ys__n37857, ys__n37858, ys__n37859,
    ys__n37860, ys__n37861, ys__n37862, ys__n37863, ys__n37864, ys__n37865,
    ys__n37866, ys__n37867, ys__n37868, ys__n37869, ys__n37870, ys__n37871,
    ys__n37872, ys__n37873, ys__n37874, ys__n37875, ys__n37876, ys__n37877,
    ys__n37878, ys__n37879, ys__n37880, ys__n37881, ys__n37882, ys__n37883,
    ys__n37884, ys__n37885, ys__n37886, ys__n37887, ys__n37888, ys__n37889,
    ys__n37890, ys__n37891, ys__n37892, ys__n37893, ys__n37894, ys__n37895,
    ys__n37896, ys__n37897, ys__n37898, ys__n37899, ys__n37900, ys__n37901,
    ys__n37902, ys__n37903, ys__n37904, ys__n37905, ys__n37906, ys__n37907,
    ys__n37908, ys__n37909, ys__n37910, ys__n37911, ys__n37912, ys__n37913,
    ys__n37914, ys__n37915, ys__n37916, ys__n37917, ys__n37918, ys__n37919,
    ys__n37920, ys__n37921, ys__n37922, ys__n37923, ys__n37924, ys__n37925,
    ys__n37926, ys__n37927, ys__n37928, ys__n37929, ys__n37930, ys__n37931,
    ys__n37932, ys__n37933, ys__n37934, ys__n37935, ys__n37936, ys__n37937,
    ys__n37938, ys__n37939, ys__n37940, ys__n37941, ys__n37942, ys__n37943,
    ys__n37944, ys__n37945, ys__n37946, ys__n37947, ys__n37948, ys__n37949,
    ys__n37950, ys__n37951, ys__n37952, ys__n37953, ys__n37954, ys__n37955,
    ys__n37956, ys__n37957, ys__n37958, ys__n37959, ys__n37960, ys__n37961,
    ys__n37962, ys__n37963, ys__n37964, ys__n37965, ys__n37966, ys__n37967,
    ys__n37968, ys__n37969, ys__n37970, ys__n37971, ys__n37972, ys__n37973,
    ys__n37974, ys__n37975, ys__n37976, ys__n37977, ys__n37978, ys__n37979,
    ys__n37980, ys__n37981, ys__n37982, ys__n37983, ys__n37984, ys__n37985,
    ys__n37986, ys__n37987, ys__n37988, ys__n37989, ys__n37990, ys__n37991,
    ys__n37992, ys__n37993, ys__n37994, ys__n37995, ys__n37996, ys__n37997,
    ys__n37998, ys__n37999, ys__n38000, ys__n38001, ys__n38002, ys__n38003,
    ys__n38004, ys__n38005, ys__n38006, ys__n38007, ys__n38008, ys__n38009,
    ys__n38010, ys__n38011, ys__n38012, ys__n38013, ys__n38014, ys__n38015,
    ys__n38016, ys__n38017, ys__n38018, ys__n38019, ys__n38020, ys__n38021,
    ys__n38022, ys__n38023, ys__n38024, ys__n38025, ys__n38026, ys__n38027,
    ys__n38028, ys__n38029, ys__n38030, ys__n38031, ys__n38032, ys__n38033,
    ys__n38034, ys__n38035, ys__n38036, ys__n38037, ys__n38038, ys__n38039,
    ys__n38040, ys__n38041, ys__n38042, ys__n38043, ys__n38044, ys__n38045,
    ys__n38046, ys__n38047, ys__n38048, ys__n38049, ys__n38050, ys__n38051,
    ys__n38052, ys__n38053, ys__n38054, ys__n38055, ys__n38056, ys__n38057,
    ys__n38058, ys__n38059, ys__n38060, ys__n38061, ys__n38062, ys__n38063,
    ys__n38064, ys__n38065, ys__n38066, ys__n38067, ys__n38068, ys__n38069,
    ys__n38070, ys__n38071, ys__n38072, ys__n38073, ys__n38074, ys__n38075,
    ys__n38076, ys__n38077, ys__n38078, ys__n38079, ys__n38080, ys__n38081,
    ys__n38082, ys__n38083, ys__n38084, ys__n38085, ys__n38086, ys__n38087,
    ys__n38088, ys__n38089, ys__n38090, ys__n38091, ys__n38092, ys__n38093,
    ys__n38094, ys__n38095, ys__n38096, ys__n38097, ys__n38098, ys__n38099,
    ys__n38100, ys__n38101, ys__n38102, ys__n38103, ys__n38104, ys__n38105,
    ys__n38106, ys__n38107, ys__n38108, ys__n38109, ys__n38110, ys__n38111,
    ys__n38112, ys__n38113, ys__n38114, ys__n38115, ys__n38116, ys__n38117,
    ys__n38118, ys__n38119, ys__n38120, ys__n38121, ys__n38122, ys__n38123,
    ys__n38124, ys__n38125, ys__n38126, ys__n38127, ys__n38128, ys__n38129,
    ys__n38130, ys__n38131, ys__n38132, ys__n38133, ys__n38134, ys__n38135,
    ys__n38136, ys__n38137, ys__n38138, ys__n38139, ys__n38140, ys__n38141,
    ys__n38142, ys__n38143, ys__n38144, ys__n38145, ys__n38146, ys__n38147,
    ys__n38148, ys__n38149, ys__n38150, ys__n38151, ys__n38152, ys__n38153,
    ys__n38154, ys__n38155, ys__n38156, ys__n38157, ys__n38158, ys__n38159,
    ys__n38160, ys__n38161, ys__n38162, ys__n38163, ys__n38164, ys__n38165,
    ys__n38166, ys__n38167, ys__n38168, ys__n38169, ys__n38170, ys__n38171,
    ys__n38172, ys__n38173, ys__n38174, ys__n38175, ys__n38176, ys__n38177,
    ys__n38178, ys__n38179, ys__n38183, ys__n38192, ys__n38193, ys__n38194,
    ys__n38195, ys__n38196, ys__n38197, ys__n38198, ys__n38199, ys__n38200,
    ys__n38201, ys__n38202, ys__n38203, ys__n38212, ys__n38215, ys__n38217,
    ys__n38219, ys__n38220, ys__n38221, ys__n38236, ys__n38237, ys__n38257,
    ys__n38259, ys__n38272, ys__n38277, ys__n38278, ys__n38279, ys__n38282,
    ys__n38283, ys__n38286, ys__n38288, ys__n38290, ys__n38291, ys__n38300,
    ys__n38304, ys__n38305, ys__n38307, ys__n38311, ys__n38315, ys__n38320,
    ys__n38323, ys__n38346, ys__n38361, ys__n38376, ys__n38378, ys__n38380,
    ys__n38382, ys__n38384, ys__n38386, ys__n38398, ys__n38407, ys__n38408,
    ys__n38413, ys__n38418, ys__n38420, ys__n38424, ys__n38427, ys__n38437,
    ys__n38438, ys__n38441, ys__n38443, ys__n38448, ys__n38449, ys__n38451,
    ys__n38473, ys__n38486, ys__n38487, ys__n38488, ys__n38489, ys__n38490,
    ys__n38491, ys__n38494, ys__n38495, ys__n38496, ys__n38497, ys__n38498,
    ys__n38499, ys__n38502, ys__n38503, ys__n38504, ys__n38505, ys__n38506,
    ys__n38507, ys__n38513, ys__n38522, ys__n38524, ys__n38526, ys__n38527,
    ys__n38528, ys__n38529, ys__n38553, ys__n38557, ys__n38561, ys__n38564,
    ys__n38565, ys__n38567, ys__n38568, ys__n38569, ys__n38585, ys__n38586,
    ys__n38587, ys__n38588, ys__n38589, ys__n38590, ys__n38591, ys__n38592,
    ys__n38593, ys__n38594, ys__n38595, ys__n38596, ys__n38597, ys__n38598,
    ys__n38599, ys__n38600, ys__n38601, ys__n38602, ys__n38603, ys__n38604,
    ys__n38605, ys__n38606, ys__n38607, ys__n38608, ys__n38609, ys__n38610,
    ys__n38611, ys__n38620, ys__n38624, ys__n38631, ys__n38649, ys__n38654,
    ys__n38670, ys__n38680, ys__n38693, ys__n38694, ys__n38695, ys__n38724,
    ys__n38776, ys__n38777, ys__n38805, ys__n38827, ys__n38828, ys__n38829,
    ys__n38830, ys__n38831, ys__n38832, ys__n38833, ys__n38834, ys__n38835,
    ys__n38836, ys__n38837, ys__n38838, ys__n38839, ys__n38840, ys__n38841,
    ys__n38842, ys__n38843, ys__n38844, ys__n38845, ys__n38846, ys__n38847,
    ys__n38848, ys__n38849, ys__n38850, ys__n38851, ys__n38852, ys__n38853,
    ys__n38854, ys__n38855, ys__n38856, ys__n38857, ys__n38858, ys__n38859,
    ys__n38861, ys__n38862, ys__n38863, ys__n38864, ys__n38865, ys__n38883,
    ys__n38885, ys__n38893, ys__n38894, ys__n38896, ys__n38897, ys__n38898,
    ys__n38902, ys__n38904, ys__n38906, ys__n38908, ys__n38910, ys__n38919,
    ys__n38922, ys__n38927, ys__n38928, ys__n38929, ys__n39167, ys__n39518,
    ys__n39520, ys__n39718, ys__n39720, ys__n39722, ys__n39724, ys__n39726,
    ys__n39728, ys__n39730, ys__n39732, ys__n39734, ys__n39736, ys__n39738,
    ys__n39740, ys__n39742, ys__n39744, ys__n39746, ys__n39748, ys__n39750,
    ys__n39752, ys__n39754, ys__n39756, ys__n39758, ys__n39760, ys__n39762,
    ys__n39764, ys__n39766, ys__n39768, ys__n39770, ys__n39772, ys__n39774,
    ys__n39776, ys__n39778, ys__n44833, ys__n44840, ys__n44842, ys__n44847,
    ys__n44849, ys__n44892, ys__n44906, ys__n44907, ys__n44908, ys__n44988,
    ys__n44989, ys__n44990, ys__n44991, ys__n44992, ys__n44993, ys__n44995,
    ys__n44996, ys__n44998, ys__n44999, ys__n45001, ys__n45002, ys__n45004,
    ys__n45005, ys__n45007, ys__n45008, ys__n45010, ys__n45011, ys__n45013,
    ys__n45014, ys__n45016, ys__n45017, ys__n45019, ys__n45020, ys__n45022,
    ys__n45023, ys__n45025, ys__n45026, ys__n45028, ys__n45029, ys__n45031,
    ys__n45032, ys__n45034, ys__n45035, ys__n45037, ys__n45038, ys__n45040,
    ys__n45041, ys__n45043, ys__n45044, ys__n45046, ys__n45047, ys__n45049,
    ys__n45050, ys__n45052, ys__n45053, ys__n45055, ys__n45056, ys__n45058,
    ys__n45059, ys__n45061, ys__n45062, ys__n45064, ys__n45065, ys__n45067,
    ys__n45068, ys__n45070, ys__n45071, ys__n45073, ys__n45074, ys__n45076,
    ys__n45077, ys__n45079, ys__n45080, ys__n45082, ys__n45083, ys__n45084,
    ys__n45085, ys__n45086, ys__n45087, ys__n45088, ys__n45089, ys__n45090,
    ys__n45091, ys__n45092, ys__n45093, ys__n45094, ys__n45095, ys__n45096,
    ys__n45097, ys__n45098, ys__n45099, ys__n45100, ys__n45101, ys__n45102,
    ys__n45103, ys__n45104, ys__n45105, ys__n45106, ys__n45107, ys__n45108,
    ys__n45109, ys__n45110, ys__n45111, ys__n45112, ys__n45113, ys__n45115,
    ys__n45116, ys__n45118, ys__n45119, ys__n45121, ys__n45122, ys__n45124,
    ys__n45125, ys__n45127, ys__n45128, ys__n45130, ys__n45131, ys__n45133,
    ys__n45134, ys__n45136, ys__n45137, ys__n45139, ys__n45140, ys__n45142,
    ys__n45143, ys__n45145, ys__n45146, ys__n45148, ys__n45149, ys__n45151,
    ys__n45152, ys__n45154, ys__n45155, ys__n45157, ys__n45158, ys__n45160,
    ys__n45161, ys__n45163, ys__n45164, ys__n45166, ys__n45167, ys__n45169,
    ys__n45170, ys__n45172, ys__n45173, ys__n45175, ys__n45176, ys__n45178,
    ys__n45179, ys__n45181, ys__n45182, ys__n45184, ys__n45185, ys__n45187,
    ys__n45188, ys__n45190, ys__n45191, ys__n45193, ys__n45194, ys__n45196,
    ys__n45197, ys__n45199, ys__n45200, ys__n45202, ys__n45203, ys__n45205,
    ys__n45206, ys__n45208, ys__n45209, ys__n45210, ys__n45211, ys__n45212,
    ys__n45214, ys__n45216, ys__n45218, ys__n45220, ys__n45222, ys__n45224,
    ys__n45226, ys__n45228, ys__n45230, ys__n45232, ys__n45234, ys__n45236,
    ys__n45238, ys__n45240, ys__n45242, ys__n45244, ys__n45246, ys__n45248,
    ys__n45250, ys__n45252, ys__n45254, ys__n45256, ys__n45258, ys__n45260,
    ys__n45262, ys__n45264, ys__n45266, ys__n45268, ys__n45270, ys__n45272,
    ys__n45274, ys__n45276, ys__n45277, ys__n45278, ys__n45279, ys__n45280,
    ys__n45281, ys__n45282, ys__n45283, ys__n45284, ys__n45285, ys__n45286,
    ys__n45287, ys__n45288, ys__n45289, ys__n45290, ys__n45291, ys__n45292,
    ys__n45293, ys__n45294, ys__n45295, ys__n45296, ys__n45297, ys__n45298,
    ys__n45299, ys__n45300, ys__n45301, ys__n45302, ys__n45303, ys__n45304,
    ys__n45305, ys__n45306, ys__n45308, ys__n45310, ys__n45312, ys__n45314,
    ys__n45316, ys__n45318, ys__n45320, ys__n45322, ys__n45324, ys__n45326,
    ys__n45328, ys__n45330, ys__n45332, ys__n45334, ys__n45336, ys__n45338,
    ys__n45340, ys__n45342, ys__n45344, ys__n45346, ys__n45348, ys__n45350,
    ys__n45352, ys__n45354, ys__n45356, ys__n45358, ys__n45360, ys__n45362,
    ys__n45364, ys__n45366, ys__n45368, ys__n45370, ys__n45371, ys__n45372,
    ys__n45373, ys__n45374, ys__n45377, ys__n45380, ys__n45382, ys__n45384,
    ys__n45386, ys__n45388, ys__n45390, ys__n45392, ys__n45394, ys__n45396,
    ys__n45398, ys__n45400, ys__n45402, ys__n45404, ys__n45406, ys__n45408,
    ys__n45410, ys__n45412, ys__n45414, ys__n45416, ys__n45418, ys__n45420,
    ys__n45422, ys__n45424, ys__n45426, ys__n45428, ys__n45430, ys__n45432,
    ys__n45434, ys__n45436, ys__n45438, ys__n45440, ys__n45441, ys__n45442,
    ys__n45443, ys__n45444, ys__n45445, ys__n45446, ys__n45447, ys__n45448,
    ys__n45449, ys__n45450, ys__n45451, ys__n45452, ys__n45453, ys__n45454,
    ys__n45455, ys__n45456, ys__n45457, ys__n45458, ys__n45459, ys__n45460,
    ys__n45461, ys__n45462, ys__n45463, ys__n45464, ys__n45465, ys__n45466,
    ys__n45467, ys__n45468, ys__n45469, ys__n45470, ys__n45472, ys__n45474,
    ys__n45476, ys__n45478, ys__n45480, ys__n45482, ys__n45484, ys__n45486,
    ys__n45488, ys__n45490, ys__n45492, ys__n45494, ys__n45496, ys__n45498,
    ys__n45500, ys__n45502, ys__n45504, ys__n45506, ys__n45508, ys__n45510,
    ys__n45512, ys__n45514, ys__n45516, ys__n45518, ys__n45520, ys__n45522,
    ys__n45524, ys__n45526, ys__n45528, ys__n45530, ys__n45532, ys__n45534,
    ys__n45535, ys__n45536, ys__n45537, ys__n45538, ys__n45541, ys__n45544,
    ys__n45546, ys__n45548, ys__n45550, ys__n45552, ys__n45554, ys__n45556,
    ys__n45558, ys__n45560, ys__n45562, ys__n45564, ys__n45566, ys__n45568,
    ys__n45570, ys__n45572, ys__n45574, ys__n45576, ys__n45578, ys__n45580,
    ys__n45582, ys__n45584, ys__n45586, ys__n45588, ys__n45590, ys__n45592,
    ys__n45594, ys__n45596, ys__n45598, ys__n45600, ys__n45602, ys__n45604,
    ys__n45605, ys__n45606, ys__n45607, ys__n45608, ys__n45609, ys__n45610,
    ys__n45611, ys__n45612, ys__n45613, ys__n45614, ys__n45615, ys__n45616,
    ys__n45617, ys__n45618, ys__n45619, ys__n45620, ys__n45621, ys__n45622,
    ys__n45623, ys__n45624, ys__n45625, ys__n45626, ys__n45627, ys__n45628,
    ys__n45629, ys__n45630, ys__n45631, ys__n45632, ys__n45633, ys__n45634,
    ys__n45636, ys__n45638, ys__n45640, ys__n45642, ys__n45644, ys__n45646,
    ys__n45648, ys__n45650, ys__n45652, ys__n45654, ys__n45656, ys__n45658,
    ys__n45660, ys__n45662, ys__n45664, ys__n45666, ys__n45668, ys__n45670,
    ys__n45672, ys__n45674, ys__n45676, ys__n45678, ys__n45680, ys__n45682,
    ys__n45684, ys__n45686, ys__n45688, ys__n45690, ys__n45692, ys__n45694,
    ys__n45696, ys__n45698, ys__n45699, ys__n45700, ys__n45701, ys__n45702,
    ys__n45704, ys__n45707, ys__n45708, ys__n45709, ys__n45710, ys__n45711,
    ys__n45712, ys__n45714, ys__n45715, ys__n45717, ys__n45718, ys__n45720,
    ys__n45721, ys__n45723, ys__n45724, ys__n45726, ys__n45727, ys__n45729,
    ys__n45730, ys__n45732, ys__n45733, ys__n45735, ys__n45736, ys__n45738,
    ys__n45739, ys__n45741, ys__n45742, ys__n45744, ys__n45745, ys__n45747,
    ys__n45748, ys__n45750, ys__n45751, ys__n45753, ys__n45754, ys__n45756,
    ys__n45757, ys__n45759, ys__n45760, ys__n45762, ys__n45763, ys__n45765,
    ys__n45766, ys__n45768, ys__n45769, ys__n45771, ys__n45772, ys__n45774,
    ys__n45775, ys__n45777, ys__n45778, ys__n45780, ys__n45781, ys__n45783,
    ys__n45784, ys__n45786, ys__n45787, ys__n45789, ys__n45790, ys__n45792,
    ys__n45793, ys__n45795, ys__n45796, ys__n45798, ys__n45799, ys__n45801,
    ys__n45802, ys__n45804, ys__n45805, ys__n45806, ys__n45807, ys__n45808,
    ys__n45809, ys__n45810, ys__n45811, ys__n45812, ys__n45813, ys__n45814,
    ys__n45815, ys__n45816, ys__n45817, ys__n45818, ys__n45819, ys__n45820,
    ys__n45821, ys__n45822, ys__n45823, ys__n45824, ys__n45825, ys__n45826,
    ys__n45827, ys__n45828, ys__n45829, ys__n45830, ys__n45831, ys__n45832,
    ys__n45833, ys__n45834, ys__n45835, ys__n45836, ys__n45838, ys__n45840,
    ys__n45842, ys__n45844, ys__n45846, ys__n45848, ys__n45850, ys__n45852,
    ys__n45854, ys__n45856, ys__n45858, ys__n45860, ys__n45862, ys__n45864,
    ys__n45866, ys__n45868, ys__n45870, ys__n45872, ys__n45874, ys__n45876,
    ys__n45878, ys__n45880, ys__n45882, ys__n45884, ys__n45886, ys__n45888,
    ys__n45890, ys__n45892, ys__n45894, ys__n45896, ys__n45898, ys__n45900,
    ys__n45901, ys__n45902, ys__n45903, ys__n45904, ys__n45905, ys__n45906,
    ys__n45907, ys__n45908, ys__n45909, ys__n45910, ys__n45911, ys__n45912,
    ys__n45913, ys__n45914, ys__n45915, ys__n45916, ys__n45917, ys__n45918,
    ys__n45919, ys__n45920, ys__n45921, ys__n45922, ys__n45923, ys__n45924,
    ys__n45925, ys__n45926, ys__n45927, ys__n45928, ys__n45929, ys__n45930,
    ys__n45931, ys__n45933, ys__n45936, ys__n45938, ys__n45940, ys__n45942,
    ys__n45944, ys__n45946, ys__n45948, ys__n45950, ys__n45952, ys__n45954,
    ys__n45956, ys__n45958, ys__n45960, ys__n45962, ys__n45964, ys__n45966,
    ys__n45968, ys__n45970, ys__n45972, ys__n45974, ys__n45976, ys__n45978,
    ys__n45980, ys__n45982, ys__n45984, ys__n45986, ys__n45988, ys__n45990,
    ys__n45992, ys__n45994, ys__n45996, ys__n45998, ys__n45999, ys__n46000,
    ys__n46001, ys__n46002, ys__n46003, ys__n46004, ys__n46005, ys__n46006,
    ys__n46007, ys__n46008, ys__n46009, ys__n46010, ys__n46011, ys__n46012,
    ys__n46013, ys__n46014, ys__n46015, ys__n46016, ys__n46017, ys__n46018,
    ys__n46019, ys__n46020, ys__n46021, ys__n46022, ys__n46023, ys__n46024,
    ys__n46025, ys__n46026, ys__n46027, ys__n46028, ys__n46029, ys__n46031,
    ys__n46034, ys__n46036, ys__n46038, ys__n46040, ys__n46042, ys__n46044,
    ys__n46046, ys__n46048, ys__n46050, ys__n46052, ys__n46054, ys__n46056,
    ys__n46058, ys__n46060, ys__n46062, ys__n46064, ys__n46066, ys__n46068,
    ys__n46070, ys__n46072, ys__n46074, ys__n46076, ys__n46078, ys__n46080,
    ys__n46082, ys__n46084, ys__n46086, ys__n46088, ys__n46090, ys__n46092,
    ys__n46094, ys__n46096, ys__n46097, ys__n46098, ys__n46099, ys__n46100,
    ys__n46101, ys__n46102, ys__n46103, ys__n46104, ys__n46105, ys__n46106,
    ys__n46107, ys__n46108, ys__n46109, ys__n46110, ys__n46111, ys__n46112,
    ys__n46113, ys__n46114, ys__n46115, ys__n46116, ys__n46117, ys__n46118,
    ys__n46119, ys__n46120, ys__n46121, ys__n46122, ys__n46123, ys__n46124,
    ys__n46125, ys__n46126, ys__n46127, ys__n46128, ys__n46130, ys__n46132,
    ys__n46134, ys__n46136, ys__n46141, ys__n46142, ys__n46150, ys__n46151,
    ys__n46152, ys__n46153, ys__n46166, ys__n46168, ys__n46169, ys__n46170,
    ys__n46171, ys__n46180, ys__n46184, ys__n46185, ys__n46186, ys__n46187,
    ys__n46198, ys__n46200, ys__n46201, ys__n46202, ys__n46203, ys__n46214,
    ys__n46216, ys__n46217, ys__n46218, ys__n46219, ys__n46230, ys__n46231,
    ys__n46238, ys__n46239, ys__n46240, ys__n46242, ys__n46244, ys__n46245,
    ys__n46247, ys__n46248, ys__n46252, ys__n46254, ys__n46256, ys__n46258,
    ys__n46260, ys__n46262, ys__n46264, ys__n46266, ys__n46268, ys__n46270,
    ys__n46272, ys__n46274, ys__n46276, ys__n46278, ys__n46280, ys__n46282,
    ys__n46284, ys__n46286, ys__n46288, ys__n46290, ys__n46292, ys__n46294,
    ys__n46296, ys__n46298, ys__n46300, ys__n46302, ys__n46304, ys__n46306,
    ys__n46308, ys__n46310, ys__n46312, ys__n46314, ys__n46315, ys__n46316,
    ys__n46317, ys__n46318, ys__n46319, ys__n46320, ys__n46321, ys__n46322,
    ys__n46323, ys__n46324, ys__n46325, ys__n46326, ys__n46327, ys__n46328,
    ys__n46329, ys__n46330, ys__n46331, ys__n46332, ys__n46333, ys__n46334,
    ys__n46335, ys__n46336, ys__n46337, ys__n46338, ys__n46339, ys__n46340,
    ys__n46341, ys__n46342, ys__n46343, ys__n46344, ys__n46345, ys__n46346,
    ys__n46348, ys__n46350, ys__n46352, ys__n46354, ys__n46356, ys__n46358,
    ys__n46360, ys__n46362, ys__n46364, ys__n46366, ys__n46368, ys__n46370,
    ys__n46372, ys__n46374, ys__n46376, ys__n46378, ys__n46380, ys__n46382,
    ys__n46384, ys__n46386, ys__n46388, ys__n46390, ys__n46392, ys__n46393,
    ys__n46394, ys__n46395, ys__n46396, ys__n46397, ys__n46398, ys__n46399,
    ys__n46400, ys__n46401, ys__n46402, ys__n46403, ys__n46404, ys__n46405,
    ys__n46406, ys__n46407, ys__n46408, ys__n46409, ys__n46410, ys__n46411,
    ys__n46412, ys__n46413, ys__n46414, ys__n46415, ys__n46416, ys__n46417,
    ys__n46418, ys__n46419, ys__n46420, ys__n46421, ys__n46422, ys__n46423,
    ys__n46428, ys__n46430, ys__n46432, ys__n46434, ys__n46436, ys__n46438,
    ys__n46440, ys__n46442, ys__n46444, ys__n46446, ys__n46448, ys__n46450,
    ys__n46452, ys__n46454, ys__n46456, ys__n46458, ys__n46460, ys__n46462,
    ys__n46464, ys__n46466, ys__n46468, ys__n46470, ys__n46472, ys__n46474,
    ys__n46476, ys__n46478, ys__n46480, ys__n46482, ys__n46484, ys__n46486,
    ys__n46488, ys__n46490, ys__n46491, ys__n46492, ys__n46493, ys__n46494,
    ys__n46495, ys__n46496, ys__n46497, ys__n46498, ys__n46499, ys__n46500,
    ys__n46501, ys__n46502, ys__n46503, ys__n46504, ys__n46505, ys__n46506,
    ys__n46507, ys__n46508, ys__n46509, ys__n46510, ys__n46511, ys__n46512,
    ys__n46513, ys__n46514, ys__n46515, ys__n46516, ys__n46517, ys__n46518,
    ys__n46519, ys__n46520, ys__n46521, ys__n46522, ys__n46524, ys__n46526,
    ys__n46528, ys__n46530, ys__n46532, ys__n46534, ys__n46536, ys__n46538,
    ys__n46540, ys__n46542, ys__n46544, ys__n46546, ys__n46548, ys__n46550,
    ys__n46552, ys__n46554, ys__n46556, ys__n46558, ys__n46560, ys__n46562,
    ys__n46564, ys__n46566, ys__n46568, ys__n46569, ys__n46570, ys__n46571,
    ys__n46572, ys__n46573, ys__n46574, ys__n46575, ys__n46576, ys__n46577,
    ys__n46578, ys__n46579, ys__n46580, ys__n46581, ys__n46582, ys__n46583,
    ys__n46584, ys__n46585, ys__n46586, ys__n46587, ys__n46588, ys__n46589,
    ys__n46590, ys__n46591, ys__n46592, ys__n46593, ys__n46594, ys__n46595,
    ys__n46596, ys__n46597, ys__n46598, ys__n46599, ys__n46604, ys__n46606,
    ys__n46608, ys__n46610, ys__n46612, ys__n46614, ys__n46616, ys__n46618,
    ys__n46620, ys__n46622, ys__n46624, ys__n46626, ys__n46628, ys__n46630,
    ys__n46632, ys__n46634, ys__n46636, ys__n46638, ys__n46640, ys__n46642,
    ys__n46644, ys__n46646, ys__n46648, ys__n46650, ys__n46652, ys__n46654,
    ys__n46656, ys__n46658, ys__n46660, ys__n46662, ys__n46664, ys__n46666,
    ys__n46667, ys__n46668, ys__n46669, ys__n46670, ys__n46671, ys__n46672,
    ys__n46673, ys__n46674, ys__n46675, ys__n46676, ys__n46677, ys__n46678,
    ys__n46679, ys__n46680, ys__n46681, ys__n46682, ys__n46683, ys__n46684,
    ys__n46685, ys__n46686, ys__n46687, ys__n46688, ys__n46689, ys__n46690,
    ys__n46691, ys__n46692, ys__n46693, ys__n46694, ys__n46695, ys__n46696,
    ys__n46697, ys__n46698, ys__n46700, ys__n46702, ys__n46704, ys__n46706,
    ys__n46708, ys__n46710, ys__n46712, ys__n46714, ys__n46716, ys__n46718,
    ys__n46720, ys__n46722, ys__n46724, ys__n46726, ys__n46728, ys__n46730,
    ys__n46732, ys__n46734, ys__n46736, ys__n46738, ys__n46740, ys__n46742,
    ys__n46744, ys__n46745, ys__n46746, ys__n46747, ys__n46748, ys__n46749,
    ys__n46750, ys__n46751, ys__n46752, ys__n46753, ys__n46754, ys__n46755,
    ys__n46756, ys__n46757, ys__n46758, ys__n46759, ys__n46760, ys__n46761,
    ys__n46762, ys__n46763, ys__n46764, ys__n46765, ys__n46766, ys__n46767,
    ys__n46768, ys__n46769, ys__n46770, ys__n46771, ys__n46772, ys__n46773,
    ys__n46774, ys__n46775, ys__n46780, ys__n46782, ys__n46784, ys__n46786,
    ys__n46788, ys__n46790, ys__n46792, ys__n46794, ys__n46796, ys__n46798,
    ys__n46800, ys__n46802, ys__n46804, ys__n46806, ys__n46808, ys__n46810,
    ys__n46812, ys__n46814, ys__n46816, ys__n46818, ys__n46820, ys__n46822,
    ys__n46824, ys__n46826, ys__n46828, ys__n46830, ys__n46832, ys__n46834,
    ys__n46836, ys__n46838, ys__n46840, ys__n46842, ys__n46843, ys__n46844,
    ys__n46845, ys__n46846, ys__n46847, ys__n46848, ys__n46849, ys__n46850,
    ys__n46851, ys__n46852, ys__n46853, ys__n46854, ys__n46855, ys__n46856,
    ys__n46857, ys__n46858, ys__n46859, ys__n46860, ys__n46861, ys__n46862,
    ys__n46863, ys__n46864, ys__n46865, ys__n46866, ys__n46867, ys__n46868,
    ys__n46869, ys__n46870, ys__n46871, ys__n46872, ys__n46873, ys__n46874,
    ys__n46876, ys__n46878, ys__n46880, ys__n46882, ys__n46884, ys__n46886,
    ys__n46888, ys__n46890, ys__n46892, ys__n46894, ys__n46896, ys__n46898,
    ys__n46900, ys__n46902, ys__n46904, ys__n46906, ys__n46908, ys__n46910,
    ys__n46912, ys__n46914, ys__n46916, ys__n46918, ys__n46920, ys__n46921,
    ys__n46922, ys__n46923, ys__n46924, ys__n46925, ys__n46926, ys__n46927,
    ys__n46928, ys__n46929, ys__n46930, ys__n46931, ys__n46932, ys__n46933,
    ys__n46934, ys__n46935, ys__n46936, ys__n46937, ys__n46938, ys__n46939,
    ys__n46940, ys__n46941, ys__n46942, ys__n46943, ys__n46944, ys__n46945,
    ys__n46946, ys__n46947, ys__n46948, ys__n46949, ys__n46950, ys__n46951,
    ys__n46954, ys__n46955, ys__n46956, ys__n46957, ys__n46958, ys__n46959,
    ys__n46960, ys__n46961, ys__n46962, ys__n46963, ys__n46964, ys__n46965,
    ys__n46966, ys__n46967, ys__n46968, ys__n46969, ys__n46970, ys__n46971,
    ys__n46972, ys__n46973, ys__n46974, ys__n46975, ys__n46976, ys__n46977,
    ys__n46978, ys__n46979, ys__n46980, ys__n46981, ys__n46982, ys__n46983,
    ys__n46984, ys__n46985, ys__n46986, ys__n46987, ys__n46988, ys__n46989,
    ys__n46990, ys__n46991, ys__n46992, ys__n46993, ys__n46994, ys__n46995,
    ys__n46996, ys__n46997, ys__n46998, ys__n46999, ys__n47000, ys__n47001,
    ys__n47002, ys__n47003, ys__n47004, ys__n47005, ys__n47006, ys__n47007,
    ys__n47008, ys__n47009, ys__n47010, ys__n47011, ys__n47012, ys__n47013,
    ys__n47014, ys__n47015, ys__n47016, ys__n47017, ys__n47018, ys__n47019,
    ys__n47020, ys__n47021, ys__n47022, ys__n47023, ys__n47024, ys__n47025,
    ys__n47026, ys__n47027, ys__n47028, ys__n47029, ys__n47030, ys__n47031,
    ys__n47032, ys__n47033, ys__n47034, ys__n47035, ys__n47036, ys__n47037,
    ys__n47038, ys__n47039, ys__n47040, ys__n47041, ys__n47074, ys__n47075,
    ys__n47076, ys__n47077, ys__n47078, ys__n47079, ys__n47080, ys__n47081,
    ys__n47082, ys__n47083, ys__n47084, ys__n47085, ys__n47086, ys__n47087,
    ys__n47088, ys__n47089, ys__n47090, ys__n47091, ys__n47092, ys__n47093,
    ys__n47094, ys__n47095, ys__n47096, ys__n47097, ys__n47098, ys__n47099,
    ys__n47100, ys__n47101, ys__n47102, ys__n47103, ys__n47104, ys__n47105,
    ys__n47106, ys__n47107, ys__n47108, ys__n47109, ys__n47110, ys__n47111,
    ys__n47112, ys__n47113, ys__n47114, ys__n47115, ys__n47116, ys__n47117,
    ys__n47118, ys__n47119, ys__n47184, ys__n47185, ys__n47186, ys__n47187,
    ys__n47188, ys__n47189, ys__n47190, ys__n47191, ys__n47192, ys__n47193,
    ys__n47194, ys__n47195, ys__n47196, ys__n47197, ys__n47198, ys__n47199,
    ys__n47200, ys__n47201, ys__n47202, ys__n47203, ys__n47204, ys__n47205,
    ys__n47206, ys__n47207, ys__n47208, ys__n47209, ys__n47210, ys__n47211,
    ys__n47212, ys__n47213, ys__n47214, ys__n47215, ys__n47216, ys__n47217,
    ys__n47218, ys__n47219, ys__n47220, ys__n47221, ys__n47222, ys__n47223,
    ys__n47224, ys__n47225, ys__n47226, ys__n47227, ys__n47228, ys__n47229,
    ys__n47230, ys__n47231, ys__n47232, ys__n47233, ys__n47234, ys__n47235,
    ys__n47236, ys__n47237, ys__n47238, ys__n47239, ys__n47240, ys__n47241,
    ys__n47242, ys__n47243, ys__n47244, ys__n47245, ys__n47246, ys__n47247,
    ys__n47248, ys__n47249, ys__n47250, ys__n47251, ys__n47252, ys__n47253,
    ys__n47254, ys__n47255, ys__n47256, ys__n47257, ys__n47258, ys__n47259,
    ys__n47260, ys__n47261, ys__n47262, ys__n47263, ys__n47264, ys__n47265,
    ys__n47266, ys__n47267, ys__n47268, ys__n47269, ys__n47270, ys__n47271,
    ys__n47272, ys__n47273, ys__n47274, ys__n47275, ys__n47276, ys__n47277,
    ys__n47278, ys__n47279, ys__n47280, ys__n47281, ys__n47282, ys__n47283,
    ys__n47284, ys__n47285, ys__n47286, ys__n47287, ys__n47288, ys__n47289,
    ys__n47290, ys__n47291, ys__n47292, ys__n47293, ys__n47294, ys__n47295,
    ys__n47296, ys__n47297, ys__n47298, ys__n47299, ys__n47300, ys__n47301,
    ys__n47302, ys__n47303, ys__n47305, ys__n47306, ys__n47307, ys__n47308,
    ys__n47309, ys__n47310, ys__n47311, ys__n47312, ys__n47313, ys__n47314,
    ys__n47315, ys__n47316, ys__n47317, ys__n47318, ys__n47319, ys__n47320,
    ys__n47321, ys__n47322, ys__n47323, ys__n47324, ys__n47325, ys__n47326,
    ys__n47327, ys__n47328, ys__n47329, ys__n47330, ys__n47331, ys__n47332,
    ys__n47333, ys__n47334, ys__n47335, ys__n47336, ys__n47337, ys__n47338,
    ys__n47339, ys__n47340, ys__n47341, ys__n47342, ys__n47343, ys__n47344,
    ys__n47345, ys__n47346, ys__n47347, ys__n47348, ys__n47349, ys__n47350,
    ys__n47351, ys__n47352, ys__n47353, ys__n47354, ys__n47355, ys__n47356,
    ys__n47357, ys__n47358, ys__n47359, ys__n47360, ys__n47361, ys__n47362,
    ys__n47363, ys__n47364, ys__n47365, ys__n47366, ys__n47367, ys__n47368,
    ys__n47369, ys__n47370, ys__n47371, ys__n47372, ys__n47373, ys__n47374,
    ys__n47375, ys__n47376, ys__n47377, ys__n47378, ys__n47379, ys__n47380,
    ys__n47381, ys__n47382, ys__n47383, ys__n47384, ys__n47385, ys__n47386,
    ys__n47387, ys__n47388, ys__n47389, ys__n47390, ys__n47391, ys__n47392,
    ys__n47393, ys__n47394, ys__n47395, ys__n47396, ys__n47397, ys__n47398,
    ys__n47399, ys__n47400, ys__n47401, ys__n47402, ys__n47403, ys__n47404,
    ys__n47405, ys__n47406, ys__n47407, ys__n47408, ys__n47409, ys__n47410,
    ys__n47411, ys__n47412, ys__n47413, ys__n47414, ys__n47415, ys__n47416,
    ys__n47417, ys__n47418, ys__n47419, ys__n47420, ys__n47421, ys__n47422,
    ys__n47423, ys__n47424, ys__n47425, ys__n47426, ys__n47427, ys__n47428,
    ys__n47429, ys__n47430, ys__n47431, ys__n47432, ys__n47433, ys__n47434,
    ys__n47435, ys__n47436, ys__n47437, ys__n47438, ys__n47439, ys__n47440,
    ys__n47441, ys__n47442, ys__n47443, ys__n47444, ys__n47445, ys__n47446,
    ys__n47447, ys__n47448, ys__n47449, ys__n47450, ys__n47451, ys__n47452,
    ys__n47453, ys__n47454, ys__n47455, ys__n47456, ys__n47457, ys__n47458,
    ys__n47459, ys__n47460, ys__n47461, ys__n47462, ys__n47463, ys__n47464,
    ys__n47465, ys__n47466, ys__n47467, ys__n47468, ys__n47469, ys__n47470,
    ys__n47471, ys__n47472, ys__n47473, ys__n47474, ys__n47475, ys__n47476,
    ys__n47477, ys__n47478, ys__n47479, ys__n47480, ys__n47481, ys__n47482,
    ys__n47483, ys__n47484, ys__n47485, ys__n47486, ys__n47487, ys__n47488,
    ys__n47489, ys__n47490, ys__n47491, ys__n47492, ys__n47493, ys__n47494,
    ys__n47495, ys__n47496, ys__n47497, ys__n47498, ys__n47499, ys__n47500,
    ys__n47501, ys__n47502, ys__n47503, ys__n47504, ys__n47505, ys__n47506,
    ys__n47507, ys__n47508, ys__n47509, ys__n47510, ys__n47511, ys__n47512,
    ys__n47513, ys__n47514, ys__n47515, ys__n47516, ys__n47517, ys__n47518,
    ys__n47519, ys__n47520, ys__n47521, ys__n47522, ys__n47523, ys__n47524,
    ys__n47525, ys__n47526, ys__n47527, ys__n47528, ys__n47529, ys__n47530,
    ys__n47531, ys__n47532, ys__n47533, ys__n47534, ys__n47535, ys__n47536,
    ys__n47537, ys__n47538, ys__n47539, ys__n47540, ys__n47541, ys__n47542,
    ys__n47543, ys__n47544, ys__n47545, ys__n47546, ys__n47547, ys__n47548,
    ys__n47549, ys__n47550, ys__n47551, ys__n47552, ys__n47553, ys__n47554,
    ys__n47555, ys__n47556, ys__n47557, ys__n47558, ys__n47559, ys__n47560,
    ys__n47561, ys__n47562, ys__n47563, ys__n47564, ys__n47565, ys__n47566,
    ys__n47567, ys__n47568, ys__n47569, ys__n47570, ys__n47571, ys__n47572,
    ys__n47573, ys__n47574, ys__n47575, ys__n47576, ys__n47577, ys__n47578,
    ys__n47579, ys__n47580, ys__n47581, ys__n47582, ys__n47583, ys__n47584,
    ys__n47585, ys__n47586, ys__n47587, ys__n47588, ys__n47589, ys__n47590,
    ys__n47591, ys__n47592, ys__n47593, ys__n47594, ys__n47595, ys__n47596,
    ys__n47597, ys__n47598, ys__n47599, ys__n47600, ys__n47601, ys__n47602,
    ys__n47603, ys__n47604, ys__n47605, ys__n47606, ys__n47607, ys__n47608,
    ys__n47609, ys__n47610, ys__n47611, ys__n47612, ys__n47613, ys__n47614,
    ys__n47615, ys__n47616, ys__n47617, ys__n47618, ys__n47619, ys__n47620,
    ys__n47621, ys__n47622, ys__n47623, ys__n47624, ys__n47625, ys__n47626,
    ys__n47627, ys__n47628, ys__n47629, ys__n47630, ys__n47631, ys__n47632,
    ys__n47633, ys__n47634, ys__n47635, ys__n47636, ys__n47637, ys__n47638,
    ys__n47639, ys__n47640, ys__n47641, ys__n47642, ys__n47643, ys__n47644,
    ys__n47645, ys__n47646, ys__n47647, ys__n47648, ys__n47649, ys__n47650,
    ys__n47651, ys__n47652, ys__n47653, ys__n47654, ys__n47655, ys__n47656,
    ys__n47657, ys__n47658, ys__n47659, ys__n47660, ys__n47661, ys__n47662,
    ys__n47663, ys__n47664, ys__n47665, ys__n47666, ys__n47667, ys__n47668,
    ys__n47669, ys__n47670, ys__n47671, ys__n47672, ys__n47673, ys__n47674,
    ys__n47675, ys__n47676, ys__n47677, ys__n47678, ys__n47679, ys__n47680,
    ys__n47681, ys__n47682, ys__n47683, ys__n47684, ys__n47685, ys__n47686,
    ys__n47687, ys__n47688, ys__n47689, ys__n47690, ys__n47691, ys__n47692,
    ys__n47693, ys__n47694, ys__n47695, ys__n47696, ys__n47697, ys__n47698,
    ys__n47699, ys__n47700, ys__n47701, ys__n47702, ys__n47703, ys__n47704,
    ys__n47705, ys__n47706, ys__n47707, ys__n47708, ys__n47709, ys__n47710,
    ys__n47711, ys__n47712, ys__n47713, ys__n47714, ys__n47715, ys__n47716,
    ys__n47717, ys__n47718, ys__n47719, ys__n47720, ys__n47721, ys__n47722,
    ys__n47723, ys__n47724, ys__n47725, ys__n47726, ys__n47727, ys__n47728,
    ys__n47729, ys__n47730, ys__n47731, ys__n47732, ys__n47733, ys__n47734,
    ys__n47735, ys__n47736, ys__n47737, ys__n47738, ys__n47739, ys__n47740,
    ys__n47741, ys__n47742, ys__n47743, ys__n47744, ys__n47745, ys__n47746,
    ys__n47747, ys__n47748, ys__n47749, ys__n47750, ys__n47751, ys__n47752,
    ys__n47753, ys__n47754, ys__n47755, ys__n47756, ys__n47757, ys__n47758,
    ys__n47759, ys__n47760, ys__n47761, ys__n47762, ys__n47763, ys__n47764,
    ys__n47765, ys__n47766, ys__n47767, ys__n47768, ys__n47769, ys__n47770,
    ys__n47771, ys__n47772, ys__n47773, ys__n47774, ys__n47775, ys__n47776,
    ys__n47777, ys__n47778, ys__n47779, ys__n47780, ys__n47781, ys__n47782,
    ys__n47783, ys__n47784, ys__n47785, ys__n47786, ys__n47787, ys__n47788,
    ys__n47789, ys__n47790, ys__n47791, ys__n47792, ys__n47793, ys__n47794,
    ys__n47795, ys__n47796, ys__n47797, ys__n47798, ys__n47799, ys__n47800,
    ys__n47801, ys__n47802, ys__n47803, ys__n47804, ys__n47805, ys__n47806,
    ys__n47807, ys__n47808, ys__n47809, ys__n47810, ys__n47811, ys__n47812,
    ys__n47813, ys__n47814, ys__n47815, ys__n47816, ys__n47817, ys__n47818,
    ys__n47819, ys__n47820, ys__n47821, ys__n47822, ys__n47823, ys__n47824,
    ys__n47825, ys__n47826, ys__n47827, ys__n47828, ys__n47829, ys__n47830,
    ys__n47831, ys__n47832, ys__n47833, ys__n47834, ys__n47835, ys__n47836,
    ys__n47837, ys__n47838, ys__n47839, ys__n47840, ys__n47841, ys__n47842,
    ys__n47843, ys__n47844, ys__n47845, ys__n47846, ys__n47847, ys__n47848,
    ys__n47849, ys__n47850, ys__n47851, ys__n47852, ys__n47853, ys__n47854,
    ys__n47855, ys__n47856, ys__n47857, ys__n47858, ys__n47859, ys__n47860,
    ys__n47861, ys__n47862, ys__n47863, ys__n47864, ys__n47865, ys__n47866,
    ys__n47867, ys__n47868, ys__n47869, ys__n47870, ys__n47871, ys__n47872,
    ys__n47873, ys__n47874, ys__n47875, ys__n47876, ys__n47877, ys__n47878,
    ys__n47879, ys__n47880, ys__n47881, ys__n47882, ys__n47883, ys__n47884,
    ys__n47885, ys__n47886, ys__n47887, ys__n47888, ys__n47889, ys__n47890,
    ys__n47891, ys__n47892, ys__n47893, ys__n47894, ys__n47895, ys__n47896,
    ys__n47897, ys__n47898, ys__n47899, ys__n47900, ys__n47901, ys__n47902,
    ys__n47903, ys__n47904, ys__n47905, ys__n47906, ys__n47907, ys__n47908,
    ys__n47909, ys__n47910, ys__n47911, ys__n47912, ys__n47913, ys__n47914,
    ys__n47915, ys__n47916, ys__n47917, ys__n47918, ys__n47919, ys__n47920,
    ys__n47921, ys__n47922, ys__n47923, ys__n47924, ys__n47925, ys__n47926,
    ys__n47927, ys__n47928, ys__n47929, ys__n47930, ys__n47931, ys__n47932,
    ys__n47933, ys__n47934, ys__n47935, ys__n47936, ys__n47937, ys__n47938,
    ys__n47939, ys__n47940, ys__n47941, ys__n47942, ys__n47943, ys__n47944,
    ys__n47945, ys__n47946, ys__n47947, ys__n47948, ys__n47949, ys__n47950,
    ys__n47951, ys__n47952, ys__n47953, ys__n47954, ys__n47955, ys__n47956,
    ys__n47957, ys__n47958, ys__n47959, ys__n47960, ys__n47961, ys__n47962,
    ys__n47963, ys__n47964, ys__n47965, ys__n47966, ys__n47967, ys__n47968,
    ys__n47969, ys__n47970, ys__n47971, ys__n47972, ys__n47973, ys__n47974,
    ys__n47975, ys__n47976, ys__n47977, ys__n47978, ys__n47979, ys__n47980,
    ys__n47981, ys__n47982, ys__n47983, ys__n47984, ys__n47985, ys__n47986,
    ys__n47987, ys__n47988, ys__n47989, ys__n47990, ys__n47991, ys__n47992,
    ys__n47993, ys__n47994, ys__n47995, ys__n47996, ys__n47997, ys__n47998,
    ys__n47999, ys__n48000, ys__n48001, ys__n48002, ys__n48003, ys__n48004,
    ys__n48005, ys__n48006, ys__n48007, ys__n48008, ys__n48009, ys__n48010,
    ys__n48011, ys__n48012, ys__n48013, ys__n48014, ys__n48015, ys__n48016,
    ys__n48017, ys__n48018, ys__n48019, ys__n48020, ys__n48021, ys__n48022,
    ys__n48023, ys__n48024, ys__n48025, ys__n48026, ys__n48027, ys__n48028,
    ys__n48029, ys__n48030, ys__n48031, ys__n48032, ys__n48033, ys__n48034,
    ys__n48035, ys__n48036, ys__n48037, ys__n48038, ys__n48039, ys__n48040,
    ys__n48041, ys__n48042, ys__n48043, ys__n48044, ys__n48045, ys__n48046,
    ys__n48047, ys__n48048, ys__n48049, ys__n48050, ys__n48051, ys__n48052,
    ys__n48053, ys__n48054, ys__n48055, ys__n48056, ys__n48057, ys__n48058,
    ys__n48059, ys__n48060, ys__n48061, ys__n48062, ys__n48063, ys__n48064,
    ys__n48065, ys__n48066, ys__n48067, ys__n48068, ys__n48069, ys__n48070,
    ys__n48071, ys__n48072, ys__n48073, ys__n48074, ys__n48075, ys__n48076,
    ys__n48077, ys__n48078, ys__n48079, ys__n48080, ys__n48081, ys__n48082,
    ys__n48083, ys__n48084, ys__n48085, ys__n48086, ys__n48087, ys__n48088,
    ys__n48089, ys__n48090, ys__n48091, ys__n48092, ys__n48093, ys__n48094,
    ys__n48095, ys__n48096, ys__n48097, ys__n48098, ys__n48099, ys__n48100,
    ys__n48101, ys__n48102, ys__n48103, ys__n48104, ys__n48105, ys__n48106,
    ys__n48107, ys__n48108, ys__n48109, ys__n48110, ys__n48111, ys__n48112,
    ys__n48113, ys__n48114, ys__n48115, ys__n48116, ys__n48117, ys__n48118,
    ys__n48119, ys__n48120, ys__n48121, ys__n48122, ys__n48123, ys__n48124,
    ys__n48125, ys__n48126, ys__n48127, ys__n48128, ys__n48129, ys__n48130,
    ys__n48131, ys__n48132, ys__n48133, ys__n48134, ys__n48135, ys__n48136,
    ys__n48137, ys__n48138, ys__n48139, ys__n48140, ys__n48141, ys__n48142,
    ys__n48143, ys__n48144, ys__n48145, ys__n48146, ys__n48147, ys__n48148,
    ys__n48149, ys__n48150, ys__n48151, ys__n48152, ys__n48153, ys__n48154,
    ys__n48155, ys__n48156, ys__n48157, ys__n48158, ys__n48159, ys__n48160,
    ys__n48161, ys__n48162, ys__n48163, ys__n48164, ys__n48165, ys__n48166,
    ys__n48167, ys__n48168, ys__n48169, ys__n48170, ys__n48171, ys__n48172,
    ys__n48173, ys__n48174, ys__n48175, ys__n48176, ys__n48177, ys__n48178,
    ys__n48179, ys__n48180, ys__n48181, ys__n48182, ys__n48183, ys__n48184,
    ys__n48185, ys__n48186, ys__n48187, ys__n48188, ys__n48189, ys__n48190,
    ys__n48191, ys__n48192, ys__n48193, ys__n48194, ys__n48195, ys__n48196,
    ys__n48197, ys__n48198, ys__n48199, ys__n48200, ys__n48201, ys__n48202,
    ys__n48203, ys__n48204, ys__n48205, ys__n48206, ys__n48207, ys__n48208,
    ys__n48209, ys__n48210, ys__n48211, ys__n48212, ys__n48213, ys__n48214,
    ys__n48215, ys__n48216, ys__n48217, ys__n48218, ys__n48219, ys__n48220,
    ys__n48221, ys__n48222, ys__n48223, ys__n48224, ys__n48225, ys__n48226,
    ys__n48227, ys__n48228, ys__n48229, ys__n48230, ys__n48231, ys__n48232,
    ys__n48233, ys__n48234, ys__n48235, ys__n48236, ys__n48237, ys__n48238,
    ys__n48239, ys__n48240, ys__n48241, ys__n48242, ys__n48243, ys__n48244,
    ys__n48245, ys__n48246, ys__n48247, ys__n48248, ys__n48249, ys__n48250,
    ys__n48251, ys__n48252, ys__n48253, ys__n48254, ys__n48255, ys__n48256,
    ys__n48257, ys__n48258, ys__n48259, ys__n48260, ys__n48261, ys__n48262,
    ys__n48263, ys__n48264, ys__n48265, ys__n48266, ys__n48267, ys__n48268,
    ys__n48269, ys__n48270, ys__n48271, ys__n48272, ys__n48273, ys__n48274,
    ys__n48275, ys__n48324, ys__n48325, ys__n48327, ys__n48330, ys__n48331,
    ys__n48332, ys__n48333, ys__n48334, ys__n48335,
    ys__n2, ys__n246, ys__n250, ys__n252, ys__n254, ys__n264, ys__n270,
    ys__n278, ys__n280, ys__n313, ys__n319, ys__n404, ys__n415, ys__n417,
    ys__n455, ys__n457, ys__n478, ys__n480, ys__n482, ys__n502, ys__n565,
    ys__n574, ys__n576, ys__n628, ys__n630, ys__n714, ys__n716, ys__n730,
    ys__n732, ys__n738, ys__n740, ys__n754, ys__n756, ys__n786, ys__n788,
    ys__n790, ys__n792, ys__n794, ys__n796, ys__n798, ys__n800, ys__n802,
    ys__n804, ys__n806, ys__n808, ys__n810, ys__n812, ys__n814, ys__n862,
    ys__n863, ys__n865, ys__n866, ys__n868, ys__n870, ys__n871, ys__n872,
    ys__n873, ys__n876, ys__n878, ys__n879, ys__n881, ys__n888, ys__n890,
    ys__n900, ys__n902, ys__n904, ys__n911, ys__n920, ys__n923, ys__n927,
    ys__n929, ys__n930, ys__n932, ys__n934, ys__n936, ys__n942, ys__n944,
    ys__n948, ys__n949, ys__n970, ys__n972, ys__n974, ys__n976, ys__n978,
    ys__n980, ys__n982, ys__n989, ys__n991, ys__n993, ys__n995, ys__n999,
    ys__n1001, ys__n1004, ys__n1007, ys__n1009, ys__n1013, ys__n1020,
    ys__n1028, ys__n1030, ys__n1031, ys__n1032, ys__n1037, ys__n1040,
    ys__n1043, ys__n1046, ys__n1047, ys__n1049, ys__n1060, ys__n1071,
    ys__n1073, ys__n1074, ys__n1075, ys__n1077, ys__n1079, ys__n1080,
    ys__n1083, ys__n1085, ys__n1087, ys__n1088, ys__n1089, ys__n1090,
    ys__n1091, ys__n1095, ys__n1103, ys__n1115, ys__n1125, ys__n1128,
    ys__n1135, ys__n1138, ys__n1141, ys__n1142, ys__n1143, ys__n1146,
    ys__n1148, ys__n1161, ys__n1163, ys__n1164, ys__n1165, ys__n1167,
    ys__n1170, ys__n1171, ys__n1183, ys__n1189, ys__n1195, ys__n1201,
    ys__n1207, ys__n1213, ys__n1219, ys__n1222, ys__n1228, ys__n1234,
    ys__n1240, ys__n1246, ys__n1252, ys__n1258, ys__n1261, ys__n1266,
    ys__n1272, ys__n1278, ys__n1284, ys__n1290, ys__n1296, ys__n1303,
    ys__n1377, ys__n1386, ys__n1445, ys__n1448, ys__n1470, ys__n1591,
    ys__n1598, ys__n1601, ys__n1616, ys__n1790, ys__n1802, ys__n1817,
    ys__n1835, ys__n1837, ys__n2152, ys__n2365, ys__n2400, ys__n2423,
    ys__n2491, ys__n2535, ys__n2536, ys__n2582, ys__n2635, ys__n2651,
    ys__n2653, ys__n2655, ys__n2674, ys__n2684, ys__n2733, ys__n2776,
    ys__n2778, ys__n2780, ys__n2782, ys__n2804, ys__n2806, ys__n2845,
    ys__n2855, ys__n3021, ys__n3024, ys__n3035, ys__n3039, ys__n3040,
    ys__n3051, ys__n3061, ys__n3068, ys__n3083, ys__n3085, ys__n3097,
    ys__n3106, ys__n3114, ys__n3115, ys__n3118, ys__n3121, ys__n3195,
    ys__n3249, ys__n3250, ys__n3252, ys__n4175, ys__n4189, ys__n4192,
    ys__n4320, ys__n4414, ys__n4521, ys__n4566, ys__n4588, ys__n4603,
    ys__n4615, ys__n4696, ys__n4764, ys__n4791, ys__n4793, ys__n4798,
    ys__n4817, ys__n4818, ys__n4820, ys__n4821, ys__n4824, ys__n4825,
    ys__n4839, ys__n4840, ys__n12455, ys__n12458, ys__n12461, ys__n12464,
    ys__n12467, ys__n12470, ys__n12473, ys__n12476, ys__n12479, ys__n12482,
    ys__n12485, ys__n12488, ys__n12491, ys__n12494, ys__n12497, ys__n12500,
    ys__n12503, ys__n12506, ys__n12509, ys__n12512, ys__n12515, ys__n12518,
    ys__n12521, ys__n12524, ys__n12527, ys__n12530, ys__n12533, ys__n12536,
    ys__n12539, ys__n12542, ys__n12545, ys__n12548, ys__n16188, ys__n16191,
    ys__n16412, ys__n16415, ys__n16424, ys__n16427, ys__n16706, ys__n16709,
    ys__n16718, ys__n16721, ys__n17692, ys__n17697, ys__n17780, ys__n18007,
    ys__n18009, ys__n18015, ys__n18019, ys__n18028, ys__n18078, ys__n18080,
    ys__n18082, ys__n18087, ys__n18088, ys__n18089, ys__n18120, ys__n18125,
    ys__n18128, ys__n18131, ys__n18133, ys__n18134, ys__n18136, ys__n18137,
    ys__n18154, ys__n18165, ys__n18166, ys__n18169, ys__n18170, ys__n18174,
    ys__n18176, ys__n18178, ys__n18210, ys__n18214, ys__n18216, ys__n18217,
    ys__n18218, ys__n18223, ys__n18227, ys__n18236, ys__n18238, ys__n18239,
    ys__n18241, ys__n18251, ys__n18268, ys__n18272, ys__n18273, ys__n18278,
    ys__n18281, ys__n18284, ys__n18287, ys__n18303, ys__n18321, ys__n18329,
    ys__n18331, ys__n18333, ys__n18335, ys__n18337, ys__n18339, ys__n18341,
    ys__n18343, ys__n18345, ys__n18347, ys__n18349, ys__n18351, ys__n18353,
    ys__n18355, ys__n18357, ys__n18360, ys__n18380, ys__n18383, ys__n18386,
    ys__n18391, ys__n18392, ys__n18394, ys__n18395, ys__n18396, ys__n18397,
    ys__n18398, ys__n18399, ys__n18400, ys__n18401, ys__n18402, ys__n18403,
    ys__n18404, ys__n18405, ys__n18406, ys__n18407, ys__n18408, ys__n18409,
    ys__n18410, ys__n18411, ys__n18412, ys__n18413, ys__n18414, ys__n18415,
    ys__n18416, ys__n18417, ys__n18418, ys__n18419, ys__n18420, ys__n18421,
    ys__n18422, ys__n18423, ys__n18424, ys__n18425, ys__n18426, ys__n18427,
    ys__n18428, ys__n18429, ys__n18430, ys__n18431, ys__n18432, ys__n18433,
    ys__n18434, ys__n18435, ys__n18436, ys__n18437, ys__n18438, ys__n18439,
    ys__n18440, ys__n18441, ys__n18442, ys__n18443, ys__n18444, ys__n18445,
    ys__n18449, ys__n18450, ys__n18452, ys__n18453, ys__n18455, ys__n18456,
    ys__n18458, ys__n18459, ys__n18461, ys__n18462, ys__n18464, ys__n18465,
    ys__n18467, ys__n18468, ys__n18470, ys__n18471, ys__n18473, ys__n18474,
    ys__n18476, ys__n18477, ys__n18479, ys__n18480, ys__n18482, ys__n18483,
    ys__n18485, ys__n18486, ys__n18488, ys__n18489, ys__n18491, ys__n18492,
    ys__n18494, ys__n18495, ys__n18497, ys__n18498, ys__n18500, ys__n18501,
    ys__n18503, ys__n18504, ys__n18506, ys__n18507, ys__n18509, ys__n18510,
    ys__n18512, ys__n18513, ys__n18515, ys__n18516, ys__n18518, ys__n18519,
    ys__n18521, ys__n18522, ys__n18524, ys__n18525, ys__n18527, ys__n18528,
    ys__n18530, ys__n18531, ys__n18533, ys__n18534, ys__n18536, ys__n18537,
    ys__n18539, ys__n18540, ys__n18542, ys__n18543, ys__n18545, ys__n18547,
    ys__n18548, ys__n18549, ys__n18550, ys__n18551, ys__n18553, ys__n18554,
    ys__n18555, ys__n18557, ys__n18559, ys__n18561, ys__n18564, ys__n18567,
    ys__n18570, ys__n18573, ys__n18576, ys__n18579, ys__n18582, ys__n18585,
    ys__n18588, ys__n18591, ys__n18594, ys__n18597, ys__n18600, ys__n18603,
    ys__n18606, ys__n18609, ys__n18612, ys__n18615, ys__n18618, ys__n18621,
    ys__n18624, ys__n18627, ys__n18629, ys__n18631, ys__n18633, ys__n18635,
    ys__n18637, ys__n18640, ys__n18643, ys__n18646, ys__n18649, ys__n18652,
    ys__n18654, ys__n18655, ys__n18657, ys__n18658, ys__n18660, ys__n18661,
    ys__n18663, ys__n18664, ys__n18666, ys__n18667, ys__n18669, ys__n18670,
    ys__n18672, ys__n18673, ys__n18675, ys__n18676, ys__n18678, ys__n18679,
    ys__n18681, ys__n18682, ys__n18684, ys__n18685, ys__n18687, ys__n18688,
    ys__n18690, ys__n18691, ys__n18693, ys__n18694, ys__n18696, ys__n18697,
    ys__n18699, ys__n18700, ys__n18702, ys__n18703, ys__n18705, ys__n18706,
    ys__n18708, ys__n18709, ys__n18711, ys__n18712, ys__n18714, ys__n18715,
    ys__n18717, ys__n18718, ys__n18720, ys__n18721, ys__n18723, ys__n18724,
    ys__n18726, ys__n18727, ys__n18729, ys__n18730, ys__n18732, ys__n18733,
    ys__n18735, ys__n18736, ys__n18738, ys__n18739, ys__n18741, ys__n18742,
    ys__n18744, ys__n18745, ys__n18747, ys__n18748, ys__n18750, ys__n18751,
    ys__n18753, ys__n18754, ys__n18757, ys__n18759, ys__n18760, ys__n18763,
    ys__n18764, ys__n18766, ys__n18768, ys__n18770, ys__n18772, ys__n18774,
    ys__n18776, ys__n18778, ys__n18780, ys__n18782, ys__n18784, ys__n18786,
    ys__n18788, ys__n18790, ys__n18792, ys__n18794, ys__n18796, ys__n18798,
    ys__n18800, ys__n18802, ys__n18804, ys__n18806, ys__n18808, ys__n18810,
    ys__n18812, ys__n18814, ys__n18816, ys__n18818, ys__n18820, ys__n18822,
    ys__n18824, ys__n18826, ys__n19149, ys__n19151, ys__n19159, ys__n19173,
    ys__n19177, ys__n19178, ys__n19183, ys__n19227, ys__n19229, ys__n19231,
    ys__n19233, ys__n19235, ys__n19239, ys__n19254, ys__n19256, ys__n19257,
    ys__n19264, ys__n19266, ys__n19878, ys__n19881, ys__n19884, ys__n19887,
    ys__n19890, ys__n19893, ys__n19896, ys__n19899, ys__n19902, ys__n19905,
    ys__n19908, ys__n19911, ys__n19914, ys__n19917, ys__n19920, ys__n19923,
    ys__n19926, ys__n19929, ys__n19932, ys__n19935, ys__n19938, ys__n19941,
    ys__n19944, ys__n19947, ys__n19950, ys__n19953, ys__n19956, ys__n19959,
    ys__n19962, ys__n19965, ys__n19968, ys__n19971, ys__n20006, ys__n20007,
    ys__n20008, ys__n20009, ys__n20010, ys__n20011, ys__n20012, ys__n20013,
    ys__n20014, ys__n20015, ys__n20016, ys__n20017, ys__n20018, ys__n20019,
    ys__n20020, ys__n20021, ys__n20022, ys__n20023, ys__n20024, ys__n20025,
    ys__n20026, ys__n20027, ys__n20028, ys__n20029, ys__n20030, ys__n20031,
    ys__n20032, ys__n20033, ys__n20034, ys__n20038, ys__n20040, ys__n20043,
    ys__n20045, ys__n20053, ys__n20059, ys__n20062, ys__n20065, ys__n20068,
    ys__n20071, ys__n20074, ys__n20077, ys__n20080, ys__n20082, ys__n20084,
    ys__n20086, ys__n20088, ys__n20090, ys__n20092, ys__n20094, ys__n20096,
    ys__n20098, ys__n20100, ys__n20102, ys__n20104, ys__n20106, ys__n20108,
    ys__n20110, ys__n20112, ys__n20114, ys__n20116, ys__n20118, ys__n20120,
    ys__n20122, ys__n20124, ys__n20126, ys__n20128, ys__n22466, ys__n22919,
    ys__n22922, ys__n22925, ys__n22928, ys__n22931, ys__n22934, ys__n22937,
    ys__n22940, ys__n22943, ys__n22946, ys__n22949, ys__n22952, ys__n22955,
    ys__n22958, ys__n22961, ys__n22964, ys__n22967, ys__n22970, ys__n22973,
    ys__n22976, ys__n22979, ys__n22982, ys__n22985, ys__n22988, ys__n22991,
    ys__n22994, ys__n22997, ys__n23000, ys__n23003, ys__n23006, ys__n23009,
    ys__n23012, ys__n23263, ys__n23264, ys__n23340, ys__n23483, ys__n23485,
    ys__n23487, ys__n23489, ys__n23491, ys__n23493, ys__n23495, ys__n23497,
    ys__n23499, ys__n23501, ys__n23503, ys__n23505, ys__n23507, ys__n23509,
    ys__n23511, ys__n23513, ys__n23515, ys__n23517, ys__n23519, ys__n23521,
    ys__n23523, ys__n23525, ys__n23527, ys__n23529, ys__n23531, ys__n23533,
    ys__n23535, ys__n23537, ys__n23539, ys__n23541, ys__n23543, ys__n23635,
    ys__n23636, ys__n23764, ys__n23795, ys__n23798, ys__n23801, ys__n23804,
    ys__n23807, ys__n23853, ys__n23865, ys__n23868, ys__n23871, ys__n23874,
    ys__n23877, ys__n23921, ys__n23933, ys__n23936, ys__n23939, ys__n23942,
    ys__n23945, ys__n24099, ys__n24101, ys__n24102, ys__n24104, ys__n24105,
    ys__n24116, ys__n24118, ys__n24120, ys__n24126, ys__n24130, ys__n24134,
    ys__n24140, ys__n24145, ys__n24149, ys__n24154, ys__n24160, ys__n24162,
    ys__n24163, ys__n24165, ys__n24166, ys__n24176, ys__n24179, ys__n24180,
    ys__n24182, ys__n24183, ys__n24185, ys__n24186, ys__n24188, ys__n24189,
    ys__n24191, ys__n24192, ys__n24194, ys__n24195, ys__n24222, ys__n24227,
    ys__n24231, ys__n24236, ys__n24240, ys__n24245, ys__n24250, ys__n24255,
    ys__n24256, ys__n24258, ys__n24259, ys__n24260, ys__n24262, ys__n24265,
    ys__n24268, ys__n24271, ys__n24272, ys__n24274, ys__n24275, ys__n24277,
    ys__n24278, ys__n24286, ys__n24289, ys__n24291, ys__n24293, ys__n24295,
    ys__n24297, ys__n24299, ys__n24301, ys__n24305, ys__n24307, ys__n24309,
    ys__n24311, ys__n24313, ys__n24315, ys__n24317, ys__n24319, ys__n24320,
    ys__n24323, ys__n24325, ys__n24327, ys__n24329, ys__n24331, ys__n24333,
    ys__n24335, ys__n24339, ys__n24341, ys__n24343, ys__n24345, ys__n24347,
    ys__n24349, ys__n24351, ys__n24353, ys__n24354, ys__n24357, ys__n24359,
    ys__n24361, ys__n24363, ys__n24365, ys__n24367, ys__n24369, ys__n24373,
    ys__n24375, ys__n24377, ys__n24379, ys__n24381, ys__n24383, ys__n24385,
    ys__n24387, ys__n24388, ys__n24392, ys__n24394, ys__n24396, ys__n24398,
    ys__n24400, ys__n24402, ys__n24404, ys__n24408, ys__n24410, ys__n24412,
    ys__n24414, ys__n24416, ys__n24418, ys__n24420, ys__n24422, ys__n24425,
    ys__n24430, ys__n24436, ys__n24440, ys__n24445, ys__n24447, ys__n24466,
    ys__n24470, ys__n24488, ys__n24499, ys__n24502, ys__n24522, ys__n24532,
    ys__n24541, ys__n24552, ys__n24570, ys__n24573, ys__n24577, ys__n24579,
    ys__n24581, ys__n24585, ys__n24604, ys__n24713, ys__n24714, ys__n24742,
    ys__n24745, ys__n24748, ys__n24751, ys__n24754, ys__n24757, ys__n24760,
    ys__n24763, ys__n24766, ys__n24769, ys__n24772, ys__n24775, ys__n24778,
    ys__n24781, ys__n24784, ys__n24787, ys__n24790, ys__n24793, ys__n24796,
    ys__n24799, ys__n24802, ys__n24805, ys__n24808, ys__n24811, ys__n24814,
    ys__n24817, ys__n24820, ys__n24823, ys__n24826, ys__n24829, ys__n24832,
    ys__n24835, ys__n24837, ys__n24839, ys__n24907, ys__n24910, ys__n24913,
    ys__n24916, ys__n24919, ys__n24922, ys__n24925, ys__n24928, ys__n24931,
    ys__n24934, ys__n24937, ys__n24940, ys__n24943, ys__n24946, ys__n24949,
    ys__n24952, ys__n24955, ys__n25294, ys__n25302, ys__n25304, ys__n25306,
    ys__n25308, ys__n25310, ys__n25385, ys__n25386, ys__n25387, ys__n25388,
    ys__n25390, ys__n25406, ys__n25421, ys__n25430, ys__n25431, ys__n25432,
    ys__n25433, ys__n25434, ys__n25435, ys__n25436, ys__n25438, ys__n25441,
    ys__n25449, ys__n25456, ys__n25461, ys__n25463, ys__n25465, ys__n25467,
    ys__n25469, ys__n25472, ys__n25486, ys__n25496, ys__n25504, ys__n25519,
    ys__n25522, ys__n25534, ys__n25550, ys__n25661, ys__n25663, ys__n25665,
    ys__n25667, ys__n25669, ys__n25671, ys__n25673, ys__n25675, ys__n25677,
    ys__n25679, ys__n25681, ys__n25683, ys__n25685, ys__n25687, ys__n25689,
    ys__n25691, ys__n25693, ys__n25695, ys__n25697, ys__n25699, ys__n25701,
    ys__n25703, ys__n25705, ys__n25707, ys__n25709, ys__n25711, ys__n25713,
    ys__n25715, ys__n25717, ys__n25719, ys__n25721, ys__n25723, ys__n25725,
    ys__n25830, ys__n25833, ys__n25836, ys__n25839, ys__n25842, ys__n25844,
    ys__n25846, ys__n25852, ys__n25957, ys__n25960, ys__n25963, ys__n25966,
    ys__n26118, ys__n26119, ys__n26120, ys__n26121, ys__n26122, ys__n26123,
    ys__n26124, ys__n26125, ys__n26126, ys__n26127, ys__n26128, ys__n26129,
    ys__n26130, ys__n26131, ys__n26132, ys__n26133, ys__n26134, ys__n26135,
    ys__n26136, ys__n26137, ys__n26138, ys__n26139, ys__n26141, ys__n26144,
    ys__n26146, ys__n26148, ys__n26150, ys__n26152, ys__n26154, ys__n26156,
    ys__n26158, ys__n26160, ys__n26220, ys__n26222, ys__n26224, ys__n26226,
    ys__n26228, ys__n26230, ys__n26232, ys__n26234, ys__n26236, ys__n26238,
    ys__n26240, ys__n26242, ys__n26244, ys__n26246, ys__n26248, ys__n26250,
    ys__n26252, ys__n26254, ys__n26256, ys__n26258, ys__n26260, ys__n26262,
    ys__n26264, ys__n26266, ys__n26268, ys__n26270, ys__n26272, ys__n26274,
    ys__n26276, ys__n26278, ys__n26282, ys__n26284, ys__n26286, ys__n26288,
    ys__n26291, ys__n26293, ys__n26294, ys__n26555, ys__n26566, ys__n26573,
    ys__n26607, ys__n26609, ys__n26611, ys__n26613, ys__n26615, ys__n26617,
    ys__n26619, ys__n26621, ys__n26623, ys__n26625, ys__n26627, ys__n26629,
    ys__n26631, ys__n26633, ys__n26635, ys__n26637, ys__n26639, ys__n26641,
    ys__n26643, ys__n26645, ys__n26647, ys__n26649, ys__n26651, ys__n26653,
    ys__n26655, ys__n26657, ys__n26659, ys__n26661, ys__n26663, ys__n26665,
    ys__n26667, ys__n26669, ys__n26671, ys__n26673, ys__n26675, ys__n26677,
    ys__n26679, ys__n26681, ys__n26683, ys__n26685, ys__n26687, ys__n26689,
    ys__n26691, ys__n26693, ys__n26695, ys__n26697, ys__n26699, ys__n26701,
    ys__n26703, ys__n26705, ys__n26707, ys__n26709, ys__n26711, ys__n26713,
    ys__n26715, ys__n26717, ys__n26719, ys__n26721, ys__n26723, ys__n26725,
    ys__n26727, ys__n26729, ys__n26731, ys__n26733, ys__n26734, ys__n26735,
    ys__n26736, ys__n26737, ys__n26738, ys__n26739, ys__n26740, ys__n26741,
    ys__n26742, ys__n26743, ys__n26744, ys__n26745, ys__n26746, ys__n26747,
    ys__n26748, ys__n26749, ys__n26750, ys__n26751, ys__n26752, ys__n26753,
    ys__n26754, ys__n26755, ys__n26756, ys__n26757, ys__n26758, ys__n26759,
    ys__n26760, ys__n26761, ys__n26762, ys__n26763, ys__n26764, ys__n26765,
    ys__n26802, ys__n26803, ys__n26804, ys__n26805, ys__n26806, ys__n26807,
    ys__n26808, ys__n26809, ys__n26810, ys__n26811, ys__n26812, ys__n26813,
    ys__n26814, ys__n26815, ys__n26816, ys__n26817, ys__n26818, ys__n26819,
    ys__n26820, ys__n26821, ys__n26822, ys__n26823, ys__n26824, ys__n26825,
    ys__n26826, ys__n26827, ys__n26828, ys__n26829, ys__n26830, ys__n26831,
    ys__n26832, ys__n26833, ys__n26834, ys__n26835, ys__n26836, ys__n26837,
    ys__n26838, ys__n26839, ys__n26840, ys__n26841, ys__n26842, ys__n26843,
    ys__n26844, ys__n26845, ys__n26846, ys__n26847, ys__n26848, ys__n26849,
    ys__n26850, ys__n26851, ys__n26852, ys__n26853, ys__n26854, ys__n26855,
    ys__n26856, ys__n26857, ys__n26858, ys__n26859, ys__n26860, ys__n26861,
    ys__n26862, ys__n26863, ys__n26864, ys__n26865, ys__n26866, ys__n26867,
    ys__n26868, ys__n26869, ys__n26870, ys__n26871, ys__n26872, ys__n26873,
    ys__n26874, ys__n26875, ys__n26876, ys__n26877, ys__n26878, ys__n26879,
    ys__n26880, ys__n26881, ys__n26882, ys__n26883, ys__n26884, ys__n26885,
    ys__n26886, ys__n26887, ys__n26888, ys__n26889, ys__n26890, ys__n26891,
    ys__n26892, ys__n26893, ys__n26894, ys__n26895, ys__n26896, ys__n26897,
    ys__n26898, ys__n26899, ys__n26900, ys__n26901, ys__n26902, ys__n26903,
    ys__n26904, ys__n26905, ys__n26906, ys__n26907, ys__n26908, ys__n26909,
    ys__n26910, ys__n26911, ys__n26912, ys__n26913, ys__n26914, ys__n26915,
    ys__n26916, ys__n26917, ys__n26918, ys__n26919, ys__n26920, ys__n26921,
    ys__n26922, ys__n26923, ys__n26924, ys__n26925, ys__n26926, ys__n26927,
    ys__n26928, ys__n26929, ys__n26930, ys__n26931, ys__n26932, ys__n26933,
    ys__n26934, ys__n26935, ys__n26936, ys__n26937, ys__n26938, ys__n26939,
    ys__n26940, ys__n26941, ys__n26942, ys__n26943, ys__n26944, ys__n26945,
    ys__n26946, ys__n26947, ys__n26948, ys__n26949, ys__n26950, ys__n26951,
    ys__n26952, ys__n26953, ys__n26954, ys__n26955, ys__n26956, ys__n26957,
    ys__n26958, ys__n26959, ys__n26960, ys__n26961, ys__n26962, ys__n26963,
    ys__n26964, ys__n26965, ys__n26966, ys__n26967, ys__n26968, ys__n26969,
    ys__n26970, ys__n26971, ys__n26972, ys__n26973, ys__n26974, ys__n26975,
    ys__n26976, ys__n26977, ys__n26978, ys__n26979, ys__n26980, ys__n26981,
    ys__n26982, ys__n26983, ys__n26984, ys__n26985, ys__n26986, ys__n26987,
    ys__n26988, ys__n26989, ys__n26990, ys__n26991, ys__n26992, ys__n26993,
    ys__n26994, ys__n26995, ys__n26996, ys__n26997, ys__n26998, ys__n26999,
    ys__n27000, ys__n27001, ys__n27002, ys__n27003, ys__n27004, ys__n27005,
    ys__n27006, ys__n27007, ys__n27008, ys__n27009, ys__n27010, ys__n27011,
    ys__n27012, ys__n27013, ys__n27014, ys__n27015, ys__n27016, ys__n27017,
    ys__n27018, ys__n27019, ys__n27020, ys__n27021, ys__n27022, ys__n27023,
    ys__n27024, ys__n27025, ys__n27026, ys__n27027, ys__n27028, ys__n27029,
    ys__n27030, ys__n27031, ys__n27032, ys__n27033, ys__n27034, ys__n27035,
    ys__n27036, ys__n27037, ys__n27038, ys__n27039, ys__n27040, ys__n27041,
    ys__n27042, ys__n27043, ys__n27044, ys__n27045, ys__n27046, ys__n27047,
    ys__n27048, ys__n27049, ys__n27050, ys__n27051, ys__n27052, ys__n27053,
    ys__n27054, ys__n27055, ys__n27056, ys__n27057, ys__n27058, ys__n27059,
    ys__n27060, ys__n27061, ys__n27062, ys__n27063, ys__n27064, ys__n27065,
    ys__n27066, ys__n27067, ys__n27068, ys__n27069, ys__n27070, ys__n27071,
    ys__n27072, ys__n27073, ys__n27074, ys__n27075, ys__n27076, ys__n27077,
    ys__n27078, ys__n27079, ys__n27080, ys__n27081, ys__n27082, ys__n27083,
    ys__n27084, ys__n27085, ys__n27086, ys__n27087, ys__n27088, ys__n27089,
    ys__n27090, ys__n27091, ys__n27092, ys__n27093, ys__n27094, ys__n27095,
    ys__n27096, ys__n27097, ys__n27098, ys__n27099, ys__n27100, ys__n27101,
    ys__n27102, ys__n27103, ys__n27104, ys__n27105, ys__n27106, ys__n27107,
    ys__n27108, ys__n27109, ys__n27110, ys__n27111, ys__n27112, ys__n27113,
    ys__n27114, ys__n27115, ys__n27116, ys__n27117, ys__n27118, ys__n27119,
    ys__n27120, ys__n27121, ys__n27122, ys__n27123, ys__n27124, ys__n27125,
    ys__n27126, ys__n27127, ys__n27128, ys__n27129, ys__n27130, ys__n27131,
    ys__n27132, ys__n27133, ys__n27134, ys__n27135, ys__n27136, ys__n27137,
    ys__n27138, ys__n27139, ys__n27140, ys__n27141, ys__n27142, ys__n27143,
    ys__n27144, ys__n27145, ys__n27146, ys__n27147, ys__n27148, ys__n27149,
    ys__n27150, ys__n27151, ys__n27152, ys__n27153, ys__n27154, ys__n27155,
    ys__n27156, ys__n27157, ys__n27158, ys__n27159, ys__n27160, ys__n27161,
    ys__n27162, ys__n27163, ys__n27164, ys__n27165, ys__n27166, ys__n27167,
    ys__n27168, ys__n27169, ys__n27170, ys__n27171, ys__n27172, ys__n27173,
    ys__n27174, ys__n27175, ys__n27176, ys__n27177, ys__n27178, ys__n27179,
    ys__n27180, ys__n27181, ys__n27182, ys__n27183, ys__n27184, ys__n27185,
    ys__n27186, ys__n27187, ys__n27188, ys__n27189, ys__n27190, ys__n27191,
    ys__n27192, ys__n27193, ys__n27194, ys__n27195, ys__n27196, ys__n27197,
    ys__n27198, ys__n27199, ys__n27200, ys__n27201, ys__n27202, ys__n27203,
    ys__n27204, ys__n27205, ys__n27206, ys__n27207, ys__n27208, ys__n27209,
    ys__n27210, ys__n27211, ys__n27212, ys__n27213, ys__n27214, ys__n27215,
    ys__n27216, ys__n27217, ys__n27218, ys__n27219, ys__n27220, ys__n27221,
    ys__n27222, ys__n27223, ys__n27224, ys__n27225, ys__n27226, ys__n27227,
    ys__n27228, ys__n27229, ys__n27230, ys__n27231, ys__n27232, ys__n27233,
    ys__n27234, ys__n27235, ys__n27236, ys__n27237, ys__n27238, ys__n27239,
    ys__n27240, ys__n27241, ys__n27242, ys__n27243, ys__n27244, ys__n27245,
    ys__n27246, ys__n27247, ys__n27248, ys__n27249, ys__n27250, ys__n27251,
    ys__n27252, ys__n27253, ys__n27254, ys__n27255, ys__n27256, ys__n27257,
    ys__n27258, ys__n27259, ys__n27260, ys__n27261, ys__n27262, ys__n27263,
    ys__n27264, ys__n27265, ys__n27266, ys__n27267, ys__n27268, ys__n27269,
    ys__n27270, ys__n27271, ys__n27272, ys__n27273, ys__n27274, ys__n27275,
    ys__n27276, ys__n27277, ys__n27278, ys__n27279, ys__n27280, ys__n27281,
    ys__n27282, ys__n27283, ys__n27284, ys__n27285, ys__n27286, ys__n27287,
    ys__n27288, ys__n27289, ys__n27290, ys__n27291, ys__n27292, ys__n27293,
    ys__n27294, ys__n27295, ys__n27296, ys__n27297, ys__n27298, ys__n27299,
    ys__n27300, ys__n27301, ys__n27302, ys__n27303, ys__n27304, ys__n27305,
    ys__n27306, ys__n27307, ys__n27308, ys__n27309, ys__n27310, ys__n27311,
    ys__n27312, ys__n27313, ys__n27314, ys__n27315, ys__n27316, ys__n27317,
    ys__n27318, ys__n27319, ys__n27320, ys__n27321, ys__n27322, ys__n27323,
    ys__n27324, ys__n27325, ys__n27326, ys__n27327, ys__n27328, ys__n27329,
    ys__n27330, ys__n27331, ys__n27332, ys__n27333, ys__n27334, ys__n27335,
    ys__n27336, ys__n27337, ys__n27338, ys__n27339, ys__n27340, ys__n27341,
    ys__n27342, ys__n27343, ys__n27344, ys__n27345, ys__n27346, ys__n27347,
    ys__n27348, ys__n27349, ys__n27350, ys__n27351, ys__n27352, ys__n27353,
    ys__n27354, ys__n27355, ys__n27356, ys__n27357, ys__n27358, ys__n27359,
    ys__n27360, ys__n27361, ys__n27362, ys__n27363, ys__n27364, ys__n27365,
    ys__n27366, ys__n27367, ys__n27368, ys__n27369, ys__n27370, ys__n27371,
    ys__n27372, ys__n27373, ys__n27374, ys__n27375, ys__n27376, ys__n27377,
    ys__n27378, ys__n27379, ys__n27380, ys__n27381, ys__n27382, ys__n27383,
    ys__n27384, ys__n27385, ys__n27386, ys__n27387, ys__n27388, ys__n27389,
    ys__n27390, ys__n27391, ys__n27392, ys__n27393, ys__n27394, ys__n27395,
    ys__n27396, ys__n27397, ys__n27398, ys__n27399, ys__n27400, ys__n27401,
    ys__n27402, ys__n27403, ys__n27404, ys__n27405, ys__n27406, ys__n27407,
    ys__n27408, ys__n27409, ys__n27410, ys__n27411, ys__n27412, ys__n27413,
    ys__n27414, ys__n27415, ys__n27416, ys__n27417, ys__n27418, ys__n27419,
    ys__n27420, ys__n27421, ys__n27422, ys__n27423, ys__n27424, ys__n27425,
    ys__n27426, ys__n27427, ys__n27428, ys__n27429, ys__n27430, ys__n27431,
    ys__n27432, ys__n27433, ys__n27434, ys__n27435, ys__n27436, ys__n27437,
    ys__n27484, ys__n27493, ys__n27504, ys__n27513, ys__n27515, ys__n27517,
    ys__n27550, ys__n27551, ys__n27598, ys__n27603, ys__n27605, ys__n27610,
    ys__n27613, ys__n27616, ys__n27619, ys__n27622, ys__n27625, ys__n27628,
    ys__n27631, ys__n27634, ys__n27637, ys__n27640, ys__n27643, ys__n27646,
    ys__n27649, ys__n27652, ys__n27655, ys__n27658, ys__n27661, ys__n27664,
    ys__n27667, ys__n27670, ys__n27673, ys__n27676, ys__n27679, ys__n27682,
    ys__n27685, ys__n27688, ys__n27691, ys__n27694, ys__n27697, ys__n27700,
    ys__n27703, ys__n27705, ys__n27706, ys__n27707, ys__n27708, ys__n27709,
    ys__n27710, ys__n27711, ys__n27712, ys__n27713, ys__n27714, ys__n27715,
    ys__n27716, ys__n27717, ys__n27718, ys__n27719, ys__n27720, ys__n27721,
    ys__n27722, ys__n27723, ys__n27724, ys__n27725, ys__n27726, ys__n27727,
    ys__n27728, ys__n27729, ys__n27730, ys__n27731, ys__n27732, ys__n27733,
    ys__n27734, ys__n27735, ys__n27736, ys__n27739, ys__n27741, ys__n28247,
    ys__n28249, ys__n28250, ys__n28251, ys__n28252, ys__n28254, ys__n28256,
    ys__n28258, ys__n28259, ys__n28261, ys__n28263, ys__n28265, ys__n28266,
    ys__n28268, ys__n28269, ys__n28270, ys__n28271, ys__n28272, ys__n28274,
    ys__n28276, ys__n28328, ys__n28330, ys__n28332, ys__n28334, ys__n28336,
    ys__n28343, ys__n28345, ys__n28347, ys__n28349, ys__n28351, ys__n28353,
    ys__n28355, ys__n28357, ys__n28359, ys__n28361, ys__n28363, ys__n28365,
    ys__n28367, ys__n28369, ys__n28371, ys__n28373, ys__n28375, ys__n28377,
    ys__n28379, ys__n28381, ys__n28383, ys__n28385, ys__n28387, ys__n28389,
    ys__n28391, ys__n28393, ys__n28395, ys__n28397, ys__n28399, ys__n28401,
    ys__n28403, ys__n28406, ys__n28409, ys__n28410, ys__n28411, ys__n28412,
    ys__n28413, ys__n28414, ys__n28415, ys__n28416, ys__n28417, ys__n28418,
    ys__n28419, ys__n28420, ys__n28421, ys__n28422, ys__n28423, ys__n28425,
    ys__n28427, ys__n28429, ys__n28431, ys__n28433, ys__n28435, ys__n28437,
    ys__n28439, ys__n28440, ys__n28441, ys__n28442, ys__n28443, ys__n28444,
    ys__n28445, ys__n28447, ys__n28448, ys__n28449, ys__n28450, ys__n28451,
    ys__n28452, ys__n28454, ys__n28456, ys__n28458, ys__n28460, ys__n28475,
    ys__n28476, ys__n28477, ys__n28478, ys__n28479, ys__n28480, ys__n28481,
    ys__n28482, ys__n28483, ys__n28484, ys__n28485, ys__n28486, ys__n28487,
    ys__n28488, ys__n28489, ys__n28490, ys__n28491, ys__n28492, ys__n28493,
    ys__n28494, ys__n28495, ys__n28496, ys__n28497, ys__n28498, ys__n28499,
    ys__n28500, ys__n28501, ys__n28502, ys__n28503, ys__n28504, ys__n28505,
    ys__n28506, ys__n28510, ys__n28513, ys__n28518, ys__n28533, ys__n28536,
    ys__n28539, ys__n28542, ys__n28545, ys__n28548, ys__n28551, ys__n28554,
    ys__n28557, ys__n28560, ys__n28563, ys__n28566, ys__n28569, ys__n28572,
    ys__n28575, ys__n28578, ys__n28581, ys__n28584, ys__n28587, ys__n28661,
    ys__n28662, ys__n28781, ys__n28782, ys__n28783, ys__n28784, ys__n28785,
    ys__n28786, ys__n28787, ys__n28788, ys__n28789, ys__n28790, ys__n28791,
    ys__n28792, ys__n28793, ys__n28794, ys__n28796, ys__n28798, ys__n28800,
    ys__n28802, ys__n28804, ys__n28806, ys__n28808, ys__n28810, ys__n28812,
    ys__n28814, ys__n28816, ys__n28818, ys__n28820, ys__n28822, ys__n28824,
    ys__n28826, ys__n28828, ys__n28830, ys__n28832, ys__n28834, ys__n28836,
    ys__n28838, ys__n28840, ys__n28842, ys__n28844, ys__n28846, ys__n28848,
    ys__n28850, ys__n28852, ys__n28854, ys__n28856, ys__n28858, ys__n29022,
    ys__n29025, ys__n29028, ys__n29031, ys__n29034, ys__n29037, ys__n29040,
    ys__n29043, ys__n29046, ys__n29049, ys__n29052, ys__n29055, ys__n29058,
    ys__n29061, ys__n29064, ys__n29067, ys__n29070, ys__n29073, ys__n29076,
    ys__n29079, ys__n29082, ys__n29085, ys__n29088, ys__n29091, ys__n29094,
    ys__n29097, ys__n29100, ys__n29103, ys__n29106, ys__n29109, ys__n29112,
    ys__n29115, ys__n29118, ys__n29122, ys__n29125, ys__n29128, ys__n29131,
    ys__n29134, ys__n29137, ys__n29140, ys__n29143, ys__n29146, ys__n29149,
    ys__n29152, ys__n29155, ys__n29158, ys__n29161, ys__n29164, ys__n29167,
    ys__n29170, ys__n29173, ys__n29176, ys__n29179, ys__n29182, ys__n29185,
    ys__n29188, ys__n29191, ys__n29194, ys__n29197, ys__n29200, ys__n29203,
    ys__n29206, ys__n29209, ys__n29212, ys__n29215, ys__n29217, ys__n29219,
    ys__n29221, ys__n29223, ys__n29225, ys__n29226, ys__n29227, ys__n29228,
    ys__n29229, ys__n29230, ys__n29231, ys__n29232, ys__n29233, ys__n29234,
    ys__n29235, ys__n29336, ys__n29339, ys__n29342, ys__n29345, ys__n29348,
    ys__n29351, ys__n29354, ys__n29357, ys__n29360, ys__n29363, ys__n29366,
    ys__n29369, ys__n29372, ys__n29375, ys__n29378, ys__n29381, ys__n29384,
    ys__n29387, ys__n29390, ys__n29393, ys__n29396, ys__n29399, ys__n29402,
    ys__n29405, ys__n29408, ys__n29411, ys__n29414, ys__n29417, ys__n29420,
    ys__n29423, ys__n29426, ys__n29429, ys__n29431, ys__n29435, ys__n29438,
    ys__n29441, ys__n29444, ys__n29447, ys__n29450, ys__n29453, ys__n29456,
    ys__n29459, ys__n29462, ys__n29465, ys__n29468, ys__n29471, ys__n29474,
    ys__n29477, ys__n29480, ys__n29483, ys__n29486, ys__n29489, ys__n29492,
    ys__n29495, ys__n29498, ys__n29501, ys__n29504, ys__n29507, ys__n29510,
    ys__n29513, ys__n29516, ys__n29519, ys__n29522, ys__n29525, ys__n29528,
    ys__n29530, ys__n29532, ys__n29534, ys__n29536, ys__n29538, ys__n29539,
    ys__n29540, ys__n29541, ys__n29542, ys__n29543, ys__n29544, ys__n29545,
    ys__n29546, ys__n29547, ys__n29548, ys__n29611, ys__n29614, ys__n29617,
    ys__n29620, ys__n29623, ys__n29626, ys__n29629, ys__n29632, ys__n29635,
    ys__n29638, ys__n29641, ys__n29644, ys__n29647, ys__n29650, ys__n29653,
    ys__n29656, ys__n29659, ys__n29662, ys__n29665, ys__n29668, ys__n29671,
    ys__n29674, ys__n29677, ys__n29680, ys__n29683, ys__n29686, ys__n29689,
    ys__n29692, ys__n29695, ys__n29698, ys__n29701, ys__n29704, ys__n29706,
    ys__n29710, ys__n29713, ys__n29716, ys__n29719, ys__n29722, ys__n29725,
    ys__n29728, ys__n29731, ys__n29734, ys__n29737, ys__n29740, ys__n29743,
    ys__n29746, ys__n29749, ys__n29752, ys__n29755, ys__n29758, ys__n29761,
    ys__n29764, ys__n29767, ys__n29770, ys__n29773, ys__n29776, ys__n29779,
    ys__n29782, ys__n29785, ys__n29788, ys__n29791, ys__n29794, ys__n29797,
    ys__n29800, ys__n29803, ys__n29805, ys__n29807, ys__n29809, ys__n29811,
    ys__n29813, ys__n29814, ys__n29815, ys__n29816, ys__n29817, ys__n29818,
    ys__n29819, ys__n29820, ys__n29821, ys__n29822, ys__n29823, ys__n29847,
    ys__n30010, ys__n30080, ys__n30081, ys__n30082, ys__n30083, ys__n30084,
    ys__n30085, ys__n30086, ys__n30087, ys__n30089, ys__n30090, ys__n30091,
    ys__n30092, ys__n30093, ys__n30094, ys__n30095, ys__n30096, ys__n30098,
    ys__n30099, ys__n30100, ys__n30101, ys__n30102, ys__n30103, ys__n30104,
    ys__n30105, ys__n30106, ys__n30107, ys__n30108, ys__n30109, ys__n30110,
    ys__n30111, ys__n30112, ys__n30113, ys__n30119, ys__n30122, ys__n30125,
    ys__n30128, ys__n30131, ys__n30134, ys__n30137, ys__n30140, ys__n30143,
    ys__n30146, ys__n30149, ys__n30152, ys__n30155, ys__n30158, ys__n30161,
    ys__n30164, ys__n30167, ys__n30170, ys__n30173, ys__n30176, ys__n30179,
    ys__n30182, ys__n30185, ys__n30188, ys__n30191, ys__n30194, ys__n30197,
    ys__n30200, ys__n30203, ys__n30206, ys__n30209, ys__n30212, ys__n30215,
    ys__n30223, ys__n30226, ys__n30235, ys__n30238, ys__n30241, ys__n30244,
    ys__n30247, ys__n30250, ys__n30253, ys__n30256, ys__n30259, ys__n30262,
    ys__n30265, ys__n30268, ys__n30271, ys__n30274, ys__n30277, ys__n30280,
    ys__n30283, ys__n30286, ys__n30289, ys__n30292, ys__n30295, ys__n30298,
    ys__n30301, ys__n30304, ys__n30307, ys__n30310, ys__n30313, ys__n30316,
    ys__n30319, ys__n30322, ys__n30325, ys__n30328, ys__n30330, ys__n30331,
    ys__n30616, ys__n30619, ys__n30622, ys__n30625, ys__n30628, ys__n30631,
    ys__n30634, ys__n30637, ys__n30640, ys__n30643, ys__n30646, ys__n30649,
    ys__n30652, ys__n30655, ys__n30658, ys__n30661, ys__n30664, ys__n30667,
    ys__n30668, ys__n30670, ys__n30797, ys__n30798, ys__n30799, ys__n30800,
    ys__n30801, ys__n30802, ys__n30803, ys__n30804, ys__n30805, ys__n30806,
    ys__n30807, ys__n30808, ys__n30809, ys__n30810, ys__n30811, ys__n30812,
    ys__n30813, ys__n30832, ys__n30833, ys__n30835, ys__n30836, ys__n30856,
    ys__n30858, ys__n30860, ys__n30864, ys__n30873, ys__n30874, ys__n30875,
    ys__n30876, ys__n30942, ys__n30943, ys__n30944, ys__n30945, ys__n30946,
    ys__n30947, ys__n30948, ys__n30949, ys__n30950, ys__n30951, ys__n30952,
    ys__n30953, ys__n30954, ys__n30955, ys__n30956, ys__n31202, ys__n31203,
    ys__n31207, ys__n31208, ys__n31209, ys__n31210, ys__n31211, ys__n31212,
    ys__n31213, ys__n31214, ys__n31215, ys__n31216, ys__n31217, ys__n31218,
    ys__n31219, ys__n31220, ys__n31221, ys__n31222, ys__n31223, ys__n31224,
    ys__n31225, ys__n31226, ys__n31227, ys__n31228, ys__n31229, ys__n31230,
    ys__n31231, ys__n31232, ys__n31233, ys__n31234, ys__n31235, ys__n31236,
    ys__n31237, ys__n31238, ys__n31326, ys__n31327, ys__n31328, ys__n31329,
    ys__n31330, ys__n31331, ys__n31332, ys__n31333, ys__n31334, ys__n31335,
    ys__n31336, ys__n31337, ys__n31338, ys__n31339, ys__n31340, ys__n31341,
    ys__n31342, ys__n31343, ys__n31344, ys__n31345, ys__n31346, ys__n31347,
    ys__n31348, ys__n31349, ys__n31350, ys__n31351, ys__n31352, ys__n31353,
    ys__n31354, ys__n31355, ys__n31356, ys__n31357, ys__n31358, ys__n31359,
    ys__n31360, ys__n31361, ys__n31362, ys__n31363, ys__n31364, ys__n31365,
    ys__n31366, ys__n31367, ys__n31368, ys__n31369, ys__n31370, ys__n31371,
    ys__n31372, ys__n31373, ys__n31374, ys__n31375, ys__n31376, ys__n31377,
    ys__n31378, ys__n31379, ys__n31380, ys__n31381, ys__n31382, ys__n31383,
    ys__n31384, ys__n31385, ys__n31386, ys__n31387, ys__n31388, ys__n31389,
    ys__n31390, ys__n31391, ys__n31392, ys__n31393, ys__n31394, ys__n31395,
    ys__n31397, ys__n31398, ys__n31399, ys__n31400, ys__n31401, ys__n31402,
    ys__n31403, ys__n31404, ys__n31405, ys__n31406, ys__n31407, ys__n31408,
    ys__n31409, ys__n31410, ys__n31411, ys__n31412, ys__n31413, ys__n31414,
    ys__n31415, ys__n31416, ys__n31417, ys__n31418, ys__n31419, ys__n31420,
    ys__n31421, ys__n31422, ys__n31423, ys__n31424, ys__n31425, ys__n31426,
    ys__n31427, ys__n31428, ys__n31429, ys__n31430, ys__n31431, ys__n31432,
    ys__n31433, ys__n31434, ys__n31435, ys__n31436, ys__n31437, ys__n31438,
    ys__n31439, ys__n31440, ys__n31441, ys__n31442, ys__n31443, ys__n31444,
    ys__n31445, ys__n31446, ys__n31447, ys__n31448, ys__n31449, ys__n31450,
    ys__n31451, ys__n31452, ys__n31453, ys__n31454, ys__n31455, ys__n31456,
    ys__n31457, ys__n31458, ys__n31459, ys__n31460, ys__n31461, ys__n31462,
    ys__n31463, ys__n31464, ys__n31465, ys__n31466, ys__n31467, ys__n31468,
    ys__n31469, ys__n31470, ys__n31471, ys__n31472, ys__n31473, ys__n31474,
    ys__n31475, ys__n31476, ys__n31477, ys__n31478, ys__n31479, ys__n31480,
    ys__n31481, ys__n31482, ys__n31483, ys__n31484, ys__n31485, ys__n31486,
    ys__n31487, ys__n31488, ys__n31489, ys__n31490, ys__n31491, ys__n31492,
    ys__n31493, ys__n31494, ys__n31495, ys__n31496, ys__n31497, ys__n31498,
    ys__n31499, ys__n31500, ys__n31501, ys__n31502, ys__n31503, ys__n31504,
    ys__n31505, ys__n31506, ys__n31507, ys__n31508, ys__n31509, ys__n31510,
    ys__n31511, ys__n31512, ys__n31513, ys__n31514, ys__n31515, ys__n31516,
    ys__n31517, ys__n31518, ys__n31519, ys__n31520, ys__n31521, ys__n31522,
    ys__n31523, ys__n31524, ys__n31525, ys__n31526, ys__n31527, ys__n31528,
    ys__n31529, ys__n31530, ys__n31531, ys__n31532, ys__n31533, ys__n31534,
    ys__n31535, ys__n31536, ys__n31537, ys__n31538, ys__n31539, ys__n31540,
    ys__n31541, ys__n31542, ys__n31543, ys__n31544, ys__n31559, ys__n31560,
    ys__n31562, ys__n31564, ys__n31567, ys__n31571, ys__n31740, ys__n31741,
    ys__n31742, ys__n31743, ys__n31744, ys__n31745, ys__n31746, ys__n31747,
    ys__n31748, ys__n31749, ys__n31750, ys__n31751, ys__n31752, ys__n31753,
    ys__n31754, ys__n31755, ys__n31756, ys__n31757, ys__n31758, ys__n31759,
    ys__n31760, ys__n31761, ys__n31762, ys__n31763, ys__n31764, ys__n31765,
    ys__n31766, ys__n31767, ys__n31768, ys__n31769, ys__n31770, ys__n31771,
    ys__n31772, ys__n31773, ys__n31774, ys__n31775, ys__n31776, ys__n31777,
    ys__n31778, ys__n31779, ys__n31780, ys__n31781, ys__n31782, ys__n31783,
    ys__n31784, ys__n31785, ys__n31786, ys__n31787, ys__n31788, ys__n31789,
    ys__n31790, ys__n31791, ys__n31792, ys__n31793, ys__n31794, ys__n31795,
    ys__n31796, ys__n31797, ys__n31798, ys__n31799, ys__n31800, ys__n31801,
    ys__n31802, ys__n31803, ys__n31804, ys__n31805, ys__n31806, ys__n31807,
    ys__n31808, ys__n31809, ys__n31810, ys__n31811, ys__n31812, ys__n31813,
    ys__n31814, ys__n31815, ys__n31816, ys__n31817, ys__n31818, ys__n31819,
    ys__n31820, ys__n31821, ys__n31822, ys__n31823, ys__n31824, ys__n31825,
    ys__n31826, ys__n31827, ys__n31828, ys__n31829, ys__n31830, ys__n31831,
    ys__n31832, ys__n31833, ys__n31834, ys__n31835, ys__n31836, ys__n31837,
    ys__n31838, ys__n31839, ys__n31840, ys__n31841, ys__n31842, ys__n31843,
    ys__n31844, ys__n31845, ys__n31846, ys__n31847, ys__n31848, ys__n31849,
    ys__n31850, ys__n31851, ys__n31852, ys__n31853, ys__n31854, ys__n31855,
    ys__n31856, ys__n31857, ys__n31858, ys__n31859, ys__n31860, ys__n31861,
    ys__n31862, ys__n31863, ys__n31864, ys__n31865, ys__n31866, ys__n31867,
    ys__n31868, ys__n31869, ys__n31870, ys__n31871, ys__n31872, ys__n31873,
    ys__n31874, ys__n31875, ys__n31876, ys__n31877, ys__n31878, ys__n31879,
    ys__n31880, ys__n31881, ys__n31882, ys__n31883, ys__n31884, ys__n31885,
    ys__n31886, ys__n31887, ys__n31888, ys__n31889, ys__n31890, ys__n31891,
    ys__n31892, ys__n31893, ys__n31894, ys__n31895, ys__n31896, ys__n31897,
    ys__n31898, ys__n31899, ys__n31900, ys__n31901, ys__n31902, ys__n31903,
    ys__n31904, ys__n31905, ys__n31906, ys__n31907, ys__n31908, ys__n31909,
    ys__n31910, ys__n31911, ys__n31912, ys__n31913, ys__n31914, ys__n31915,
    ys__n31916, ys__n31917, ys__n31918, ys__n31919, ys__n31920, ys__n31921,
    ys__n31922, ys__n31923, ys__n31924, ys__n31925, ys__n31926, ys__n31927,
    ys__n31928, ys__n31929, ys__n31930, ys__n31931, ys__n31932, ys__n31933,
    ys__n31934, ys__n31935, ys__n31936, ys__n31937, ys__n31938, ys__n31939,
    ys__n31940, ys__n31941, ys__n31942, ys__n31943, ys__n31944, ys__n31945,
    ys__n31946, ys__n31947, ys__n31948, ys__n31949, ys__n31950, ys__n31953,
    ys__n31954, ys__n31955, ys__n31965, ys__n31971, ys__n31973, ys__n31975,
    ys__n31976, ys__n31978, ys__n31979, ys__n31984, ys__n31986, ys__n31988,
    ys__n31990, ys__n31992, ys__n31994, ys__n31996, ys__n31998, ys__n32000,
    ys__n32002, ys__n32004, ys__n32006, ys__n32007, ys__n32008, ys__n32010,
    ys__n32012, ys__n32014, ys__n32016, ys__n32018, ys__n32022, ys__n32023,
    ys__n32024, ys__n32025, ys__n32026, ys__n32027, ys__n32028, ys__n32029,
    ys__n32030, ys__n32031, ys__n32032, ys__n32033, ys__n32034, ys__n32035,
    ys__n32036, ys__n32037, ys__n32038, ys__n32039, ys__n32040, ys__n32041,
    ys__n32042, ys__n32043, ys__n32044, ys__n32045, ys__n32046, ys__n32047,
    ys__n32048, ys__n32049, ys__n32050, ys__n32051, ys__n32052, ys__n32053,
    ys__n32054, ys__n32055, ys__n32056, ys__n32057, ys__n32058, ys__n32059,
    ys__n32060, ys__n32061, ys__n32062, ys__n32063, ys__n32064, ys__n32065,
    ys__n32066, ys__n32067, ys__n32068, ys__n32069, ys__n32070, ys__n32071,
    ys__n32072, ys__n32073, ys__n32074, ys__n32075, ys__n32076, ys__n32077,
    ys__n32078, ys__n32079, ys__n32080, ys__n32081, ys__n32082, ys__n32083,
    ys__n32084, ys__n32085, ys__n32086, ys__n32087, ys__n32088, ys__n32124,
    ys__n32125, ys__n32126, ys__n32127, ys__n32128, ys__n32129, ys__n32130,
    ys__n32131, ys__n32132, ys__n32133, ys__n32134, ys__n32135, ys__n32136,
    ys__n32137, ys__n32138, ys__n32139, ys__n32140, ys__n32141, ys__n32142,
    ys__n32143, ys__n32144, ys__n32145, ys__n32146, ys__n32147, ys__n32148,
    ys__n32149, ys__n32150, ys__n32151, ys__n32152, ys__n32153, ys__n32154,
    ys__n32155, ys__n32158, ys__n32159, ys__n32160, ys__n32161, ys__n32162,
    ys__n32163, ys__n32164, ys__n32165, ys__n32166, ys__n32167, ys__n32168,
    ys__n32169, ys__n32170, ys__n32171, ys__n32172, ys__n32173, ys__n32174,
    ys__n32175, ys__n32176, ys__n32177, ys__n32178, ys__n32179, ys__n32180,
    ys__n32181, ys__n32182, ys__n32183, ys__n32184, ys__n32185, ys__n32186,
    ys__n32187, ys__n32188, ys__n32189, ys__n32190, ys__n32191, ys__n32192,
    ys__n32193, ys__n32194, ys__n32195, ys__n32196, ys__n32197, ys__n32198,
    ys__n32199, ys__n32200, ys__n32201, ys__n32202, ys__n32203, ys__n32204,
    ys__n32205, ys__n32206, ys__n32207, ys__n32208, ys__n32209, ys__n32210,
    ys__n32211, ys__n32212, ys__n32213, ys__n32214, ys__n32215, ys__n32216,
    ys__n32217, ys__n32218, ys__n32219, ys__n32220, ys__n32221, ys__n32222,
    ys__n32223, ys__n32224, ys__n32225, ys__n32226, ys__n32227, ys__n32228,
    ys__n32229, ys__n32230, ys__n32231, ys__n32232, ys__n32233, ys__n32234,
    ys__n32235, ys__n32236, ys__n32237, ys__n32238, ys__n32239, ys__n32240,
    ys__n32241, ys__n32242, ys__n32243, ys__n32244, ys__n32245, ys__n32246,
    ys__n32247, ys__n32248, ys__n32249, ys__n32250, ys__n32251, ys__n32252,
    ys__n32253, ys__n32254, ys__n32255, ys__n32256, ys__n32257, ys__n32258,
    ys__n32259, ys__n32260, ys__n32261, ys__n32262, ys__n32263, ys__n32264,
    ys__n32265, ys__n32266, ys__n32267, ys__n32268, ys__n32269, ys__n32270,
    ys__n32271, ys__n32272, ys__n32273, ys__n32274, ys__n32275, ys__n32276,
    ys__n32277, ys__n32278, ys__n32279, ys__n32280, ys__n32281, ys__n32282,
    ys__n32283, ys__n32284, ys__n32285, ys__n32286, ys__n32287, ys__n32288,
    ys__n32289, ys__n32290, ys__n32291, ys__n32292, ys__n32293, ys__n32294,
    ys__n32295, ys__n32296, ys__n32297, ys__n32298, ys__n32299, ys__n32300,
    ys__n32301, ys__n32302, ys__n32303, ys__n32304, ys__n32305, ys__n32306,
    ys__n32307, ys__n32308, ys__n32309, ys__n32310, ys__n32311, ys__n32312,
    ys__n32313, ys__n32314, ys__n32315, ys__n32316, ys__n32317, ys__n32318,
    ys__n32319, ys__n32320, ys__n32321, ys__n32322, ys__n32323, ys__n32324,
    ys__n32325, ys__n32326, ys__n32327, ys__n32328, ys__n32329, ys__n32330,
    ys__n32331, ys__n32332, ys__n32333, ys__n32334, ys__n32335, ys__n32336,
    ys__n32337, ys__n32338, ys__n32339, ys__n32340, ys__n32341, ys__n32342,
    ys__n32343, ys__n32344, ys__n32345, ys__n32346, ys__n32347, ys__n32348,
    ys__n32349, ys__n32350, ys__n32351, ys__n32352, ys__n32353, ys__n32354,
    ys__n32355, ys__n32356, ys__n32357, ys__n32358, ys__n32359, ys__n32360,
    ys__n32361, ys__n32362, ys__n32363, ys__n32364, ys__n32365, ys__n32366,
    ys__n32367, ys__n32368, ys__n32369, ys__n32370, ys__n32371, ys__n32372,
    ys__n32373, ys__n32374, ys__n32375, ys__n32376, ys__n32377, ys__n32378,
    ys__n32379, ys__n32380, ys__n32381, ys__n32382, ys__n32383, ys__n32384,
    ys__n32385, ys__n32386, ys__n32387, ys__n32388, ys__n32389, ys__n32390,
    ys__n32391, ys__n32392, ys__n32393, ys__n32394, ys__n32395, ys__n32396,
    ys__n32397, ys__n32398, ys__n32399, ys__n32400, ys__n32401, ys__n32402,
    ys__n32403, ys__n32404, ys__n32405, ys__n32406, ys__n32407, ys__n32408,
    ys__n32409, ys__n32410, ys__n32411, ys__n32412, ys__n32413, ys__n32414,
    ys__n32415, ys__n32416, ys__n32417, ys__n32418, ys__n32419, ys__n32420,
    ys__n32421, ys__n32422, ys__n32423, ys__n32424, ys__n32425, ys__n32426,
    ys__n32427, ys__n32428, ys__n32429, ys__n32430, ys__n32431, ys__n32432,
    ys__n32433, ys__n32434, ys__n32435, ys__n32436, ys__n32437, ys__n32438,
    ys__n32439, ys__n32440, ys__n32441, ys__n32442, ys__n32443, ys__n32444,
    ys__n32445, ys__n32446, ys__n32447, ys__n32448, ys__n32449, ys__n32450,
    ys__n32451, ys__n32452, ys__n32453, ys__n32454, ys__n32455, ys__n32456,
    ys__n32457, ys__n32458, ys__n32459, ys__n32460, ys__n32461, ys__n32462,
    ys__n32463, ys__n32464, ys__n32465, ys__n32466, ys__n32467, ys__n32468,
    ys__n32469, ys__n32470, ys__n32471, ys__n32472, ys__n32473, ys__n32474,
    ys__n32475, ys__n32476, ys__n32477, ys__n32478, ys__n32479, ys__n32480,
    ys__n32481, ys__n32482, ys__n32483, ys__n32484, ys__n32485, ys__n32486,
    ys__n32487, ys__n32488, ys__n32489, ys__n32490, ys__n32491, ys__n32492,
    ys__n32493, ys__n32494, ys__n32495, ys__n32496, ys__n32497, ys__n32498,
    ys__n32499, ys__n32500, ys__n32501, ys__n32502, ys__n32503, ys__n32504,
    ys__n32505, ys__n32506, ys__n32507, ys__n32508, ys__n32509, ys__n32510,
    ys__n32511, ys__n32512, ys__n32513, ys__n32514, ys__n32515, ys__n32516,
    ys__n32517, ys__n32518, ys__n32519, ys__n32520, ys__n32521, ys__n32522,
    ys__n32523, ys__n32524, ys__n32525, ys__n32526, ys__n32527, ys__n32528,
    ys__n32529, ys__n32530, ys__n32531, ys__n32532, ys__n32533, ys__n32534,
    ys__n32535, ys__n32536, ys__n32537, ys__n32538, ys__n32539, ys__n32540,
    ys__n32541, ys__n32542, ys__n32543, ys__n32544, ys__n32545, ys__n32546,
    ys__n32547, ys__n32548, ys__n32549, ys__n32550, ys__n32551, ys__n32552,
    ys__n32553, ys__n32554, ys__n32555, ys__n32556, ys__n32557, ys__n32558,
    ys__n32559, ys__n32560, ys__n32561, ys__n32562, ys__n32563, ys__n32564,
    ys__n32565, ys__n32566, ys__n32567, ys__n32568, ys__n32569, ys__n32570,
    ys__n32571, ys__n32572, ys__n32573, ys__n32574, ys__n32575, ys__n32576,
    ys__n32577, ys__n32578, ys__n32579, ys__n32580, ys__n32581, ys__n32582,
    ys__n32583, ys__n32584, ys__n32585, ys__n32586, ys__n32587, ys__n32588,
    ys__n32589, ys__n32590, ys__n32591, ys__n32592, ys__n32593, ys__n32594,
    ys__n32595, ys__n32596, ys__n32597, ys__n32598, ys__n32599, ys__n32600,
    ys__n32601, ys__n32602, ys__n32603, ys__n32604, ys__n32605, ys__n32606,
    ys__n32607, ys__n32608, ys__n32609, ys__n32610, ys__n32611, ys__n32612,
    ys__n32613, ys__n32614, ys__n32615, ys__n32616, ys__n32617, ys__n32618,
    ys__n32619, ys__n32620, ys__n32621, ys__n32622, ys__n32623, ys__n32624,
    ys__n32625, ys__n32626, ys__n32627, ys__n32628, ys__n32629, ys__n32630,
    ys__n32631, ys__n32632, ys__n32633, ys__n32634, ys__n32635, ys__n32636,
    ys__n32637, ys__n32638, ys__n32639, ys__n32640, ys__n32641, ys__n32642,
    ys__n32643, ys__n32644, ys__n32645, ys__n32646, ys__n32647, ys__n32648,
    ys__n32649, ys__n32650, ys__n32651, ys__n32652, ys__n32653, ys__n32654,
    ys__n32655, ys__n32656, ys__n32657, ys__n32658, ys__n32659, ys__n32660,
    ys__n32661, ys__n32662, ys__n32663, ys__n32664, ys__n32665, ys__n32666,
    ys__n32667, ys__n32668, ys__n32669, ys__n32670, ys__n32671, ys__n32672,
    ys__n32673, ys__n32674, ys__n32675, ys__n32676, ys__n32677, ys__n32678,
    ys__n32679, ys__n32680, ys__n32681, ys__n32682, ys__n32683, ys__n32684,
    ys__n32685, ys__n32686, ys__n32687, ys__n32688, ys__n32689, ys__n32690,
    ys__n32691, ys__n32692, ys__n32693, ys__n32694, ys__n32695, ys__n32696,
    ys__n32697, ys__n32698, ys__n32699, ys__n32700, ys__n32701, ys__n32702,
    ys__n32703, ys__n32704, ys__n32705, ys__n32706, ys__n32707, ys__n32708,
    ys__n32709, ys__n32710, ys__n32711, ys__n32712, ys__n32713, ys__n32714,
    ys__n32715, ys__n32716, ys__n32717, ys__n32718, ys__n32719, ys__n32720,
    ys__n32721, ys__n32722, ys__n32723, ys__n32724, ys__n32725, ys__n32726,
    ys__n32727, ys__n32728, ys__n32729, ys__n32730, ys__n32731, ys__n32732,
    ys__n32733, ys__n32734, ys__n32735, ys__n32736, ys__n32737, ys__n32738,
    ys__n32739, ys__n32740, ys__n32741, ys__n32742, ys__n32743, ys__n32744,
    ys__n32745, ys__n32746, ys__n32747, ys__n32748, ys__n32749, ys__n32750,
    ys__n32751, ys__n32752, ys__n32753, ys__n32754, ys__n32755, ys__n32756,
    ys__n32757, ys__n32758, ys__n32759, ys__n32760, ys__n32761, ys__n32762,
    ys__n32763, ys__n32764, ys__n32765, ys__n32766, ys__n32767, ys__n32768,
    ys__n32769, ys__n32770, ys__n32771, ys__n32772, ys__n32773, ys__n32774,
    ys__n32775, ys__n32776, ys__n32777, ys__n32778, ys__n32779, ys__n32780,
    ys__n32781, ys__n32782, ys__n32783, ys__n32784, ys__n32785, ys__n32786,
    ys__n32787, ys__n32788, ys__n32789, ys__n32790, ys__n32791, ys__n32792,
    ys__n32793, ys__n32794, ys__n32795, ys__n32796, ys__n32797, ys__n32798,
    ys__n32799, ys__n32800, ys__n32801, ys__n32802, ys__n32803, ys__n32804,
    ys__n32805, ys__n32806, ys__n32807, ys__n32808, ys__n32809, ys__n32810,
    ys__n32811, ys__n32812, ys__n32813, ys__n32814, ys__n32815, ys__n32816,
    ys__n32817, ys__n32818, ys__n32819, ys__n32820, ys__n32821, ys__n32822,
    ys__n32823, ys__n32824, ys__n32825, ys__n32826, ys__n32827, ys__n32828,
    ys__n32829, ys__n32830, ys__n32831, ys__n32832, ys__n32833, ys__n32834,
    ys__n32835, ys__n32836, ys__n32837, ys__n32838, ys__n32839, ys__n32840,
    ys__n32841, ys__n32842, ys__n32843, ys__n32844, ys__n32845, ys__n32846,
    ys__n32847, ys__n32848, ys__n32849, ys__n32850, ys__n32851, ys__n32852,
    ys__n32853, ys__n32854, ys__n32855, ys__n32856, ys__n32857, ys__n32858,
    ys__n32859, ys__n32860, ys__n32861, ys__n32862, ys__n32863, ys__n32864,
    ys__n32865, ys__n32866, ys__n32867, ys__n32868, ys__n32869, ys__n32870,
    ys__n32871, ys__n32872, ys__n32873, ys__n32874, ys__n32875, ys__n32876,
    ys__n32877, ys__n32878, ys__n32879, ys__n32880, ys__n32881, ys__n32882,
    ys__n32883, ys__n32884, ys__n32885, ys__n32886, ys__n32887, ys__n32888,
    ys__n32889, ys__n32890, ys__n32891, ys__n32892, ys__n32893, ys__n32894,
    ys__n32895, ys__n32896, ys__n32897, ys__n32898, ys__n32899, ys__n32900,
    ys__n32901, ys__n32902, ys__n32903, ys__n32904, ys__n32905, ys__n32906,
    ys__n32907, ys__n32908, ys__n32909, ys__n32910, ys__n32911, ys__n32912,
    ys__n32913, ys__n32914, ys__n32915, ys__n32916, ys__n32917, ys__n32918,
    ys__n32919, ys__n32920, ys__n32921, ys__n32922, ys__n32923, ys__n32924,
    ys__n32925, ys__n32926, ys__n32927, ys__n32928, ys__n32929, ys__n32930,
    ys__n32931, ys__n32932, ys__n32933, ys__n32934, ys__n32935, ys__n32936,
    ys__n32937, ys__n32938, ys__n32939, ys__n32940, ys__n32941, ys__n32942,
    ys__n32943, ys__n32944, ys__n32945, ys__n32946, ys__n32947, ys__n32948,
    ys__n32949, ys__n32950, ys__n32951, ys__n32952, ys__n32953, ys__n32954,
    ys__n32955, ys__n32956, ys__n32957, ys__n32958, ys__n32959, ys__n32960,
    ys__n32961, ys__n32962, ys__n32963, ys__n32964, ys__n32965, ys__n32966,
    ys__n32967, ys__n32968, ys__n32969, ys__n32970, ys__n32971, ys__n32972,
    ys__n32973, ys__n32974, ys__n32975, ys__n32976, ys__n32977, ys__n32978,
    ys__n32979, ys__n32980, ys__n32981, ys__n32982, ys__n32983, ys__n32984,
    ys__n32985, ys__n32986, ys__n32987, ys__n32988, ys__n32989, ys__n32990,
    ys__n32991, ys__n32992, ys__n32993, ys__n32994, ys__n32995, ys__n32996,
    ys__n32997, ys__n32998, ys__n33007, ys__n33008, ys__n33009, ys__n33014,
    ys__n33015, ys__n33016, ys__n33017, ys__n33018, ys__n33019, ys__n33020,
    ys__n33021, ys__n33022, ys__n33023, ys__n33024, ys__n33025, ys__n33026,
    ys__n33027, ys__n33028, ys__n33029, ys__n33030, ys__n33031, ys__n33032,
    ys__n33033, ys__n33034, ys__n33035, ys__n33036, ys__n33037, ys__n33038,
    ys__n33039, ys__n33040, ys__n33041, ys__n33042, ys__n33043, ys__n33044,
    ys__n33045, ys__n33046, ys__n33047, ys__n33048, ys__n33049, ys__n33050,
    ys__n33051, ys__n33052, ys__n33053, ys__n33054, ys__n33055, ys__n33056,
    ys__n33058, ys__n33059, ys__n33060, ys__n33061, ys__n33062, ys__n33063,
    ys__n33064, ys__n33065, ys__n33066, ys__n33067, ys__n33068, ys__n33069,
    ys__n33070, ys__n33071, ys__n33072, ys__n33073, ys__n33074, ys__n33075,
    ys__n33076, ys__n33077, ys__n33078, ys__n33079, ys__n33080, ys__n33081,
    ys__n33082, ys__n33083, ys__n33084, ys__n33085, ys__n33086, ys__n33087,
    ys__n33088, ys__n33089, ys__n33090, ys__n33091, ys__n33092, ys__n33093,
    ys__n33094, ys__n33095, ys__n33096, ys__n33097, ys__n33098, ys__n33099,
    ys__n33100, ys__n33101, ys__n33102, ys__n33103, ys__n33104, ys__n33105,
    ys__n33106, ys__n33107, ys__n33108, ys__n33109, ys__n33110, ys__n33111,
    ys__n33178, ys__n33179, ys__n33180, ys__n33181, ys__n33182, ys__n33183,
    ys__n33184, ys__n33185, ys__n33186, ys__n33187, ys__n33188, ys__n33189,
    ys__n33190, ys__n33191, ys__n33192, ys__n33193, ys__n33194, ys__n33195,
    ys__n33196, ys__n33197, ys__n33198, ys__n33199, ys__n33200, ys__n33201,
    ys__n33202, ys__n33203, ys__n33204, ys__n33205, ys__n33206, ys__n33207,
    ys__n33208, ys__n33209, ys__n33211, ys__n33317, ys__n33324, ys__n33329,
    ys__n33331, ys__n33333, ys__n33335, ys__n33337, ys__n33339, ys__n33357,
    ys__n33366, ys__n33414, ys__n33420, ys__n33437, ys__n33438, ys__n33439,
    ys__n33453, ys__n33454, ys__n33455, ys__n33456, ys__n33457, ys__n33513,
    ys__n33514, ys__n33515, ys__n33521, ys__n33535, ys__n34952, ys__n34953,
    ys__n34962, ys__n35052, ys__n35144, ys__n35146, ys__n35148, ys__n35150,
    ys__n35152, ys__n35154, ys__n35156, ys__n35158, ys__n35160, ys__n35162,
    ys__n35164, ys__n35166, ys__n35168, ys__n35170, ys__n35172, ys__n35174,
    ys__n35176, ys__n35178, ys__n35180, ys__n35182, ys__n35184, ys__n35186,
    ys__n35188, ys__n35190, ys__n35192, ys__n35194, ys__n35196, ys__n35198,
    ys__n35200, ys__n35202, ys__n35204, ys__n35206, ys__n35402, ys__n35404,
    ys__n35406, ys__n35408, ys__n35410, ys__n35412, ys__n35425, ys__n35705,
    ys__n35706, ys__n35708, ys__n35710, ys__n35712, ys__n35714, ys__n35716,
    ys__n37676, ys__n37687, ys__n37695, ys__n37697, ys__n37699, ys__n37702,
    ys__n37703, ys__n37707, ys__n37714, ys__n37731, ys__n37732, ys__n37733,
    ys__n37738, ys__n37739, ys__n37741, ys__n37742, ys__n38180, ys__n38182,
    ys__n38184, ys__n38185, ys__n38186, ys__n38188, ys__n38191, ys__n38205,
    ys__n38207, ys__n38209, ys__n38211, ys__n38213, ys__n38214, ys__n38216,
    ys__n38218, ys__n38222, ys__n38224, ys__n38246, ys__n38247, ys__n38248,
    ys__n38250, ys__n38252, ys__n38263, ys__n38266, ys__n38281, ys__n38285,
    ys__n38287, ys__n38289, ys__n38292, ys__n38294, ys__n38296, ys__n38303,
    ys__n38325, ys__n38326, ys__n38327, ys__n38328, ys__n38330, ys__n38331,
    ys__n38332, ys__n38334, ys__n38336, ys__n38337, ys__n38338, ys__n38339,
    ys__n38340, ys__n38341, ys__n38342, ys__n38343, ys__n38344, ys__n38345,
    ys__n38347, ys__n38349, ys__n38351, ys__n38352, ys__n38353, ys__n38354,
    ys__n38355, ys__n38356, ys__n38357, ys__n38359, ys__n38360, ys__n38362,
    ys__n38364, ys__n38365, ys__n38366, ys__n38367, ys__n38368, ys__n38369,
    ys__n38370, ys__n38371, ys__n38372, ys__n38373, ys__n38374, ys__n38375,
    ys__n38377, ys__n38379, ys__n38381, ys__n38383, ys__n38385, ys__n38387,
    ys__n38388, ys__n38389, ys__n38390, ys__n38391, ys__n38392, ys__n38393,
    ys__n38394, ys__n38396, ys__n38397, ys__n38417, ys__n38453, ys__n38456,
    ys__n38508, ys__n38509, ys__n38510, ys__n38515, ys__n38518, ys__n38520,
    ys__n38521, ys__n38523, ys__n38525, ys__n38552, ys__n38555, ys__n38556,
    ys__n38563, ys__n38566, ys__n38615, ys__n38623, ys__n38628, ys__n38633,
    ys__n38650, ys__n38662, ys__n38668, ys__n38669, ys__n38672, ys__n38674,
    ys__n38677, ys__n38689, ys__n38742, ys__n38768, ys__n38795, ys__n38799,
    ys__n38801, ys__n38884, ys__n38886, ys__n38887, ys__n38900, ys__n38912,
    ys__n38913, ys__n38914, ys__n38915, ys__n38917, ys__n38923, ys__n38925,
    ys__n38930, ys__n39392, ys__n39393, ys__n39395, ys__n39396, ys__n39397,
    ys__n39398, ys__n39399, ys__n39400, ys__n39401, ys__n39402, ys__n39403,
    ys__n39404, ys__n39405, ys__n39406, ys__n39407, ys__n39408, ys__n39409,
    ys__n39410, ys__n39411, ys__n39412, ys__n39413, ys__n39414, ys__n39415,
    ys__n39416, ys__n39417, ys__n39418, ys__n40052, ys__n42129, ys__n42153,
    ys__n42189, ys__n42194, ys__n42229, ys__n42234, ys__n42270, ys__n42275,
    ys__n42311, ys__n42316, ys__n42352, ys__n42357, ys__n42393, ys__n42398,
    ys__n42434, ys__n42439, ys__n42488, ys__n42493, ys__n42541, ys__n42546,
    ys__n42594, ys__n42599, ys__n42647, ys__n42652, ys__n42701, ys__n42706,
    ys__n42755, ys__n42760, ys__n42809, ys__n42814, ys__n42863, ys__n42868,
    ys__n42917, ys__n42922, ys__n42971, ys__n42976, ys__n43025, ys__n43030,
    ys__n43079, ys__n43084, ys__n43133, ys__n43138, ys__n43187, ys__n43192,
    ys__n43241, ys__n43246, ys__n43295, ys__n43300, ys__n43349, ys__n43354,
    ys__n43403, ys__n43408, ys__n43457, ys__n43462, ys__n43511, ys__n43516,
    ys__n43565, ys__n43570, ys__n43619, ys__n43624, ys__n43673, ys__n43678,
    ys__n43727, ys__n43732, ys__n43781, ys__n43786, ys__n43835, ys__n43840,
    ys__n43889, ys__n43894, ys__n43932, ys__n43937, ys__n43975, ys__n43980,
    ys__n44018, ys__n44023, ys__n44048, ys__n44053, ys__n44089, ys__n44094,
    ys__n44119, ys__n44122, ys__n44136, ys__n44139, ys__n44155, ys__n44160,
    ys__n44183, ys__n44186, ys__n44189, ys__n44192, ys__n44195, ys__n44198,
    ys__n44205, ys__n44213, ys__n44216, ys__n44219, ys__n44836, ys__n44838,
    ys__n44841, ys__n44843, ys__n44844, ys__n44845, ys__n44846, ys__n44848,
    ys__n44850, ys__n44851, ys__n44852, ys__n44853, ys__n44854, ys__n44855,
    ys__n44858, ys__n44948, ys__n44949, ys__n44950, ys__n44952, ys__n44953,
    ys__n44954, ys__n44955, ys__n44956, ys__n44957, ys__n44958, ys__n44959,
    ys__n44960, ys__n44961, ys__n44962, ys__n44963, ys__n44964, ys__n44965,
    ys__n44966, ys__n44967, ys__n44968, ys__n44969, ys__n44970, ys__n44971,
    ys__n44972, ys__n44973, ys__n44974, ys__n44975, ys__n44976, ys__n44977,
    ys__n44978, ys__n44979, ys__n44980, ys__n44981, ys__n44982, ys__n44983,
    ys__n44985, ys__n44987, ys__n46131, ys__n46133, ys__n46135, ys__n46137,
    ys__n46143, ys__n46146, ys__n46154, ys__n46155, ys__n46158, ys__n46159,
    ys__n46162, ys__n46163, ys__n46172, ys__n46173, ys__n46176, ys__n46179,
    ys__n46188, ys__n46189, ys__n46192, ys__n46195, ys__n46204, ys__n46205,
    ys__n46208, ys__n46211, ys__n46220, ys__n46221, ys__n46224, ys__n46227,
    ys__n46233, ys__n46234, ys__n48339, ys__n48340, ys__n48341, ys__n48342,
    ys__n48343, ys__n48344, ys__n48348, ys__n48349, ys__n48350, ys__n48351,
    ys__n48352, ys__n48353, ys__n48354, ys__n48355, ys__n48356, ys__n48357,
    ys__n48358, ys__n48359, ys__n48360, ys__n48361, ys__n48362  );
  input  ys__n14, ys__n16, ys__n22, ys__n24, ys__n26, ys__n28, ys__n30,
    ys__n32, ys__n34, ys__n36, ys__n38, ys__n40, ys__n42, ys__n44, ys__n46,
    ys__n48, ys__n50, ys__n52, ys__n54, ys__n56, ys__n58, ys__n60, ys__n62,
    ys__n66, ys__n70, ys__n72, ys__n74, ys__n76, ys__n78, ys__n80, ys__n82,
    ys__n84, ys__n86, ys__n88, ys__n90, ys__n96, ys__n98, ys__n100,
    ys__n108, ys__n110, ys__n112, ys__n114, ys__n116, ys__n118, ys__n120,
    ys__n122, ys__n124, ys__n126, ys__n128, ys__n130, ys__n132, ys__n134,
    ys__n136, ys__n138, ys__n140, ys__n142, ys__n148, ys__n150, ys__n152,
    ys__n156, ys__n158, ys__n160, ys__n162, ys__n164, ys__n166, ys__n168,
    ys__n170, ys__n172, ys__n174, ys__n176, ys__n178, ys__n182, ys__n184,
    ys__n186, ys__n190, ys__n192, ys__n194, ys__n196, ys__n198, ys__n202,
    ys__n204, ys__n206, ys__n208, ys__n210, ys__n212, ys__n214, ys__n216,
    ys__n218, ys__n220, ys__n222, ys__n226, ys__n232, ys__n238, ys__n240,
    ys__n242, ys__n244, ys__n248, ys__n256, ys__n258, ys__n262, ys__n290,
    ys__n294, ys__n296, ys__n298, ys__n300, ys__n302, ys__n304, ys__n306,
    ys__n308, ys__n310, ys__n312, ys__n314, ys__n316, ys__n318, ys__n326,
    ys__n328, ys__n330, ys__n332, ys__n336, ys__n338, ys__n340, ys__n342,
    ys__n344, ys__n346, ys__n348, ys__n350, ys__n352, ys__n354, ys__n356,
    ys__n358, ys__n360, ys__n362, ys__n364, ys__n366, ys__n368, ys__n370,
    ys__n372, ys__n374, ys__n376, ys__n378, ys__n380, ys__n382, ys__n384,
    ys__n386, ys__n392, ys__n394, ys__n396, ys__n398, ys__n402, ys__n408,
    ys__n414, ys__n416, ys__n418, ys__n420, ys__n422, ys__n424, ys__n426,
    ys__n428, ys__n430, ys__n432, ys__n434, ys__n436, ys__n438, ys__n440,
    ys__n442, ys__n444, ys__n446, ys__n448, ys__n450, ys__n452, ys__n454,
    ys__n456, ys__n464, ys__n488, ys__n490, ys__n500, ys__n504, ys__n512,
    ys__n514, ys__n516, ys__n518, ys__n520, ys__n522, ys__n524, ys__n526,
    ys__n528, ys__n530, ys__n532, ys__n536, ys__n538, ys__n544, ys__n546,
    ys__n548, ys__n550, ys__n556, ys__n558, ys__n562, ys__n564, ys__n566,
    ys__n568, ys__n570, ys__n572, ys__n580, ys__n582, ys__n584, ys__n586,
    ys__n588, ys__n598, ys__n600, ys__n602, ys__n604, ys__n606, ys__n608,
    ys__n610, ys__n612, ys__n614, ys__n616, ys__n618, ys__n620, ys__n622,
    ys__n624, ys__n626, ys__n632, ys__n634, ys__n636, ys__n638, ys__n640,
    ys__n642, ys__n644, ys__n646, ys__n648, ys__n650, ys__n652, ys__n654,
    ys__n656, ys__n658, ys__n660, ys__n662, ys__n664, ys__n666, ys__n668,
    ys__n670, ys__n672, ys__n674, ys__n676, ys__n678, ys__n680, ys__n682,
    ys__n684, ys__n686, ys__n688, ys__n690, ys__n692, ys__n694, ys__n696,
    ys__n698, ys__n700, ys__n702, ys__n704, ys__n706, ys__n708, ys__n710,
    ys__n712, ys__n718, ys__n720, ys__n722, ys__n724, ys__n726, ys__n728,
    ys__n736, ys__n742, ys__n744, ys__n746, ys__n748, ys__n750, ys__n752,
    ys__n758, ys__n760, ys__n762, ys__n764, ys__n766, ys__n768, ys__n770,
    ys__n772, ys__n774, ys__n776, ys__n778, ys__n780, ys__n782, ys__n784,
    ys__n816, ys__n818, ys__n820, ys__n822, ys__n824, ys__n826, ys__n828,
    ys__n830, ys__n832, ys__n834, ys__n836, ys__n838, ys__n840, ys__n842,
    ys__n844, ys__n846, ys__n848, ys__n850, ys__n852, ys__n854, ys__n856,
    ys__n858, ys__n860, ys__n874, ys__n889, ys__n935, ys__n1029, ys__n1036,
    ys__n1038, ys__n1048, ys__n1072, ys__n1076, ys__n1078, ys__n1084,
    ys__n1094, ys__n1098, ys__n1099, ys__n1106, ys__n1107, ys__n1109,
    ys__n1110, ys__n1116, ys__n1117, ys__n1119, ys__n1120, ys__n1129,
    ys__n1147, ys__n1151, ys__n1153, ys__n1154, ys__n1156, ys__n1157,
    ys__n1301, ys__n1309, ys__n1489, ys__n1490, ys__n1492, ys__n1493,
    ys__n1495, ys__n1496, ys__n1498, ys__n1499, ys__n1502, ys__n1503,
    ys__n1505, ys__n1506, ys__n1508, ys__n1509, ys__n1511, ys__n1535,
    ys__n2024, ys__n2233, ys__n2239, ys__n2245, ys__n2247, ys__n2251,
    ys__n2276, ys__n2282, ys__n2306, ys__n2308, ys__n2312, ys__n2427,
    ys__n2429, ys__n2433, ys__n2644, ys__n2652, ys__n2693, ys__n2716,
    ys__n2779, ys__n2830, ys__n2924, ys__n3214, ys__n4168, ys__n4176,
    ys__n4177, ys__n4184, ys__n4185, ys__n4190, ys__n4291, ys__n4292,
    ys__n4294, ys__n4296, ys__n4297, ys__n4299, ys__n4300, ys__n4305,
    ys__n4340, ys__n4448, ys__n4449, ys__n4451, ys__n4452, ys__n4454,
    ys__n4455, ys__n4457, ys__n4458, ys__n4460, ys__n4461, ys__n4465,
    ys__n4478, ys__n4480, ys__n4488, ys__n4494, ys__n4496, ys__n4613,
    ys__n4625, ys__n4627, ys__n4688, ys__n4698, ys__n4736, ys__n4744,
    ys__n4746, ys__n4750, ys__n4751, ys__n4753, ys__n4754, ys__n4756,
    ys__n4757, ys__n4759, ys__n4761, ys__n4783, ys__n4784, ys__n4810,
    ys__n4826, ys__n4832, ys__n4833, ys__n4836, ys__n4837, ys__n6112,
    ys__n6113, ys__n6115, ys__n6118, ys__n6119, ys__n6120, ys__n6121,
    ys__n6123, ys__n6124, ys__n6126, ys__n6127, ys__n6129, ys__n6130,
    ys__n6133, ys__n6134, ys__n17803, ys__n17804, ys__n17806, ys__n17807,
    ys__n17809, ys__n17810, ys__n17812, ys__n17813, ys__n17815, ys__n17816,
    ys__n17818, ys__n17819, ys__n17821, ys__n17822, ys__n17824, ys__n17825,
    ys__n17827, ys__n17828, ys__n17830, ys__n17831, ys__n17833, ys__n17834,
    ys__n17836, ys__n17837, ys__n17839, ys__n17840, ys__n17842, ys__n17843,
    ys__n17845, ys__n17846, ys__n17848, ys__n17849, ys__n17866, ys__n17867,
    ys__n17869, ys__n17870, ys__n17872, ys__n17873, ys__n17875, ys__n17876,
    ys__n17878, ys__n17879, ys__n17881, ys__n17882, ys__n17884, ys__n17885,
    ys__n17887, ys__n17888, ys__n17890, ys__n17891, ys__n17893, ys__n17894,
    ys__n17896, ys__n17897, ys__n17899, ys__n17900, ys__n17902, ys__n17903,
    ys__n17905, ys__n17906, ys__n17908, ys__n17909, ys__n17911, ys__n17912,
    ys__n17941, ys__n17943, ys__n18041, ys__n18043, ys__n18045, ys__n18047,
    ys__n18049, ys__n18051, ys__n18053, ys__n18055, ys__n18057, ys__n18059,
    ys__n18061, ys__n18063, ys__n18065, ys__n18067, ys__n18070, ys__n18071,
    ys__n18090, ys__n18101, ys__n18105, ys__n18106, ys__n18109, ys__n18111,
    ys__n18112, ys__n18114, ys__n18116, ys__n18118, ys__n18121, ys__n18122,
    ys__n18124, ys__n18143, ys__n18149, ys__n18150, ys__n18156, ys__n18173,
    ys__n18208, ys__n18226, ys__n18229, ys__n18231, ys__n18240, ys__n18242,
    ys__n18243, ys__n18270, ys__n18271, ys__n18277, ys__n18280, ys__n18283,
    ys__n18286, ys__n18317, ys__n18378, ys__n18381, ys__n18384, ys__n18389,
    ys__n18393, ys__n18448, ys__n18451, ys__n18454, ys__n18457, ys__n18460,
    ys__n18463, ys__n18466, ys__n18469, ys__n18472, ys__n18475, ys__n18478,
    ys__n18481, ys__n18484, ys__n18487, ys__n18490, ys__n18493, ys__n18496,
    ys__n18499, ys__n18502, ys__n18505, ys__n18508, ys__n18511, ys__n18514,
    ys__n18517, ys__n18520, ys__n18523, ys__n18526, ys__n18529, ys__n18532,
    ys__n18535, ys__n18538, ys__n18541, ys__n18544, ys__n18546, ys__n18556,
    ys__n18558, ys__n18560, ys__n18562, ys__n18565, ys__n18568, ys__n18569,
    ys__n18571, ys__n18572, ys__n18574, ys__n18575, ys__n18577, ys__n18578,
    ys__n18580, ys__n18581, ys__n18583, ys__n18584, ys__n18586, ys__n18587,
    ys__n18589, ys__n18590, ys__n18592, ys__n18593, ys__n18595, ys__n18596,
    ys__n18598, ys__n18599, ys__n18601, ys__n18602, ys__n18604, ys__n18605,
    ys__n18607, ys__n18608, ys__n18610, ys__n18611, ys__n18613, ys__n18614,
    ys__n18616, ys__n18617, ys__n18619, ys__n18620, ys__n18622, ys__n18623,
    ys__n18625, ys__n18626, ys__n18628, ys__n18630, ys__n18632, ys__n18634,
    ys__n18636, ys__n18638, ys__n18639, ys__n18641, ys__n18642, ys__n18644,
    ys__n18645, ys__n18647, ys__n18650, ys__n18651, ys__n18749, ys__n18752,
    ys__n18755, ys__n18758, ys__n18761, ys__n18762, ys__n18765, ys__n18767,
    ys__n18769, ys__n18771, ys__n18773, ys__n18775, ys__n18777, ys__n18779,
    ys__n18781, ys__n18783, ys__n18785, ys__n18787, ys__n18789, ys__n18791,
    ys__n18793, ys__n18795, ys__n18797, ys__n18799, ys__n18801, ys__n18803,
    ys__n18805, ys__n18807, ys__n18809, ys__n18811, ys__n18813, ys__n18815,
    ys__n18817, ys__n18819, ys__n18821, ys__n18823, ys__n18825, ys__n18827,
    ys__n18829, ys__n18831, ys__n18833, ys__n18835, ys__n18837, ys__n18839,
    ys__n18841, ys__n18843, ys__n18845, ys__n18847, ys__n18849, ys__n18851,
    ys__n18853, ys__n18855, ys__n18857, ys__n18859, ys__n18861, ys__n18863,
    ys__n18865, ys__n18867, ys__n18869, ys__n18871, ys__n18873, ys__n18875,
    ys__n18877, ys__n18879, ys__n18881, ys__n18883, ys__n18885, ys__n18887,
    ys__n18889, ys__n18891, ys__n18956, ys__n18957, ys__n18958, ys__n18959,
    ys__n18960, ys__n18961, ys__n18962, ys__n18963, ys__n18964, ys__n18965,
    ys__n18966, ys__n18967, ys__n18968, ys__n18969, ys__n18970, ys__n18971,
    ys__n18972, ys__n18973, ys__n18974, ys__n18975, ys__n18976, ys__n18977,
    ys__n18978, ys__n18979, ys__n18980, ys__n18981, ys__n18982, ys__n18983,
    ys__n18984, ys__n18985, ys__n18986, ys__n18987, ys__n18989, ys__n18991,
    ys__n18993, ys__n18995, ys__n18997, ys__n18999, ys__n19001, ys__n19003,
    ys__n19005, ys__n19007, ys__n19009, ys__n19011, ys__n19013, ys__n19015,
    ys__n19017, ys__n19019, ys__n19021, ys__n19023, ys__n19025, ys__n19027,
    ys__n19029, ys__n19031, ys__n19033, ys__n19035, ys__n19037, ys__n19039,
    ys__n19041, ys__n19043, ys__n19045, ys__n19047, ys__n19049, ys__n19051,
    ys__n19116, ys__n19117, ys__n19118, ys__n19119, ys__n19120, ys__n19121,
    ys__n19122, ys__n19123, ys__n19124, ys__n19125, ys__n19126, ys__n19127,
    ys__n19128, ys__n19129, ys__n19130, ys__n19131, ys__n19132, ys__n19133,
    ys__n19134, ys__n19135, ys__n19136, ys__n19137, ys__n19138, ys__n19139,
    ys__n19140, ys__n19141, ys__n19142, ys__n19143, ys__n19144, ys__n19145,
    ys__n19146, ys__n19147, ys__n19156, ys__n19157, ys__n19166, ys__n19171,
    ys__n19203, ys__n19215, ys__n19245, ys__n19251, ys__n19253, ys__n19259,
    ys__n19261, ys__n19263, ys__n19843, ys__n19844, ys__n19845, ys__n19846,
    ys__n19847, ys__n19848, ys__n19849, ys__n19850, ys__n19851, ys__n19852,
    ys__n19853, ys__n19854, ys__n19855, ys__n19856, ys__n19857, ys__n19858,
    ys__n19859, ys__n19860, ys__n19861, ys__n19862, ys__n19863, ys__n19864,
    ys__n19865, ys__n19866, ys__n19867, ys__n19868, ys__n19869, ys__n19870,
    ys__n19871, ys__n19872, ys__n19873, ys__n19874, ys__n19875, ys__n19972,
    ys__n19973, ys__n19974, ys__n19975, ys__n19976, ys__n19977, ys__n19978,
    ys__n19979, ys__n19980, ys__n19981, ys__n19982, ys__n19983, ys__n19984,
    ys__n19985, ys__n19986, ys__n19987, ys__n19988, ys__n19989, ys__n19990,
    ys__n19991, ys__n19992, ys__n19993, ys__n19994, ys__n19995, ys__n19996,
    ys__n19997, ys__n19998, ys__n19999, ys__n20000, ys__n20001, ys__n20002,
    ys__n20003, ys__n20004, ys__n20035, ys__n20058, ys__n20061, ys__n20064,
    ys__n20067, ys__n20070, ys__n20073, ys__n20076, ys__n20079, ys__n20138,
    ys__n20140, ys__n20142, ys__n20144, ys__n20146, ys__n20148, ys__n20150,
    ys__n20152, ys__n20186, ys__n20188, ys__n20190, ys__n20192, ys__n20194,
    ys__n20196, ys__n20198, ys__n20200, ys__n20202, ys__n20204, ys__n20206,
    ys__n20208, ys__n20210, ys__n20212, ys__n20214, ys__n20216, ys__n20273,
    ys__n20279, ys__n20280, ys__n20540, ys__n20542, ys__n20544, ys__n20546,
    ys__n20548, ys__n20550, ys__n20552, ys__n20554, ys__n20556, ys__n20558,
    ys__n20560, ys__n20562, ys__n20564, ys__n20566, ys__n20568, ys__n20570,
    ys__n20572, ys__n20574, ys__n20576, ys__n20578, ys__n20580, ys__n20582,
    ys__n20584, ys__n20586, ys__n20588, ys__n20590, ys__n20592, ys__n20594,
    ys__n20596, ys__n20598, ys__n20600, ys__n20602, ys__n20604, ys__n20606,
    ys__n20608, ys__n20610, ys__n20612, ys__n20614, ys__n20616, ys__n20618,
    ys__n20620, ys__n20622, ys__n20624, ys__n20626, ys__n20628, ys__n20630,
    ys__n20632, ys__n20634, ys__n20636, ys__n20638, ys__n20640, ys__n20642,
    ys__n20644, ys__n20646, ys__n20648, ys__n20650, ys__n20652, ys__n20654,
    ys__n20656, ys__n20658, ys__n20660, ys__n20662, ys__n20664, ys__n20666,
    ys__n20668, ys__n20670, ys__n20672, ys__n20674, ys__n20676, ys__n20678,
    ys__n20680, ys__n20682, ys__n20684, ys__n20686, ys__n20688, ys__n20690,
    ys__n20692, ys__n20694, ys__n20696, ys__n20698, ys__n20700, ys__n20702,
    ys__n20704, ys__n20706, ys__n20708, ys__n20710, ys__n20712, ys__n20714,
    ys__n20716, ys__n20718, ys__n20720, ys__n20722, ys__n20724, ys__n20726,
    ys__n20728, ys__n20730, ys__n20732, ys__n20734, ys__n20736, ys__n20738,
    ys__n20740, ys__n20742, ys__n20744, ys__n20746, ys__n20748, ys__n20750,
    ys__n20752, ys__n20754, ys__n20756, ys__n20758, ys__n20760, ys__n20762,
    ys__n20764, ys__n20766, ys__n20768, ys__n20770, ys__n20772, ys__n20774,
    ys__n20776, ys__n20778, ys__n20780, ys__n20782, ys__n20784, ys__n20786,
    ys__n20788, ys__n20790, ys__n20792, ys__n20794, ys__n20796, ys__n20798,
    ys__n20800, ys__n20802, ys__n20804, ys__n20806, ys__n20808, ys__n20810,
    ys__n20812, ys__n20814, ys__n20816, ys__n20818, ys__n20820, ys__n20822,
    ys__n20824, ys__n20826, ys__n20828, ys__n20830, ys__n20832, ys__n20834,
    ys__n20836, ys__n20838, ys__n20840, ys__n20842, ys__n20844, ys__n20846,
    ys__n20848, ys__n20850, ys__n20852, ys__n20854, ys__n20856, ys__n20858,
    ys__n20860, ys__n20862, ys__n20864, ys__n20866, ys__n20868, ys__n20870,
    ys__n20872, ys__n20874, ys__n20876, ys__n20878, ys__n20880, ys__n20882,
    ys__n20884, ys__n20886, ys__n20888, ys__n20890, ys__n20892, ys__n20894,
    ys__n20896, ys__n20898, ys__n20900, ys__n20902, ys__n20904, ys__n20906,
    ys__n20908, ys__n20910, ys__n20912, ys__n20914, ys__n20916, ys__n20918,
    ys__n20920, ys__n20922, ys__n20924, ys__n20925, ys__n20926, ys__n20927,
    ys__n20928, ys__n20929, ys__n20930, ys__n20931, ys__n20932, ys__n20933,
    ys__n20934, ys__n20935, ys__n20936, ys__n20937, ys__n20938, ys__n20939,
    ys__n20940, ys__n20941, ys__n20942, ys__n20943, ys__n20944, ys__n20945,
    ys__n20946, ys__n20947, ys__n20948, ys__n20949, ys__n20950, ys__n20951,
    ys__n20952, ys__n20953, ys__n20954, ys__n20955, ys__n20956, ys__n20958,
    ys__n20960, ys__n20962, ys__n20964, ys__n20966, ys__n20968, ys__n20970,
    ys__n20972, ys__n20974, ys__n20976, ys__n20978, ys__n20980, ys__n20982,
    ys__n20984, ys__n20986, ys__n20988, ys__n20990, ys__n20992, ys__n20994,
    ys__n20996, ys__n20998, ys__n21000, ys__n21002, ys__n21004, ys__n21006,
    ys__n21008, ys__n21010, ys__n21012, ys__n21014, ys__n21016, ys__n21018,
    ys__n21020, ys__n21022, ys__n21024, ys__n21026, ys__n21028, ys__n21030,
    ys__n21032, ys__n21034, ys__n21036, ys__n21038, ys__n21040, ys__n21042,
    ys__n21044, ys__n21046, ys__n21048, ys__n21050, ys__n21052, ys__n21054,
    ys__n21056, ys__n21058, ys__n21060, ys__n21062, ys__n21064, ys__n21066,
    ys__n21068, ys__n21070, ys__n21072, ys__n21074, ys__n21076, ys__n21078,
    ys__n21080, ys__n21082, ys__n21084, ys__n21086, ys__n21088, ys__n21090,
    ys__n21092, ys__n21094, ys__n21096, ys__n21098, ys__n21100, ys__n21102,
    ys__n21104, ys__n21106, ys__n21108, ys__n21110, ys__n21112, ys__n21114,
    ys__n21116, ys__n21118, ys__n21120, ys__n21122, ys__n21124, ys__n21126,
    ys__n21128, ys__n21130, ys__n21132, ys__n21134, ys__n21136, ys__n21138,
    ys__n21140, ys__n21142, ys__n21144, ys__n21146, ys__n21148, ys__n21150,
    ys__n21152, ys__n21154, ys__n21156, ys__n21158, ys__n21160, ys__n21162,
    ys__n21164, ys__n21166, ys__n21168, ys__n21170, ys__n21172, ys__n21174,
    ys__n21176, ys__n21178, ys__n21180, ys__n21182, ys__n21184, ys__n21186,
    ys__n21188, ys__n21190, ys__n21192, ys__n21194, ys__n21196, ys__n21198,
    ys__n21200, ys__n21202, ys__n21204, ys__n21206, ys__n21208, ys__n21210,
    ys__n21212, ys__n21214, ys__n21216, ys__n21218, ys__n21220, ys__n21222,
    ys__n21224, ys__n21226, ys__n21228, ys__n21230, ys__n21232, ys__n21234,
    ys__n21236, ys__n21238, ys__n21240, ys__n21242, ys__n21244, ys__n21246,
    ys__n21248, ys__n21250, ys__n21252, ys__n21254, ys__n21256, ys__n21258,
    ys__n21260, ys__n21262, ys__n21264, ys__n21266, ys__n21268, ys__n21270,
    ys__n21272, ys__n21274, ys__n21276, ys__n21278, ys__n21280, ys__n21282,
    ys__n21284, ys__n21286, ys__n21288, ys__n21290, ys__n21292, ys__n21294,
    ys__n21296, ys__n21298, ys__n21300, ys__n21302, ys__n21304, ys__n21306,
    ys__n21308, ys__n21310, ys__n21312, ys__n21314, ys__n21316, ys__n21318,
    ys__n21320, ys__n21322, ys__n21324, ys__n21326, ys__n21328, ys__n21330,
    ys__n21332, ys__n21334, ys__n21336, ys__n21338, ys__n21340, ys__n21342,
    ys__n21344, ys__n21346, ys__n21348, ys__n21350, ys__n21352, ys__n21354,
    ys__n21356, ys__n21358, ys__n21360, ys__n21362, ys__n21364, ys__n21366,
    ys__n21368, ys__n21370, ys__n21372, ys__n21374, ys__n21376, ys__n21378,
    ys__n21380, ys__n21382, ys__n21384, ys__n21386, ys__n21388, ys__n21390,
    ys__n21392, ys__n21394, ys__n21396, ys__n21398, ys__n21400, ys__n21402,
    ys__n21404, ys__n21405, ys__n21406, ys__n21407, ys__n21408, ys__n21409,
    ys__n21410, ys__n21411, ys__n21412, ys__n21413, ys__n21414, ys__n21415,
    ys__n21416, ys__n21417, ys__n21418, ys__n21419, ys__n21420, ys__n21421,
    ys__n21422, ys__n21423, ys__n21424, ys__n21425, ys__n21426, ys__n21427,
    ys__n21428, ys__n21429, ys__n21430, ys__n21431, ys__n21432, ys__n21433,
    ys__n21434, ys__n21435, ys__n21500, ys__n21502, ys__n21504, ys__n21506,
    ys__n21508, ys__n21510, ys__n21512, ys__n21514, ys__n21516, ys__n21518,
    ys__n21520, ys__n21522, ys__n21524, ys__n21526, ys__n21528, ys__n21530,
    ys__n21532, ys__n21534, ys__n21536, ys__n21538, ys__n21540, ys__n21542,
    ys__n21544, ys__n21546, ys__n21548, ys__n21550, ys__n21552, ys__n21554,
    ys__n21556, ys__n21558, ys__n21560, ys__n21562, ys__n21564, ys__n21566,
    ys__n21568, ys__n21570, ys__n21572, ys__n21574, ys__n21576, ys__n21578,
    ys__n21580, ys__n21582, ys__n21584, ys__n21586, ys__n21588, ys__n21590,
    ys__n21592, ys__n21594, ys__n21596, ys__n21598, ys__n21600, ys__n21602,
    ys__n21604, ys__n21606, ys__n21608, ys__n21610, ys__n21612, ys__n21614,
    ys__n21616, ys__n21618, ys__n21620, ys__n21622, ys__n21624, ys__n21626,
    ys__n21628, ys__n21630, ys__n21632, ys__n21634, ys__n21636, ys__n21638,
    ys__n21640, ys__n21642, ys__n21644, ys__n21646, ys__n21648, ys__n21650,
    ys__n21652, ys__n21654, ys__n21656, ys__n21658, ys__n21660, ys__n21662,
    ys__n21664, ys__n21666, ys__n21668, ys__n21670, ys__n21672, ys__n21674,
    ys__n21676, ys__n21678, ys__n21680, ys__n21682, ys__n21684, ys__n21686,
    ys__n21688, ys__n21690, ys__n21692, ys__n21694, ys__n21696, ys__n21698,
    ys__n21700, ys__n21702, ys__n21704, ys__n21706, ys__n21708, ys__n21710,
    ys__n21712, ys__n21714, ys__n21716, ys__n21718, ys__n21720, ys__n21722,
    ys__n21724, ys__n21726, ys__n21728, ys__n21730, ys__n21732, ys__n21734,
    ys__n21736, ys__n21738, ys__n21740, ys__n21742, ys__n21744, ys__n21746,
    ys__n21748, ys__n21750, ys__n21752, ys__n21754, ys__n21756, ys__n21758,
    ys__n21760, ys__n21762, ys__n21764, ys__n21766, ys__n21768, ys__n21770,
    ys__n21772, ys__n21774, ys__n21776, ys__n21778, ys__n21780, ys__n21782,
    ys__n21784, ys__n21786, ys__n21788, ys__n21790, ys__n21792, ys__n21794,
    ys__n21796, ys__n21798, ys__n21800, ys__n21802, ys__n21804, ys__n21806,
    ys__n21808, ys__n21810, ys__n21812, ys__n21814, ys__n21816, ys__n21818,
    ys__n21820, ys__n21822, ys__n21824, ys__n21826, ys__n21828, ys__n21830,
    ys__n21832, ys__n21834, ys__n21836, ys__n21838, ys__n21840, ys__n21842,
    ys__n21844, ys__n21846, ys__n21848, ys__n21850, ys__n21852, ys__n21854,
    ys__n21856, ys__n21858, ys__n21860, ys__n21862, ys__n21864, ys__n21866,
    ys__n21868, ys__n21870, ys__n21872, ys__n21874, ys__n21876, ys__n21878,
    ys__n21880, ys__n21882, ys__n21884, ys__n21886, ys__n21888, ys__n21890,
    ys__n21892, ys__n21894, ys__n21896, ys__n21898, ys__n21900, ys__n21902,
    ys__n21904, ys__n21906, ys__n21908, ys__n21910, ys__n21912, ys__n21914,
    ys__n21916, ys__n21918, ys__n21920, ys__n21922, ys__n21924, ys__n21926,
    ys__n21928, ys__n21930, ys__n21932, ys__n21934, ys__n21936, ys__n21938,
    ys__n21940, ys__n21942, ys__n21944, ys__n21946, ys__n21948, ys__n21949,
    ys__n21950, ys__n21951, ys__n21952, ys__n21953, ys__n21954, ys__n21955,
    ys__n21956, ys__n21957, ys__n21958, ys__n21959, ys__n21960, ys__n21961,
    ys__n21962, ys__n21963, ys__n21964, ys__n21965, ys__n21966, ys__n21967,
    ys__n21968, ys__n21969, ys__n21970, ys__n21971, ys__n21972, ys__n21973,
    ys__n21974, ys__n21975, ys__n21976, ys__n21977, ys__n21978, ys__n21979,
    ys__n21980, ys__n21982, ys__n21984, ys__n21986, ys__n21988, ys__n21990,
    ys__n21992, ys__n21994, ys__n21996, ys__n21998, ys__n22000, ys__n22002,
    ys__n22004, ys__n22006, ys__n22008, ys__n22010, ys__n22012, ys__n22014,
    ys__n22016, ys__n22018, ys__n22020, ys__n22022, ys__n22024, ys__n22026,
    ys__n22028, ys__n22030, ys__n22032, ys__n22034, ys__n22036, ys__n22038,
    ys__n22040, ys__n22042, ys__n22044, ys__n22046, ys__n22048, ys__n22050,
    ys__n22052, ys__n22054, ys__n22056, ys__n22058, ys__n22060, ys__n22062,
    ys__n22064, ys__n22066, ys__n22068, ys__n22070, ys__n22072, ys__n22074,
    ys__n22076, ys__n22078, ys__n22080, ys__n22082, ys__n22084, ys__n22086,
    ys__n22088, ys__n22090, ys__n22092, ys__n22094, ys__n22096, ys__n22098,
    ys__n22100, ys__n22102, ys__n22104, ys__n22106, ys__n22108, ys__n22110,
    ys__n22112, ys__n22114, ys__n22116, ys__n22118, ys__n22120, ys__n22122,
    ys__n22124, ys__n22126, ys__n22128, ys__n22130, ys__n22132, ys__n22134,
    ys__n22136, ys__n22138, ys__n22140, ys__n22142, ys__n22144, ys__n22146,
    ys__n22148, ys__n22150, ys__n22152, ys__n22154, ys__n22156, ys__n22158,
    ys__n22160, ys__n22162, ys__n22164, ys__n22166, ys__n22168, ys__n22170,
    ys__n22172, ys__n22174, ys__n22176, ys__n22178, ys__n22180, ys__n22182,
    ys__n22184, ys__n22186, ys__n22188, ys__n22190, ys__n22192, ys__n22194,
    ys__n22196, ys__n22198, ys__n22200, ys__n22202, ys__n22204, ys__n22206,
    ys__n22208, ys__n22210, ys__n22212, ys__n22214, ys__n22216, ys__n22218,
    ys__n22220, ys__n22222, ys__n22224, ys__n22226, ys__n22228, ys__n22230,
    ys__n22232, ys__n22234, ys__n22236, ys__n22238, ys__n22240, ys__n22242,
    ys__n22244, ys__n22246, ys__n22248, ys__n22250, ys__n22252, ys__n22254,
    ys__n22256, ys__n22258, ys__n22260, ys__n22262, ys__n22264, ys__n22266,
    ys__n22268, ys__n22270, ys__n22272, ys__n22274, ys__n22276, ys__n22278,
    ys__n22280, ys__n22282, ys__n22284, ys__n22286, ys__n22288, ys__n22290,
    ys__n22292, ys__n22294, ys__n22296, ys__n22298, ys__n22300, ys__n22302,
    ys__n22304, ys__n22306, ys__n22308, ys__n22310, ys__n22312, ys__n22314,
    ys__n22316, ys__n22318, ys__n22320, ys__n22322, ys__n22324, ys__n22326,
    ys__n22328, ys__n22330, ys__n22332, ys__n22334, ys__n22336, ys__n22338,
    ys__n22340, ys__n22342, ys__n22344, ys__n22346, ys__n22348, ys__n22350,
    ys__n22352, ys__n22354, ys__n22356, ys__n22358, ys__n22360, ys__n22362,
    ys__n22364, ys__n22366, ys__n22368, ys__n22370, ys__n22372, ys__n22374,
    ys__n22376, ys__n22378, ys__n22380, ys__n22382, ys__n22384, ys__n22386,
    ys__n22388, ys__n22390, ys__n22392, ys__n22394, ys__n22396, ys__n22398,
    ys__n22400, ys__n22402, ys__n22404, ys__n22406, ys__n22408, ys__n22410,
    ys__n22412, ys__n22414, ys__n22416, ys__n22418, ys__n22420, ys__n22422,
    ys__n22424, ys__n22426, ys__n22428, ys__n22429, ys__n22430, ys__n22431,
    ys__n22432, ys__n22433, ys__n22434, ys__n22435, ys__n22436, ys__n22437,
    ys__n22438, ys__n22439, ys__n22440, ys__n22441, ys__n22442, ys__n22443,
    ys__n22444, ys__n22445, ys__n22446, ys__n22447, ys__n22448, ys__n22449,
    ys__n22450, ys__n22451, ys__n22452, ys__n22453, ys__n22454, ys__n22455,
    ys__n22456, ys__n22457, ys__n22458, ys__n22459, ys__n22464, ys__n22465,
    ys__n22564, ys__n22566, ys__n22568, ys__n22570, ys__n22572, ys__n22574,
    ys__n22576, ys__n22578, ys__n22580, ys__n22582, ys__n22584, ys__n22586,
    ys__n22588, ys__n22590, ys__n22592, ys__n22594, ys__n22596, ys__n22598,
    ys__n22600, ys__n22602, ys__n22604, ys__n22606, ys__n22608, ys__n22610,
    ys__n22612, ys__n22614, ys__n22616, ys__n22618, ys__n22620, ys__n22622,
    ys__n22624, ys__n22626, ys__n22630, ys__n22632, ys__n22634, ys__n22636,
    ys__n22640, ys__n22642, ys__n22644, ys__n22646, ys__n22648, ys__n22650,
    ys__n22652, ys__n22654, ys__n22668, ys__n22670, ys__n22673, ys__n22675,
    ys__n22677, ys__n22679, ys__n22681, ys__n22683, ys__n22685, ys__n22687,
    ys__n22689, ys__n22715, ys__n22717, ys__n22719, ys__n22721, ys__n22723,
    ys__n22725, ys__n22727, ys__n22729, ys__n22731, ys__n22733, ys__n22735,
    ys__n22737, ys__n22739, ys__n22741, ys__n22743, ys__n22745, ys__n22747,
    ys__n22749, ys__n22751, ys__n22753, ys__n22755, ys__n22757, ys__n22759,
    ys__n22761, ys__n22763, ys__n22765, ys__n22767, ys__n22769, ys__n22771,
    ys__n22773, ys__n22775, ys__n22777, ys__n22779, ys__n22781, ys__n22783,
    ys__n22785, ys__n22787, ys__n22789, ys__n22792, ys__n22794, ys__n22799,
    ys__n22818, ys__n22820, ys__n22822, ys__n22824, ys__n22826, ys__n22828,
    ys__n22830, ys__n22832, ys__n22834, ys__n22836, ys__n22838, ys__n22840,
    ys__n22842, ys__n22844, ys__n22846, ys__n22848, ys__n22850, ys__n22852,
    ys__n22854, ys__n22856, ys__n22858, ys__n22860, ys__n22862, ys__n22864,
    ys__n22866, ys__n22868, ys__n22870, ys__n22872, ys__n22874, ys__n22876,
    ys__n22878, ys__n22880, ys__n22882, ys__n22884, ys__n22885, ys__n22886,
    ys__n22887, ys__n22888, ys__n22889, ys__n22890, ys__n22891, ys__n22892,
    ys__n22893, ys__n22894, ys__n22895, ys__n22896, ys__n22897, ys__n22898,
    ys__n22899, ys__n22900, ys__n22901, ys__n22902, ys__n22903, ys__n22904,
    ys__n22905, ys__n22906, ys__n22907, ys__n22908, ys__n22909, ys__n22910,
    ys__n22911, ys__n22912, ys__n22913, ys__n22914, ys__n22915, ys__n22916,
    ys__n22918, ys__n22921, ys__n22924, ys__n22927, ys__n22930, ys__n22933,
    ys__n22936, ys__n22939, ys__n22942, ys__n22945, ys__n22948, ys__n22951,
    ys__n22954, ys__n22957, ys__n22960, ys__n22963, ys__n22966, ys__n22969,
    ys__n22972, ys__n22975, ys__n22978, ys__n22981, ys__n22984, ys__n22987,
    ys__n22990, ys__n22993, ys__n22996, ys__n22999, ys__n23002, ys__n23005,
    ys__n23008, ys__n23011, ys__n23014, ys__n23016, ys__n23018, ys__n23020,
    ys__n23022, ys__n23024, ys__n23026, ys__n23028, ys__n23030, ys__n23032,
    ys__n23034, ys__n23036, ys__n23038, ys__n23040, ys__n23042, ys__n23044,
    ys__n23046, ys__n23048, ys__n23050, ys__n23052, ys__n23054, ys__n23056,
    ys__n23058, ys__n23060, ys__n23062, ys__n23064, ys__n23066, ys__n23068,
    ys__n23070, ys__n23072, ys__n23074, ys__n23076, ys__n23077, ys__n23078,
    ys__n23079, ys__n23080, ys__n23081, ys__n23082, ys__n23083, ys__n23084,
    ys__n23085, ys__n23086, ys__n23087, ys__n23088, ys__n23089, ys__n23090,
    ys__n23091, ys__n23092, ys__n23093, ys__n23094, ys__n23095, ys__n23096,
    ys__n23097, ys__n23098, ys__n23099, ys__n23100, ys__n23101, ys__n23102,
    ys__n23103, ys__n23104, ys__n23105, ys__n23106, ys__n23107, ys__n23108,
    ys__n23111, ys__n23114, ys__n23117, ys__n23120, ys__n23123, ys__n23126,
    ys__n23129, ys__n23132, ys__n23135, ys__n23138, ys__n23141, ys__n23144,
    ys__n23147, ys__n23150, ys__n23153, ys__n23156, ys__n23159, ys__n23162,
    ys__n23165, ys__n23168, ys__n23171, ys__n23174, ys__n23177, ys__n23180,
    ys__n23183, ys__n23186, ys__n23189, ys__n23192, ys__n23195, ys__n23198,
    ys__n23203, ys__n23205, ys__n23207, ys__n23209, ys__n23211, ys__n23213,
    ys__n23215, ys__n23217, ys__n23219, ys__n23221, ys__n23223, ys__n23225,
    ys__n23227, ys__n23229, ys__n23231, ys__n23233, ys__n23235, ys__n23237,
    ys__n23239, ys__n23241, ys__n23243, ys__n23245, ys__n23247, ys__n23249,
    ys__n23251, ys__n23253, ys__n23255, ys__n23257, ys__n23259, ys__n23261,
    ys__n23269, ys__n23271, ys__n23272, ys__n23274, ys__n23276, ys__n23278,
    ys__n23280, ys__n23282, ys__n23284, ys__n23286, ys__n23288, ys__n23290,
    ys__n23292, ys__n23294, ys__n23296, ys__n23298, ys__n23300, ys__n23302,
    ys__n23304, ys__n23306, ys__n23308, ys__n23310, ys__n23312, ys__n23314,
    ys__n23316, ys__n23318, ys__n23320, ys__n23322, ys__n23324, ys__n23326,
    ys__n23328, ys__n23330, ys__n23332, ys__n23335, ys__n23339, ys__n23480,
    ys__n23548, ys__n23550, ys__n23552, ys__n23554, ys__n23556, ys__n23558,
    ys__n23560, ys__n23562, ys__n23564, ys__n23566, ys__n23568, ys__n23570,
    ys__n23572, ys__n23574, ys__n23627, ys__n23629, ys__n23641, ys__n23644,
    ys__n23645, ys__n23647, ys__n23650, ys__n23652, ys__n23655, ys__n23658,
    ys__n23661, ys__n23663, ys__n23705, ys__n23706, ys__n23707, ys__n23708,
    ys__n23709, ys__n23710, ys__n23711, ys__n23712, ys__n23713, ys__n23714,
    ys__n23715, ys__n23717, ys__n23729, ys__n23730, ys__n23763, ys__n23818,
    ys__n23819, ys__n23820, ys__n23821, ys__n23822, ys__n23834, ys__n23836,
    ys__n23838, ys__n23840, ys__n23842, ys__n23850, ys__n23888, ys__n23889,
    ys__n23890, ys__n23891, ys__n23892, ys__n23904, ys__n23906, ys__n23908,
    ys__n23910, ys__n23912, ys__n23956, ys__n23957, ys__n23958, ys__n23959,
    ys__n23960, ys__n23977, ys__n23979, ys__n23981, ys__n23983, ys__n23985,
    ys__n24106, ys__n24107, ys__n24108, ys__n24112, ys__n24123, ys__n24124,
    ys__n24131, ys__n24143, ys__n24158, ys__n24167, ys__n24168, ys__n24177,
    ys__n24197, ys__n24199, ys__n24201, ys__n24203, ys__n24205, ys__n24207,
    ys__n24209, ys__n24211, ys__n24213, ys__n24215, ys__n24217, ys__n24219,
    ys__n24228, ys__n24233, ys__n24235, ys__n24243, ys__n24248, ys__n24279,
    ys__n24280, ys__n24303, ys__n24306, ys__n24308, ys__n24310, ys__n24312,
    ys__n24314, ys__n24316, ys__n24318, ys__n24337, ys__n24340, ys__n24342,
    ys__n24344, ys__n24346, ys__n24348, ys__n24350, ys__n24352, ys__n24371,
    ys__n24374, ys__n24376, ys__n24378, ys__n24380, ys__n24382, ys__n24384,
    ys__n24386, ys__n24389, ys__n24406, ys__n24409, ys__n24411, ys__n24413,
    ys__n24415, ys__n24417, ys__n24419, ys__n24421, ys__n24427, ys__n24433,
    ys__n24434, ys__n24461, ys__n24463, ys__n24464, ys__n24483, ys__n24485,
    ys__n24506, ys__n24519, ys__n24567, ys__n24575, ys__n24578, ys__n24590,
    ys__n24591, ys__n24615, ys__n24616, ys__n24617, ys__n24618, ys__n24619,
    ys__n24620, ys__n24621, ys__n24622, ys__n24623, ys__n24624, ys__n24625,
    ys__n24626, ys__n24627, ys__n24628, ys__n24629, ys__n24630, ys__n24631,
    ys__n24632, ys__n24633, ys__n24634, ys__n24635, ys__n24636, ys__n24637,
    ys__n24638, ys__n24639, ys__n24640, ys__n24641, ys__n24642, ys__n24643,
    ys__n24644, ys__n24645, ys__n24646, ys__n24647, ys__n24648, ys__n24649,
    ys__n24650, ys__n24651, ys__n24652, ys__n24653, ys__n24654, ys__n24655,
    ys__n24656, ys__n24657, ys__n24658, ys__n24659, ys__n24660, ys__n24661,
    ys__n24662, ys__n24663, ys__n24664, ys__n24665, ys__n24666, ys__n24667,
    ys__n24668, ys__n24669, ys__n24670, ys__n24671, ys__n24672, ys__n24673,
    ys__n24674, ys__n24675, ys__n24677, ys__n24679, ys__n24681, ys__n24683,
    ys__n24684, ys__n24685, ys__n24686, ys__n24687, ys__n24688, ys__n24689,
    ys__n24690, ys__n24691, ys__n24692, ys__n24693, ys__n24694, ys__n24695,
    ys__n24696, ys__n24697, ys__n24698, ys__n24699, ys__n24700, ys__n24701,
    ys__n24702, ys__n24703, ys__n24704, ys__n24705, ys__n24706, ys__n24707,
    ys__n24708, ys__n24709, ys__n24710, ys__n24711, ys__n24712, ys__n24741,
    ys__n24744, ys__n24747, ys__n24750, ys__n24753, ys__n24756, ys__n24759,
    ys__n24762, ys__n24765, ys__n24768, ys__n24771, ys__n24774, ys__n24777,
    ys__n24780, ys__n24783, ys__n24786, ys__n24789, ys__n24792, ys__n24795,
    ys__n24798, ys__n24801, ys__n24804, ys__n24807, ys__n24810, ys__n24813,
    ys__n24816, ys__n24819, ys__n24822, ys__n24825, ys__n24828, ys__n24831,
    ys__n24834, ys__n25292, ys__n25300, ys__n25381, ys__n25382, ys__n25383,
    ys__n25384, ys__n25470, ys__n25564, ys__n25567, ys__n25570, ys__n25573,
    ys__n25576, ys__n25579, ys__n25582, ys__n25585, ys__n25588, ys__n25591,
    ys__n25594, ys__n25597, ys__n25600, ys__n25603, ys__n25606, ys__n25609,
    ys__n25612, ys__n25615, ys__n25618, ys__n25621, ys__n25624, ys__n25627,
    ys__n25630, ys__n25633, ys__n25636, ys__n25639, ys__n25642, ys__n25645,
    ys__n25648, ys__n25651, ys__n25654, ys__n25657, ys__n25727, ys__n25730,
    ys__n25733, ys__n25736, ys__n25853, ys__n25856, ys__n25859, ys__n25862,
    ys__n25980, ys__n25984, ys__n25987, ys__n25990, ys__n25993, ys__n25996,
    ys__n25999, ys__n26002, ys__n26005, ys__n26008, ys__n26011, ys__n26014,
    ys__n26017, ys__n26020, ys__n26023, ys__n26026, ys__n26029, ys__n26032,
    ys__n26035, ys__n26038, ys__n26041, ys__n26044, ys__n26047, ys__n26050,
    ys__n26053, ys__n26056, ys__n26059, ys__n26062, ys__n26065, ys__n26068,
    ys__n26071, ys__n26074, ys__n26143, ys__n26145, ys__n26147, ys__n26149,
    ys__n26151, ys__n26153, ys__n26155, ys__n26157, ys__n26159, ys__n26161,
    ys__n26162, ys__n26164, ys__n26166, ys__n26168, ys__n26170, ys__n26172,
    ys__n26174, ys__n26176, ys__n26178, ys__n26180, ys__n26182, ys__n26184,
    ys__n26186, ys__n26188, ys__n26190, ys__n26192, ys__n26194, ys__n26196,
    ys__n26198, ys__n26200, ys__n26202, ys__n26204, ys__n26206, ys__n26208,
    ys__n26210, ys__n26212, ys__n26214, ys__n26216, ys__n26218, ys__n26279,
    ys__n26285, ys__n26359, ys__n26362, ys__n26425, ys__n26428, ys__n26431,
    ys__n26434, ys__n26437, ys__n26440, ys__n26443, ys__n26446, ys__n26449,
    ys__n26452, ys__n26455, ys__n26460, ys__n26463, ys__n26466, ys__n26469,
    ys__n26472, ys__n26475, ys__n26478, ys__n26481, ys__n26484, ys__n26487,
    ys__n26490, ys__n26493, ys__n26496, ys__n26499, ys__n26502, ys__n26505,
    ys__n26508, ys__n26511, ys__n26514, ys__n26517, ys__n26552, ys__n26553,
    ys__n26554, ys__n26556, ys__n26557, ys__n26558, ys__n26559, ys__n26560,
    ys__n26561, ys__n26562, ys__n26563, ys__n26564, ys__n26565, ys__n26567,
    ys__n26568, ys__n26569, ys__n26570, ys__n26571, ys__n26572, ys__n26766,
    ys__n26768, ys__n26770, ys__n26772, ys__n27479, ys__n27481, ys__n27485,
    ys__n27488, ys__n27496, ys__n27498, ys__n27499, ys__n27507, ys__n27509,
    ys__n27510, ys__n27518, ys__n27520, ys__n27607, ys__n27608, ys__n27611,
    ys__n27612, ys__n27614, ys__n27615, ys__n27617, ys__n27618, ys__n27620,
    ys__n27621, ys__n27623, ys__n27624, ys__n27626, ys__n27627, ys__n27629,
    ys__n27630, ys__n27632, ys__n27633, ys__n27635, ys__n27636, ys__n27638,
    ys__n27639, ys__n27641, ys__n27642, ys__n27644, ys__n27645, ys__n27647,
    ys__n27648, ys__n27650, ys__n27651, ys__n27653, ys__n27654, ys__n27656,
    ys__n27657, ys__n27659, ys__n27660, ys__n27662, ys__n27663, ys__n27665,
    ys__n27666, ys__n27668, ys__n27669, ys__n27671, ys__n27672, ys__n27674,
    ys__n27675, ys__n27677, ys__n27678, ys__n27680, ys__n27681, ys__n27683,
    ys__n27684, ys__n27686, ys__n27687, ys__n27689, ys__n27690, ys__n27692,
    ys__n27693, ys__n27695, ys__n27696, ys__n27698, ys__n27699, ys__n27701,
    ys__n27702, ys__n27737, ys__n27738, ys__n27740, ys__n27743, ys__n27747,
    ys__n27750, ys__n27753, ys__n27756, ys__n27759, ys__n27762, ys__n27765,
    ys__n27768, ys__n27771, ys__n27774, ys__n27777, ys__n27780, ys__n27783,
    ys__n27786, ys__n27789, ys__n27792, ys__n27795, ys__n27798, ys__n27801,
    ys__n27804, ys__n27807, ys__n27810, ys__n27813, ys__n27816, ys__n27819,
    ys__n27822, ys__n27825, ys__n27828, ys__n27831, ys__n27834, ys__n27837,
    ys__n27855, ys__n27857, ys__n27859, ys__n27861, ys__n27863, ys__n27865,
    ys__n27867, ys__n27869, ys__n27871, ys__n27873, ys__n27875, ys__n27877,
    ys__n27879, ys__n27881, ys__n27883, ys__n27885, ys__n28015, ys__n28016,
    ys__n28017, ys__n28018, ys__n28019, ys__n28020, ys__n28021, ys__n28022,
    ys__n28023, ys__n28024, ys__n28025, ys__n28026, ys__n28027, ys__n28028,
    ys__n28029, ys__n28030, ys__n28243, ys__n28287, ys__n28288, ys__n28290,
    ys__n28292, ys__n28294, ys__n28296, ys__n28424, ys__n28426, ys__n28428,
    ys__n28430, ys__n28432, ys__n28434, ys__n28436, ys__n28438, ys__n28446,
    ys__n28453, ys__n28455, ys__n28457, ys__n28459, ys__n28462, ys__n28464,
    ys__n28466, ys__n28468, ys__n28470, ys__n28472, ys__n28632, ys__n28633,
    ys__n28634, ys__n28635, ys__n28636, ys__n28637, ys__n28638, ys__n28639,
    ys__n28640, ys__n28641, ys__n28718, ys__n28719, ys__n28720, ys__n28859,
    ys__n28863, ys__n28866, ys__n28869, ys__n28872, ys__n28875, ys__n28878,
    ys__n28881, ys__n28884, ys__n28887, ys__n28890, ys__n28893, ys__n28896,
    ys__n28899, ys__n28902, ys__n28905, ys__n28908, ys__n28911, ys__n28914,
    ys__n28917, ys__n28920, ys__n28923, ys__n28926, ys__n28929, ys__n28932,
    ys__n28935, ys__n28938, ys__n28941, ys__n28944, ys__n28947, ys__n28950,
    ys__n28953, ys__n29117, ys__n29119, ys__n29120, ys__n29121, ys__n29123,
    ys__n29124, ys__n29126, ys__n29127, ys__n29129, ys__n29130, ys__n29132,
    ys__n29133, ys__n29135, ys__n29136, ys__n29138, ys__n29139, ys__n29141,
    ys__n29142, ys__n29144, ys__n29145, ys__n29147, ys__n29148, ys__n29150,
    ys__n29151, ys__n29153, ys__n29154, ys__n29156, ys__n29157, ys__n29159,
    ys__n29160, ys__n29162, ys__n29163, ys__n29165, ys__n29166, ys__n29168,
    ys__n29169, ys__n29171, ys__n29172, ys__n29174, ys__n29175, ys__n29177,
    ys__n29178, ys__n29180, ys__n29181, ys__n29183, ys__n29184, ys__n29186,
    ys__n29187, ys__n29189, ys__n29190, ys__n29192, ys__n29193, ys__n29195,
    ys__n29196, ys__n29198, ys__n29199, ys__n29201, ys__n29202, ys__n29204,
    ys__n29205, ys__n29207, ys__n29208, ys__n29210, ys__n29211, ys__n29213,
    ys__n29214, ys__n29218, ys__n29220, ys__n29224, ys__n29237, ys__n29240,
    ys__n29242, ys__n29244, ys__n29246, ys__n29248, ys__n29250, ys__n29252,
    ys__n29254, ys__n29256, ys__n29258, ys__n29260, ys__n29262, ys__n29264,
    ys__n29266, ys__n29268, ys__n29270, ys__n29272, ys__n29274, ys__n29276,
    ys__n29278, ys__n29280, ys__n29282, ys__n29284, ys__n29286, ys__n29288,
    ys__n29290, ys__n29292, ys__n29294, ys__n29296, ys__n29298, ys__n29300,
    ys__n29432, ys__n29433, ys__n29434, ys__n29436, ys__n29437, ys__n29439,
    ys__n29440, ys__n29442, ys__n29443, ys__n29445, ys__n29446, ys__n29448,
    ys__n29449, ys__n29451, ys__n29452, ys__n29454, ys__n29455, ys__n29457,
    ys__n29458, ys__n29460, ys__n29461, ys__n29463, ys__n29464, ys__n29466,
    ys__n29467, ys__n29469, ys__n29470, ys__n29472, ys__n29473, ys__n29475,
    ys__n29476, ys__n29478, ys__n29479, ys__n29481, ys__n29482, ys__n29484,
    ys__n29485, ys__n29487, ys__n29488, ys__n29490, ys__n29491, ys__n29493,
    ys__n29494, ys__n29496, ys__n29497, ys__n29499, ys__n29500, ys__n29502,
    ys__n29503, ys__n29505, ys__n29506, ys__n29508, ys__n29509, ys__n29511,
    ys__n29512, ys__n29514, ys__n29515, ys__n29517, ys__n29518, ys__n29520,
    ys__n29521, ys__n29523, ys__n29524, ys__n29526, ys__n29527, ys__n29531,
    ys__n29533, ys__n29537, ys__n29550, ys__n29552, ys__n29553, ys__n29554,
    ys__n29555, ys__n29556, ys__n29557, ys__n29558, ys__n29559, ys__n29560,
    ys__n29561, ys__n29562, ys__n29563, ys__n29564, ys__n29565, ys__n29566,
    ys__n29567, ys__n29568, ys__n29569, ys__n29570, ys__n29571, ys__n29572,
    ys__n29573, ys__n29574, ys__n29575, ys__n29576, ys__n29577, ys__n29578,
    ys__n29579, ys__n29580, ys__n29581, ys__n29582, ys__n29583, ys__n29584,
    ys__n29585, ys__n29586, ys__n29587, ys__n29588, ys__n29589, ys__n29590,
    ys__n29591, ys__n29592, ys__n29593, ys__n29594, ys__n29595, ys__n29596,
    ys__n29597, ys__n29598, ys__n29599, ys__n29600, ys__n29601, ys__n29602,
    ys__n29603, ys__n29604, ys__n29605, ys__n29606, ys__n29607, ys__n29608,
    ys__n29707, ys__n29708, ys__n29709, ys__n29711, ys__n29712, ys__n29714,
    ys__n29715, ys__n29717, ys__n29718, ys__n29720, ys__n29721, ys__n29723,
    ys__n29724, ys__n29726, ys__n29727, ys__n29729, ys__n29730, ys__n29732,
    ys__n29733, ys__n29735, ys__n29736, ys__n29738, ys__n29739, ys__n29741,
    ys__n29742, ys__n29744, ys__n29745, ys__n29747, ys__n29748, ys__n29750,
    ys__n29751, ys__n29753, ys__n29754, ys__n29756, ys__n29757, ys__n29759,
    ys__n29760, ys__n29762, ys__n29763, ys__n29765, ys__n29766, ys__n29768,
    ys__n29769, ys__n29771, ys__n29772, ys__n29774, ys__n29775, ys__n29777,
    ys__n29778, ys__n29780, ys__n29781, ys__n29783, ys__n29784, ys__n29786,
    ys__n29787, ys__n29789, ys__n29790, ys__n29792, ys__n29793, ys__n29795,
    ys__n29796, ys__n29798, ys__n29799, ys__n29801, ys__n29802, ys__n29806,
    ys__n29808, ys__n29812, ys__n29846, ys__n29880, ys__n29881, ys__n29883,
    ys__n29884, ys__n29885, ys__n29886, ys__n29887, ys__n29888, ys__n29889,
    ys__n29890, ys__n29891, ys__n29892, ys__n29893, ys__n29894, ys__n29895,
    ys__n29896, ys__n29897, ys__n29898, ys__n29899, ys__n29900, ys__n29901,
    ys__n29902, ys__n29903, ys__n29904, ys__n29905, ys__n29906, ys__n29907,
    ys__n29908, ys__n29909, ys__n29910, ys__n29911, ys__n29912, ys__n29913,
    ys__n30011, ys__n30014, ys__n30016, ys__n30018, ys__n30020, ys__n30022,
    ys__n30024, ys__n30026, ys__n30028, ys__n30030, ys__n30032, ys__n30034,
    ys__n30036, ys__n30038, ys__n30040, ys__n30042, ys__n30044, ys__n30046,
    ys__n30048, ys__n30050, ys__n30052, ys__n30054, ys__n30056, ys__n30058,
    ys__n30060, ys__n30062, ys__n30064, ys__n30066, ys__n30068, ys__n30070,
    ys__n30072, ys__n30074, ys__n30214, ys__n30216, ys__n30217, ys__n30219,
    ys__n30220, ys__n30225, ys__n30230, ys__n30232, ys__n30333, ys__n30334,
    ys__n30553, ys__n30815, ys__n30816, ys__n30818, ys__n30819, ys__n30820,
    ys__n30837, ys__n30861, ys__n30862, ys__n30863, ys__n30865, ys__n30867,
    ys__n30869, ys__n30871, ys__n30877, ys__n30879, ys__n30881, ys__n30883,
    ys__n30885, ys__n30887, ys__n30889, ys__n30891, ys__n30893, ys__n30895,
    ys__n30897, ys__n30899, ys__n30901, ys__n30903, ys__n30905, ys__n30907,
    ys__n30909, ys__n30911, ys__n30913, ys__n30915, ys__n30917, ys__n30919,
    ys__n30921, ys__n30923, ys__n30925, ys__n30927, ys__n30929, ys__n30931,
    ys__n30933, ys__n30935, ys__n30937, ys__n30939, ys__n30941, ys__n30957,
    ys__n30960, ys__n30961, ys__n30962, ys__n30974, ys__n31031, ys__n33212,
    ys__n33214, ys__n33216, ys__n33218, ys__n33220, ys__n33222, ys__n33259,
    ys__n33261, ys__n33263, ys__n33265, ys__n33267, ys__n33269, ys__n33272,
    ys__n33274, ys__n33276, ys__n33278, ys__n33300, ys__n33309, ys__n33311,
    ys__n33313, ys__n33318, ys__n33320, ys__n33328, ys__n33330, ys__n33332,
    ys__n33334, ys__n33336, ys__n33338, ys__n33340, ys__n33342, ys__n33350,
    ys__n33352, ys__n33359, ys__n33364, ys__n33370, ys__n33375, ys__n33380,
    ys__n33384, ys__n33386, ys__n33389, ys__n33394, ys__n33396, ys__n33398,
    ys__n33403, ys__n33407, ys__n33409, ys__n33411, ys__n33423, ys__n33431,
    ys__n33442, ys__n33451, ys__n33464, ys__n33469, ys__n33471, ys__n33473,
    ys__n33475, ys__n33479, ys__n33481, ys__n33488, ys__n33491, ys__n33493,
    ys__n33495, ys__n33497, ys__n33499, ys__n33509, ys__n33511, ys__n33522,
    ys__n33532, ys__n33541, ys__n33545, ys__n33548, ys__n33552, ys__n33558,
    ys__n33563, ys__n33564, ys__n33566, ys__n33568, ys__n33570, ys__n33572,
    ys__n33574, ys__n33576, ys__n33579, ys__n33581, ys__n33614, ys__n33632,
    ys__n33634, ys__n33636, ys__n33638, ys__n33640, ys__n33642, ys__n33644,
    ys__n33646, ys__n33648, ys__n33650, ys__n33652, ys__n33654, ys__n33656,
    ys__n33658, ys__n33660, ys__n33662, ys__n33664, ys__n33666, ys__n33668,
    ys__n33670, ys__n33672, ys__n33674, ys__n33676, ys__n33678, ys__n33681,
    ys__n33683, ys__n33685, ys__n33687, ys__n33689, ys__n33691, ys__n33693,
    ys__n33695, ys__n33697, ys__n33699, ys__n33701, ys__n33703, ys__n33705,
    ys__n33707, ys__n33709, ys__n33711, ys__n33713, ys__n33715, ys__n33717,
    ys__n33719, ys__n33721, ys__n33723, ys__n33725, ys__n33727, ys__n33729,
    ys__n33731, ys__n33733, ys__n33735, ys__n33737, ys__n33739, ys__n33741,
    ys__n33743, ys__n33745, ys__n33747, ys__n33749, ys__n34666, ys__n34668,
    ys__n34670, ys__n34672, ys__n34674, ys__n34676, ys__n34678, ys__n34680,
    ys__n34682, ys__n34684, ys__n34686, ys__n34688, ys__n34690, ys__n34692,
    ys__n34694, ys__n34696, ys__n34698, ys__n34700, ys__n34702, ys__n34704,
    ys__n34706, ys__n34708, ys__n34710, ys__n34712, ys__n34714, ys__n34716,
    ys__n34718, ys__n34720, ys__n34722, ys__n34724, ys__n34726, ys__n34728,
    ys__n34730, ys__n34732, ys__n34734, ys__n34736, ys__n34738, ys__n34740,
    ys__n34742, ys__n34744, ys__n34746, ys__n34748, ys__n34750, ys__n34752,
    ys__n34754, ys__n34756, ys__n34758, ys__n34760, ys__n34762, ys__n34764,
    ys__n34766, ys__n34768, ys__n34770, ys__n34772, ys__n34774, ys__n34776,
    ys__n34778, ys__n34780, ys__n34782, ys__n34784, ys__n34786, ys__n34788,
    ys__n34790, ys__n34792, ys__n34794, ys__n34796, ys__n34798, ys__n34800,
    ys__n34802, ys__n34804, ys__n34806, ys__n34808, ys__n34810, ys__n34812,
    ys__n34814, ys__n34816, ys__n34818, ys__n34820, ys__n34822, ys__n34824,
    ys__n34826, ys__n34828, ys__n34830, ys__n34832, ys__n34834, ys__n34836,
    ys__n34838, ys__n34840, ys__n34842, ys__n34844, ys__n34846, ys__n34848,
    ys__n34850, ys__n34852, ys__n34854, ys__n34856, ys__n34858, ys__n34860,
    ys__n34862, ys__n34864, ys__n34866, ys__n34868, ys__n34870, ys__n34872,
    ys__n34874, ys__n34876, ys__n34878, ys__n34880, ys__n34882, ys__n34884,
    ys__n34886, ys__n34888, ys__n34890, ys__n34892, ys__n34894, ys__n34896,
    ys__n34898, ys__n34900, ys__n34902, ys__n34904, ys__n34906, ys__n34908,
    ys__n34910, ys__n34912, ys__n34914, ys__n34916, ys__n34918, ys__n34920,
    ys__n34922, ys__n34924, ys__n34926, ys__n34928, ys__n34930, ys__n34932,
    ys__n34934, ys__n34936, ys__n34938, ys__n34940, ys__n34942, ys__n34944,
    ys__n34946, ys__n34948, ys__n34950, ys__n34959, ys__n34966, ys__n34972,
    ys__n34976, ys__n34978, ys__n34984, ys__n34988, ys__n34990, ys__n34996,
    ys__n35000, ys__n35002, ys__n35008, ys__n35012, ys__n35014, ys__n35020,
    ys__n35024, ys__n35026, ys__n35028, ys__n35031, ys__n35033, ys__n35035,
    ys__n35037, ys__n35039, ys__n35041, ys__n35047, ys__n35049, ys__n35057,
    ys__n35059, ys__n35065, ys__n35076, ys__n35078, ys__n35080, ys__n35082,
    ys__n35084, ys__n35086, ys__n35088, ys__n35090, ys__n35092, ys__n35094,
    ys__n35096, ys__n35098, ys__n35102, ys__n35104, ys__n35106, ys__n35108,
    ys__n35110, ys__n35112, ys__n35114, ys__n35116, ys__n35118, ys__n35120,
    ys__n35122, ys__n35124, ys__n35413, ys__n35415, ys__n35417, ys__n35419,
    ys__n35421, ys__n35423, ys__n35426, ys__n35704, ys__n35717, ys__n35719,
    ys__n35721, ys__n35723, ys__n35725, ys__n35727, ys__n37668, ys__n37669,
    ys__n37670, ys__n37671, ys__n37672, ys__n37673, ys__n37674, ys__n37675,
    ys__n37678, ys__n37679, ys__n37682, ys__n37692, ys__n37694, ys__n37696,
    ys__n37710, ys__n37712, ys__n37713, ys__n37743, ys__n37744, ys__n37745,
    ys__n37746, ys__n37747, ys__n37748, ys__n37749, ys__n37750, ys__n37751,
    ys__n37752, ys__n37753, ys__n37754, ys__n37755, ys__n37756, ys__n37757,
    ys__n37758, ys__n37759, ys__n37760, ys__n37761, ys__n37762, ys__n37763,
    ys__n37764, ys__n37765, ys__n37766, ys__n37767, ys__n37768, ys__n37769,
    ys__n37770, ys__n37771, ys__n37772, ys__n37773, ys__n37774, ys__n37775,
    ys__n37776, ys__n37777, ys__n37778, ys__n37779, ys__n37780, ys__n37781,
    ys__n37782, ys__n37783, ys__n37784, ys__n37785, ys__n37786, ys__n37787,
    ys__n37788, ys__n37789, ys__n37790, ys__n37791, ys__n37792, ys__n37793,
    ys__n37794, ys__n37795, ys__n37796, ys__n37797, ys__n37798, ys__n37799,
    ys__n37800, ys__n37801, ys__n37802, ys__n37803, ys__n37804, ys__n37805,
    ys__n37806, ys__n37807, ys__n37808, ys__n37809, ys__n37810, ys__n37811,
    ys__n37812, ys__n37813, ys__n37814, ys__n37815, ys__n37816, ys__n37817,
    ys__n37818, ys__n37819, ys__n37820, ys__n37821, ys__n37822, ys__n37823,
    ys__n37824, ys__n37825, ys__n37826, ys__n37827, ys__n37828, ys__n37829,
    ys__n37830, ys__n37831, ys__n37832, ys__n37833, ys__n37834, ys__n37835,
    ys__n37836, ys__n37837, ys__n37838, ys__n37839, ys__n37840, ys__n37841,
    ys__n37842, ys__n37843, ys__n37844, ys__n37845, ys__n37846, ys__n37847,
    ys__n37848, ys__n37849, ys__n37850, ys__n37851, ys__n37852, ys__n37853,
    ys__n37854, ys__n37855, ys__n37856, ys__n37857, ys__n37858, ys__n37859,
    ys__n37860, ys__n37861, ys__n37862, ys__n37863, ys__n37864, ys__n37865,
    ys__n37866, ys__n37867, ys__n37868, ys__n37869, ys__n37870, ys__n37871,
    ys__n37872, ys__n37873, ys__n37874, ys__n37875, ys__n37876, ys__n37877,
    ys__n37878, ys__n37879, ys__n37880, ys__n37881, ys__n37882, ys__n37883,
    ys__n37884, ys__n37885, ys__n37886, ys__n37887, ys__n37888, ys__n37889,
    ys__n37890, ys__n37891, ys__n37892, ys__n37893, ys__n37894, ys__n37895,
    ys__n37896, ys__n37897, ys__n37898, ys__n37899, ys__n37900, ys__n37901,
    ys__n37902, ys__n37903, ys__n37904, ys__n37905, ys__n37906, ys__n37907,
    ys__n37908, ys__n37909, ys__n37910, ys__n37911, ys__n37912, ys__n37913,
    ys__n37914, ys__n37915, ys__n37916, ys__n37917, ys__n37918, ys__n37919,
    ys__n37920, ys__n37921, ys__n37922, ys__n37923, ys__n37924, ys__n37925,
    ys__n37926, ys__n37927, ys__n37928, ys__n37929, ys__n37930, ys__n37931,
    ys__n37932, ys__n37933, ys__n37934, ys__n37935, ys__n37936, ys__n37937,
    ys__n37938, ys__n37939, ys__n37940, ys__n37941, ys__n37942, ys__n37943,
    ys__n37944, ys__n37945, ys__n37946, ys__n37947, ys__n37948, ys__n37949,
    ys__n37950, ys__n37951, ys__n37952, ys__n37953, ys__n37954, ys__n37955,
    ys__n37956, ys__n37957, ys__n37958, ys__n37959, ys__n37960, ys__n37961,
    ys__n37962, ys__n37963, ys__n37964, ys__n37965, ys__n37966, ys__n37967,
    ys__n37968, ys__n37969, ys__n37970, ys__n37971, ys__n37972, ys__n37973,
    ys__n37974, ys__n37975, ys__n37976, ys__n37977, ys__n37978, ys__n37979,
    ys__n37980, ys__n37981, ys__n37982, ys__n37983, ys__n37984, ys__n37985,
    ys__n37986, ys__n37987, ys__n37988, ys__n37989, ys__n37990, ys__n37991,
    ys__n37992, ys__n37993, ys__n37994, ys__n37995, ys__n37996, ys__n37997,
    ys__n37998, ys__n37999, ys__n38000, ys__n38001, ys__n38002, ys__n38003,
    ys__n38004, ys__n38005, ys__n38006, ys__n38007, ys__n38008, ys__n38009,
    ys__n38010, ys__n38011, ys__n38012, ys__n38013, ys__n38014, ys__n38015,
    ys__n38016, ys__n38017, ys__n38018, ys__n38019, ys__n38020, ys__n38021,
    ys__n38022, ys__n38023, ys__n38024, ys__n38025, ys__n38026, ys__n38027,
    ys__n38028, ys__n38029, ys__n38030, ys__n38031, ys__n38032, ys__n38033,
    ys__n38034, ys__n38035, ys__n38036, ys__n38037, ys__n38038, ys__n38039,
    ys__n38040, ys__n38041, ys__n38042, ys__n38043, ys__n38044, ys__n38045,
    ys__n38046, ys__n38047, ys__n38048, ys__n38049, ys__n38050, ys__n38051,
    ys__n38052, ys__n38053, ys__n38054, ys__n38055, ys__n38056, ys__n38057,
    ys__n38058, ys__n38059, ys__n38060, ys__n38061, ys__n38062, ys__n38063,
    ys__n38064, ys__n38065, ys__n38066, ys__n38067, ys__n38068, ys__n38069,
    ys__n38070, ys__n38071, ys__n38072, ys__n38073, ys__n38074, ys__n38075,
    ys__n38076, ys__n38077, ys__n38078, ys__n38079, ys__n38080, ys__n38081,
    ys__n38082, ys__n38083, ys__n38084, ys__n38085, ys__n38086, ys__n38087,
    ys__n38088, ys__n38089, ys__n38090, ys__n38091, ys__n38092, ys__n38093,
    ys__n38094, ys__n38095, ys__n38096, ys__n38097, ys__n38098, ys__n38099,
    ys__n38100, ys__n38101, ys__n38102, ys__n38103, ys__n38104, ys__n38105,
    ys__n38106, ys__n38107, ys__n38108, ys__n38109, ys__n38110, ys__n38111,
    ys__n38112, ys__n38113, ys__n38114, ys__n38115, ys__n38116, ys__n38117,
    ys__n38118, ys__n38119, ys__n38120, ys__n38121, ys__n38122, ys__n38123,
    ys__n38124, ys__n38125, ys__n38126, ys__n38127, ys__n38128, ys__n38129,
    ys__n38130, ys__n38131, ys__n38132, ys__n38133, ys__n38134, ys__n38135,
    ys__n38136, ys__n38137, ys__n38138, ys__n38139, ys__n38140, ys__n38141,
    ys__n38142, ys__n38143, ys__n38144, ys__n38145, ys__n38146, ys__n38147,
    ys__n38148, ys__n38149, ys__n38150, ys__n38151, ys__n38152, ys__n38153,
    ys__n38154, ys__n38155, ys__n38156, ys__n38157, ys__n38158, ys__n38159,
    ys__n38160, ys__n38161, ys__n38162, ys__n38163, ys__n38164, ys__n38165,
    ys__n38166, ys__n38167, ys__n38168, ys__n38169, ys__n38170, ys__n38171,
    ys__n38172, ys__n38173, ys__n38174, ys__n38175, ys__n38176, ys__n38177,
    ys__n38178, ys__n38179, ys__n38183, ys__n38192, ys__n38193, ys__n38194,
    ys__n38195, ys__n38196, ys__n38197, ys__n38198, ys__n38199, ys__n38200,
    ys__n38201, ys__n38202, ys__n38203, ys__n38212, ys__n38215, ys__n38217,
    ys__n38219, ys__n38220, ys__n38221, ys__n38236, ys__n38237, ys__n38257,
    ys__n38259, ys__n38272, ys__n38277, ys__n38278, ys__n38279, ys__n38282,
    ys__n38283, ys__n38286, ys__n38288, ys__n38290, ys__n38291, ys__n38300,
    ys__n38304, ys__n38305, ys__n38307, ys__n38311, ys__n38315, ys__n38320,
    ys__n38323, ys__n38346, ys__n38361, ys__n38376, ys__n38378, ys__n38380,
    ys__n38382, ys__n38384, ys__n38386, ys__n38398, ys__n38407, ys__n38408,
    ys__n38413, ys__n38418, ys__n38420, ys__n38424, ys__n38427, ys__n38437,
    ys__n38438, ys__n38441, ys__n38443, ys__n38448, ys__n38449, ys__n38451,
    ys__n38473, ys__n38486, ys__n38487, ys__n38488, ys__n38489, ys__n38490,
    ys__n38491, ys__n38494, ys__n38495, ys__n38496, ys__n38497, ys__n38498,
    ys__n38499, ys__n38502, ys__n38503, ys__n38504, ys__n38505, ys__n38506,
    ys__n38507, ys__n38513, ys__n38522, ys__n38524, ys__n38526, ys__n38527,
    ys__n38528, ys__n38529, ys__n38553, ys__n38557, ys__n38561, ys__n38564,
    ys__n38565, ys__n38567, ys__n38568, ys__n38569, ys__n38585, ys__n38586,
    ys__n38587, ys__n38588, ys__n38589, ys__n38590, ys__n38591, ys__n38592,
    ys__n38593, ys__n38594, ys__n38595, ys__n38596, ys__n38597, ys__n38598,
    ys__n38599, ys__n38600, ys__n38601, ys__n38602, ys__n38603, ys__n38604,
    ys__n38605, ys__n38606, ys__n38607, ys__n38608, ys__n38609, ys__n38610,
    ys__n38611, ys__n38620, ys__n38624, ys__n38631, ys__n38649, ys__n38654,
    ys__n38670, ys__n38680, ys__n38693, ys__n38694, ys__n38695, ys__n38724,
    ys__n38776, ys__n38777, ys__n38805, ys__n38827, ys__n38828, ys__n38829,
    ys__n38830, ys__n38831, ys__n38832, ys__n38833, ys__n38834, ys__n38835,
    ys__n38836, ys__n38837, ys__n38838, ys__n38839, ys__n38840, ys__n38841,
    ys__n38842, ys__n38843, ys__n38844, ys__n38845, ys__n38846, ys__n38847,
    ys__n38848, ys__n38849, ys__n38850, ys__n38851, ys__n38852, ys__n38853,
    ys__n38854, ys__n38855, ys__n38856, ys__n38857, ys__n38858, ys__n38859,
    ys__n38861, ys__n38862, ys__n38863, ys__n38864, ys__n38865, ys__n38883,
    ys__n38885, ys__n38893, ys__n38894, ys__n38896, ys__n38897, ys__n38898,
    ys__n38902, ys__n38904, ys__n38906, ys__n38908, ys__n38910, ys__n38919,
    ys__n38922, ys__n38927, ys__n38928, ys__n38929, ys__n39167, ys__n39518,
    ys__n39520, ys__n39718, ys__n39720, ys__n39722, ys__n39724, ys__n39726,
    ys__n39728, ys__n39730, ys__n39732, ys__n39734, ys__n39736, ys__n39738,
    ys__n39740, ys__n39742, ys__n39744, ys__n39746, ys__n39748, ys__n39750,
    ys__n39752, ys__n39754, ys__n39756, ys__n39758, ys__n39760, ys__n39762,
    ys__n39764, ys__n39766, ys__n39768, ys__n39770, ys__n39772, ys__n39774,
    ys__n39776, ys__n39778, ys__n44833, ys__n44840, ys__n44842, ys__n44847,
    ys__n44849, ys__n44892, ys__n44906, ys__n44907, ys__n44908, ys__n44988,
    ys__n44989, ys__n44990, ys__n44991, ys__n44992, ys__n44993, ys__n44995,
    ys__n44996, ys__n44998, ys__n44999, ys__n45001, ys__n45002, ys__n45004,
    ys__n45005, ys__n45007, ys__n45008, ys__n45010, ys__n45011, ys__n45013,
    ys__n45014, ys__n45016, ys__n45017, ys__n45019, ys__n45020, ys__n45022,
    ys__n45023, ys__n45025, ys__n45026, ys__n45028, ys__n45029, ys__n45031,
    ys__n45032, ys__n45034, ys__n45035, ys__n45037, ys__n45038, ys__n45040,
    ys__n45041, ys__n45043, ys__n45044, ys__n45046, ys__n45047, ys__n45049,
    ys__n45050, ys__n45052, ys__n45053, ys__n45055, ys__n45056, ys__n45058,
    ys__n45059, ys__n45061, ys__n45062, ys__n45064, ys__n45065, ys__n45067,
    ys__n45068, ys__n45070, ys__n45071, ys__n45073, ys__n45074, ys__n45076,
    ys__n45077, ys__n45079, ys__n45080, ys__n45082, ys__n45083, ys__n45084,
    ys__n45085, ys__n45086, ys__n45087, ys__n45088, ys__n45089, ys__n45090,
    ys__n45091, ys__n45092, ys__n45093, ys__n45094, ys__n45095, ys__n45096,
    ys__n45097, ys__n45098, ys__n45099, ys__n45100, ys__n45101, ys__n45102,
    ys__n45103, ys__n45104, ys__n45105, ys__n45106, ys__n45107, ys__n45108,
    ys__n45109, ys__n45110, ys__n45111, ys__n45112, ys__n45113, ys__n45115,
    ys__n45116, ys__n45118, ys__n45119, ys__n45121, ys__n45122, ys__n45124,
    ys__n45125, ys__n45127, ys__n45128, ys__n45130, ys__n45131, ys__n45133,
    ys__n45134, ys__n45136, ys__n45137, ys__n45139, ys__n45140, ys__n45142,
    ys__n45143, ys__n45145, ys__n45146, ys__n45148, ys__n45149, ys__n45151,
    ys__n45152, ys__n45154, ys__n45155, ys__n45157, ys__n45158, ys__n45160,
    ys__n45161, ys__n45163, ys__n45164, ys__n45166, ys__n45167, ys__n45169,
    ys__n45170, ys__n45172, ys__n45173, ys__n45175, ys__n45176, ys__n45178,
    ys__n45179, ys__n45181, ys__n45182, ys__n45184, ys__n45185, ys__n45187,
    ys__n45188, ys__n45190, ys__n45191, ys__n45193, ys__n45194, ys__n45196,
    ys__n45197, ys__n45199, ys__n45200, ys__n45202, ys__n45203, ys__n45205,
    ys__n45206, ys__n45208, ys__n45209, ys__n45210, ys__n45211, ys__n45212,
    ys__n45214, ys__n45216, ys__n45218, ys__n45220, ys__n45222, ys__n45224,
    ys__n45226, ys__n45228, ys__n45230, ys__n45232, ys__n45234, ys__n45236,
    ys__n45238, ys__n45240, ys__n45242, ys__n45244, ys__n45246, ys__n45248,
    ys__n45250, ys__n45252, ys__n45254, ys__n45256, ys__n45258, ys__n45260,
    ys__n45262, ys__n45264, ys__n45266, ys__n45268, ys__n45270, ys__n45272,
    ys__n45274, ys__n45276, ys__n45277, ys__n45278, ys__n45279, ys__n45280,
    ys__n45281, ys__n45282, ys__n45283, ys__n45284, ys__n45285, ys__n45286,
    ys__n45287, ys__n45288, ys__n45289, ys__n45290, ys__n45291, ys__n45292,
    ys__n45293, ys__n45294, ys__n45295, ys__n45296, ys__n45297, ys__n45298,
    ys__n45299, ys__n45300, ys__n45301, ys__n45302, ys__n45303, ys__n45304,
    ys__n45305, ys__n45306, ys__n45308, ys__n45310, ys__n45312, ys__n45314,
    ys__n45316, ys__n45318, ys__n45320, ys__n45322, ys__n45324, ys__n45326,
    ys__n45328, ys__n45330, ys__n45332, ys__n45334, ys__n45336, ys__n45338,
    ys__n45340, ys__n45342, ys__n45344, ys__n45346, ys__n45348, ys__n45350,
    ys__n45352, ys__n45354, ys__n45356, ys__n45358, ys__n45360, ys__n45362,
    ys__n45364, ys__n45366, ys__n45368, ys__n45370, ys__n45371, ys__n45372,
    ys__n45373, ys__n45374, ys__n45377, ys__n45380, ys__n45382, ys__n45384,
    ys__n45386, ys__n45388, ys__n45390, ys__n45392, ys__n45394, ys__n45396,
    ys__n45398, ys__n45400, ys__n45402, ys__n45404, ys__n45406, ys__n45408,
    ys__n45410, ys__n45412, ys__n45414, ys__n45416, ys__n45418, ys__n45420,
    ys__n45422, ys__n45424, ys__n45426, ys__n45428, ys__n45430, ys__n45432,
    ys__n45434, ys__n45436, ys__n45438, ys__n45440, ys__n45441, ys__n45442,
    ys__n45443, ys__n45444, ys__n45445, ys__n45446, ys__n45447, ys__n45448,
    ys__n45449, ys__n45450, ys__n45451, ys__n45452, ys__n45453, ys__n45454,
    ys__n45455, ys__n45456, ys__n45457, ys__n45458, ys__n45459, ys__n45460,
    ys__n45461, ys__n45462, ys__n45463, ys__n45464, ys__n45465, ys__n45466,
    ys__n45467, ys__n45468, ys__n45469, ys__n45470, ys__n45472, ys__n45474,
    ys__n45476, ys__n45478, ys__n45480, ys__n45482, ys__n45484, ys__n45486,
    ys__n45488, ys__n45490, ys__n45492, ys__n45494, ys__n45496, ys__n45498,
    ys__n45500, ys__n45502, ys__n45504, ys__n45506, ys__n45508, ys__n45510,
    ys__n45512, ys__n45514, ys__n45516, ys__n45518, ys__n45520, ys__n45522,
    ys__n45524, ys__n45526, ys__n45528, ys__n45530, ys__n45532, ys__n45534,
    ys__n45535, ys__n45536, ys__n45537, ys__n45538, ys__n45541, ys__n45544,
    ys__n45546, ys__n45548, ys__n45550, ys__n45552, ys__n45554, ys__n45556,
    ys__n45558, ys__n45560, ys__n45562, ys__n45564, ys__n45566, ys__n45568,
    ys__n45570, ys__n45572, ys__n45574, ys__n45576, ys__n45578, ys__n45580,
    ys__n45582, ys__n45584, ys__n45586, ys__n45588, ys__n45590, ys__n45592,
    ys__n45594, ys__n45596, ys__n45598, ys__n45600, ys__n45602, ys__n45604,
    ys__n45605, ys__n45606, ys__n45607, ys__n45608, ys__n45609, ys__n45610,
    ys__n45611, ys__n45612, ys__n45613, ys__n45614, ys__n45615, ys__n45616,
    ys__n45617, ys__n45618, ys__n45619, ys__n45620, ys__n45621, ys__n45622,
    ys__n45623, ys__n45624, ys__n45625, ys__n45626, ys__n45627, ys__n45628,
    ys__n45629, ys__n45630, ys__n45631, ys__n45632, ys__n45633, ys__n45634,
    ys__n45636, ys__n45638, ys__n45640, ys__n45642, ys__n45644, ys__n45646,
    ys__n45648, ys__n45650, ys__n45652, ys__n45654, ys__n45656, ys__n45658,
    ys__n45660, ys__n45662, ys__n45664, ys__n45666, ys__n45668, ys__n45670,
    ys__n45672, ys__n45674, ys__n45676, ys__n45678, ys__n45680, ys__n45682,
    ys__n45684, ys__n45686, ys__n45688, ys__n45690, ys__n45692, ys__n45694,
    ys__n45696, ys__n45698, ys__n45699, ys__n45700, ys__n45701, ys__n45702,
    ys__n45704, ys__n45707, ys__n45708, ys__n45709, ys__n45710, ys__n45711,
    ys__n45712, ys__n45714, ys__n45715, ys__n45717, ys__n45718, ys__n45720,
    ys__n45721, ys__n45723, ys__n45724, ys__n45726, ys__n45727, ys__n45729,
    ys__n45730, ys__n45732, ys__n45733, ys__n45735, ys__n45736, ys__n45738,
    ys__n45739, ys__n45741, ys__n45742, ys__n45744, ys__n45745, ys__n45747,
    ys__n45748, ys__n45750, ys__n45751, ys__n45753, ys__n45754, ys__n45756,
    ys__n45757, ys__n45759, ys__n45760, ys__n45762, ys__n45763, ys__n45765,
    ys__n45766, ys__n45768, ys__n45769, ys__n45771, ys__n45772, ys__n45774,
    ys__n45775, ys__n45777, ys__n45778, ys__n45780, ys__n45781, ys__n45783,
    ys__n45784, ys__n45786, ys__n45787, ys__n45789, ys__n45790, ys__n45792,
    ys__n45793, ys__n45795, ys__n45796, ys__n45798, ys__n45799, ys__n45801,
    ys__n45802, ys__n45804, ys__n45805, ys__n45806, ys__n45807, ys__n45808,
    ys__n45809, ys__n45810, ys__n45811, ys__n45812, ys__n45813, ys__n45814,
    ys__n45815, ys__n45816, ys__n45817, ys__n45818, ys__n45819, ys__n45820,
    ys__n45821, ys__n45822, ys__n45823, ys__n45824, ys__n45825, ys__n45826,
    ys__n45827, ys__n45828, ys__n45829, ys__n45830, ys__n45831, ys__n45832,
    ys__n45833, ys__n45834, ys__n45835, ys__n45836, ys__n45838, ys__n45840,
    ys__n45842, ys__n45844, ys__n45846, ys__n45848, ys__n45850, ys__n45852,
    ys__n45854, ys__n45856, ys__n45858, ys__n45860, ys__n45862, ys__n45864,
    ys__n45866, ys__n45868, ys__n45870, ys__n45872, ys__n45874, ys__n45876,
    ys__n45878, ys__n45880, ys__n45882, ys__n45884, ys__n45886, ys__n45888,
    ys__n45890, ys__n45892, ys__n45894, ys__n45896, ys__n45898, ys__n45900,
    ys__n45901, ys__n45902, ys__n45903, ys__n45904, ys__n45905, ys__n45906,
    ys__n45907, ys__n45908, ys__n45909, ys__n45910, ys__n45911, ys__n45912,
    ys__n45913, ys__n45914, ys__n45915, ys__n45916, ys__n45917, ys__n45918,
    ys__n45919, ys__n45920, ys__n45921, ys__n45922, ys__n45923, ys__n45924,
    ys__n45925, ys__n45926, ys__n45927, ys__n45928, ys__n45929, ys__n45930,
    ys__n45931, ys__n45933, ys__n45936, ys__n45938, ys__n45940, ys__n45942,
    ys__n45944, ys__n45946, ys__n45948, ys__n45950, ys__n45952, ys__n45954,
    ys__n45956, ys__n45958, ys__n45960, ys__n45962, ys__n45964, ys__n45966,
    ys__n45968, ys__n45970, ys__n45972, ys__n45974, ys__n45976, ys__n45978,
    ys__n45980, ys__n45982, ys__n45984, ys__n45986, ys__n45988, ys__n45990,
    ys__n45992, ys__n45994, ys__n45996, ys__n45998, ys__n45999, ys__n46000,
    ys__n46001, ys__n46002, ys__n46003, ys__n46004, ys__n46005, ys__n46006,
    ys__n46007, ys__n46008, ys__n46009, ys__n46010, ys__n46011, ys__n46012,
    ys__n46013, ys__n46014, ys__n46015, ys__n46016, ys__n46017, ys__n46018,
    ys__n46019, ys__n46020, ys__n46021, ys__n46022, ys__n46023, ys__n46024,
    ys__n46025, ys__n46026, ys__n46027, ys__n46028, ys__n46029, ys__n46031,
    ys__n46034, ys__n46036, ys__n46038, ys__n46040, ys__n46042, ys__n46044,
    ys__n46046, ys__n46048, ys__n46050, ys__n46052, ys__n46054, ys__n46056,
    ys__n46058, ys__n46060, ys__n46062, ys__n46064, ys__n46066, ys__n46068,
    ys__n46070, ys__n46072, ys__n46074, ys__n46076, ys__n46078, ys__n46080,
    ys__n46082, ys__n46084, ys__n46086, ys__n46088, ys__n46090, ys__n46092,
    ys__n46094, ys__n46096, ys__n46097, ys__n46098, ys__n46099, ys__n46100,
    ys__n46101, ys__n46102, ys__n46103, ys__n46104, ys__n46105, ys__n46106,
    ys__n46107, ys__n46108, ys__n46109, ys__n46110, ys__n46111, ys__n46112,
    ys__n46113, ys__n46114, ys__n46115, ys__n46116, ys__n46117, ys__n46118,
    ys__n46119, ys__n46120, ys__n46121, ys__n46122, ys__n46123, ys__n46124,
    ys__n46125, ys__n46126, ys__n46127, ys__n46128, ys__n46130, ys__n46132,
    ys__n46134, ys__n46136, ys__n46141, ys__n46142, ys__n46150, ys__n46151,
    ys__n46152, ys__n46153, ys__n46166, ys__n46168, ys__n46169, ys__n46170,
    ys__n46171, ys__n46180, ys__n46184, ys__n46185, ys__n46186, ys__n46187,
    ys__n46198, ys__n46200, ys__n46201, ys__n46202, ys__n46203, ys__n46214,
    ys__n46216, ys__n46217, ys__n46218, ys__n46219, ys__n46230, ys__n46231,
    ys__n46238, ys__n46239, ys__n46240, ys__n46242, ys__n46244, ys__n46245,
    ys__n46247, ys__n46248, ys__n46252, ys__n46254, ys__n46256, ys__n46258,
    ys__n46260, ys__n46262, ys__n46264, ys__n46266, ys__n46268, ys__n46270,
    ys__n46272, ys__n46274, ys__n46276, ys__n46278, ys__n46280, ys__n46282,
    ys__n46284, ys__n46286, ys__n46288, ys__n46290, ys__n46292, ys__n46294,
    ys__n46296, ys__n46298, ys__n46300, ys__n46302, ys__n46304, ys__n46306,
    ys__n46308, ys__n46310, ys__n46312, ys__n46314, ys__n46315, ys__n46316,
    ys__n46317, ys__n46318, ys__n46319, ys__n46320, ys__n46321, ys__n46322,
    ys__n46323, ys__n46324, ys__n46325, ys__n46326, ys__n46327, ys__n46328,
    ys__n46329, ys__n46330, ys__n46331, ys__n46332, ys__n46333, ys__n46334,
    ys__n46335, ys__n46336, ys__n46337, ys__n46338, ys__n46339, ys__n46340,
    ys__n46341, ys__n46342, ys__n46343, ys__n46344, ys__n46345, ys__n46346,
    ys__n46348, ys__n46350, ys__n46352, ys__n46354, ys__n46356, ys__n46358,
    ys__n46360, ys__n46362, ys__n46364, ys__n46366, ys__n46368, ys__n46370,
    ys__n46372, ys__n46374, ys__n46376, ys__n46378, ys__n46380, ys__n46382,
    ys__n46384, ys__n46386, ys__n46388, ys__n46390, ys__n46392, ys__n46393,
    ys__n46394, ys__n46395, ys__n46396, ys__n46397, ys__n46398, ys__n46399,
    ys__n46400, ys__n46401, ys__n46402, ys__n46403, ys__n46404, ys__n46405,
    ys__n46406, ys__n46407, ys__n46408, ys__n46409, ys__n46410, ys__n46411,
    ys__n46412, ys__n46413, ys__n46414, ys__n46415, ys__n46416, ys__n46417,
    ys__n46418, ys__n46419, ys__n46420, ys__n46421, ys__n46422, ys__n46423,
    ys__n46428, ys__n46430, ys__n46432, ys__n46434, ys__n46436, ys__n46438,
    ys__n46440, ys__n46442, ys__n46444, ys__n46446, ys__n46448, ys__n46450,
    ys__n46452, ys__n46454, ys__n46456, ys__n46458, ys__n46460, ys__n46462,
    ys__n46464, ys__n46466, ys__n46468, ys__n46470, ys__n46472, ys__n46474,
    ys__n46476, ys__n46478, ys__n46480, ys__n46482, ys__n46484, ys__n46486,
    ys__n46488, ys__n46490, ys__n46491, ys__n46492, ys__n46493, ys__n46494,
    ys__n46495, ys__n46496, ys__n46497, ys__n46498, ys__n46499, ys__n46500,
    ys__n46501, ys__n46502, ys__n46503, ys__n46504, ys__n46505, ys__n46506,
    ys__n46507, ys__n46508, ys__n46509, ys__n46510, ys__n46511, ys__n46512,
    ys__n46513, ys__n46514, ys__n46515, ys__n46516, ys__n46517, ys__n46518,
    ys__n46519, ys__n46520, ys__n46521, ys__n46522, ys__n46524, ys__n46526,
    ys__n46528, ys__n46530, ys__n46532, ys__n46534, ys__n46536, ys__n46538,
    ys__n46540, ys__n46542, ys__n46544, ys__n46546, ys__n46548, ys__n46550,
    ys__n46552, ys__n46554, ys__n46556, ys__n46558, ys__n46560, ys__n46562,
    ys__n46564, ys__n46566, ys__n46568, ys__n46569, ys__n46570, ys__n46571,
    ys__n46572, ys__n46573, ys__n46574, ys__n46575, ys__n46576, ys__n46577,
    ys__n46578, ys__n46579, ys__n46580, ys__n46581, ys__n46582, ys__n46583,
    ys__n46584, ys__n46585, ys__n46586, ys__n46587, ys__n46588, ys__n46589,
    ys__n46590, ys__n46591, ys__n46592, ys__n46593, ys__n46594, ys__n46595,
    ys__n46596, ys__n46597, ys__n46598, ys__n46599, ys__n46604, ys__n46606,
    ys__n46608, ys__n46610, ys__n46612, ys__n46614, ys__n46616, ys__n46618,
    ys__n46620, ys__n46622, ys__n46624, ys__n46626, ys__n46628, ys__n46630,
    ys__n46632, ys__n46634, ys__n46636, ys__n46638, ys__n46640, ys__n46642,
    ys__n46644, ys__n46646, ys__n46648, ys__n46650, ys__n46652, ys__n46654,
    ys__n46656, ys__n46658, ys__n46660, ys__n46662, ys__n46664, ys__n46666,
    ys__n46667, ys__n46668, ys__n46669, ys__n46670, ys__n46671, ys__n46672,
    ys__n46673, ys__n46674, ys__n46675, ys__n46676, ys__n46677, ys__n46678,
    ys__n46679, ys__n46680, ys__n46681, ys__n46682, ys__n46683, ys__n46684,
    ys__n46685, ys__n46686, ys__n46687, ys__n46688, ys__n46689, ys__n46690,
    ys__n46691, ys__n46692, ys__n46693, ys__n46694, ys__n46695, ys__n46696,
    ys__n46697, ys__n46698, ys__n46700, ys__n46702, ys__n46704, ys__n46706,
    ys__n46708, ys__n46710, ys__n46712, ys__n46714, ys__n46716, ys__n46718,
    ys__n46720, ys__n46722, ys__n46724, ys__n46726, ys__n46728, ys__n46730,
    ys__n46732, ys__n46734, ys__n46736, ys__n46738, ys__n46740, ys__n46742,
    ys__n46744, ys__n46745, ys__n46746, ys__n46747, ys__n46748, ys__n46749,
    ys__n46750, ys__n46751, ys__n46752, ys__n46753, ys__n46754, ys__n46755,
    ys__n46756, ys__n46757, ys__n46758, ys__n46759, ys__n46760, ys__n46761,
    ys__n46762, ys__n46763, ys__n46764, ys__n46765, ys__n46766, ys__n46767,
    ys__n46768, ys__n46769, ys__n46770, ys__n46771, ys__n46772, ys__n46773,
    ys__n46774, ys__n46775, ys__n46780, ys__n46782, ys__n46784, ys__n46786,
    ys__n46788, ys__n46790, ys__n46792, ys__n46794, ys__n46796, ys__n46798,
    ys__n46800, ys__n46802, ys__n46804, ys__n46806, ys__n46808, ys__n46810,
    ys__n46812, ys__n46814, ys__n46816, ys__n46818, ys__n46820, ys__n46822,
    ys__n46824, ys__n46826, ys__n46828, ys__n46830, ys__n46832, ys__n46834,
    ys__n46836, ys__n46838, ys__n46840, ys__n46842, ys__n46843, ys__n46844,
    ys__n46845, ys__n46846, ys__n46847, ys__n46848, ys__n46849, ys__n46850,
    ys__n46851, ys__n46852, ys__n46853, ys__n46854, ys__n46855, ys__n46856,
    ys__n46857, ys__n46858, ys__n46859, ys__n46860, ys__n46861, ys__n46862,
    ys__n46863, ys__n46864, ys__n46865, ys__n46866, ys__n46867, ys__n46868,
    ys__n46869, ys__n46870, ys__n46871, ys__n46872, ys__n46873, ys__n46874,
    ys__n46876, ys__n46878, ys__n46880, ys__n46882, ys__n46884, ys__n46886,
    ys__n46888, ys__n46890, ys__n46892, ys__n46894, ys__n46896, ys__n46898,
    ys__n46900, ys__n46902, ys__n46904, ys__n46906, ys__n46908, ys__n46910,
    ys__n46912, ys__n46914, ys__n46916, ys__n46918, ys__n46920, ys__n46921,
    ys__n46922, ys__n46923, ys__n46924, ys__n46925, ys__n46926, ys__n46927,
    ys__n46928, ys__n46929, ys__n46930, ys__n46931, ys__n46932, ys__n46933,
    ys__n46934, ys__n46935, ys__n46936, ys__n46937, ys__n46938, ys__n46939,
    ys__n46940, ys__n46941, ys__n46942, ys__n46943, ys__n46944, ys__n46945,
    ys__n46946, ys__n46947, ys__n46948, ys__n46949, ys__n46950, ys__n46951,
    ys__n46954, ys__n46955, ys__n46956, ys__n46957, ys__n46958, ys__n46959,
    ys__n46960, ys__n46961, ys__n46962, ys__n46963, ys__n46964, ys__n46965,
    ys__n46966, ys__n46967, ys__n46968, ys__n46969, ys__n46970, ys__n46971,
    ys__n46972, ys__n46973, ys__n46974, ys__n46975, ys__n46976, ys__n46977,
    ys__n46978, ys__n46979, ys__n46980, ys__n46981, ys__n46982, ys__n46983,
    ys__n46984, ys__n46985, ys__n46986, ys__n46987, ys__n46988, ys__n46989,
    ys__n46990, ys__n46991, ys__n46992, ys__n46993, ys__n46994, ys__n46995,
    ys__n46996, ys__n46997, ys__n46998, ys__n46999, ys__n47000, ys__n47001,
    ys__n47002, ys__n47003, ys__n47004, ys__n47005, ys__n47006, ys__n47007,
    ys__n47008, ys__n47009, ys__n47010, ys__n47011, ys__n47012, ys__n47013,
    ys__n47014, ys__n47015, ys__n47016, ys__n47017, ys__n47018, ys__n47019,
    ys__n47020, ys__n47021, ys__n47022, ys__n47023, ys__n47024, ys__n47025,
    ys__n47026, ys__n47027, ys__n47028, ys__n47029, ys__n47030, ys__n47031,
    ys__n47032, ys__n47033, ys__n47034, ys__n47035, ys__n47036, ys__n47037,
    ys__n47038, ys__n47039, ys__n47040, ys__n47041, ys__n47074, ys__n47075,
    ys__n47076, ys__n47077, ys__n47078, ys__n47079, ys__n47080, ys__n47081,
    ys__n47082, ys__n47083, ys__n47084, ys__n47085, ys__n47086, ys__n47087,
    ys__n47088, ys__n47089, ys__n47090, ys__n47091, ys__n47092, ys__n47093,
    ys__n47094, ys__n47095, ys__n47096, ys__n47097, ys__n47098, ys__n47099,
    ys__n47100, ys__n47101, ys__n47102, ys__n47103, ys__n47104, ys__n47105,
    ys__n47106, ys__n47107, ys__n47108, ys__n47109, ys__n47110, ys__n47111,
    ys__n47112, ys__n47113, ys__n47114, ys__n47115, ys__n47116, ys__n47117,
    ys__n47118, ys__n47119, ys__n47184, ys__n47185, ys__n47186, ys__n47187,
    ys__n47188, ys__n47189, ys__n47190, ys__n47191, ys__n47192, ys__n47193,
    ys__n47194, ys__n47195, ys__n47196, ys__n47197, ys__n47198, ys__n47199,
    ys__n47200, ys__n47201, ys__n47202, ys__n47203, ys__n47204, ys__n47205,
    ys__n47206, ys__n47207, ys__n47208, ys__n47209, ys__n47210, ys__n47211,
    ys__n47212, ys__n47213, ys__n47214, ys__n47215, ys__n47216, ys__n47217,
    ys__n47218, ys__n47219, ys__n47220, ys__n47221, ys__n47222, ys__n47223,
    ys__n47224, ys__n47225, ys__n47226, ys__n47227, ys__n47228, ys__n47229,
    ys__n47230, ys__n47231, ys__n47232, ys__n47233, ys__n47234, ys__n47235,
    ys__n47236, ys__n47237, ys__n47238, ys__n47239, ys__n47240, ys__n47241,
    ys__n47242, ys__n47243, ys__n47244, ys__n47245, ys__n47246, ys__n47247,
    ys__n47248, ys__n47249, ys__n47250, ys__n47251, ys__n47252, ys__n47253,
    ys__n47254, ys__n47255, ys__n47256, ys__n47257, ys__n47258, ys__n47259,
    ys__n47260, ys__n47261, ys__n47262, ys__n47263, ys__n47264, ys__n47265,
    ys__n47266, ys__n47267, ys__n47268, ys__n47269, ys__n47270, ys__n47271,
    ys__n47272, ys__n47273, ys__n47274, ys__n47275, ys__n47276, ys__n47277,
    ys__n47278, ys__n47279, ys__n47280, ys__n47281, ys__n47282, ys__n47283,
    ys__n47284, ys__n47285, ys__n47286, ys__n47287, ys__n47288, ys__n47289,
    ys__n47290, ys__n47291, ys__n47292, ys__n47293, ys__n47294, ys__n47295,
    ys__n47296, ys__n47297, ys__n47298, ys__n47299, ys__n47300, ys__n47301,
    ys__n47302, ys__n47303, ys__n47305, ys__n47306, ys__n47307, ys__n47308,
    ys__n47309, ys__n47310, ys__n47311, ys__n47312, ys__n47313, ys__n47314,
    ys__n47315, ys__n47316, ys__n47317, ys__n47318, ys__n47319, ys__n47320,
    ys__n47321, ys__n47322, ys__n47323, ys__n47324, ys__n47325, ys__n47326,
    ys__n47327, ys__n47328, ys__n47329, ys__n47330, ys__n47331, ys__n47332,
    ys__n47333, ys__n47334, ys__n47335, ys__n47336, ys__n47337, ys__n47338,
    ys__n47339, ys__n47340, ys__n47341, ys__n47342, ys__n47343, ys__n47344,
    ys__n47345, ys__n47346, ys__n47347, ys__n47348, ys__n47349, ys__n47350,
    ys__n47351, ys__n47352, ys__n47353, ys__n47354, ys__n47355, ys__n47356,
    ys__n47357, ys__n47358, ys__n47359, ys__n47360, ys__n47361, ys__n47362,
    ys__n47363, ys__n47364, ys__n47365, ys__n47366, ys__n47367, ys__n47368,
    ys__n47369, ys__n47370, ys__n47371, ys__n47372, ys__n47373, ys__n47374,
    ys__n47375, ys__n47376, ys__n47377, ys__n47378, ys__n47379, ys__n47380,
    ys__n47381, ys__n47382, ys__n47383, ys__n47384, ys__n47385, ys__n47386,
    ys__n47387, ys__n47388, ys__n47389, ys__n47390, ys__n47391, ys__n47392,
    ys__n47393, ys__n47394, ys__n47395, ys__n47396, ys__n47397, ys__n47398,
    ys__n47399, ys__n47400, ys__n47401, ys__n47402, ys__n47403, ys__n47404,
    ys__n47405, ys__n47406, ys__n47407, ys__n47408, ys__n47409, ys__n47410,
    ys__n47411, ys__n47412, ys__n47413, ys__n47414, ys__n47415, ys__n47416,
    ys__n47417, ys__n47418, ys__n47419, ys__n47420, ys__n47421, ys__n47422,
    ys__n47423, ys__n47424, ys__n47425, ys__n47426, ys__n47427, ys__n47428,
    ys__n47429, ys__n47430, ys__n47431, ys__n47432, ys__n47433, ys__n47434,
    ys__n47435, ys__n47436, ys__n47437, ys__n47438, ys__n47439, ys__n47440,
    ys__n47441, ys__n47442, ys__n47443, ys__n47444, ys__n47445, ys__n47446,
    ys__n47447, ys__n47448, ys__n47449, ys__n47450, ys__n47451, ys__n47452,
    ys__n47453, ys__n47454, ys__n47455, ys__n47456, ys__n47457, ys__n47458,
    ys__n47459, ys__n47460, ys__n47461, ys__n47462, ys__n47463, ys__n47464,
    ys__n47465, ys__n47466, ys__n47467, ys__n47468, ys__n47469, ys__n47470,
    ys__n47471, ys__n47472, ys__n47473, ys__n47474, ys__n47475, ys__n47476,
    ys__n47477, ys__n47478, ys__n47479, ys__n47480, ys__n47481, ys__n47482,
    ys__n47483, ys__n47484, ys__n47485, ys__n47486, ys__n47487, ys__n47488,
    ys__n47489, ys__n47490, ys__n47491, ys__n47492, ys__n47493, ys__n47494,
    ys__n47495, ys__n47496, ys__n47497, ys__n47498, ys__n47499, ys__n47500,
    ys__n47501, ys__n47502, ys__n47503, ys__n47504, ys__n47505, ys__n47506,
    ys__n47507, ys__n47508, ys__n47509, ys__n47510, ys__n47511, ys__n47512,
    ys__n47513, ys__n47514, ys__n47515, ys__n47516, ys__n47517, ys__n47518,
    ys__n47519, ys__n47520, ys__n47521, ys__n47522, ys__n47523, ys__n47524,
    ys__n47525, ys__n47526, ys__n47527, ys__n47528, ys__n47529, ys__n47530,
    ys__n47531, ys__n47532, ys__n47533, ys__n47534, ys__n47535, ys__n47536,
    ys__n47537, ys__n47538, ys__n47539, ys__n47540, ys__n47541, ys__n47542,
    ys__n47543, ys__n47544, ys__n47545, ys__n47546, ys__n47547, ys__n47548,
    ys__n47549, ys__n47550, ys__n47551, ys__n47552, ys__n47553, ys__n47554,
    ys__n47555, ys__n47556, ys__n47557, ys__n47558, ys__n47559, ys__n47560,
    ys__n47561, ys__n47562, ys__n47563, ys__n47564, ys__n47565, ys__n47566,
    ys__n47567, ys__n47568, ys__n47569, ys__n47570, ys__n47571, ys__n47572,
    ys__n47573, ys__n47574, ys__n47575, ys__n47576, ys__n47577, ys__n47578,
    ys__n47579, ys__n47580, ys__n47581, ys__n47582, ys__n47583, ys__n47584,
    ys__n47585, ys__n47586, ys__n47587, ys__n47588, ys__n47589, ys__n47590,
    ys__n47591, ys__n47592, ys__n47593, ys__n47594, ys__n47595, ys__n47596,
    ys__n47597, ys__n47598, ys__n47599, ys__n47600, ys__n47601, ys__n47602,
    ys__n47603, ys__n47604, ys__n47605, ys__n47606, ys__n47607, ys__n47608,
    ys__n47609, ys__n47610, ys__n47611, ys__n47612, ys__n47613, ys__n47614,
    ys__n47615, ys__n47616, ys__n47617, ys__n47618, ys__n47619, ys__n47620,
    ys__n47621, ys__n47622, ys__n47623, ys__n47624, ys__n47625, ys__n47626,
    ys__n47627, ys__n47628, ys__n47629, ys__n47630, ys__n47631, ys__n47632,
    ys__n47633, ys__n47634, ys__n47635, ys__n47636, ys__n47637, ys__n47638,
    ys__n47639, ys__n47640, ys__n47641, ys__n47642, ys__n47643, ys__n47644,
    ys__n47645, ys__n47646, ys__n47647, ys__n47648, ys__n47649, ys__n47650,
    ys__n47651, ys__n47652, ys__n47653, ys__n47654, ys__n47655, ys__n47656,
    ys__n47657, ys__n47658, ys__n47659, ys__n47660, ys__n47661, ys__n47662,
    ys__n47663, ys__n47664, ys__n47665, ys__n47666, ys__n47667, ys__n47668,
    ys__n47669, ys__n47670, ys__n47671, ys__n47672, ys__n47673, ys__n47674,
    ys__n47675, ys__n47676, ys__n47677, ys__n47678, ys__n47679, ys__n47680,
    ys__n47681, ys__n47682, ys__n47683, ys__n47684, ys__n47685, ys__n47686,
    ys__n47687, ys__n47688, ys__n47689, ys__n47690, ys__n47691, ys__n47692,
    ys__n47693, ys__n47694, ys__n47695, ys__n47696, ys__n47697, ys__n47698,
    ys__n47699, ys__n47700, ys__n47701, ys__n47702, ys__n47703, ys__n47704,
    ys__n47705, ys__n47706, ys__n47707, ys__n47708, ys__n47709, ys__n47710,
    ys__n47711, ys__n47712, ys__n47713, ys__n47714, ys__n47715, ys__n47716,
    ys__n47717, ys__n47718, ys__n47719, ys__n47720, ys__n47721, ys__n47722,
    ys__n47723, ys__n47724, ys__n47725, ys__n47726, ys__n47727, ys__n47728,
    ys__n47729, ys__n47730, ys__n47731, ys__n47732, ys__n47733, ys__n47734,
    ys__n47735, ys__n47736, ys__n47737, ys__n47738, ys__n47739, ys__n47740,
    ys__n47741, ys__n47742, ys__n47743, ys__n47744, ys__n47745, ys__n47746,
    ys__n47747, ys__n47748, ys__n47749, ys__n47750, ys__n47751, ys__n47752,
    ys__n47753, ys__n47754, ys__n47755, ys__n47756, ys__n47757, ys__n47758,
    ys__n47759, ys__n47760, ys__n47761, ys__n47762, ys__n47763, ys__n47764,
    ys__n47765, ys__n47766, ys__n47767, ys__n47768, ys__n47769, ys__n47770,
    ys__n47771, ys__n47772, ys__n47773, ys__n47774, ys__n47775, ys__n47776,
    ys__n47777, ys__n47778, ys__n47779, ys__n47780, ys__n47781, ys__n47782,
    ys__n47783, ys__n47784, ys__n47785, ys__n47786, ys__n47787, ys__n47788,
    ys__n47789, ys__n47790, ys__n47791, ys__n47792, ys__n47793, ys__n47794,
    ys__n47795, ys__n47796, ys__n47797, ys__n47798, ys__n47799, ys__n47800,
    ys__n47801, ys__n47802, ys__n47803, ys__n47804, ys__n47805, ys__n47806,
    ys__n47807, ys__n47808, ys__n47809, ys__n47810, ys__n47811, ys__n47812,
    ys__n47813, ys__n47814, ys__n47815, ys__n47816, ys__n47817, ys__n47818,
    ys__n47819, ys__n47820, ys__n47821, ys__n47822, ys__n47823, ys__n47824,
    ys__n47825, ys__n47826, ys__n47827, ys__n47828, ys__n47829, ys__n47830,
    ys__n47831, ys__n47832, ys__n47833, ys__n47834, ys__n47835, ys__n47836,
    ys__n47837, ys__n47838, ys__n47839, ys__n47840, ys__n47841, ys__n47842,
    ys__n47843, ys__n47844, ys__n47845, ys__n47846, ys__n47847, ys__n47848,
    ys__n47849, ys__n47850, ys__n47851, ys__n47852, ys__n47853, ys__n47854,
    ys__n47855, ys__n47856, ys__n47857, ys__n47858, ys__n47859, ys__n47860,
    ys__n47861, ys__n47862, ys__n47863, ys__n47864, ys__n47865, ys__n47866,
    ys__n47867, ys__n47868, ys__n47869, ys__n47870, ys__n47871, ys__n47872,
    ys__n47873, ys__n47874, ys__n47875, ys__n47876, ys__n47877, ys__n47878,
    ys__n47879, ys__n47880, ys__n47881, ys__n47882, ys__n47883, ys__n47884,
    ys__n47885, ys__n47886, ys__n47887, ys__n47888, ys__n47889, ys__n47890,
    ys__n47891, ys__n47892, ys__n47893, ys__n47894, ys__n47895, ys__n47896,
    ys__n47897, ys__n47898, ys__n47899, ys__n47900, ys__n47901, ys__n47902,
    ys__n47903, ys__n47904, ys__n47905, ys__n47906, ys__n47907, ys__n47908,
    ys__n47909, ys__n47910, ys__n47911, ys__n47912, ys__n47913, ys__n47914,
    ys__n47915, ys__n47916, ys__n47917, ys__n47918, ys__n47919, ys__n47920,
    ys__n47921, ys__n47922, ys__n47923, ys__n47924, ys__n47925, ys__n47926,
    ys__n47927, ys__n47928, ys__n47929, ys__n47930, ys__n47931, ys__n47932,
    ys__n47933, ys__n47934, ys__n47935, ys__n47936, ys__n47937, ys__n47938,
    ys__n47939, ys__n47940, ys__n47941, ys__n47942, ys__n47943, ys__n47944,
    ys__n47945, ys__n47946, ys__n47947, ys__n47948, ys__n47949, ys__n47950,
    ys__n47951, ys__n47952, ys__n47953, ys__n47954, ys__n47955, ys__n47956,
    ys__n47957, ys__n47958, ys__n47959, ys__n47960, ys__n47961, ys__n47962,
    ys__n47963, ys__n47964, ys__n47965, ys__n47966, ys__n47967, ys__n47968,
    ys__n47969, ys__n47970, ys__n47971, ys__n47972, ys__n47973, ys__n47974,
    ys__n47975, ys__n47976, ys__n47977, ys__n47978, ys__n47979, ys__n47980,
    ys__n47981, ys__n47982, ys__n47983, ys__n47984, ys__n47985, ys__n47986,
    ys__n47987, ys__n47988, ys__n47989, ys__n47990, ys__n47991, ys__n47992,
    ys__n47993, ys__n47994, ys__n47995, ys__n47996, ys__n47997, ys__n47998,
    ys__n47999, ys__n48000, ys__n48001, ys__n48002, ys__n48003, ys__n48004,
    ys__n48005, ys__n48006, ys__n48007, ys__n48008, ys__n48009, ys__n48010,
    ys__n48011, ys__n48012, ys__n48013, ys__n48014, ys__n48015, ys__n48016,
    ys__n48017, ys__n48018, ys__n48019, ys__n48020, ys__n48021, ys__n48022,
    ys__n48023, ys__n48024, ys__n48025, ys__n48026, ys__n48027, ys__n48028,
    ys__n48029, ys__n48030, ys__n48031, ys__n48032, ys__n48033, ys__n48034,
    ys__n48035, ys__n48036, ys__n48037, ys__n48038, ys__n48039, ys__n48040,
    ys__n48041, ys__n48042, ys__n48043, ys__n48044, ys__n48045, ys__n48046,
    ys__n48047, ys__n48048, ys__n48049, ys__n48050, ys__n48051, ys__n48052,
    ys__n48053, ys__n48054, ys__n48055, ys__n48056, ys__n48057, ys__n48058,
    ys__n48059, ys__n48060, ys__n48061, ys__n48062, ys__n48063, ys__n48064,
    ys__n48065, ys__n48066, ys__n48067, ys__n48068, ys__n48069, ys__n48070,
    ys__n48071, ys__n48072, ys__n48073, ys__n48074, ys__n48075, ys__n48076,
    ys__n48077, ys__n48078, ys__n48079, ys__n48080, ys__n48081, ys__n48082,
    ys__n48083, ys__n48084, ys__n48085, ys__n48086, ys__n48087, ys__n48088,
    ys__n48089, ys__n48090, ys__n48091, ys__n48092, ys__n48093, ys__n48094,
    ys__n48095, ys__n48096, ys__n48097, ys__n48098, ys__n48099, ys__n48100,
    ys__n48101, ys__n48102, ys__n48103, ys__n48104, ys__n48105, ys__n48106,
    ys__n48107, ys__n48108, ys__n48109, ys__n48110, ys__n48111, ys__n48112,
    ys__n48113, ys__n48114, ys__n48115, ys__n48116, ys__n48117, ys__n48118,
    ys__n48119, ys__n48120, ys__n48121, ys__n48122, ys__n48123, ys__n48124,
    ys__n48125, ys__n48126, ys__n48127, ys__n48128, ys__n48129, ys__n48130,
    ys__n48131, ys__n48132, ys__n48133, ys__n48134, ys__n48135, ys__n48136,
    ys__n48137, ys__n48138, ys__n48139, ys__n48140, ys__n48141, ys__n48142,
    ys__n48143, ys__n48144, ys__n48145, ys__n48146, ys__n48147, ys__n48148,
    ys__n48149, ys__n48150, ys__n48151, ys__n48152, ys__n48153, ys__n48154,
    ys__n48155, ys__n48156, ys__n48157, ys__n48158, ys__n48159, ys__n48160,
    ys__n48161, ys__n48162, ys__n48163, ys__n48164, ys__n48165, ys__n48166,
    ys__n48167, ys__n48168, ys__n48169, ys__n48170, ys__n48171, ys__n48172,
    ys__n48173, ys__n48174, ys__n48175, ys__n48176, ys__n48177, ys__n48178,
    ys__n48179, ys__n48180, ys__n48181, ys__n48182, ys__n48183, ys__n48184,
    ys__n48185, ys__n48186, ys__n48187, ys__n48188, ys__n48189, ys__n48190,
    ys__n48191, ys__n48192, ys__n48193, ys__n48194, ys__n48195, ys__n48196,
    ys__n48197, ys__n48198, ys__n48199, ys__n48200, ys__n48201, ys__n48202,
    ys__n48203, ys__n48204, ys__n48205, ys__n48206, ys__n48207, ys__n48208,
    ys__n48209, ys__n48210, ys__n48211, ys__n48212, ys__n48213, ys__n48214,
    ys__n48215, ys__n48216, ys__n48217, ys__n48218, ys__n48219, ys__n48220,
    ys__n48221, ys__n48222, ys__n48223, ys__n48224, ys__n48225, ys__n48226,
    ys__n48227, ys__n48228, ys__n48229, ys__n48230, ys__n48231, ys__n48232,
    ys__n48233, ys__n48234, ys__n48235, ys__n48236, ys__n48237, ys__n48238,
    ys__n48239, ys__n48240, ys__n48241, ys__n48242, ys__n48243, ys__n48244,
    ys__n48245, ys__n48246, ys__n48247, ys__n48248, ys__n48249, ys__n48250,
    ys__n48251, ys__n48252, ys__n48253, ys__n48254, ys__n48255, ys__n48256,
    ys__n48257, ys__n48258, ys__n48259, ys__n48260, ys__n48261, ys__n48262,
    ys__n48263, ys__n48264, ys__n48265, ys__n48266, ys__n48267, ys__n48268,
    ys__n48269, ys__n48270, ys__n48271, ys__n48272, ys__n48273, ys__n48274,
    ys__n48275, ys__n48324, ys__n48325, ys__n48327, ys__n48330, ys__n48331,
    ys__n48332, ys__n48333, ys__n48334, ys__n48335;
  output ys__n2, ys__n246, ys__n250, ys__n252, ys__n254, ys__n264, ys__n270,
    ys__n278, ys__n280, ys__n313, ys__n319, ys__n404, ys__n415, ys__n417,
    ys__n455, ys__n457, ys__n478, ys__n480, ys__n482, ys__n502, ys__n565,
    ys__n574, ys__n576, ys__n628, ys__n630, ys__n714, ys__n716, ys__n730,
    ys__n732, ys__n738, ys__n740, ys__n754, ys__n756, ys__n786, ys__n788,
    ys__n790, ys__n792, ys__n794, ys__n796, ys__n798, ys__n800, ys__n802,
    ys__n804, ys__n806, ys__n808, ys__n810, ys__n812, ys__n814, ys__n862,
    ys__n863, ys__n865, ys__n866, ys__n868, ys__n870, ys__n871, ys__n872,
    ys__n873, ys__n876, ys__n878, ys__n879, ys__n881, ys__n888, ys__n890,
    ys__n900, ys__n902, ys__n904, ys__n911, ys__n920, ys__n923, ys__n927,
    ys__n929, ys__n930, ys__n932, ys__n934, ys__n936, ys__n942, ys__n944,
    ys__n948, ys__n949, ys__n970, ys__n972, ys__n974, ys__n976, ys__n978,
    ys__n980, ys__n982, ys__n989, ys__n991, ys__n993, ys__n995, ys__n999,
    ys__n1001, ys__n1004, ys__n1007, ys__n1009, ys__n1013, ys__n1020,
    ys__n1028, ys__n1030, ys__n1031, ys__n1032, ys__n1037, ys__n1040,
    ys__n1043, ys__n1046, ys__n1047, ys__n1049, ys__n1060, ys__n1071,
    ys__n1073, ys__n1074, ys__n1075, ys__n1077, ys__n1079, ys__n1080,
    ys__n1083, ys__n1085, ys__n1087, ys__n1088, ys__n1089, ys__n1090,
    ys__n1091, ys__n1095, ys__n1103, ys__n1115, ys__n1125, ys__n1128,
    ys__n1135, ys__n1138, ys__n1141, ys__n1142, ys__n1143, ys__n1146,
    ys__n1148, ys__n1161, ys__n1163, ys__n1164, ys__n1165, ys__n1167,
    ys__n1170, ys__n1171, ys__n1183, ys__n1189, ys__n1195, ys__n1201,
    ys__n1207, ys__n1213, ys__n1219, ys__n1222, ys__n1228, ys__n1234,
    ys__n1240, ys__n1246, ys__n1252, ys__n1258, ys__n1261, ys__n1266,
    ys__n1272, ys__n1278, ys__n1284, ys__n1290, ys__n1296, ys__n1303,
    ys__n1377, ys__n1386, ys__n1445, ys__n1448, ys__n1470, ys__n1591,
    ys__n1598, ys__n1601, ys__n1616, ys__n1790, ys__n1802, ys__n1817,
    ys__n1835, ys__n1837, ys__n2152, ys__n2365, ys__n2400, ys__n2423,
    ys__n2491, ys__n2535, ys__n2536, ys__n2582, ys__n2635, ys__n2651,
    ys__n2653, ys__n2655, ys__n2674, ys__n2684, ys__n2733, ys__n2776,
    ys__n2778, ys__n2780, ys__n2782, ys__n2804, ys__n2806, ys__n2845,
    ys__n2855, ys__n3021, ys__n3024, ys__n3035, ys__n3039, ys__n3040,
    ys__n3051, ys__n3061, ys__n3068, ys__n3083, ys__n3085, ys__n3097,
    ys__n3106, ys__n3114, ys__n3115, ys__n3118, ys__n3121, ys__n3195,
    ys__n3249, ys__n3250, ys__n3252, ys__n4175, ys__n4189, ys__n4192,
    ys__n4320, ys__n4414, ys__n4521, ys__n4566, ys__n4588, ys__n4603,
    ys__n4615, ys__n4696, ys__n4764, ys__n4791, ys__n4793, ys__n4798,
    ys__n4817, ys__n4818, ys__n4820, ys__n4821, ys__n4824, ys__n4825,
    ys__n4839, ys__n4840, ys__n12455, ys__n12458, ys__n12461, ys__n12464,
    ys__n12467, ys__n12470, ys__n12473, ys__n12476, ys__n12479, ys__n12482,
    ys__n12485, ys__n12488, ys__n12491, ys__n12494, ys__n12497, ys__n12500,
    ys__n12503, ys__n12506, ys__n12509, ys__n12512, ys__n12515, ys__n12518,
    ys__n12521, ys__n12524, ys__n12527, ys__n12530, ys__n12533, ys__n12536,
    ys__n12539, ys__n12542, ys__n12545, ys__n12548, ys__n16188, ys__n16191,
    ys__n16412, ys__n16415, ys__n16424, ys__n16427, ys__n16706, ys__n16709,
    ys__n16718, ys__n16721, ys__n17692, ys__n17697, ys__n17780, ys__n18007,
    ys__n18009, ys__n18015, ys__n18019, ys__n18028, ys__n18078, ys__n18080,
    ys__n18082, ys__n18087, ys__n18088, ys__n18089, ys__n18120, ys__n18125,
    ys__n18128, ys__n18131, ys__n18133, ys__n18134, ys__n18136, ys__n18137,
    ys__n18154, ys__n18165, ys__n18166, ys__n18169, ys__n18170, ys__n18174,
    ys__n18176, ys__n18178, ys__n18210, ys__n18214, ys__n18216, ys__n18217,
    ys__n18218, ys__n18223, ys__n18227, ys__n18236, ys__n18238, ys__n18239,
    ys__n18241, ys__n18251, ys__n18268, ys__n18272, ys__n18273, ys__n18278,
    ys__n18281, ys__n18284, ys__n18287, ys__n18303, ys__n18321, ys__n18329,
    ys__n18331, ys__n18333, ys__n18335, ys__n18337, ys__n18339, ys__n18341,
    ys__n18343, ys__n18345, ys__n18347, ys__n18349, ys__n18351, ys__n18353,
    ys__n18355, ys__n18357, ys__n18360, ys__n18380, ys__n18383, ys__n18386,
    ys__n18391, ys__n18392, ys__n18394, ys__n18395, ys__n18396, ys__n18397,
    ys__n18398, ys__n18399, ys__n18400, ys__n18401, ys__n18402, ys__n18403,
    ys__n18404, ys__n18405, ys__n18406, ys__n18407, ys__n18408, ys__n18409,
    ys__n18410, ys__n18411, ys__n18412, ys__n18413, ys__n18414, ys__n18415,
    ys__n18416, ys__n18417, ys__n18418, ys__n18419, ys__n18420, ys__n18421,
    ys__n18422, ys__n18423, ys__n18424, ys__n18425, ys__n18426, ys__n18427,
    ys__n18428, ys__n18429, ys__n18430, ys__n18431, ys__n18432, ys__n18433,
    ys__n18434, ys__n18435, ys__n18436, ys__n18437, ys__n18438, ys__n18439,
    ys__n18440, ys__n18441, ys__n18442, ys__n18443, ys__n18444, ys__n18445,
    ys__n18449, ys__n18450, ys__n18452, ys__n18453, ys__n18455, ys__n18456,
    ys__n18458, ys__n18459, ys__n18461, ys__n18462, ys__n18464, ys__n18465,
    ys__n18467, ys__n18468, ys__n18470, ys__n18471, ys__n18473, ys__n18474,
    ys__n18476, ys__n18477, ys__n18479, ys__n18480, ys__n18482, ys__n18483,
    ys__n18485, ys__n18486, ys__n18488, ys__n18489, ys__n18491, ys__n18492,
    ys__n18494, ys__n18495, ys__n18497, ys__n18498, ys__n18500, ys__n18501,
    ys__n18503, ys__n18504, ys__n18506, ys__n18507, ys__n18509, ys__n18510,
    ys__n18512, ys__n18513, ys__n18515, ys__n18516, ys__n18518, ys__n18519,
    ys__n18521, ys__n18522, ys__n18524, ys__n18525, ys__n18527, ys__n18528,
    ys__n18530, ys__n18531, ys__n18533, ys__n18534, ys__n18536, ys__n18537,
    ys__n18539, ys__n18540, ys__n18542, ys__n18543, ys__n18545, ys__n18547,
    ys__n18548, ys__n18549, ys__n18550, ys__n18551, ys__n18553, ys__n18554,
    ys__n18555, ys__n18557, ys__n18559, ys__n18561, ys__n18564, ys__n18567,
    ys__n18570, ys__n18573, ys__n18576, ys__n18579, ys__n18582, ys__n18585,
    ys__n18588, ys__n18591, ys__n18594, ys__n18597, ys__n18600, ys__n18603,
    ys__n18606, ys__n18609, ys__n18612, ys__n18615, ys__n18618, ys__n18621,
    ys__n18624, ys__n18627, ys__n18629, ys__n18631, ys__n18633, ys__n18635,
    ys__n18637, ys__n18640, ys__n18643, ys__n18646, ys__n18649, ys__n18652,
    ys__n18654, ys__n18655, ys__n18657, ys__n18658, ys__n18660, ys__n18661,
    ys__n18663, ys__n18664, ys__n18666, ys__n18667, ys__n18669, ys__n18670,
    ys__n18672, ys__n18673, ys__n18675, ys__n18676, ys__n18678, ys__n18679,
    ys__n18681, ys__n18682, ys__n18684, ys__n18685, ys__n18687, ys__n18688,
    ys__n18690, ys__n18691, ys__n18693, ys__n18694, ys__n18696, ys__n18697,
    ys__n18699, ys__n18700, ys__n18702, ys__n18703, ys__n18705, ys__n18706,
    ys__n18708, ys__n18709, ys__n18711, ys__n18712, ys__n18714, ys__n18715,
    ys__n18717, ys__n18718, ys__n18720, ys__n18721, ys__n18723, ys__n18724,
    ys__n18726, ys__n18727, ys__n18729, ys__n18730, ys__n18732, ys__n18733,
    ys__n18735, ys__n18736, ys__n18738, ys__n18739, ys__n18741, ys__n18742,
    ys__n18744, ys__n18745, ys__n18747, ys__n18748, ys__n18750, ys__n18751,
    ys__n18753, ys__n18754, ys__n18757, ys__n18759, ys__n18760, ys__n18763,
    ys__n18764, ys__n18766, ys__n18768, ys__n18770, ys__n18772, ys__n18774,
    ys__n18776, ys__n18778, ys__n18780, ys__n18782, ys__n18784, ys__n18786,
    ys__n18788, ys__n18790, ys__n18792, ys__n18794, ys__n18796, ys__n18798,
    ys__n18800, ys__n18802, ys__n18804, ys__n18806, ys__n18808, ys__n18810,
    ys__n18812, ys__n18814, ys__n18816, ys__n18818, ys__n18820, ys__n18822,
    ys__n18824, ys__n18826, ys__n19149, ys__n19151, ys__n19159, ys__n19173,
    ys__n19177, ys__n19178, ys__n19183, ys__n19227, ys__n19229, ys__n19231,
    ys__n19233, ys__n19235, ys__n19239, ys__n19254, ys__n19256, ys__n19257,
    ys__n19264, ys__n19266, ys__n19878, ys__n19881, ys__n19884, ys__n19887,
    ys__n19890, ys__n19893, ys__n19896, ys__n19899, ys__n19902, ys__n19905,
    ys__n19908, ys__n19911, ys__n19914, ys__n19917, ys__n19920, ys__n19923,
    ys__n19926, ys__n19929, ys__n19932, ys__n19935, ys__n19938, ys__n19941,
    ys__n19944, ys__n19947, ys__n19950, ys__n19953, ys__n19956, ys__n19959,
    ys__n19962, ys__n19965, ys__n19968, ys__n19971, ys__n20006, ys__n20007,
    ys__n20008, ys__n20009, ys__n20010, ys__n20011, ys__n20012, ys__n20013,
    ys__n20014, ys__n20015, ys__n20016, ys__n20017, ys__n20018, ys__n20019,
    ys__n20020, ys__n20021, ys__n20022, ys__n20023, ys__n20024, ys__n20025,
    ys__n20026, ys__n20027, ys__n20028, ys__n20029, ys__n20030, ys__n20031,
    ys__n20032, ys__n20033, ys__n20034, ys__n20038, ys__n20040, ys__n20043,
    ys__n20045, ys__n20053, ys__n20059, ys__n20062, ys__n20065, ys__n20068,
    ys__n20071, ys__n20074, ys__n20077, ys__n20080, ys__n20082, ys__n20084,
    ys__n20086, ys__n20088, ys__n20090, ys__n20092, ys__n20094, ys__n20096,
    ys__n20098, ys__n20100, ys__n20102, ys__n20104, ys__n20106, ys__n20108,
    ys__n20110, ys__n20112, ys__n20114, ys__n20116, ys__n20118, ys__n20120,
    ys__n20122, ys__n20124, ys__n20126, ys__n20128, ys__n22466, ys__n22919,
    ys__n22922, ys__n22925, ys__n22928, ys__n22931, ys__n22934, ys__n22937,
    ys__n22940, ys__n22943, ys__n22946, ys__n22949, ys__n22952, ys__n22955,
    ys__n22958, ys__n22961, ys__n22964, ys__n22967, ys__n22970, ys__n22973,
    ys__n22976, ys__n22979, ys__n22982, ys__n22985, ys__n22988, ys__n22991,
    ys__n22994, ys__n22997, ys__n23000, ys__n23003, ys__n23006, ys__n23009,
    ys__n23012, ys__n23263, ys__n23264, ys__n23340, ys__n23483, ys__n23485,
    ys__n23487, ys__n23489, ys__n23491, ys__n23493, ys__n23495, ys__n23497,
    ys__n23499, ys__n23501, ys__n23503, ys__n23505, ys__n23507, ys__n23509,
    ys__n23511, ys__n23513, ys__n23515, ys__n23517, ys__n23519, ys__n23521,
    ys__n23523, ys__n23525, ys__n23527, ys__n23529, ys__n23531, ys__n23533,
    ys__n23535, ys__n23537, ys__n23539, ys__n23541, ys__n23543, ys__n23635,
    ys__n23636, ys__n23764, ys__n23795, ys__n23798, ys__n23801, ys__n23804,
    ys__n23807, ys__n23853, ys__n23865, ys__n23868, ys__n23871, ys__n23874,
    ys__n23877, ys__n23921, ys__n23933, ys__n23936, ys__n23939, ys__n23942,
    ys__n23945, ys__n24099, ys__n24101, ys__n24102, ys__n24104, ys__n24105,
    ys__n24116, ys__n24118, ys__n24120, ys__n24126, ys__n24130, ys__n24134,
    ys__n24140, ys__n24145, ys__n24149, ys__n24154, ys__n24160, ys__n24162,
    ys__n24163, ys__n24165, ys__n24166, ys__n24176, ys__n24179, ys__n24180,
    ys__n24182, ys__n24183, ys__n24185, ys__n24186, ys__n24188, ys__n24189,
    ys__n24191, ys__n24192, ys__n24194, ys__n24195, ys__n24222, ys__n24227,
    ys__n24231, ys__n24236, ys__n24240, ys__n24245, ys__n24250, ys__n24255,
    ys__n24256, ys__n24258, ys__n24259, ys__n24260, ys__n24262, ys__n24265,
    ys__n24268, ys__n24271, ys__n24272, ys__n24274, ys__n24275, ys__n24277,
    ys__n24278, ys__n24286, ys__n24289, ys__n24291, ys__n24293, ys__n24295,
    ys__n24297, ys__n24299, ys__n24301, ys__n24305, ys__n24307, ys__n24309,
    ys__n24311, ys__n24313, ys__n24315, ys__n24317, ys__n24319, ys__n24320,
    ys__n24323, ys__n24325, ys__n24327, ys__n24329, ys__n24331, ys__n24333,
    ys__n24335, ys__n24339, ys__n24341, ys__n24343, ys__n24345, ys__n24347,
    ys__n24349, ys__n24351, ys__n24353, ys__n24354, ys__n24357, ys__n24359,
    ys__n24361, ys__n24363, ys__n24365, ys__n24367, ys__n24369, ys__n24373,
    ys__n24375, ys__n24377, ys__n24379, ys__n24381, ys__n24383, ys__n24385,
    ys__n24387, ys__n24388, ys__n24392, ys__n24394, ys__n24396, ys__n24398,
    ys__n24400, ys__n24402, ys__n24404, ys__n24408, ys__n24410, ys__n24412,
    ys__n24414, ys__n24416, ys__n24418, ys__n24420, ys__n24422, ys__n24425,
    ys__n24430, ys__n24436, ys__n24440, ys__n24445, ys__n24447, ys__n24466,
    ys__n24470, ys__n24488, ys__n24499, ys__n24502, ys__n24522, ys__n24532,
    ys__n24541, ys__n24552, ys__n24570, ys__n24573, ys__n24577, ys__n24579,
    ys__n24581, ys__n24585, ys__n24604, ys__n24713, ys__n24714, ys__n24742,
    ys__n24745, ys__n24748, ys__n24751, ys__n24754, ys__n24757, ys__n24760,
    ys__n24763, ys__n24766, ys__n24769, ys__n24772, ys__n24775, ys__n24778,
    ys__n24781, ys__n24784, ys__n24787, ys__n24790, ys__n24793, ys__n24796,
    ys__n24799, ys__n24802, ys__n24805, ys__n24808, ys__n24811, ys__n24814,
    ys__n24817, ys__n24820, ys__n24823, ys__n24826, ys__n24829, ys__n24832,
    ys__n24835, ys__n24837, ys__n24839, ys__n24907, ys__n24910, ys__n24913,
    ys__n24916, ys__n24919, ys__n24922, ys__n24925, ys__n24928, ys__n24931,
    ys__n24934, ys__n24937, ys__n24940, ys__n24943, ys__n24946, ys__n24949,
    ys__n24952, ys__n24955, ys__n25294, ys__n25302, ys__n25304, ys__n25306,
    ys__n25308, ys__n25310, ys__n25385, ys__n25386, ys__n25387, ys__n25388,
    ys__n25390, ys__n25406, ys__n25421, ys__n25430, ys__n25431, ys__n25432,
    ys__n25433, ys__n25434, ys__n25435, ys__n25436, ys__n25438, ys__n25441,
    ys__n25449, ys__n25456, ys__n25461, ys__n25463, ys__n25465, ys__n25467,
    ys__n25469, ys__n25472, ys__n25486, ys__n25496, ys__n25504, ys__n25519,
    ys__n25522, ys__n25534, ys__n25550, ys__n25661, ys__n25663, ys__n25665,
    ys__n25667, ys__n25669, ys__n25671, ys__n25673, ys__n25675, ys__n25677,
    ys__n25679, ys__n25681, ys__n25683, ys__n25685, ys__n25687, ys__n25689,
    ys__n25691, ys__n25693, ys__n25695, ys__n25697, ys__n25699, ys__n25701,
    ys__n25703, ys__n25705, ys__n25707, ys__n25709, ys__n25711, ys__n25713,
    ys__n25715, ys__n25717, ys__n25719, ys__n25721, ys__n25723, ys__n25725,
    ys__n25830, ys__n25833, ys__n25836, ys__n25839, ys__n25842, ys__n25844,
    ys__n25846, ys__n25852, ys__n25957, ys__n25960, ys__n25963, ys__n25966,
    ys__n26118, ys__n26119, ys__n26120, ys__n26121, ys__n26122, ys__n26123,
    ys__n26124, ys__n26125, ys__n26126, ys__n26127, ys__n26128, ys__n26129,
    ys__n26130, ys__n26131, ys__n26132, ys__n26133, ys__n26134, ys__n26135,
    ys__n26136, ys__n26137, ys__n26138, ys__n26139, ys__n26141, ys__n26144,
    ys__n26146, ys__n26148, ys__n26150, ys__n26152, ys__n26154, ys__n26156,
    ys__n26158, ys__n26160, ys__n26220, ys__n26222, ys__n26224, ys__n26226,
    ys__n26228, ys__n26230, ys__n26232, ys__n26234, ys__n26236, ys__n26238,
    ys__n26240, ys__n26242, ys__n26244, ys__n26246, ys__n26248, ys__n26250,
    ys__n26252, ys__n26254, ys__n26256, ys__n26258, ys__n26260, ys__n26262,
    ys__n26264, ys__n26266, ys__n26268, ys__n26270, ys__n26272, ys__n26274,
    ys__n26276, ys__n26278, ys__n26282, ys__n26284, ys__n26286, ys__n26288,
    ys__n26291, ys__n26293, ys__n26294, ys__n26555, ys__n26566, ys__n26573,
    ys__n26607, ys__n26609, ys__n26611, ys__n26613, ys__n26615, ys__n26617,
    ys__n26619, ys__n26621, ys__n26623, ys__n26625, ys__n26627, ys__n26629,
    ys__n26631, ys__n26633, ys__n26635, ys__n26637, ys__n26639, ys__n26641,
    ys__n26643, ys__n26645, ys__n26647, ys__n26649, ys__n26651, ys__n26653,
    ys__n26655, ys__n26657, ys__n26659, ys__n26661, ys__n26663, ys__n26665,
    ys__n26667, ys__n26669, ys__n26671, ys__n26673, ys__n26675, ys__n26677,
    ys__n26679, ys__n26681, ys__n26683, ys__n26685, ys__n26687, ys__n26689,
    ys__n26691, ys__n26693, ys__n26695, ys__n26697, ys__n26699, ys__n26701,
    ys__n26703, ys__n26705, ys__n26707, ys__n26709, ys__n26711, ys__n26713,
    ys__n26715, ys__n26717, ys__n26719, ys__n26721, ys__n26723, ys__n26725,
    ys__n26727, ys__n26729, ys__n26731, ys__n26733, ys__n26734, ys__n26735,
    ys__n26736, ys__n26737, ys__n26738, ys__n26739, ys__n26740, ys__n26741,
    ys__n26742, ys__n26743, ys__n26744, ys__n26745, ys__n26746, ys__n26747,
    ys__n26748, ys__n26749, ys__n26750, ys__n26751, ys__n26752, ys__n26753,
    ys__n26754, ys__n26755, ys__n26756, ys__n26757, ys__n26758, ys__n26759,
    ys__n26760, ys__n26761, ys__n26762, ys__n26763, ys__n26764, ys__n26765,
    ys__n26802, ys__n26803, ys__n26804, ys__n26805, ys__n26806, ys__n26807,
    ys__n26808, ys__n26809, ys__n26810, ys__n26811, ys__n26812, ys__n26813,
    ys__n26814, ys__n26815, ys__n26816, ys__n26817, ys__n26818, ys__n26819,
    ys__n26820, ys__n26821, ys__n26822, ys__n26823, ys__n26824, ys__n26825,
    ys__n26826, ys__n26827, ys__n26828, ys__n26829, ys__n26830, ys__n26831,
    ys__n26832, ys__n26833, ys__n26834, ys__n26835, ys__n26836, ys__n26837,
    ys__n26838, ys__n26839, ys__n26840, ys__n26841, ys__n26842, ys__n26843,
    ys__n26844, ys__n26845, ys__n26846, ys__n26847, ys__n26848, ys__n26849,
    ys__n26850, ys__n26851, ys__n26852, ys__n26853, ys__n26854, ys__n26855,
    ys__n26856, ys__n26857, ys__n26858, ys__n26859, ys__n26860, ys__n26861,
    ys__n26862, ys__n26863, ys__n26864, ys__n26865, ys__n26866, ys__n26867,
    ys__n26868, ys__n26869, ys__n26870, ys__n26871, ys__n26872, ys__n26873,
    ys__n26874, ys__n26875, ys__n26876, ys__n26877, ys__n26878, ys__n26879,
    ys__n26880, ys__n26881, ys__n26882, ys__n26883, ys__n26884, ys__n26885,
    ys__n26886, ys__n26887, ys__n26888, ys__n26889, ys__n26890, ys__n26891,
    ys__n26892, ys__n26893, ys__n26894, ys__n26895, ys__n26896, ys__n26897,
    ys__n26898, ys__n26899, ys__n26900, ys__n26901, ys__n26902, ys__n26903,
    ys__n26904, ys__n26905, ys__n26906, ys__n26907, ys__n26908, ys__n26909,
    ys__n26910, ys__n26911, ys__n26912, ys__n26913, ys__n26914, ys__n26915,
    ys__n26916, ys__n26917, ys__n26918, ys__n26919, ys__n26920, ys__n26921,
    ys__n26922, ys__n26923, ys__n26924, ys__n26925, ys__n26926, ys__n26927,
    ys__n26928, ys__n26929, ys__n26930, ys__n26931, ys__n26932, ys__n26933,
    ys__n26934, ys__n26935, ys__n26936, ys__n26937, ys__n26938, ys__n26939,
    ys__n26940, ys__n26941, ys__n26942, ys__n26943, ys__n26944, ys__n26945,
    ys__n26946, ys__n26947, ys__n26948, ys__n26949, ys__n26950, ys__n26951,
    ys__n26952, ys__n26953, ys__n26954, ys__n26955, ys__n26956, ys__n26957,
    ys__n26958, ys__n26959, ys__n26960, ys__n26961, ys__n26962, ys__n26963,
    ys__n26964, ys__n26965, ys__n26966, ys__n26967, ys__n26968, ys__n26969,
    ys__n26970, ys__n26971, ys__n26972, ys__n26973, ys__n26974, ys__n26975,
    ys__n26976, ys__n26977, ys__n26978, ys__n26979, ys__n26980, ys__n26981,
    ys__n26982, ys__n26983, ys__n26984, ys__n26985, ys__n26986, ys__n26987,
    ys__n26988, ys__n26989, ys__n26990, ys__n26991, ys__n26992, ys__n26993,
    ys__n26994, ys__n26995, ys__n26996, ys__n26997, ys__n26998, ys__n26999,
    ys__n27000, ys__n27001, ys__n27002, ys__n27003, ys__n27004, ys__n27005,
    ys__n27006, ys__n27007, ys__n27008, ys__n27009, ys__n27010, ys__n27011,
    ys__n27012, ys__n27013, ys__n27014, ys__n27015, ys__n27016, ys__n27017,
    ys__n27018, ys__n27019, ys__n27020, ys__n27021, ys__n27022, ys__n27023,
    ys__n27024, ys__n27025, ys__n27026, ys__n27027, ys__n27028, ys__n27029,
    ys__n27030, ys__n27031, ys__n27032, ys__n27033, ys__n27034, ys__n27035,
    ys__n27036, ys__n27037, ys__n27038, ys__n27039, ys__n27040, ys__n27041,
    ys__n27042, ys__n27043, ys__n27044, ys__n27045, ys__n27046, ys__n27047,
    ys__n27048, ys__n27049, ys__n27050, ys__n27051, ys__n27052, ys__n27053,
    ys__n27054, ys__n27055, ys__n27056, ys__n27057, ys__n27058, ys__n27059,
    ys__n27060, ys__n27061, ys__n27062, ys__n27063, ys__n27064, ys__n27065,
    ys__n27066, ys__n27067, ys__n27068, ys__n27069, ys__n27070, ys__n27071,
    ys__n27072, ys__n27073, ys__n27074, ys__n27075, ys__n27076, ys__n27077,
    ys__n27078, ys__n27079, ys__n27080, ys__n27081, ys__n27082, ys__n27083,
    ys__n27084, ys__n27085, ys__n27086, ys__n27087, ys__n27088, ys__n27089,
    ys__n27090, ys__n27091, ys__n27092, ys__n27093, ys__n27094, ys__n27095,
    ys__n27096, ys__n27097, ys__n27098, ys__n27099, ys__n27100, ys__n27101,
    ys__n27102, ys__n27103, ys__n27104, ys__n27105, ys__n27106, ys__n27107,
    ys__n27108, ys__n27109, ys__n27110, ys__n27111, ys__n27112, ys__n27113,
    ys__n27114, ys__n27115, ys__n27116, ys__n27117, ys__n27118, ys__n27119,
    ys__n27120, ys__n27121, ys__n27122, ys__n27123, ys__n27124, ys__n27125,
    ys__n27126, ys__n27127, ys__n27128, ys__n27129, ys__n27130, ys__n27131,
    ys__n27132, ys__n27133, ys__n27134, ys__n27135, ys__n27136, ys__n27137,
    ys__n27138, ys__n27139, ys__n27140, ys__n27141, ys__n27142, ys__n27143,
    ys__n27144, ys__n27145, ys__n27146, ys__n27147, ys__n27148, ys__n27149,
    ys__n27150, ys__n27151, ys__n27152, ys__n27153, ys__n27154, ys__n27155,
    ys__n27156, ys__n27157, ys__n27158, ys__n27159, ys__n27160, ys__n27161,
    ys__n27162, ys__n27163, ys__n27164, ys__n27165, ys__n27166, ys__n27167,
    ys__n27168, ys__n27169, ys__n27170, ys__n27171, ys__n27172, ys__n27173,
    ys__n27174, ys__n27175, ys__n27176, ys__n27177, ys__n27178, ys__n27179,
    ys__n27180, ys__n27181, ys__n27182, ys__n27183, ys__n27184, ys__n27185,
    ys__n27186, ys__n27187, ys__n27188, ys__n27189, ys__n27190, ys__n27191,
    ys__n27192, ys__n27193, ys__n27194, ys__n27195, ys__n27196, ys__n27197,
    ys__n27198, ys__n27199, ys__n27200, ys__n27201, ys__n27202, ys__n27203,
    ys__n27204, ys__n27205, ys__n27206, ys__n27207, ys__n27208, ys__n27209,
    ys__n27210, ys__n27211, ys__n27212, ys__n27213, ys__n27214, ys__n27215,
    ys__n27216, ys__n27217, ys__n27218, ys__n27219, ys__n27220, ys__n27221,
    ys__n27222, ys__n27223, ys__n27224, ys__n27225, ys__n27226, ys__n27227,
    ys__n27228, ys__n27229, ys__n27230, ys__n27231, ys__n27232, ys__n27233,
    ys__n27234, ys__n27235, ys__n27236, ys__n27237, ys__n27238, ys__n27239,
    ys__n27240, ys__n27241, ys__n27242, ys__n27243, ys__n27244, ys__n27245,
    ys__n27246, ys__n27247, ys__n27248, ys__n27249, ys__n27250, ys__n27251,
    ys__n27252, ys__n27253, ys__n27254, ys__n27255, ys__n27256, ys__n27257,
    ys__n27258, ys__n27259, ys__n27260, ys__n27261, ys__n27262, ys__n27263,
    ys__n27264, ys__n27265, ys__n27266, ys__n27267, ys__n27268, ys__n27269,
    ys__n27270, ys__n27271, ys__n27272, ys__n27273, ys__n27274, ys__n27275,
    ys__n27276, ys__n27277, ys__n27278, ys__n27279, ys__n27280, ys__n27281,
    ys__n27282, ys__n27283, ys__n27284, ys__n27285, ys__n27286, ys__n27287,
    ys__n27288, ys__n27289, ys__n27290, ys__n27291, ys__n27292, ys__n27293,
    ys__n27294, ys__n27295, ys__n27296, ys__n27297, ys__n27298, ys__n27299,
    ys__n27300, ys__n27301, ys__n27302, ys__n27303, ys__n27304, ys__n27305,
    ys__n27306, ys__n27307, ys__n27308, ys__n27309, ys__n27310, ys__n27311,
    ys__n27312, ys__n27313, ys__n27314, ys__n27315, ys__n27316, ys__n27317,
    ys__n27318, ys__n27319, ys__n27320, ys__n27321, ys__n27322, ys__n27323,
    ys__n27324, ys__n27325, ys__n27326, ys__n27327, ys__n27328, ys__n27329,
    ys__n27330, ys__n27331, ys__n27332, ys__n27333, ys__n27334, ys__n27335,
    ys__n27336, ys__n27337, ys__n27338, ys__n27339, ys__n27340, ys__n27341,
    ys__n27342, ys__n27343, ys__n27344, ys__n27345, ys__n27346, ys__n27347,
    ys__n27348, ys__n27349, ys__n27350, ys__n27351, ys__n27352, ys__n27353,
    ys__n27354, ys__n27355, ys__n27356, ys__n27357, ys__n27358, ys__n27359,
    ys__n27360, ys__n27361, ys__n27362, ys__n27363, ys__n27364, ys__n27365,
    ys__n27366, ys__n27367, ys__n27368, ys__n27369, ys__n27370, ys__n27371,
    ys__n27372, ys__n27373, ys__n27374, ys__n27375, ys__n27376, ys__n27377,
    ys__n27378, ys__n27379, ys__n27380, ys__n27381, ys__n27382, ys__n27383,
    ys__n27384, ys__n27385, ys__n27386, ys__n27387, ys__n27388, ys__n27389,
    ys__n27390, ys__n27391, ys__n27392, ys__n27393, ys__n27394, ys__n27395,
    ys__n27396, ys__n27397, ys__n27398, ys__n27399, ys__n27400, ys__n27401,
    ys__n27402, ys__n27403, ys__n27404, ys__n27405, ys__n27406, ys__n27407,
    ys__n27408, ys__n27409, ys__n27410, ys__n27411, ys__n27412, ys__n27413,
    ys__n27414, ys__n27415, ys__n27416, ys__n27417, ys__n27418, ys__n27419,
    ys__n27420, ys__n27421, ys__n27422, ys__n27423, ys__n27424, ys__n27425,
    ys__n27426, ys__n27427, ys__n27428, ys__n27429, ys__n27430, ys__n27431,
    ys__n27432, ys__n27433, ys__n27434, ys__n27435, ys__n27436, ys__n27437,
    ys__n27484, ys__n27493, ys__n27504, ys__n27513, ys__n27515, ys__n27517,
    ys__n27550, ys__n27551, ys__n27598, ys__n27603, ys__n27605, ys__n27610,
    ys__n27613, ys__n27616, ys__n27619, ys__n27622, ys__n27625, ys__n27628,
    ys__n27631, ys__n27634, ys__n27637, ys__n27640, ys__n27643, ys__n27646,
    ys__n27649, ys__n27652, ys__n27655, ys__n27658, ys__n27661, ys__n27664,
    ys__n27667, ys__n27670, ys__n27673, ys__n27676, ys__n27679, ys__n27682,
    ys__n27685, ys__n27688, ys__n27691, ys__n27694, ys__n27697, ys__n27700,
    ys__n27703, ys__n27705, ys__n27706, ys__n27707, ys__n27708, ys__n27709,
    ys__n27710, ys__n27711, ys__n27712, ys__n27713, ys__n27714, ys__n27715,
    ys__n27716, ys__n27717, ys__n27718, ys__n27719, ys__n27720, ys__n27721,
    ys__n27722, ys__n27723, ys__n27724, ys__n27725, ys__n27726, ys__n27727,
    ys__n27728, ys__n27729, ys__n27730, ys__n27731, ys__n27732, ys__n27733,
    ys__n27734, ys__n27735, ys__n27736, ys__n27739, ys__n27741, ys__n28247,
    ys__n28249, ys__n28250, ys__n28251, ys__n28252, ys__n28254, ys__n28256,
    ys__n28258, ys__n28259, ys__n28261, ys__n28263, ys__n28265, ys__n28266,
    ys__n28268, ys__n28269, ys__n28270, ys__n28271, ys__n28272, ys__n28274,
    ys__n28276, ys__n28328, ys__n28330, ys__n28332, ys__n28334, ys__n28336,
    ys__n28343, ys__n28345, ys__n28347, ys__n28349, ys__n28351, ys__n28353,
    ys__n28355, ys__n28357, ys__n28359, ys__n28361, ys__n28363, ys__n28365,
    ys__n28367, ys__n28369, ys__n28371, ys__n28373, ys__n28375, ys__n28377,
    ys__n28379, ys__n28381, ys__n28383, ys__n28385, ys__n28387, ys__n28389,
    ys__n28391, ys__n28393, ys__n28395, ys__n28397, ys__n28399, ys__n28401,
    ys__n28403, ys__n28406, ys__n28409, ys__n28410, ys__n28411, ys__n28412,
    ys__n28413, ys__n28414, ys__n28415, ys__n28416, ys__n28417, ys__n28418,
    ys__n28419, ys__n28420, ys__n28421, ys__n28422, ys__n28423, ys__n28425,
    ys__n28427, ys__n28429, ys__n28431, ys__n28433, ys__n28435, ys__n28437,
    ys__n28439, ys__n28440, ys__n28441, ys__n28442, ys__n28443, ys__n28444,
    ys__n28445, ys__n28447, ys__n28448, ys__n28449, ys__n28450, ys__n28451,
    ys__n28452, ys__n28454, ys__n28456, ys__n28458, ys__n28460, ys__n28475,
    ys__n28476, ys__n28477, ys__n28478, ys__n28479, ys__n28480, ys__n28481,
    ys__n28482, ys__n28483, ys__n28484, ys__n28485, ys__n28486, ys__n28487,
    ys__n28488, ys__n28489, ys__n28490, ys__n28491, ys__n28492, ys__n28493,
    ys__n28494, ys__n28495, ys__n28496, ys__n28497, ys__n28498, ys__n28499,
    ys__n28500, ys__n28501, ys__n28502, ys__n28503, ys__n28504, ys__n28505,
    ys__n28506, ys__n28510, ys__n28513, ys__n28518, ys__n28533, ys__n28536,
    ys__n28539, ys__n28542, ys__n28545, ys__n28548, ys__n28551, ys__n28554,
    ys__n28557, ys__n28560, ys__n28563, ys__n28566, ys__n28569, ys__n28572,
    ys__n28575, ys__n28578, ys__n28581, ys__n28584, ys__n28587, ys__n28661,
    ys__n28662, ys__n28781, ys__n28782, ys__n28783, ys__n28784, ys__n28785,
    ys__n28786, ys__n28787, ys__n28788, ys__n28789, ys__n28790, ys__n28791,
    ys__n28792, ys__n28793, ys__n28794, ys__n28796, ys__n28798, ys__n28800,
    ys__n28802, ys__n28804, ys__n28806, ys__n28808, ys__n28810, ys__n28812,
    ys__n28814, ys__n28816, ys__n28818, ys__n28820, ys__n28822, ys__n28824,
    ys__n28826, ys__n28828, ys__n28830, ys__n28832, ys__n28834, ys__n28836,
    ys__n28838, ys__n28840, ys__n28842, ys__n28844, ys__n28846, ys__n28848,
    ys__n28850, ys__n28852, ys__n28854, ys__n28856, ys__n28858, ys__n29022,
    ys__n29025, ys__n29028, ys__n29031, ys__n29034, ys__n29037, ys__n29040,
    ys__n29043, ys__n29046, ys__n29049, ys__n29052, ys__n29055, ys__n29058,
    ys__n29061, ys__n29064, ys__n29067, ys__n29070, ys__n29073, ys__n29076,
    ys__n29079, ys__n29082, ys__n29085, ys__n29088, ys__n29091, ys__n29094,
    ys__n29097, ys__n29100, ys__n29103, ys__n29106, ys__n29109, ys__n29112,
    ys__n29115, ys__n29118, ys__n29122, ys__n29125, ys__n29128, ys__n29131,
    ys__n29134, ys__n29137, ys__n29140, ys__n29143, ys__n29146, ys__n29149,
    ys__n29152, ys__n29155, ys__n29158, ys__n29161, ys__n29164, ys__n29167,
    ys__n29170, ys__n29173, ys__n29176, ys__n29179, ys__n29182, ys__n29185,
    ys__n29188, ys__n29191, ys__n29194, ys__n29197, ys__n29200, ys__n29203,
    ys__n29206, ys__n29209, ys__n29212, ys__n29215, ys__n29217, ys__n29219,
    ys__n29221, ys__n29223, ys__n29225, ys__n29226, ys__n29227, ys__n29228,
    ys__n29229, ys__n29230, ys__n29231, ys__n29232, ys__n29233, ys__n29234,
    ys__n29235, ys__n29336, ys__n29339, ys__n29342, ys__n29345, ys__n29348,
    ys__n29351, ys__n29354, ys__n29357, ys__n29360, ys__n29363, ys__n29366,
    ys__n29369, ys__n29372, ys__n29375, ys__n29378, ys__n29381, ys__n29384,
    ys__n29387, ys__n29390, ys__n29393, ys__n29396, ys__n29399, ys__n29402,
    ys__n29405, ys__n29408, ys__n29411, ys__n29414, ys__n29417, ys__n29420,
    ys__n29423, ys__n29426, ys__n29429, ys__n29431, ys__n29435, ys__n29438,
    ys__n29441, ys__n29444, ys__n29447, ys__n29450, ys__n29453, ys__n29456,
    ys__n29459, ys__n29462, ys__n29465, ys__n29468, ys__n29471, ys__n29474,
    ys__n29477, ys__n29480, ys__n29483, ys__n29486, ys__n29489, ys__n29492,
    ys__n29495, ys__n29498, ys__n29501, ys__n29504, ys__n29507, ys__n29510,
    ys__n29513, ys__n29516, ys__n29519, ys__n29522, ys__n29525, ys__n29528,
    ys__n29530, ys__n29532, ys__n29534, ys__n29536, ys__n29538, ys__n29539,
    ys__n29540, ys__n29541, ys__n29542, ys__n29543, ys__n29544, ys__n29545,
    ys__n29546, ys__n29547, ys__n29548, ys__n29611, ys__n29614, ys__n29617,
    ys__n29620, ys__n29623, ys__n29626, ys__n29629, ys__n29632, ys__n29635,
    ys__n29638, ys__n29641, ys__n29644, ys__n29647, ys__n29650, ys__n29653,
    ys__n29656, ys__n29659, ys__n29662, ys__n29665, ys__n29668, ys__n29671,
    ys__n29674, ys__n29677, ys__n29680, ys__n29683, ys__n29686, ys__n29689,
    ys__n29692, ys__n29695, ys__n29698, ys__n29701, ys__n29704, ys__n29706,
    ys__n29710, ys__n29713, ys__n29716, ys__n29719, ys__n29722, ys__n29725,
    ys__n29728, ys__n29731, ys__n29734, ys__n29737, ys__n29740, ys__n29743,
    ys__n29746, ys__n29749, ys__n29752, ys__n29755, ys__n29758, ys__n29761,
    ys__n29764, ys__n29767, ys__n29770, ys__n29773, ys__n29776, ys__n29779,
    ys__n29782, ys__n29785, ys__n29788, ys__n29791, ys__n29794, ys__n29797,
    ys__n29800, ys__n29803, ys__n29805, ys__n29807, ys__n29809, ys__n29811,
    ys__n29813, ys__n29814, ys__n29815, ys__n29816, ys__n29817, ys__n29818,
    ys__n29819, ys__n29820, ys__n29821, ys__n29822, ys__n29823, ys__n29847,
    ys__n30010, ys__n30080, ys__n30081, ys__n30082, ys__n30083, ys__n30084,
    ys__n30085, ys__n30086, ys__n30087, ys__n30089, ys__n30090, ys__n30091,
    ys__n30092, ys__n30093, ys__n30094, ys__n30095, ys__n30096, ys__n30098,
    ys__n30099, ys__n30100, ys__n30101, ys__n30102, ys__n30103, ys__n30104,
    ys__n30105, ys__n30106, ys__n30107, ys__n30108, ys__n30109, ys__n30110,
    ys__n30111, ys__n30112, ys__n30113, ys__n30119, ys__n30122, ys__n30125,
    ys__n30128, ys__n30131, ys__n30134, ys__n30137, ys__n30140, ys__n30143,
    ys__n30146, ys__n30149, ys__n30152, ys__n30155, ys__n30158, ys__n30161,
    ys__n30164, ys__n30167, ys__n30170, ys__n30173, ys__n30176, ys__n30179,
    ys__n30182, ys__n30185, ys__n30188, ys__n30191, ys__n30194, ys__n30197,
    ys__n30200, ys__n30203, ys__n30206, ys__n30209, ys__n30212, ys__n30215,
    ys__n30223, ys__n30226, ys__n30235, ys__n30238, ys__n30241, ys__n30244,
    ys__n30247, ys__n30250, ys__n30253, ys__n30256, ys__n30259, ys__n30262,
    ys__n30265, ys__n30268, ys__n30271, ys__n30274, ys__n30277, ys__n30280,
    ys__n30283, ys__n30286, ys__n30289, ys__n30292, ys__n30295, ys__n30298,
    ys__n30301, ys__n30304, ys__n30307, ys__n30310, ys__n30313, ys__n30316,
    ys__n30319, ys__n30322, ys__n30325, ys__n30328, ys__n30330, ys__n30331,
    ys__n30616, ys__n30619, ys__n30622, ys__n30625, ys__n30628, ys__n30631,
    ys__n30634, ys__n30637, ys__n30640, ys__n30643, ys__n30646, ys__n30649,
    ys__n30652, ys__n30655, ys__n30658, ys__n30661, ys__n30664, ys__n30667,
    ys__n30668, ys__n30670, ys__n30797, ys__n30798, ys__n30799, ys__n30800,
    ys__n30801, ys__n30802, ys__n30803, ys__n30804, ys__n30805, ys__n30806,
    ys__n30807, ys__n30808, ys__n30809, ys__n30810, ys__n30811, ys__n30812,
    ys__n30813, ys__n30832, ys__n30833, ys__n30835, ys__n30836, ys__n30856,
    ys__n30858, ys__n30860, ys__n30864, ys__n30873, ys__n30874, ys__n30875,
    ys__n30876, ys__n30942, ys__n30943, ys__n30944, ys__n30945, ys__n30946,
    ys__n30947, ys__n30948, ys__n30949, ys__n30950, ys__n30951, ys__n30952,
    ys__n30953, ys__n30954, ys__n30955, ys__n30956, ys__n31202, ys__n31203,
    ys__n31207, ys__n31208, ys__n31209, ys__n31210, ys__n31211, ys__n31212,
    ys__n31213, ys__n31214, ys__n31215, ys__n31216, ys__n31217, ys__n31218,
    ys__n31219, ys__n31220, ys__n31221, ys__n31222, ys__n31223, ys__n31224,
    ys__n31225, ys__n31226, ys__n31227, ys__n31228, ys__n31229, ys__n31230,
    ys__n31231, ys__n31232, ys__n31233, ys__n31234, ys__n31235, ys__n31236,
    ys__n31237, ys__n31238, ys__n31326, ys__n31327, ys__n31328, ys__n31329,
    ys__n31330, ys__n31331, ys__n31332, ys__n31333, ys__n31334, ys__n31335,
    ys__n31336, ys__n31337, ys__n31338, ys__n31339, ys__n31340, ys__n31341,
    ys__n31342, ys__n31343, ys__n31344, ys__n31345, ys__n31346, ys__n31347,
    ys__n31348, ys__n31349, ys__n31350, ys__n31351, ys__n31352, ys__n31353,
    ys__n31354, ys__n31355, ys__n31356, ys__n31357, ys__n31358, ys__n31359,
    ys__n31360, ys__n31361, ys__n31362, ys__n31363, ys__n31364, ys__n31365,
    ys__n31366, ys__n31367, ys__n31368, ys__n31369, ys__n31370, ys__n31371,
    ys__n31372, ys__n31373, ys__n31374, ys__n31375, ys__n31376, ys__n31377,
    ys__n31378, ys__n31379, ys__n31380, ys__n31381, ys__n31382, ys__n31383,
    ys__n31384, ys__n31385, ys__n31386, ys__n31387, ys__n31388, ys__n31389,
    ys__n31390, ys__n31391, ys__n31392, ys__n31393, ys__n31394, ys__n31395,
    ys__n31397, ys__n31398, ys__n31399, ys__n31400, ys__n31401, ys__n31402,
    ys__n31403, ys__n31404, ys__n31405, ys__n31406, ys__n31407, ys__n31408,
    ys__n31409, ys__n31410, ys__n31411, ys__n31412, ys__n31413, ys__n31414,
    ys__n31415, ys__n31416, ys__n31417, ys__n31418, ys__n31419, ys__n31420,
    ys__n31421, ys__n31422, ys__n31423, ys__n31424, ys__n31425, ys__n31426,
    ys__n31427, ys__n31428, ys__n31429, ys__n31430, ys__n31431, ys__n31432,
    ys__n31433, ys__n31434, ys__n31435, ys__n31436, ys__n31437, ys__n31438,
    ys__n31439, ys__n31440, ys__n31441, ys__n31442, ys__n31443, ys__n31444,
    ys__n31445, ys__n31446, ys__n31447, ys__n31448, ys__n31449, ys__n31450,
    ys__n31451, ys__n31452, ys__n31453, ys__n31454, ys__n31455, ys__n31456,
    ys__n31457, ys__n31458, ys__n31459, ys__n31460, ys__n31461, ys__n31462,
    ys__n31463, ys__n31464, ys__n31465, ys__n31466, ys__n31467, ys__n31468,
    ys__n31469, ys__n31470, ys__n31471, ys__n31472, ys__n31473, ys__n31474,
    ys__n31475, ys__n31476, ys__n31477, ys__n31478, ys__n31479, ys__n31480,
    ys__n31481, ys__n31482, ys__n31483, ys__n31484, ys__n31485, ys__n31486,
    ys__n31487, ys__n31488, ys__n31489, ys__n31490, ys__n31491, ys__n31492,
    ys__n31493, ys__n31494, ys__n31495, ys__n31496, ys__n31497, ys__n31498,
    ys__n31499, ys__n31500, ys__n31501, ys__n31502, ys__n31503, ys__n31504,
    ys__n31505, ys__n31506, ys__n31507, ys__n31508, ys__n31509, ys__n31510,
    ys__n31511, ys__n31512, ys__n31513, ys__n31514, ys__n31515, ys__n31516,
    ys__n31517, ys__n31518, ys__n31519, ys__n31520, ys__n31521, ys__n31522,
    ys__n31523, ys__n31524, ys__n31525, ys__n31526, ys__n31527, ys__n31528,
    ys__n31529, ys__n31530, ys__n31531, ys__n31532, ys__n31533, ys__n31534,
    ys__n31535, ys__n31536, ys__n31537, ys__n31538, ys__n31539, ys__n31540,
    ys__n31541, ys__n31542, ys__n31543, ys__n31544, ys__n31559, ys__n31560,
    ys__n31562, ys__n31564, ys__n31567, ys__n31571, ys__n31740, ys__n31741,
    ys__n31742, ys__n31743, ys__n31744, ys__n31745, ys__n31746, ys__n31747,
    ys__n31748, ys__n31749, ys__n31750, ys__n31751, ys__n31752, ys__n31753,
    ys__n31754, ys__n31755, ys__n31756, ys__n31757, ys__n31758, ys__n31759,
    ys__n31760, ys__n31761, ys__n31762, ys__n31763, ys__n31764, ys__n31765,
    ys__n31766, ys__n31767, ys__n31768, ys__n31769, ys__n31770, ys__n31771,
    ys__n31772, ys__n31773, ys__n31774, ys__n31775, ys__n31776, ys__n31777,
    ys__n31778, ys__n31779, ys__n31780, ys__n31781, ys__n31782, ys__n31783,
    ys__n31784, ys__n31785, ys__n31786, ys__n31787, ys__n31788, ys__n31789,
    ys__n31790, ys__n31791, ys__n31792, ys__n31793, ys__n31794, ys__n31795,
    ys__n31796, ys__n31797, ys__n31798, ys__n31799, ys__n31800, ys__n31801,
    ys__n31802, ys__n31803, ys__n31804, ys__n31805, ys__n31806, ys__n31807,
    ys__n31808, ys__n31809, ys__n31810, ys__n31811, ys__n31812, ys__n31813,
    ys__n31814, ys__n31815, ys__n31816, ys__n31817, ys__n31818, ys__n31819,
    ys__n31820, ys__n31821, ys__n31822, ys__n31823, ys__n31824, ys__n31825,
    ys__n31826, ys__n31827, ys__n31828, ys__n31829, ys__n31830, ys__n31831,
    ys__n31832, ys__n31833, ys__n31834, ys__n31835, ys__n31836, ys__n31837,
    ys__n31838, ys__n31839, ys__n31840, ys__n31841, ys__n31842, ys__n31843,
    ys__n31844, ys__n31845, ys__n31846, ys__n31847, ys__n31848, ys__n31849,
    ys__n31850, ys__n31851, ys__n31852, ys__n31853, ys__n31854, ys__n31855,
    ys__n31856, ys__n31857, ys__n31858, ys__n31859, ys__n31860, ys__n31861,
    ys__n31862, ys__n31863, ys__n31864, ys__n31865, ys__n31866, ys__n31867,
    ys__n31868, ys__n31869, ys__n31870, ys__n31871, ys__n31872, ys__n31873,
    ys__n31874, ys__n31875, ys__n31876, ys__n31877, ys__n31878, ys__n31879,
    ys__n31880, ys__n31881, ys__n31882, ys__n31883, ys__n31884, ys__n31885,
    ys__n31886, ys__n31887, ys__n31888, ys__n31889, ys__n31890, ys__n31891,
    ys__n31892, ys__n31893, ys__n31894, ys__n31895, ys__n31896, ys__n31897,
    ys__n31898, ys__n31899, ys__n31900, ys__n31901, ys__n31902, ys__n31903,
    ys__n31904, ys__n31905, ys__n31906, ys__n31907, ys__n31908, ys__n31909,
    ys__n31910, ys__n31911, ys__n31912, ys__n31913, ys__n31914, ys__n31915,
    ys__n31916, ys__n31917, ys__n31918, ys__n31919, ys__n31920, ys__n31921,
    ys__n31922, ys__n31923, ys__n31924, ys__n31925, ys__n31926, ys__n31927,
    ys__n31928, ys__n31929, ys__n31930, ys__n31931, ys__n31932, ys__n31933,
    ys__n31934, ys__n31935, ys__n31936, ys__n31937, ys__n31938, ys__n31939,
    ys__n31940, ys__n31941, ys__n31942, ys__n31943, ys__n31944, ys__n31945,
    ys__n31946, ys__n31947, ys__n31948, ys__n31949, ys__n31950, ys__n31953,
    ys__n31954, ys__n31955, ys__n31965, ys__n31971, ys__n31973, ys__n31975,
    ys__n31976, ys__n31978, ys__n31979, ys__n31984, ys__n31986, ys__n31988,
    ys__n31990, ys__n31992, ys__n31994, ys__n31996, ys__n31998, ys__n32000,
    ys__n32002, ys__n32004, ys__n32006, ys__n32007, ys__n32008, ys__n32010,
    ys__n32012, ys__n32014, ys__n32016, ys__n32018, ys__n32022, ys__n32023,
    ys__n32024, ys__n32025, ys__n32026, ys__n32027, ys__n32028, ys__n32029,
    ys__n32030, ys__n32031, ys__n32032, ys__n32033, ys__n32034, ys__n32035,
    ys__n32036, ys__n32037, ys__n32038, ys__n32039, ys__n32040, ys__n32041,
    ys__n32042, ys__n32043, ys__n32044, ys__n32045, ys__n32046, ys__n32047,
    ys__n32048, ys__n32049, ys__n32050, ys__n32051, ys__n32052, ys__n32053,
    ys__n32054, ys__n32055, ys__n32056, ys__n32057, ys__n32058, ys__n32059,
    ys__n32060, ys__n32061, ys__n32062, ys__n32063, ys__n32064, ys__n32065,
    ys__n32066, ys__n32067, ys__n32068, ys__n32069, ys__n32070, ys__n32071,
    ys__n32072, ys__n32073, ys__n32074, ys__n32075, ys__n32076, ys__n32077,
    ys__n32078, ys__n32079, ys__n32080, ys__n32081, ys__n32082, ys__n32083,
    ys__n32084, ys__n32085, ys__n32086, ys__n32087, ys__n32088, ys__n32124,
    ys__n32125, ys__n32126, ys__n32127, ys__n32128, ys__n32129, ys__n32130,
    ys__n32131, ys__n32132, ys__n32133, ys__n32134, ys__n32135, ys__n32136,
    ys__n32137, ys__n32138, ys__n32139, ys__n32140, ys__n32141, ys__n32142,
    ys__n32143, ys__n32144, ys__n32145, ys__n32146, ys__n32147, ys__n32148,
    ys__n32149, ys__n32150, ys__n32151, ys__n32152, ys__n32153, ys__n32154,
    ys__n32155, ys__n32158, ys__n32159, ys__n32160, ys__n32161, ys__n32162,
    ys__n32163, ys__n32164, ys__n32165, ys__n32166, ys__n32167, ys__n32168,
    ys__n32169, ys__n32170, ys__n32171, ys__n32172, ys__n32173, ys__n32174,
    ys__n32175, ys__n32176, ys__n32177, ys__n32178, ys__n32179, ys__n32180,
    ys__n32181, ys__n32182, ys__n32183, ys__n32184, ys__n32185, ys__n32186,
    ys__n32187, ys__n32188, ys__n32189, ys__n32190, ys__n32191, ys__n32192,
    ys__n32193, ys__n32194, ys__n32195, ys__n32196, ys__n32197, ys__n32198,
    ys__n32199, ys__n32200, ys__n32201, ys__n32202, ys__n32203, ys__n32204,
    ys__n32205, ys__n32206, ys__n32207, ys__n32208, ys__n32209, ys__n32210,
    ys__n32211, ys__n32212, ys__n32213, ys__n32214, ys__n32215, ys__n32216,
    ys__n32217, ys__n32218, ys__n32219, ys__n32220, ys__n32221, ys__n32222,
    ys__n32223, ys__n32224, ys__n32225, ys__n32226, ys__n32227, ys__n32228,
    ys__n32229, ys__n32230, ys__n32231, ys__n32232, ys__n32233, ys__n32234,
    ys__n32235, ys__n32236, ys__n32237, ys__n32238, ys__n32239, ys__n32240,
    ys__n32241, ys__n32242, ys__n32243, ys__n32244, ys__n32245, ys__n32246,
    ys__n32247, ys__n32248, ys__n32249, ys__n32250, ys__n32251, ys__n32252,
    ys__n32253, ys__n32254, ys__n32255, ys__n32256, ys__n32257, ys__n32258,
    ys__n32259, ys__n32260, ys__n32261, ys__n32262, ys__n32263, ys__n32264,
    ys__n32265, ys__n32266, ys__n32267, ys__n32268, ys__n32269, ys__n32270,
    ys__n32271, ys__n32272, ys__n32273, ys__n32274, ys__n32275, ys__n32276,
    ys__n32277, ys__n32278, ys__n32279, ys__n32280, ys__n32281, ys__n32282,
    ys__n32283, ys__n32284, ys__n32285, ys__n32286, ys__n32287, ys__n32288,
    ys__n32289, ys__n32290, ys__n32291, ys__n32292, ys__n32293, ys__n32294,
    ys__n32295, ys__n32296, ys__n32297, ys__n32298, ys__n32299, ys__n32300,
    ys__n32301, ys__n32302, ys__n32303, ys__n32304, ys__n32305, ys__n32306,
    ys__n32307, ys__n32308, ys__n32309, ys__n32310, ys__n32311, ys__n32312,
    ys__n32313, ys__n32314, ys__n32315, ys__n32316, ys__n32317, ys__n32318,
    ys__n32319, ys__n32320, ys__n32321, ys__n32322, ys__n32323, ys__n32324,
    ys__n32325, ys__n32326, ys__n32327, ys__n32328, ys__n32329, ys__n32330,
    ys__n32331, ys__n32332, ys__n32333, ys__n32334, ys__n32335, ys__n32336,
    ys__n32337, ys__n32338, ys__n32339, ys__n32340, ys__n32341, ys__n32342,
    ys__n32343, ys__n32344, ys__n32345, ys__n32346, ys__n32347, ys__n32348,
    ys__n32349, ys__n32350, ys__n32351, ys__n32352, ys__n32353, ys__n32354,
    ys__n32355, ys__n32356, ys__n32357, ys__n32358, ys__n32359, ys__n32360,
    ys__n32361, ys__n32362, ys__n32363, ys__n32364, ys__n32365, ys__n32366,
    ys__n32367, ys__n32368, ys__n32369, ys__n32370, ys__n32371, ys__n32372,
    ys__n32373, ys__n32374, ys__n32375, ys__n32376, ys__n32377, ys__n32378,
    ys__n32379, ys__n32380, ys__n32381, ys__n32382, ys__n32383, ys__n32384,
    ys__n32385, ys__n32386, ys__n32387, ys__n32388, ys__n32389, ys__n32390,
    ys__n32391, ys__n32392, ys__n32393, ys__n32394, ys__n32395, ys__n32396,
    ys__n32397, ys__n32398, ys__n32399, ys__n32400, ys__n32401, ys__n32402,
    ys__n32403, ys__n32404, ys__n32405, ys__n32406, ys__n32407, ys__n32408,
    ys__n32409, ys__n32410, ys__n32411, ys__n32412, ys__n32413, ys__n32414,
    ys__n32415, ys__n32416, ys__n32417, ys__n32418, ys__n32419, ys__n32420,
    ys__n32421, ys__n32422, ys__n32423, ys__n32424, ys__n32425, ys__n32426,
    ys__n32427, ys__n32428, ys__n32429, ys__n32430, ys__n32431, ys__n32432,
    ys__n32433, ys__n32434, ys__n32435, ys__n32436, ys__n32437, ys__n32438,
    ys__n32439, ys__n32440, ys__n32441, ys__n32442, ys__n32443, ys__n32444,
    ys__n32445, ys__n32446, ys__n32447, ys__n32448, ys__n32449, ys__n32450,
    ys__n32451, ys__n32452, ys__n32453, ys__n32454, ys__n32455, ys__n32456,
    ys__n32457, ys__n32458, ys__n32459, ys__n32460, ys__n32461, ys__n32462,
    ys__n32463, ys__n32464, ys__n32465, ys__n32466, ys__n32467, ys__n32468,
    ys__n32469, ys__n32470, ys__n32471, ys__n32472, ys__n32473, ys__n32474,
    ys__n32475, ys__n32476, ys__n32477, ys__n32478, ys__n32479, ys__n32480,
    ys__n32481, ys__n32482, ys__n32483, ys__n32484, ys__n32485, ys__n32486,
    ys__n32487, ys__n32488, ys__n32489, ys__n32490, ys__n32491, ys__n32492,
    ys__n32493, ys__n32494, ys__n32495, ys__n32496, ys__n32497, ys__n32498,
    ys__n32499, ys__n32500, ys__n32501, ys__n32502, ys__n32503, ys__n32504,
    ys__n32505, ys__n32506, ys__n32507, ys__n32508, ys__n32509, ys__n32510,
    ys__n32511, ys__n32512, ys__n32513, ys__n32514, ys__n32515, ys__n32516,
    ys__n32517, ys__n32518, ys__n32519, ys__n32520, ys__n32521, ys__n32522,
    ys__n32523, ys__n32524, ys__n32525, ys__n32526, ys__n32527, ys__n32528,
    ys__n32529, ys__n32530, ys__n32531, ys__n32532, ys__n32533, ys__n32534,
    ys__n32535, ys__n32536, ys__n32537, ys__n32538, ys__n32539, ys__n32540,
    ys__n32541, ys__n32542, ys__n32543, ys__n32544, ys__n32545, ys__n32546,
    ys__n32547, ys__n32548, ys__n32549, ys__n32550, ys__n32551, ys__n32552,
    ys__n32553, ys__n32554, ys__n32555, ys__n32556, ys__n32557, ys__n32558,
    ys__n32559, ys__n32560, ys__n32561, ys__n32562, ys__n32563, ys__n32564,
    ys__n32565, ys__n32566, ys__n32567, ys__n32568, ys__n32569, ys__n32570,
    ys__n32571, ys__n32572, ys__n32573, ys__n32574, ys__n32575, ys__n32576,
    ys__n32577, ys__n32578, ys__n32579, ys__n32580, ys__n32581, ys__n32582,
    ys__n32583, ys__n32584, ys__n32585, ys__n32586, ys__n32587, ys__n32588,
    ys__n32589, ys__n32590, ys__n32591, ys__n32592, ys__n32593, ys__n32594,
    ys__n32595, ys__n32596, ys__n32597, ys__n32598, ys__n32599, ys__n32600,
    ys__n32601, ys__n32602, ys__n32603, ys__n32604, ys__n32605, ys__n32606,
    ys__n32607, ys__n32608, ys__n32609, ys__n32610, ys__n32611, ys__n32612,
    ys__n32613, ys__n32614, ys__n32615, ys__n32616, ys__n32617, ys__n32618,
    ys__n32619, ys__n32620, ys__n32621, ys__n32622, ys__n32623, ys__n32624,
    ys__n32625, ys__n32626, ys__n32627, ys__n32628, ys__n32629, ys__n32630,
    ys__n32631, ys__n32632, ys__n32633, ys__n32634, ys__n32635, ys__n32636,
    ys__n32637, ys__n32638, ys__n32639, ys__n32640, ys__n32641, ys__n32642,
    ys__n32643, ys__n32644, ys__n32645, ys__n32646, ys__n32647, ys__n32648,
    ys__n32649, ys__n32650, ys__n32651, ys__n32652, ys__n32653, ys__n32654,
    ys__n32655, ys__n32656, ys__n32657, ys__n32658, ys__n32659, ys__n32660,
    ys__n32661, ys__n32662, ys__n32663, ys__n32664, ys__n32665, ys__n32666,
    ys__n32667, ys__n32668, ys__n32669, ys__n32670, ys__n32671, ys__n32672,
    ys__n32673, ys__n32674, ys__n32675, ys__n32676, ys__n32677, ys__n32678,
    ys__n32679, ys__n32680, ys__n32681, ys__n32682, ys__n32683, ys__n32684,
    ys__n32685, ys__n32686, ys__n32687, ys__n32688, ys__n32689, ys__n32690,
    ys__n32691, ys__n32692, ys__n32693, ys__n32694, ys__n32695, ys__n32696,
    ys__n32697, ys__n32698, ys__n32699, ys__n32700, ys__n32701, ys__n32702,
    ys__n32703, ys__n32704, ys__n32705, ys__n32706, ys__n32707, ys__n32708,
    ys__n32709, ys__n32710, ys__n32711, ys__n32712, ys__n32713, ys__n32714,
    ys__n32715, ys__n32716, ys__n32717, ys__n32718, ys__n32719, ys__n32720,
    ys__n32721, ys__n32722, ys__n32723, ys__n32724, ys__n32725, ys__n32726,
    ys__n32727, ys__n32728, ys__n32729, ys__n32730, ys__n32731, ys__n32732,
    ys__n32733, ys__n32734, ys__n32735, ys__n32736, ys__n32737, ys__n32738,
    ys__n32739, ys__n32740, ys__n32741, ys__n32742, ys__n32743, ys__n32744,
    ys__n32745, ys__n32746, ys__n32747, ys__n32748, ys__n32749, ys__n32750,
    ys__n32751, ys__n32752, ys__n32753, ys__n32754, ys__n32755, ys__n32756,
    ys__n32757, ys__n32758, ys__n32759, ys__n32760, ys__n32761, ys__n32762,
    ys__n32763, ys__n32764, ys__n32765, ys__n32766, ys__n32767, ys__n32768,
    ys__n32769, ys__n32770, ys__n32771, ys__n32772, ys__n32773, ys__n32774,
    ys__n32775, ys__n32776, ys__n32777, ys__n32778, ys__n32779, ys__n32780,
    ys__n32781, ys__n32782, ys__n32783, ys__n32784, ys__n32785, ys__n32786,
    ys__n32787, ys__n32788, ys__n32789, ys__n32790, ys__n32791, ys__n32792,
    ys__n32793, ys__n32794, ys__n32795, ys__n32796, ys__n32797, ys__n32798,
    ys__n32799, ys__n32800, ys__n32801, ys__n32802, ys__n32803, ys__n32804,
    ys__n32805, ys__n32806, ys__n32807, ys__n32808, ys__n32809, ys__n32810,
    ys__n32811, ys__n32812, ys__n32813, ys__n32814, ys__n32815, ys__n32816,
    ys__n32817, ys__n32818, ys__n32819, ys__n32820, ys__n32821, ys__n32822,
    ys__n32823, ys__n32824, ys__n32825, ys__n32826, ys__n32827, ys__n32828,
    ys__n32829, ys__n32830, ys__n32831, ys__n32832, ys__n32833, ys__n32834,
    ys__n32835, ys__n32836, ys__n32837, ys__n32838, ys__n32839, ys__n32840,
    ys__n32841, ys__n32842, ys__n32843, ys__n32844, ys__n32845, ys__n32846,
    ys__n32847, ys__n32848, ys__n32849, ys__n32850, ys__n32851, ys__n32852,
    ys__n32853, ys__n32854, ys__n32855, ys__n32856, ys__n32857, ys__n32858,
    ys__n32859, ys__n32860, ys__n32861, ys__n32862, ys__n32863, ys__n32864,
    ys__n32865, ys__n32866, ys__n32867, ys__n32868, ys__n32869, ys__n32870,
    ys__n32871, ys__n32872, ys__n32873, ys__n32874, ys__n32875, ys__n32876,
    ys__n32877, ys__n32878, ys__n32879, ys__n32880, ys__n32881, ys__n32882,
    ys__n32883, ys__n32884, ys__n32885, ys__n32886, ys__n32887, ys__n32888,
    ys__n32889, ys__n32890, ys__n32891, ys__n32892, ys__n32893, ys__n32894,
    ys__n32895, ys__n32896, ys__n32897, ys__n32898, ys__n32899, ys__n32900,
    ys__n32901, ys__n32902, ys__n32903, ys__n32904, ys__n32905, ys__n32906,
    ys__n32907, ys__n32908, ys__n32909, ys__n32910, ys__n32911, ys__n32912,
    ys__n32913, ys__n32914, ys__n32915, ys__n32916, ys__n32917, ys__n32918,
    ys__n32919, ys__n32920, ys__n32921, ys__n32922, ys__n32923, ys__n32924,
    ys__n32925, ys__n32926, ys__n32927, ys__n32928, ys__n32929, ys__n32930,
    ys__n32931, ys__n32932, ys__n32933, ys__n32934, ys__n32935, ys__n32936,
    ys__n32937, ys__n32938, ys__n32939, ys__n32940, ys__n32941, ys__n32942,
    ys__n32943, ys__n32944, ys__n32945, ys__n32946, ys__n32947, ys__n32948,
    ys__n32949, ys__n32950, ys__n32951, ys__n32952, ys__n32953, ys__n32954,
    ys__n32955, ys__n32956, ys__n32957, ys__n32958, ys__n32959, ys__n32960,
    ys__n32961, ys__n32962, ys__n32963, ys__n32964, ys__n32965, ys__n32966,
    ys__n32967, ys__n32968, ys__n32969, ys__n32970, ys__n32971, ys__n32972,
    ys__n32973, ys__n32974, ys__n32975, ys__n32976, ys__n32977, ys__n32978,
    ys__n32979, ys__n32980, ys__n32981, ys__n32982, ys__n32983, ys__n32984,
    ys__n32985, ys__n32986, ys__n32987, ys__n32988, ys__n32989, ys__n32990,
    ys__n32991, ys__n32992, ys__n32993, ys__n32994, ys__n32995, ys__n32996,
    ys__n32997, ys__n32998, ys__n33007, ys__n33008, ys__n33009, ys__n33014,
    ys__n33015, ys__n33016, ys__n33017, ys__n33018, ys__n33019, ys__n33020,
    ys__n33021, ys__n33022, ys__n33023, ys__n33024, ys__n33025, ys__n33026,
    ys__n33027, ys__n33028, ys__n33029, ys__n33030, ys__n33031, ys__n33032,
    ys__n33033, ys__n33034, ys__n33035, ys__n33036, ys__n33037, ys__n33038,
    ys__n33039, ys__n33040, ys__n33041, ys__n33042, ys__n33043, ys__n33044,
    ys__n33045, ys__n33046, ys__n33047, ys__n33048, ys__n33049, ys__n33050,
    ys__n33051, ys__n33052, ys__n33053, ys__n33054, ys__n33055, ys__n33056,
    ys__n33058, ys__n33059, ys__n33060, ys__n33061, ys__n33062, ys__n33063,
    ys__n33064, ys__n33065, ys__n33066, ys__n33067, ys__n33068, ys__n33069,
    ys__n33070, ys__n33071, ys__n33072, ys__n33073, ys__n33074, ys__n33075,
    ys__n33076, ys__n33077, ys__n33078, ys__n33079, ys__n33080, ys__n33081,
    ys__n33082, ys__n33083, ys__n33084, ys__n33085, ys__n33086, ys__n33087,
    ys__n33088, ys__n33089, ys__n33090, ys__n33091, ys__n33092, ys__n33093,
    ys__n33094, ys__n33095, ys__n33096, ys__n33097, ys__n33098, ys__n33099,
    ys__n33100, ys__n33101, ys__n33102, ys__n33103, ys__n33104, ys__n33105,
    ys__n33106, ys__n33107, ys__n33108, ys__n33109, ys__n33110, ys__n33111,
    ys__n33178, ys__n33179, ys__n33180, ys__n33181, ys__n33182, ys__n33183,
    ys__n33184, ys__n33185, ys__n33186, ys__n33187, ys__n33188, ys__n33189,
    ys__n33190, ys__n33191, ys__n33192, ys__n33193, ys__n33194, ys__n33195,
    ys__n33196, ys__n33197, ys__n33198, ys__n33199, ys__n33200, ys__n33201,
    ys__n33202, ys__n33203, ys__n33204, ys__n33205, ys__n33206, ys__n33207,
    ys__n33208, ys__n33209, ys__n33211, ys__n33317, ys__n33324, ys__n33329,
    ys__n33331, ys__n33333, ys__n33335, ys__n33337, ys__n33339, ys__n33357,
    ys__n33366, ys__n33414, ys__n33420, ys__n33437, ys__n33438, ys__n33439,
    ys__n33453, ys__n33454, ys__n33455, ys__n33456, ys__n33457, ys__n33513,
    ys__n33514, ys__n33515, ys__n33521, ys__n33535, ys__n34952, ys__n34953,
    ys__n34962, ys__n35052, ys__n35144, ys__n35146, ys__n35148, ys__n35150,
    ys__n35152, ys__n35154, ys__n35156, ys__n35158, ys__n35160, ys__n35162,
    ys__n35164, ys__n35166, ys__n35168, ys__n35170, ys__n35172, ys__n35174,
    ys__n35176, ys__n35178, ys__n35180, ys__n35182, ys__n35184, ys__n35186,
    ys__n35188, ys__n35190, ys__n35192, ys__n35194, ys__n35196, ys__n35198,
    ys__n35200, ys__n35202, ys__n35204, ys__n35206, ys__n35402, ys__n35404,
    ys__n35406, ys__n35408, ys__n35410, ys__n35412, ys__n35425, ys__n35705,
    ys__n35706, ys__n35708, ys__n35710, ys__n35712, ys__n35714, ys__n35716,
    ys__n37676, ys__n37687, ys__n37695, ys__n37697, ys__n37699, ys__n37702,
    ys__n37703, ys__n37707, ys__n37714, ys__n37731, ys__n37732, ys__n37733,
    ys__n37738, ys__n37739, ys__n37741, ys__n37742, ys__n38180, ys__n38182,
    ys__n38184, ys__n38185, ys__n38186, ys__n38188, ys__n38191, ys__n38205,
    ys__n38207, ys__n38209, ys__n38211, ys__n38213, ys__n38214, ys__n38216,
    ys__n38218, ys__n38222, ys__n38224, ys__n38246, ys__n38247, ys__n38248,
    ys__n38250, ys__n38252, ys__n38263, ys__n38266, ys__n38281, ys__n38285,
    ys__n38287, ys__n38289, ys__n38292, ys__n38294, ys__n38296, ys__n38303,
    ys__n38325, ys__n38326, ys__n38327, ys__n38328, ys__n38330, ys__n38331,
    ys__n38332, ys__n38334, ys__n38336, ys__n38337, ys__n38338, ys__n38339,
    ys__n38340, ys__n38341, ys__n38342, ys__n38343, ys__n38344, ys__n38345,
    ys__n38347, ys__n38349, ys__n38351, ys__n38352, ys__n38353, ys__n38354,
    ys__n38355, ys__n38356, ys__n38357, ys__n38359, ys__n38360, ys__n38362,
    ys__n38364, ys__n38365, ys__n38366, ys__n38367, ys__n38368, ys__n38369,
    ys__n38370, ys__n38371, ys__n38372, ys__n38373, ys__n38374, ys__n38375,
    ys__n38377, ys__n38379, ys__n38381, ys__n38383, ys__n38385, ys__n38387,
    ys__n38388, ys__n38389, ys__n38390, ys__n38391, ys__n38392, ys__n38393,
    ys__n38394, ys__n38396, ys__n38397, ys__n38417, ys__n38453, ys__n38456,
    ys__n38508, ys__n38509, ys__n38510, ys__n38515, ys__n38518, ys__n38520,
    ys__n38521, ys__n38523, ys__n38525, ys__n38552, ys__n38555, ys__n38556,
    ys__n38563, ys__n38566, ys__n38615, ys__n38623, ys__n38628, ys__n38633,
    ys__n38650, ys__n38662, ys__n38668, ys__n38669, ys__n38672, ys__n38674,
    ys__n38677, ys__n38689, ys__n38742, ys__n38768, ys__n38795, ys__n38799,
    ys__n38801, ys__n38884, ys__n38886, ys__n38887, ys__n38900, ys__n38912,
    ys__n38913, ys__n38914, ys__n38915, ys__n38917, ys__n38923, ys__n38925,
    ys__n38930, ys__n39392, ys__n39393, ys__n39395, ys__n39396, ys__n39397,
    ys__n39398, ys__n39399, ys__n39400, ys__n39401, ys__n39402, ys__n39403,
    ys__n39404, ys__n39405, ys__n39406, ys__n39407, ys__n39408, ys__n39409,
    ys__n39410, ys__n39411, ys__n39412, ys__n39413, ys__n39414, ys__n39415,
    ys__n39416, ys__n39417, ys__n39418, ys__n40052, ys__n42129, ys__n42153,
    ys__n42189, ys__n42194, ys__n42229, ys__n42234, ys__n42270, ys__n42275,
    ys__n42311, ys__n42316, ys__n42352, ys__n42357, ys__n42393, ys__n42398,
    ys__n42434, ys__n42439, ys__n42488, ys__n42493, ys__n42541, ys__n42546,
    ys__n42594, ys__n42599, ys__n42647, ys__n42652, ys__n42701, ys__n42706,
    ys__n42755, ys__n42760, ys__n42809, ys__n42814, ys__n42863, ys__n42868,
    ys__n42917, ys__n42922, ys__n42971, ys__n42976, ys__n43025, ys__n43030,
    ys__n43079, ys__n43084, ys__n43133, ys__n43138, ys__n43187, ys__n43192,
    ys__n43241, ys__n43246, ys__n43295, ys__n43300, ys__n43349, ys__n43354,
    ys__n43403, ys__n43408, ys__n43457, ys__n43462, ys__n43511, ys__n43516,
    ys__n43565, ys__n43570, ys__n43619, ys__n43624, ys__n43673, ys__n43678,
    ys__n43727, ys__n43732, ys__n43781, ys__n43786, ys__n43835, ys__n43840,
    ys__n43889, ys__n43894, ys__n43932, ys__n43937, ys__n43975, ys__n43980,
    ys__n44018, ys__n44023, ys__n44048, ys__n44053, ys__n44089, ys__n44094,
    ys__n44119, ys__n44122, ys__n44136, ys__n44139, ys__n44155, ys__n44160,
    ys__n44183, ys__n44186, ys__n44189, ys__n44192, ys__n44195, ys__n44198,
    ys__n44205, ys__n44213, ys__n44216, ys__n44219, ys__n44836, ys__n44838,
    ys__n44841, ys__n44843, ys__n44844, ys__n44845, ys__n44846, ys__n44848,
    ys__n44850, ys__n44851, ys__n44852, ys__n44853, ys__n44854, ys__n44855,
    ys__n44858, ys__n44948, ys__n44949, ys__n44950, ys__n44952, ys__n44953,
    ys__n44954, ys__n44955, ys__n44956, ys__n44957, ys__n44958, ys__n44959,
    ys__n44960, ys__n44961, ys__n44962, ys__n44963, ys__n44964, ys__n44965,
    ys__n44966, ys__n44967, ys__n44968, ys__n44969, ys__n44970, ys__n44971,
    ys__n44972, ys__n44973, ys__n44974, ys__n44975, ys__n44976, ys__n44977,
    ys__n44978, ys__n44979, ys__n44980, ys__n44981, ys__n44982, ys__n44983,
    ys__n44985, ys__n44987, ys__n46131, ys__n46133, ys__n46135, ys__n46137,
    ys__n46143, ys__n46146, ys__n46154, ys__n46155, ys__n46158, ys__n46159,
    ys__n46162, ys__n46163, ys__n46172, ys__n46173, ys__n46176, ys__n46179,
    ys__n46188, ys__n46189, ys__n46192, ys__n46195, ys__n46204, ys__n46205,
    ys__n46208, ys__n46211, ys__n46220, ys__n46221, ys__n46224, ys__n46227,
    ys__n46233, ys__n46234, ys__n48339, ys__n48340, ys__n48341, ys__n48342,
    ys__n48343, ys__n48344, ys__n48348, ys__n48349, ys__n48350, ys__n48351,
    ys__n48352, ys__n48353, ys__n48354, ys__n48355, ys__n48356, ys__n48357,
    ys__n48358, ys__n48359, ys__n48360, ys__n48361, ys__n48362;
  wire new_new_n98__, new_new_n99__, new_new_n101__, new_new_n102__,
    new_new_n104__, new_new_n105__, new_new_n107__, new_new_n108__,
    new_new_n110__, new_new_n111__, new_new_n113__, new_new_n114__,
    new_new_n116__, new_new_n117__, new_new_n119__, new_new_n120__,
    new_new_n122__, new_new_n123__, new_new_n125__, new_new_n126__,
    new_new_n128__, new_new_n129__, new_new_n131__, new_new_n132__,
    new_new_n134__, new_new_n135__, new_new_n137__, new_new_n138__,
    new_new_n140__, new_new_n141__, new_new_n143__, new_new_n144__,
    new_new_n146__, new_new_n147__, new_new_n149__, new_new_n150__,
    new_new_n152__, new_new_n153__, new_new_n155__, new_new_n156__,
    new_new_n158__, new_new_n159__, new_new_n161__, new_new_n162__,
    new_new_n164__, new_new_n165__, new_new_n167__, new_new_n168__,
    new_new_n170__, new_new_n171__, new_new_n173__, new_new_n174__,
    new_new_n176__, new_new_n177__, new_new_n179__, new_new_n180__,
    new_new_n182__, new_new_n183__, new_new_n185__, new_new_n186__,
    new_new_n188__, new_new_n189__, new_new_n191__, new_new_n192__,
    new_new_n98_5_, new_new_n99_5_, new_new_n101_5_, new_new_n102_5_,
    new_new_n104_5_, new_new_n105_5_, new_new_n107_5_, new_new_n108_5_,
    new_new_n110_5_, new_new_n111_5_, new_new_n113_5_, new_new_n114_5_,
    new_new_n116_5_, new_new_n117_5_, new_new_n119_5_, new_new_n120_5_,
    new_new_n122_5_, new_new_n123_5_, new_new_n125_5_, new_new_n126_5_,
    new_new_n128_5_, new_new_n129_5_, new_new_n131_5_, new_new_n132_5_,
    new_new_n134_5_, new_new_n135_5_, new_new_n137_5_, new_new_n138_5_,
    new_new_n140_5_, new_new_n141_5_, new_new_n143_5_, new_new_n144_5_,
    new_new_n146_5_, new_new_n147_5_, new_new_n149_5_, new_new_n150_5_,
    new_new_n152_5_, new_new_n153_5_, new_new_n155_5_, new_new_n156_5_,
    new_new_n158_5_, new_new_n159_5_, new_new_n161_5_, new_new_n162_5_,
    new_new_n164_5_, new_new_n165_5_, new_new_n167_5_, new_new_n168_5_,
    new_new_n170_5_, new_new_n171_5_, new_new_n173_5_, new_new_n174_5_,
    new_new_n176_5_, new_new_n177_5_, new_new_n179_5_, new_new_n180_5_,
    new_new_n182_5_, new_new_n183_5_, new_new_n185_5_, new_new_n186_5_,
    new_new_n188_5_, new_new_n189_5_, new_new_n191_5_, new_new_n192_5_,
    new_new_n10398__, new_new_n10399__, new_new_n10400__, new_new_n10401__,
    new_new_n10402__, new_new_n10403__, new_new_n10404__, new_new_n10405__,
    new_new_n10406__, new_new_n10407__, new_new_n10408__, new_new_n10409__,
    new_new_n10410__, new_new_n10411__, new_new_n10412__, new_new_n10413__,
    new_new_n10414__, new_new_n10415__, new_new_n10416__, new_new_n10417__,
    new_new_n10418__, new_new_n10419__, new_new_n10420__, new_new_n10421__,
    new_new_n10422__, new_new_n10423__, new_new_n10424__, new_new_n10425__,
    new_new_n10426__, new_new_n10427__, new_new_n10428__, new_new_n10429__,
    new_new_n10430__, new_new_n10431__, new_new_n10432__, new_new_n10433__,
    new_new_n10434__, new_new_n10435__, new_new_n10436__, new_new_n10437__,
    new_new_n10438__, new_new_n10439__, new_new_n10440__, new_new_n10441__,
    new_new_n10442__, new_new_n10443__, new_new_n10444__, new_new_n10445__,
    new_new_n10446__, new_new_n10447__, new_new_n10448__, new_new_n10449__,
    new_new_n10450__, new_new_n10451__, new_new_n10452__, new_new_n10453__,
    new_new_n10454__, new_new_n10455__, new_new_n10456__, new_new_n10457__,
    new_new_n10458__, new_new_n10459__, new_new_n10460__, new_new_n10461__,
    new_new_n10462__, new_new_n10463__, new_new_n10464__, new_new_n10465__,
    new_new_n10466__, new_new_n10467__, new_new_n10468__, new_new_n10469__,
    new_new_n10470__, new_new_n10471__, new_new_n10472__, new_new_n10473__,
    new_new_n10474__, new_new_n10475__, new_new_n10476__, new_new_n10477__,
    new_new_n10478__, new_new_n10479__, new_new_n10480__, new_new_n10481__,
    new_new_n10482__, new_new_n10483__, new_new_n10484__, new_new_n10485__,
    new_new_n10486__, new_new_n10487__, new_new_n10488__, new_new_n10489__,
    new_new_n10490__, new_new_n10491__, new_new_n10492__, new_new_n10493__,
    new_new_n10494__, new_new_n10495__, new_new_n10496__, new_new_n10497__,
    new_new_n10498__, new_new_n10499__, new_new_n10500__, new_new_n10501__,
    new_new_n10502__, new_new_n10503__, new_new_n10504__, new_new_n10505__,
    new_new_n10506__, new_new_n10507__, new_new_n10508__, new_new_n10509__,
    new_new_n10510__, new_new_n10511__, new_new_n10512__, new_new_n10513__,
    new_new_n10514__, new_new_n10515__, new_new_n10516__, new_new_n10517__,
    new_new_n10518__, new_new_n10519__, new_new_n10520__, new_new_n10521__,
    new_new_n10522__, new_new_n10523__, new_new_n10524__, new_new_n10525__,
    new_new_n10526__, new_new_n10527__, new_new_n10528__, new_new_n10529__,
    new_new_n10530__, new_new_n10531__, new_new_n10532__, new_new_n10533__,
    new_new_n10534__, new_new_n10535__, new_new_n10536__, new_new_n10537__,
    new_new_n10538__, new_new_n10539__, new_new_n10540__, new_new_n10541__,
    new_new_n10542__, new_new_n10543__, new_new_n10544__, new_new_n10545__,
    new_new_n10546__, new_new_n10547__, new_new_n10548__, new_new_n10549__,
    new_new_n10550__, new_new_n10551__, new_new_n10552__, new_new_n10553__,
    new_new_n10554__, new_new_n10555__, new_new_n10556__, new_new_n10557__,
    new_new_n10558__, new_new_n10559__, new_new_n10560__, new_new_n10561__,
    new_new_n10562__, new_new_n10563__, new_new_n10564__, new_new_n10565__,
    new_new_n10566__, new_new_n10567__, new_new_n10568__, new_new_n10569__,
    new_new_n10570__, new_new_n10571__, new_new_n10572__, new_new_n10573__,
    new_new_n10574__, new_new_n10575__, new_new_n10576__, new_new_n10577__,
    new_new_n10578__, new_new_n10579__, new_new_n10580__, new_new_n10581__,
    new_new_n10582__, new_new_n10583__, new_new_n10584__, new_new_n10585__,
    new_new_n10586__, new_new_n10587__, new_new_n10588__, new_new_n10589__,
    new_new_n10590__, new_new_n10591__, new_new_n10592__, new_new_n10593__,
    new_new_n10594__, new_new_n10595__, new_new_n10596__, new_new_n10597__,
    new_new_n10598__, new_new_n10599__, new_new_n10600__, new_new_n10601__,
    new_new_n10602__, new_new_n10603__, new_new_n10604__, new_new_n10605__,
    new_new_n10607__, new_new_n10608__, new_new_n10609__, new_new_n10610__,
    new_new_n10611__, new_new_n10612__, new_new_n10613__, new_new_n10615__,
    new_new_n10616__, new_new_n10618__, new_new_n10619__, new_new_n10620__,
    new_new_n10621__, new_new_n10622__, new_new_n10624__, new_new_n10625__,
    new_new_n10626__, new_new_n10627__, new_new_n10628__, new_new_n10629__,
    new_new_n10630__, new_new_n10631__, new_new_n10632__, new_new_n10633__,
    new_new_n10634__, new_new_n10635__, new_new_n10636__, new_new_n10637__,
    new_new_n10638__, new_new_n10639__, new_new_n10640__, new_new_n10641__,
    new_new_n10642__, new_new_n10643__, new_new_n10644__, new_new_n10645__,
    new_new_n10646__, new_new_n10647__, new_new_n10648__, new_new_n10649__,
    new_new_n10650__, new_new_n10651__, new_new_n10652__, new_new_n10653__,
    new_new_n10654__, new_new_n10655__, new_new_n10656__, new_new_n10657__,
    new_new_n10658__, new_new_n10659__, new_new_n10660__, new_new_n10661__,
    new_new_n10662__, new_new_n10663__, new_new_n10664__, new_new_n10665__,
    new_new_n10666__, new_new_n10667__, new_new_n10668__, new_new_n10669__,
    new_new_n10670__, new_new_n10671__, new_new_n10672__, new_new_n10673__,
    new_new_n10674__, new_new_n10675__, new_new_n10676__, new_new_n10677__,
    new_new_n10678__, new_new_n10679__, new_new_n10680__, new_new_n10681__,
    new_new_n10682__, new_new_n10683__, new_new_n10684__, new_new_n10685__,
    new_new_n10686__, new_new_n10687__, new_new_n10688__, new_new_n10689__,
    new_new_n10690__, new_new_n10691__, new_new_n10692__, new_new_n10693__,
    new_new_n10694__, new_new_n10695__, new_new_n10696__, new_new_n10697__,
    new_new_n10698__, new_new_n10699__, new_new_n10700__, new_new_n10701__,
    new_new_n10702__, new_new_n10703__, new_new_n10704__, new_new_n10705__,
    new_new_n10706__, new_new_n10707__, new_new_n10708__, new_new_n10709__,
    new_new_n10710__, new_new_n10711__, new_new_n10712__, new_new_n10713__,
    new_new_n10714__, new_new_n10715__, new_new_n10716__, new_new_n10717__,
    new_new_n10718__, new_new_n10719__, new_new_n10720__, new_new_n10721__,
    new_new_n10722__, new_new_n10723__, new_new_n10724__, new_new_n10725__,
    new_new_n10726__, new_new_n10727__, new_new_n10728__, new_new_n10729__,
    new_new_n10730__, new_new_n10731__, new_new_n10732__, new_new_n10733__,
    new_new_n10734__, new_new_n10735__, new_new_n10736__, new_new_n10737__,
    new_new_n10738__, new_new_n10739__, new_new_n10740__, new_new_n10741__,
    new_new_n10742__, new_new_n10743__, new_new_n10744__, new_new_n10745__,
    new_new_n10746__, new_new_n10747__, new_new_n10748__, new_new_n10749__,
    new_new_n10750__, new_new_n10751__, new_new_n10752__, new_new_n10753__,
    new_new_n10754__, new_new_n10755__, new_new_n10756__, new_new_n10757__,
    new_new_n10758__, new_new_n10759__, new_new_n10760__, new_new_n10761__,
    new_new_n10762__, new_new_n10763__, new_new_n10764__, new_new_n10765__,
    new_new_n10766__, new_new_n10767__, new_new_n10768__, new_new_n10769__,
    new_new_n10770__, new_new_n10771__, new_new_n10772__, new_new_n10773__,
    new_new_n10774__, new_new_n10775__, new_new_n10776__, new_new_n10777__,
    new_new_n10778__, new_new_n10779__, new_new_n10780__, new_new_n10781__,
    new_new_n10782__, new_new_n10783__, new_new_n10784__, new_new_n10785__,
    new_new_n10786__, new_new_n10787__, new_new_n10788__, new_new_n10789__,
    new_new_n10790__, new_new_n10791__, new_new_n10792__, new_new_n10793__,
    new_new_n10794__, new_new_n10795__, new_new_n10796__, new_new_n10797__,
    new_new_n10798__, new_new_n10799__, new_new_n10800__, new_new_n10801__,
    new_new_n10802__, new_new_n10803__, new_new_n10804__, new_new_n10805__,
    new_new_n10806__, new_new_n10807__, new_new_n10808__, new_new_n10809__,
    new_new_n10810__, new_new_n10811__, new_new_n10812__, new_new_n10813__,
    new_new_n10814__, new_new_n10815__, new_new_n10816__, new_new_n10817__,
    new_new_n10818__, new_new_n10819__, new_new_n10820__, new_new_n10821__,
    new_new_n10822__, new_new_n10823__, new_new_n10824__, new_new_n10825__,
    new_new_n10826__, new_new_n10827__, new_new_n10830__, new_new_n10831__,
    new_new_n10832__, new_new_n10834__, new_new_n10835__, new_new_n10836__,
    new_new_n10837__, new_new_n10838__, new_new_n10839__, new_new_n10840__,
    new_new_n10841__, new_new_n10842__, new_new_n10843__, new_new_n10845__,
    new_new_n10846__, new_new_n10847__, new_new_n10848__, new_new_n10849__,
    new_new_n10850__, new_new_n10851__, new_new_n10852__, new_new_n10853__,
    new_new_n10854__, new_new_n10855__, new_new_n10856__, new_new_n10858__,
    new_new_n10859__, new_new_n10860__, new_new_n10861__, new_new_n10862__,
    new_new_n10863__, new_new_n10864__, new_new_n10865__, new_new_n10866__,
    new_new_n10868__, new_new_n10869__, new_new_n10870__, new_new_n10871__,
    new_new_n10872__, new_new_n10874__, new_new_n10875__, new_new_n10876__,
    new_new_n10878__, new_new_n10879__, new_new_n10880__, new_new_n10881__,
    new_new_n10882__, new_new_n10883__, new_new_n10884__, new_new_n10885__,
    new_new_n10886__, new_new_n10887__, new_new_n10888__, new_new_n10890__,
    new_new_n10891__, new_new_n10892__, new_new_n10893__, new_new_n10894__,
    new_new_n10895__, new_new_n10896__, new_new_n10897__, new_new_n10898__,
    new_new_n10899__, new_new_n10900__, new_new_n10901__, new_new_n10902__,
    new_new_n10903__, new_new_n10904__, new_new_n10905__, new_new_n10906__,
    new_new_n10907__, new_new_n10908__, new_new_n10909__, new_new_n10911__,
    new_new_n10912__, new_new_n10913__, new_new_n10914__, new_new_n10915__,
    new_new_n10916__, new_new_n10917__, new_new_n10918__, new_new_n10919__,
    new_new_n10920__, new_new_n10921__, new_new_n10922__, new_new_n10923__,
    new_new_n10924__, new_new_n10925__, new_new_n10926__, new_new_n10927__,
    new_new_n10928__, new_new_n10929__, new_new_n10930__, new_new_n10931__,
    new_new_n10932__, new_new_n10933__, new_new_n10934__, new_new_n10935__,
    new_new_n10936__, new_new_n10937__, new_new_n10938__, new_new_n10939__,
    new_new_n10941__, new_new_n10942__, new_new_n10943__, new_new_n10944__,
    new_new_n10945__, new_new_n10947__, new_new_n10948__, new_new_n10949__,
    new_new_n10950__, new_new_n10951__, new_new_n10952__, new_new_n10953__,
    new_new_n10954__, new_new_n10955__, new_new_n10956__, new_new_n10957__,
    new_new_n10958__, new_new_n10959__, new_new_n10960__, new_new_n10961__,
    new_new_n10962__, new_new_n10963__, new_new_n10964__, new_new_n10965__,
    new_new_n10967__, new_new_n10970__, new_new_n10971__, new_new_n10972__,
    new_new_n10973__, new_new_n10974__, new_new_n10975__, new_new_n10976__,
    new_new_n10977__, new_new_n10978__, new_new_n10979__, new_new_n10980__,
    new_new_n10982__, new_new_n10983__, new_new_n10984__, new_new_n10986__,
    new_new_n10987__, new_new_n10988__, new_new_n10989__, new_new_n10990__,
    new_new_n10991__, new_new_n10992__, new_new_n10993__, new_new_n10994__,
    new_new_n10995__, new_new_n10996__, new_new_n10997__, new_new_n10998__,
    new_new_n10999__, new_new_n11000__, new_new_n11001__, new_new_n11002__,
    new_new_n11003__, new_new_n11004__, new_new_n11005__, new_new_n11006__,
    new_new_n11008__, new_new_n11009__, new_new_n11010__, new_new_n11011__,
    new_new_n11012__, new_new_n11013__, new_new_n11014__, new_new_n11015__,
    new_new_n11016__, new_new_n11017__, new_new_n11018__, new_new_n11019__,
    new_new_n11020__, new_new_n11021__, new_new_n11022__, new_new_n11023__,
    new_new_n11024__, new_new_n11025__, new_new_n11026__, new_new_n11028__,
    new_new_n11029__, new_new_n11030__, new_new_n11031__, new_new_n11032__,
    new_new_n11033__, new_new_n11034__, new_new_n11035__, new_new_n11036__,
    new_new_n11038__, new_new_n11039__, new_new_n11040__, new_new_n11041__,
    new_new_n11042__, new_new_n11043__, new_new_n11044__, new_new_n11045__,
    new_new_n11046__, new_new_n11047__, new_new_n11048__, new_new_n11049__,
    new_new_n11050__, new_new_n11051__, new_new_n11052__, new_new_n11053__,
    new_new_n11054__, new_new_n11055__, new_new_n11056__, new_new_n11057__,
    new_new_n11058__, new_new_n11059__, new_new_n11060__, new_new_n11061__,
    new_new_n11063__, new_new_n11064__, new_new_n11065__, new_new_n11066__,
    new_new_n11067__, new_new_n11068__, new_new_n11069__, new_new_n11070__,
    new_new_n11071__, new_new_n11072__, new_new_n11073__, new_new_n11074__,
    new_new_n11075__, new_new_n11076__, new_new_n11077__, new_new_n11078__,
    new_new_n11079__, new_new_n11080__, new_new_n11081__, new_new_n11082__,
    new_new_n11083__, new_new_n11084__, new_new_n11085__, new_new_n11086__,
    new_new_n11087__, new_new_n11088__, new_new_n11089__, new_new_n11090__,
    new_new_n11091__, new_new_n11092__, new_new_n11093__, new_new_n11094__,
    new_new_n11095__, new_new_n11096__, new_new_n11097__, new_new_n11098__,
    new_new_n11099__, new_new_n11100__, new_new_n11101__, new_new_n11102__,
    new_new_n11103__, new_new_n11104__, new_new_n11105__, new_new_n11106__,
    new_new_n11107__, new_new_n11108__, new_new_n11109__, new_new_n11111__,
    new_new_n11112__, new_new_n11114__, new_new_n11115__, new_new_n11116__,
    new_new_n11117__, new_new_n11119__, new_new_n11120__, new_new_n11121__,
    new_new_n11122__, new_new_n11124__, new_new_n11125__, new_new_n11126__,
    new_new_n11127__, new_new_n11128__, new_new_n11129__, new_new_n11130__,
    new_new_n11131__, new_new_n11132__, new_new_n11133__, new_new_n11134__,
    new_new_n11135__, new_new_n11137__, new_new_n11138__, new_new_n11140__,
    new_new_n11141__, new_new_n11142__, new_new_n11143__, new_new_n11144__,
    new_new_n11145__, new_new_n11146__, new_new_n11147__, new_new_n11148__,
    new_new_n11149__, new_new_n11150__, new_new_n11151__, new_new_n11152__,
    new_new_n11153__, new_new_n11154__, new_new_n11155__, new_new_n11157__,
    new_new_n11158__, new_new_n11159__, new_new_n11160__, new_new_n11161__,
    new_new_n11163__, new_new_n11164__, new_new_n11165__, new_new_n11166__,
    new_new_n11167__, new_new_n11168__, new_new_n11169__, new_new_n11170__,
    new_new_n11171__, new_new_n11172__, new_new_n11173__, new_new_n11174__,
    new_new_n11175__, new_new_n11176__, new_new_n11177__, new_new_n11178__,
    new_new_n11179__, new_new_n11180__, new_new_n11181__, new_new_n11182__,
    new_new_n11183__, new_new_n11184__, new_new_n11185__, new_new_n11186__,
    new_new_n11187__, new_new_n11188__, new_new_n11189__, new_new_n11190__,
    new_new_n11191__, new_new_n11192__, new_new_n11193__, new_new_n11194__,
    new_new_n11195__, new_new_n11196__, new_new_n11197__, new_new_n11198__,
    new_new_n11199__, new_new_n11200__, new_new_n11201__, new_new_n11202__,
    new_new_n11203__, new_new_n11204__, new_new_n11205__, new_new_n11206__,
    new_new_n11207__, new_new_n11208__, new_new_n11209__, new_new_n11210__,
    new_new_n11211__, new_new_n11212__, new_new_n11213__, new_new_n11214__,
    new_new_n11215__, new_new_n11216__, new_new_n11217__, new_new_n11218__,
    new_new_n11219__, new_new_n11220__, new_new_n11221__, new_new_n11222__,
    new_new_n11223__, new_new_n11224__, new_new_n11225__, new_new_n11226__,
    new_new_n11227__, new_new_n11228__, new_new_n11229__, new_new_n11230__,
    new_new_n11231__, new_new_n11232__, new_new_n11233__, new_new_n11234__,
    new_new_n11235__, new_new_n11236__, new_new_n11237__, new_new_n11238__,
    new_new_n11239__, new_new_n11240__, new_new_n11241__, new_new_n11242__,
    new_new_n11243__, new_new_n11244__, new_new_n11245__, new_new_n11246__,
    new_new_n11247__, new_new_n11248__, new_new_n11249__, new_new_n11250__,
    new_new_n11251__, new_new_n11252__, new_new_n11253__, new_new_n11254__,
    new_new_n11255__, new_new_n11256__, new_new_n11257__, new_new_n11258__,
    new_new_n11259__, new_new_n11260__, new_new_n11261__, new_new_n11262__,
    new_new_n11263__, new_new_n11264__, new_new_n11265__, new_new_n11266__,
    new_new_n11267__, new_new_n11268__, new_new_n11269__, new_new_n11270__,
    new_new_n11271__, new_new_n11272__, new_new_n11273__, new_new_n11274__,
    new_new_n11275__, new_new_n11276__, new_new_n11277__, new_new_n11278__,
    new_new_n11279__, new_new_n11280__, new_new_n11281__, new_new_n11282__,
    new_new_n11283__, new_new_n11284__, new_new_n11285__, new_new_n11286__,
    new_new_n11287__, new_new_n11288__, new_new_n11289__, new_new_n11290__,
    new_new_n11291__, new_new_n11292__, new_new_n11293__, new_new_n11294__,
    new_new_n11295__, new_new_n11296__, new_new_n11297__, new_new_n11298__,
    new_new_n11299__, new_new_n11300__, new_new_n11301__, new_new_n11302__,
    new_new_n11303__, new_new_n11304__, new_new_n11305__, new_new_n11306__,
    new_new_n11307__, new_new_n11308__, new_new_n11309__, new_new_n11311__,
    new_new_n11312__, new_new_n11313__, new_new_n11314__, new_new_n11315__,
    new_new_n11316__, new_new_n11317__, new_new_n11318__, new_new_n11319__,
    new_new_n11320__, new_new_n11321__, new_new_n11322__, new_new_n11323__,
    new_new_n11324__, new_new_n11325__, new_new_n11326__, new_new_n11327__,
    new_new_n11328__, new_new_n11329__, new_new_n11330__, new_new_n11331__,
    new_new_n11332__, new_new_n11333__, new_new_n11334__, new_new_n11335__,
    new_new_n11336__, new_new_n11337__, new_new_n11338__, new_new_n11339__,
    new_new_n11340__, new_new_n11341__, new_new_n11342__, new_new_n11343__,
    new_new_n11344__, new_new_n11345__, new_new_n11346__, new_new_n11347__,
    new_new_n11348__, new_new_n11349__, new_new_n11350__, new_new_n11351__,
    new_new_n11352__, new_new_n11353__, new_new_n11354__, new_new_n11355__,
    new_new_n11356__, new_new_n11357__, new_new_n11358__, new_new_n11359__,
    new_new_n11360__, new_new_n11361__, new_new_n11362__, new_new_n11363__,
    new_new_n11364__, new_new_n11365__, new_new_n11366__, new_new_n11367__,
    new_new_n11368__, new_new_n11369__, new_new_n11370__, new_new_n11371__,
    new_new_n11372__, new_new_n11373__, new_new_n11374__, new_new_n11375__,
    new_new_n11376__, new_new_n11377__, new_new_n11378__, new_new_n11379__,
    new_new_n11380__, new_new_n11381__, new_new_n11382__, new_new_n11383__,
    new_new_n11384__, new_new_n11385__, new_new_n11386__, new_new_n11387__,
    new_new_n11388__, new_new_n11389__, new_new_n11390__, new_new_n11391__,
    new_new_n11392__, new_new_n11393__, new_new_n11394__, new_new_n11395__,
    new_new_n11396__, new_new_n11397__, new_new_n11398__, new_new_n11399__,
    new_new_n11400__, new_new_n11401__, new_new_n11402__, new_new_n11403__,
    new_new_n11404__, new_new_n11405__, new_new_n11406__, new_new_n11407__,
    new_new_n11408__, new_new_n11409__, new_new_n11410__, new_new_n11411__,
    new_new_n11412__, new_new_n11413__, new_new_n11414__, new_new_n11415__,
    new_new_n11416__, new_new_n11417__, new_new_n11418__, new_new_n11419__,
    new_new_n11420__, new_new_n11421__, new_new_n11422__, new_new_n11423__,
    new_new_n11424__, new_new_n11425__, new_new_n11426__, new_new_n11427__,
    new_new_n11428__, new_new_n11429__, new_new_n11430__, new_new_n11431__,
    new_new_n11432__, new_new_n11433__, new_new_n11434__, new_new_n11435__,
    new_new_n11436__, new_new_n11437__, new_new_n11438__, new_new_n11439__,
    new_new_n11440__, new_new_n11441__, new_new_n11442__, new_new_n11443__,
    new_new_n11444__, new_new_n11445__, new_new_n11446__, new_new_n11447__,
    new_new_n11448__, new_new_n11449__, new_new_n11450__, new_new_n11451__,
    new_new_n11452__, new_new_n11453__, new_new_n11454__, new_new_n11455__,
    new_new_n11456__, new_new_n11457__, new_new_n11458__, new_new_n11459__,
    new_new_n11460__, new_new_n11461__, new_new_n11462__, new_new_n11463__,
    new_new_n11464__, new_new_n11465__, new_new_n11466__, new_new_n11467__,
    new_new_n11468__, new_new_n11469__, new_new_n11470__, new_new_n11471__,
    new_new_n11472__, new_new_n11473__, new_new_n11474__, new_new_n11475__,
    new_new_n11476__, new_new_n11477__, new_new_n11478__, new_new_n11479__,
    new_new_n11480__, new_new_n11481__, new_new_n11482__, new_new_n11483__,
    new_new_n11484__, new_new_n11485__, new_new_n11486__, new_new_n11487__,
    new_new_n11488__, new_new_n11489__, new_new_n11490__, new_new_n11491__,
    new_new_n11492__, new_new_n11493__, new_new_n11494__, new_new_n11495__,
    new_new_n11496__, new_new_n11497__, new_new_n11498__, new_new_n11499__,
    new_new_n11500__, new_new_n11501__, new_new_n11502__, new_new_n11503__,
    new_new_n11504__, new_new_n11505__, new_new_n11506__, new_new_n11507__,
    new_new_n11508__, new_new_n11509__, new_new_n11510__, new_new_n11511__,
    new_new_n11512__, new_new_n11513__, new_new_n11514__, new_new_n11515__,
    new_new_n11516__, new_new_n11517__, new_new_n11518__, new_new_n11519__,
    new_new_n11520__, new_new_n11521__, new_new_n11522__, new_new_n11523__,
    new_new_n11524__, new_new_n11525__, new_new_n11526__, new_new_n11527__,
    new_new_n11528__, new_new_n11529__, new_new_n11530__, new_new_n11531__,
    new_new_n11532__, new_new_n11533__, new_new_n11534__, new_new_n11535__,
    new_new_n11536__, new_new_n11537__, new_new_n11538__, new_new_n11539__,
    new_new_n11540__, new_new_n11541__, new_new_n11542__, new_new_n11543__,
    new_new_n11544__, new_new_n11545__, new_new_n11546__, new_new_n11547__,
    new_new_n11548__, new_new_n11549__, new_new_n11550__, new_new_n11551__,
    new_new_n11552__, new_new_n11553__, new_new_n11554__, new_new_n11555__,
    new_new_n11556__, new_new_n11557__, new_new_n11558__, new_new_n11559__,
    new_new_n11560__, new_new_n11561__, new_new_n11562__, new_new_n11563__,
    new_new_n11564__, new_new_n11565__, new_new_n11566__, new_new_n11567__,
    new_new_n11568__, new_new_n11569__, new_new_n11570__, new_new_n11571__,
    new_new_n11572__, new_new_n11573__, new_new_n11574__, new_new_n11575__,
    new_new_n11576__, new_new_n11577__, new_new_n11578__, new_new_n11579__,
    new_new_n11580__, new_new_n11581__, new_new_n11582__, new_new_n11583__,
    new_new_n11584__, new_new_n11585__, new_new_n11586__, new_new_n11587__,
    new_new_n11588__, new_new_n11589__, new_new_n11590__, new_new_n11591__,
    new_new_n11592__, new_new_n11593__, new_new_n11594__, new_new_n11595__,
    new_new_n11596__, new_new_n11597__, new_new_n11598__, new_new_n11599__,
    new_new_n11600__, new_new_n11601__, new_new_n11602__, new_new_n11603__,
    new_new_n11604__, new_new_n11605__, new_new_n11606__, new_new_n11607__,
    new_new_n11608__, new_new_n11609__, new_new_n11610__, new_new_n11611__,
    new_new_n11612__, new_new_n11613__, new_new_n11614__, new_new_n11615__,
    new_new_n11616__, new_new_n11617__, new_new_n11618__, new_new_n11619__,
    new_new_n11620__, new_new_n11621__, new_new_n11622__, new_new_n11623__,
    new_new_n11624__, new_new_n11625__, new_new_n11626__, new_new_n11627__,
    new_new_n11628__, new_new_n11629__, new_new_n11630__, new_new_n11631__,
    new_new_n11632__, new_new_n11633__, new_new_n11634__, new_new_n11635__,
    new_new_n11636__, new_new_n11637__, new_new_n11638__, new_new_n11639__,
    new_new_n11640__, new_new_n11641__, new_new_n11642__, new_new_n11643__,
    new_new_n11644__, new_new_n11645__, new_new_n11646__, new_new_n11647__,
    new_new_n11648__, new_new_n11649__, new_new_n11650__, new_new_n11651__,
    new_new_n11653__, new_new_n11654__, new_new_n11655__, new_new_n11656__,
    new_new_n11657__, new_new_n11658__, new_new_n11659__, new_new_n11660__,
    new_new_n11661__, new_new_n11662__, new_new_n11663__, new_new_n11664__,
    new_new_n11665__, new_new_n11666__, new_new_n11667__, new_new_n11668__,
    new_new_n11669__, new_new_n11671__, new_new_n11672__, new_new_n11673__,
    new_new_n11674__, new_new_n11675__, new_new_n11676__, new_new_n11677__,
    new_new_n11678__, new_new_n11679__, new_new_n11680__, new_new_n11681__,
    new_new_n11682__, new_new_n11683__, new_new_n11684__, new_new_n11685__,
    new_new_n11686__, new_new_n11687__, new_new_n11688__, new_new_n11689__,
    new_new_n11690__, new_new_n11691__, new_new_n11692__, new_new_n11693__,
    new_new_n11694__, new_new_n11695__, new_new_n11696__, new_new_n11697__,
    new_new_n11698__, new_new_n11699__, new_new_n11700__, new_new_n11701__,
    new_new_n11702__, new_new_n11703__, new_new_n11704__, new_new_n11705__,
    new_new_n11706__, new_new_n11708__, new_new_n11709__, new_new_n11710__,
    new_new_n11711__, new_new_n11712__, new_new_n11713__, new_new_n11714__,
    new_new_n11715__, new_new_n11716__, new_new_n11717__, new_new_n11719__,
    new_new_n11720__, new_new_n11721__, new_new_n11722__, new_new_n11723__,
    new_new_n11724__, new_new_n11725__, new_new_n11726__, new_new_n11727__,
    new_new_n11728__, new_new_n11729__, new_new_n11730__, new_new_n11731__,
    new_new_n11732__, new_new_n11733__, new_new_n11735__, new_new_n11736__,
    new_new_n11737__, new_new_n11739__, new_new_n11740__, new_new_n11741__,
    new_new_n11743__, new_new_n11745__, new_new_n11746__, new_new_n11747__,
    new_new_n11748__, new_new_n11750__, new_new_n11751__, new_new_n11752__,
    new_new_n11753__, new_new_n11754__, new_new_n11756__, new_new_n11757__,
    new_new_n11758__, new_new_n11759__, new_new_n11760__, new_new_n11761__,
    new_new_n11762__, new_new_n11763__, new_new_n11764__, new_new_n11765__,
    new_new_n11766__, new_new_n11767__, new_new_n11768__, new_new_n11769__,
    new_new_n11771__, new_new_n11772__, new_new_n11773__, new_new_n11774__,
    new_new_n11775__, new_new_n11776__, new_new_n11777__, new_new_n11778__,
    new_new_n11779__, new_new_n11781__, new_new_n11782__, new_new_n11783__,
    new_new_n11784__, new_new_n11785__, new_new_n11786__, new_new_n11787__,
    new_new_n11789__, new_new_n11791__, new_new_n11792__, new_new_n11793__,
    new_new_n11794__, new_new_n11795__, new_new_n11796__, new_new_n11797__,
    new_new_n11798__, new_new_n11799__, new_new_n11800__, new_new_n11801__,
    new_new_n11802__, new_new_n11803__, new_new_n11804__, new_new_n11806__,
    new_new_n11807__, new_new_n11808__, new_new_n11809__, new_new_n11810__,
    new_new_n11811__, new_new_n11812__, new_new_n11814__, new_new_n11815__,
    new_new_n11816__, new_new_n11817__, new_new_n11819__, new_new_n11820__,
    new_new_n11821__, new_new_n11822__, new_new_n11823__, new_new_n11824__,
    new_new_n11826__, new_new_n11828__, new_new_n11829__, new_new_n11830__,
    new_new_n11831__, new_new_n11832__, new_new_n11833__, new_new_n11834__,
    new_new_n11836__, new_new_n11837__, new_new_n11838__, new_new_n11840__,
    new_new_n11841__, new_new_n11842__, new_new_n11843__, new_new_n11844__,
    new_new_n11845__, new_new_n11846__, new_new_n11848__, new_new_n11849__,
    new_new_n11851__, new_new_n11852__, new_new_n11853__, new_new_n11854__,
    new_new_n11856__, new_new_n11857__, new_new_n11858__, new_new_n11859__,
    new_new_n11860__, new_new_n11861__, new_new_n11863__, new_new_n11865__,
    new_new_n11866__, new_new_n11867__, new_new_n11868__, new_new_n11869__,
    new_new_n11871__, new_new_n11872__, new_new_n11873__, new_new_n11874__,
    new_new_n11876__, new_new_n11877__, new_new_n11878__, new_new_n11879__,
    new_new_n11881__, new_new_n11882__, new_new_n11883__, new_new_n11884__,
    new_new_n11885__, new_new_n11886__, new_new_n11888__, new_new_n11890__,
    new_new_n11891__, new_new_n11892__, new_new_n11893__, new_new_n11894__,
    new_new_n11896__, new_new_n11897__, new_new_n11898__, new_new_n11899__,
    new_new_n11901__, new_new_n11902__, new_new_n11903__, new_new_n11904__,
    new_new_n11906__, new_new_n11907__, new_new_n11908__, new_new_n11909__,
    new_new_n11910__, new_new_n11911__, new_new_n11913__, new_new_n11915__,
    new_new_n11916__, new_new_n11917__, new_new_n11918__, new_new_n11919__,
    new_new_n11921__, new_new_n11922__, new_new_n11923__, new_new_n11924__,
    new_new_n11926__, new_new_n11927__, new_new_n11928__, new_new_n11929__,
    new_new_n11931__, new_new_n11932__, new_new_n11933__, new_new_n11934__,
    new_new_n11935__, new_new_n11936__, new_new_n11938__, new_new_n11940__,
    new_new_n11941__, new_new_n11942__, new_new_n11943__, new_new_n11944__,
    new_new_n11946__, new_new_n11947__, new_new_n11948__, new_new_n11949__,
    new_new_n11951__, new_new_n11952__, new_new_n11953__, new_new_n11954__,
    new_new_n11956__, new_new_n11957__, new_new_n11958__, new_new_n11959__,
    new_new_n11960__, new_new_n11961__, new_new_n11963__, new_new_n11965__,
    new_new_n11966__, new_new_n11967__, new_new_n11968__, new_new_n11969__,
    new_new_n11971__, new_new_n11972__, new_new_n11973__, new_new_n11974__,
    new_new_n11976__, new_new_n11977__, new_new_n11978__, new_new_n11979__,
    new_new_n11981__, new_new_n11982__, new_new_n11983__, new_new_n11984__,
    new_new_n11985__, new_new_n11986__, new_new_n11988__, new_new_n11990__,
    new_new_n11991__, new_new_n11992__, new_new_n11993__, new_new_n11994__,
    new_new_n11996__, new_new_n11997__, new_new_n11998__, new_new_n11999__,
    new_new_n12001__, new_new_n12002__, new_new_n12003__, new_new_n12004__,
    new_new_n12006__, new_new_n12007__, new_new_n12008__, new_new_n12009__,
    new_new_n12010__, new_new_n12011__, new_new_n12013__, new_new_n12015__,
    new_new_n12016__, new_new_n12017__, new_new_n12018__, new_new_n12019__,
    new_new_n12021__, new_new_n12022__, new_new_n12023__, new_new_n12024__,
    new_new_n12026__, new_new_n12027__, new_new_n12028__, new_new_n12029__,
    new_new_n12031__, new_new_n12032__, new_new_n12033__, new_new_n12034__,
    new_new_n12035__, new_new_n12036__, new_new_n12038__, new_new_n12040__,
    new_new_n12041__, new_new_n12042__, new_new_n12043__, new_new_n12044__,
    new_new_n12046__, new_new_n12047__, new_new_n12048__, new_new_n12049__,
    new_new_n12051__, new_new_n12053__, new_new_n12054__, new_new_n12055__,
    new_new_n12056__, new_new_n12057__, new_new_n12058__, new_new_n12059__,
    new_new_n12060__, new_new_n12061__, new_new_n12062__, new_new_n12063__,
    new_new_n12064__, new_new_n12065__, new_new_n12067__, new_new_n12068__,
    new_new_n12069__, new_new_n12070__, new_new_n12072__, new_new_n12073__,
    new_new_n12074__, new_new_n12075__, new_new_n12076__, new_new_n12077__,
    new_new_n12078__, new_new_n12079__, new_new_n12080__, new_new_n12081__,
    new_new_n12082__, new_new_n12083__, new_new_n12084__, new_new_n12085__,
    new_new_n12086__, new_new_n12087__, new_new_n12088__, new_new_n12089__,
    new_new_n12090__, new_new_n12092__, new_new_n12093__, new_new_n12094__,
    new_new_n12095__, new_new_n12096__, new_new_n12097__, new_new_n12098__,
    new_new_n12099__, new_new_n12100__, new_new_n12101__, new_new_n12102__,
    new_new_n12103__, new_new_n12104__, new_new_n12105__, new_new_n12106__,
    new_new_n12108__, new_new_n12111__, new_new_n12112__, new_new_n12113__,
    new_new_n12114__, new_new_n12115__, new_new_n12116__, new_new_n12117__,
    new_new_n12118__, new_new_n12119__, new_new_n12120__, new_new_n12121__,
    new_new_n12122__, new_new_n12124__, new_new_n12125__, new_new_n12126__,
    new_new_n12127__, new_new_n12129__, new_new_n12130__, new_new_n12131__,
    new_new_n12132__, new_new_n12133__, new_new_n12134__, new_new_n12135__,
    new_new_n12136__, new_new_n12137__, new_new_n12138__, new_new_n12140__,
    new_new_n12141__, new_new_n12142__, new_new_n12143__, new_new_n12144__,
    new_new_n12146__, new_new_n12148__, new_new_n12149__, new_new_n12150__,
    new_new_n12151__, new_new_n12152__, new_new_n12153__, new_new_n12154__,
    new_new_n12155__, new_new_n12156__, new_new_n12157__, new_new_n12159__,
    new_new_n12160__, new_new_n12161__, new_new_n12162__, new_new_n12163__,
    new_new_n12164__, new_new_n12165__, new_new_n12166__, new_new_n12167__,
    new_new_n12168__, new_new_n12170__, new_new_n12171__, new_new_n12172__,
    new_new_n12173__, new_new_n12174__, new_new_n12175__, new_new_n12176__,
    new_new_n12177__, new_new_n12178__, new_new_n12179__, new_new_n12181__,
    new_new_n12182__, new_new_n12183__, new_new_n12184__, new_new_n12185__,
    new_new_n12186__, new_new_n12187__, new_new_n12188__, new_new_n12189__,
    new_new_n12190__, new_new_n12192__, new_new_n12193__, new_new_n12194__,
    new_new_n12195__, new_new_n12196__, new_new_n12197__, new_new_n12198__,
    new_new_n12199__, new_new_n12200__, new_new_n12201__, new_new_n12203__,
    new_new_n12204__, new_new_n12205__, new_new_n12206__, new_new_n12207__,
    new_new_n12208__, new_new_n12209__, new_new_n12210__, new_new_n12211__,
    new_new_n12212__, new_new_n12214__, new_new_n12215__, new_new_n12216__,
    new_new_n12217__, new_new_n12218__, new_new_n12219__, new_new_n12221__,
    new_new_n12222__, new_new_n12223__, new_new_n12224__, new_new_n12225__,
    new_new_n12226__, new_new_n12227__, new_new_n12228__, new_new_n12232__,
    new_new_n12234__, new_new_n12235__, new_new_n12236__, new_new_n12237__,
    new_new_n12238__, new_new_n12240__, new_new_n12241__, new_new_n12242__,
    new_new_n12243__, new_new_n12244__, new_new_n12245__, new_new_n12246__,
    new_new_n12247__, new_new_n12248__, new_new_n12249__, new_new_n12250__,
    new_new_n12251__, new_new_n12252__, new_new_n12253__, new_new_n12254__,
    new_new_n12255__, new_new_n12256__, new_new_n12257__, new_new_n12259__,
    new_new_n12260__, new_new_n12261__, new_new_n12262__, new_new_n12263__,
    new_new_n12264__, new_new_n12265__, new_new_n12266__, new_new_n12267__,
    new_new_n12268__, new_new_n12269__, new_new_n12270__, new_new_n12271__,
    new_new_n12272__, new_new_n12273__, new_new_n12274__, new_new_n12275__,
    new_new_n12276__, new_new_n12277__, new_new_n12278__, new_new_n12279__,
    new_new_n12280__, new_new_n12281__, new_new_n12282__, new_new_n12283__,
    new_new_n12284__, new_new_n12285__, new_new_n12286__, new_new_n12287__,
    new_new_n12289__, new_new_n12291__, new_new_n12292__, new_new_n12293__,
    new_new_n12294__, new_new_n12297__, new_new_n12298__, new_new_n12300__,
    new_new_n12303__, new_new_n12304__, new_new_n12305__, new_new_n12306__,
    new_new_n12307__, new_new_n12308__, new_new_n12309__, new_new_n12310__,
    new_new_n12312__, new_new_n12313__, new_new_n12314__, new_new_n12315__,
    new_new_n12316__, new_new_n12317__, new_new_n12318__, new_new_n12319__,
    new_new_n12320__, new_new_n12321__, new_new_n12322__, new_new_n12323__,
    new_new_n12324__, new_new_n12325__, new_new_n12326__, new_new_n12327__,
    new_new_n12328__, new_new_n12329__, new_new_n12331__, new_new_n12332__,
    new_new_n12333__, new_new_n12336__, new_new_n12337__, new_new_n12338__,
    new_new_n12339__, new_new_n12340__, new_new_n12341__, new_new_n12342__,
    new_new_n12343__, new_new_n12344__, new_new_n12345__, new_new_n12346__,
    new_new_n12347__, new_new_n12348__, new_new_n12349__, new_new_n12350__,
    new_new_n12351__, new_new_n12352__, new_new_n12354__, new_new_n12355__,
    new_new_n12356__, new_new_n12357__, new_new_n12358__, new_new_n12359__,
    new_new_n12360__, new_new_n12361__, new_new_n12362__, new_new_n12363__,
    new_new_n12364__, new_new_n12365__, new_new_n12366__, new_new_n12368__,
    new_new_n12369__, new_new_n12370__, new_new_n12371__, new_new_n12373__,
    new_new_n12374__, new_new_n12375__, new_new_n12377__, new_new_n12378__,
    new_new_n12379__, new_new_n12380__, new_new_n12382__, new_new_n12383__,
    new_new_n12385__, new_new_n12386__, new_new_n12388__, new_new_n12389__,
    new_new_n12391__, new_new_n12392__, new_new_n12393__, new_new_n12394__,
    new_new_n12395__, new_new_n12396__, new_new_n12397__, new_new_n12400__,
    new_new_n12401__, new_new_n12403__, new_new_n12404__, new_new_n12406__,
    new_new_n12407__, new_new_n12408__, new_new_n12410__, new_new_n12411__,
    new_new_n12413__, new_new_n12414__, new_new_n12416__, new_new_n12417__,
    new_new_n12419__, new_new_n12420__, new_new_n12422__, new_new_n12423__,
    new_new_n12425__, new_new_n12426__, new_new_n12428__, new_new_n12429__,
    new_new_n12430__, new_new_n12431__, new_new_n12432__, new_new_n12434__,
    new_new_n12439__, new_new_n12443__, new_new_n12447__, new_new_n12448__,
    new_new_n12450__, new_new_n12451__, new_new_n12452__, new_new_n12453__,
    new_new_n12455__, new_new_n12456__, new_new_n12458__, new_new_n12459__,
    new_new_n12460__, new_new_n12461__, new_new_n12472__, new_new_n12473__,
    new_new_n12475__, new_new_n12476__, new_new_n12477__, new_new_n12483__,
    new_new_n12484__, new_new_n12485__, new_new_n12486__, new_new_n12488__,
    new_new_n12489__, new_new_n12490__, new_new_n12491__, new_new_n12492__,
    new_new_n12494__, new_new_n12495__, new_new_n12496__, new_new_n12497__,
    new_new_n12498__, new_new_n12499__, new_new_n12500__, new_new_n12501__,
    new_new_n12502__, new_new_n12503__, new_new_n12505__, new_new_n12507__,
    new_new_n12509__, new_new_n12510__, new_new_n12517__, new_new_n12518__,
    new_new_n12519__, new_new_n12521__, new_new_n12526__, new_new_n12528__,
    new_new_n12553__, new_new_n12555__, new_new_n12556__, new_new_n12557__,
    new_new_n12558__, new_new_n12559__, new_new_n12560__, new_new_n12562__,
    new_new_n12564__, new_new_n12565__, new_new_n12566__, new_new_n12567__,
    new_new_n12568__, new_new_n12569__, new_new_n12573__, new_new_n12574__,
    new_new_n12575__, new_new_n12579__, new_new_n12580__, new_new_n12581__,
    new_new_n12582__, new_new_n12583__, new_new_n12584__, new_new_n12585__,
    new_new_n12586__, new_new_n12588__, new_new_n12589__, new_new_n12592__,
    new_new_n12593__, new_new_n12594__, new_new_n12595__, new_new_n12596__,
    new_new_n12597__, new_new_n12598__, new_new_n12599__, new_new_n12600__,
    new_new_n12601__, new_new_n12602__, new_new_n12603__, new_new_n12604__,
    new_new_n12605__, new_new_n12606__, new_new_n12607__, new_new_n12608__,
    new_new_n12610__, new_new_n12612__, new_new_n12613__, new_new_n12614__,
    new_new_n12615__, new_new_n12616__, new_new_n12617__, new_new_n12618__,
    new_new_n12619__, new_new_n12620__, new_new_n12621__, new_new_n12622__,
    new_new_n12623__, new_new_n12624__, new_new_n12625__, new_new_n12626__,
    new_new_n12627__, new_new_n12629__, new_new_n12631__, new_new_n12633__,
    new_new_n12635__, new_new_n12637__, new_new_n12638__, new_new_n12639__,
    new_new_n12640__, new_new_n12641__, new_new_n12642__, new_new_n12643__,
    new_new_n12644__, new_new_n12645__, new_new_n12646__, new_new_n12647__,
    new_new_n12648__, new_new_n12649__, new_new_n12650__, new_new_n12651__,
    new_new_n12652__, new_new_n12653__, new_new_n12654__, new_new_n12655__,
    new_new_n12656__, new_new_n12657__, new_new_n12658__, new_new_n12659__,
    new_new_n12660__, new_new_n12661__, new_new_n12662__, new_new_n12663__,
    new_new_n12664__, new_new_n12665__, new_new_n12666__, new_new_n12667__,
    new_new_n12668__, new_new_n12669__, new_new_n12670__, new_new_n12671__,
    new_new_n12672__, new_new_n12673__, new_new_n12674__, new_new_n12675__,
    new_new_n12676__, new_new_n12677__, new_new_n12678__, new_new_n12679__,
    new_new_n12680__, new_new_n12681__, new_new_n12682__, new_new_n12683__,
    new_new_n12684__, new_new_n12685__, new_new_n12686__, new_new_n12687__,
    new_new_n12688__, new_new_n12689__, new_new_n12690__, new_new_n12691__,
    new_new_n12692__, new_new_n12693__, new_new_n12694__, new_new_n12695__,
    new_new_n12696__, new_new_n12697__, new_new_n12698__, new_new_n12699__,
    new_new_n12700__, new_new_n12701__, new_new_n12702__, new_new_n12703__,
    new_new_n12704__, new_new_n12705__, new_new_n12706__, new_new_n12707__,
    new_new_n12708__, new_new_n12709__, new_new_n12710__, new_new_n12711__,
    new_new_n12712__, new_new_n12713__, new_new_n12714__, new_new_n12715__,
    new_new_n12716__, new_new_n12717__, new_new_n12718__, new_new_n12719__,
    new_new_n12720__, new_new_n12721__, new_new_n12722__, new_new_n12723__,
    new_new_n12724__, new_new_n12725__, new_new_n12726__, new_new_n12727__,
    new_new_n12728__, new_new_n12729__, new_new_n12730__, new_new_n12731__,
    new_new_n12732__, new_new_n12733__, new_new_n12734__, new_new_n12735__,
    new_new_n12736__, new_new_n12737__, new_new_n12738__, new_new_n12739__,
    new_new_n12740__, new_new_n12741__, new_new_n12742__, new_new_n12743__,
    new_new_n12744__, new_new_n12745__, new_new_n12746__, new_new_n12747__,
    new_new_n12748__, new_new_n12749__, new_new_n12750__, new_new_n12751__,
    new_new_n12752__, new_new_n12753__, new_new_n12754__, new_new_n12755__,
    new_new_n12756__, new_new_n12757__, new_new_n12758__, new_new_n12759__,
    new_new_n12760__, new_new_n12761__, new_new_n12762__, new_new_n12763__,
    new_new_n12764__, new_new_n12765__, new_new_n12766__, new_new_n12767__,
    new_new_n12768__, new_new_n12769__, new_new_n12770__, new_new_n12771__,
    new_new_n12772__, new_new_n12773__, new_new_n12774__, new_new_n12775__,
    new_new_n12776__, new_new_n12777__, new_new_n12778__, new_new_n12779__,
    new_new_n12780__, new_new_n12781__, new_new_n12782__, new_new_n12783__,
    new_new_n12784__, new_new_n12785__, new_new_n12786__, new_new_n12787__,
    new_new_n12788__, new_new_n12789__, new_new_n12790__, new_new_n12791__,
    new_new_n12792__, new_new_n12793__, new_new_n12794__, new_new_n12795__,
    new_new_n12796__, new_new_n12797__, new_new_n12798__, new_new_n12799__,
    new_new_n12800__, new_new_n12801__, new_new_n12802__, new_new_n12803__,
    new_new_n12804__, new_new_n12805__, new_new_n12806__, new_new_n12807__,
    new_new_n12808__, new_new_n12809__, new_new_n12810__, new_new_n12811__,
    new_new_n12812__, new_new_n12813__, new_new_n12814__, new_new_n12815__,
    new_new_n12816__, new_new_n12817__, new_new_n12818__, new_new_n12819__,
    new_new_n12820__, new_new_n12821__, new_new_n12822__, new_new_n12823__,
    new_new_n12824__, new_new_n12825__, new_new_n12826__, new_new_n12827__,
    new_new_n12828__, new_new_n12829__, new_new_n12830__, new_new_n12831__,
    new_new_n12832__, new_new_n12833__, new_new_n12834__, new_new_n12835__,
    new_new_n12836__, new_new_n12837__, new_new_n12838__, new_new_n12839__,
    new_new_n12840__, new_new_n12841__, new_new_n12842__, new_new_n12843__,
    new_new_n12844__, new_new_n12845__, new_new_n12846__, new_new_n12847__,
    new_new_n12848__, new_new_n12849__, new_new_n12850__, new_new_n12851__,
    new_new_n12852__, new_new_n12853__, new_new_n12854__, new_new_n12855__,
    new_new_n12856__, new_new_n12857__, new_new_n12858__, new_new_n12859__,
    new_new_n12860__, new_new_n12861__, new_new_n12862__, new_new_n12863__,
    new_new_n12864__, new_new_n12865__, new_new_n12866__, new_new_n12867__,
    new_new_n12868__, new_new_n12869__, new_new_n12870__, new_new_n12871__,
    new_new_n12872__, new_new_n12873__, new_new_n12874__, new_new_n12875__,
    new_new_n12876__, new_new_n12877__, new_new_n12878__, new_new_n12879__,
    new_new_n12880__, new_new_n12881__, new_new_n12882__, new_new_n12883__,
    new_new_n12884__, new_new_n12885__, new_new_n12886__, new_new_n12887__,
    new_new_n12888__, new_new_n12889__, new_new_n12890__, new_new_n12891__,
    new_new_n12892__, new_new_n12893__, new_new_n12894__, new_new_n12895__,
    new_new_n12896__, new_new_n12897__, new_new_n12898__, new_new_n12899__,
    new_new_n12900__, new_new_n12901__, new_new_n12902__, new_new_n12903__,
    new_new_n12904__, new_new_n12905__, new_new_n12906__, new_new_n12907__,
    new_new_n12908__, new_new_n12909__, new_new_n12910__, new_new_n12911__,
    new_new_n12912__, new_new_n12913__, new_new_n12914__, new_new_n12915__,
    new_new_n12916__, new_new_n12917__, new_new_n12918__, new_new_n12919__,
    new_new_n12920__, new_new_n12921__, new_new_n12922__, new_new_n12923__,
    new_new_n12924__, new_new_n12925__, new_new_n12926__, new_new_n12927__,
    new_new_n12928__, new_new_n12929__, new_new_n12930__, new_new_n12931__,
    new_new_n12932__, new_new_n12933__, new_new_n12934__, new_new_n12935__,
    new_new_n12936__, new_new_n12937__, new_new_n12938__, new_new_n12939__,
    new_new_n12940__, new_new_n12941__, new_new_n12942__, new_new_n12943__,
    new_new_n12944__, new_new_n12945__, new_new_n12946__, new_new_n12947__,
    new_new_n12948__, new_new_n12949__, new_new_n12950__, new_new_n12951__,
    new_new_n12952__, new_new_n12953__, new_new_n12954__, new_new_n12955__,
    new_new_n12956__, new_new_n12957__, new_new_n12958__, new_new_n12959__,
    new_new_n12960__, new_new_n12961__, new_new_n12962__, new_new_n12963__,
    new_new_n12964__, new_new_n12965__, new_new_n12966__, new_new_n12967__,
    new_new_n12968__, new_new_n12969__, new_new_n12970__, new_new_n12971__,
    new_new_n12972__, new_new_n12973__, new_new_n12974__, new_new_n12975__,
    new_new_n12976__, new_new_n12977__, new_new_n12978__, new_new_n12979__,
    new_new_n12980__, new_new_n12981__, new_new_n12982__, new_new_n12983__,
    new_new_n12984__, new_new_n12985__, new_new_n12986__, new_new_n12987__,
    new_new_n12988__, new_new_n12989__, new_new_n12990__, new_new_n12991__,
    new_new_n12992__, new_new_n12993__, new_new_n12994__, new_new_n12995__,
    new_new_n12996__, new_new_n12997__, new_new_n12998__, new_new_n12999__,
    new_new_n13000__, new_new_n13001__, new_new_n13002__, new_new_n13003__,
    new_new_n13004__, new_new_n13005__, new_new_n13006__, new_new_n13007__,
    new_new_n13008__, new_new_n13009__, new_new_n13010__, new_new_n13011__,
    new_new_n13012__, new_new_n13013__, new_new_n13014__, new_new_n13015__,
    new_new_n13016__, new_new_n13017__, new_new_n13018__, new_new_n13019__,
    new_new_n13020__, new_new_n13021__, new_new_n13022__, new_new_n13023__,
    new_new_n13024__, new_new_n13025__, new_new_n13026__, new_new_n13027__,
    new_new_n13028__, new_new_n13029__, new_new_n13030__, new_new_n13031__,
    new_new_n13032__, new_new_n13033__, new_new_n13034__, new_new_n13035__,
    new_new_n13036__, new_new_n13037__, new_new_n13038__, new_new_n13039__,
    new_new_n13040__, new_new_n13041__, new_new_n13042__, new_new_n13043__,
    new_new_n13044__, new_new_n13045__, new_new_n13046__, new_new_n13047__,
    new_new_n13048__, new_new_n13049__, new_new_n13050__, new_new_n13051__,
    new_new_n13052__, new_new_n13053__, new_new_n13054__, new_new_n13055__,
    new_new_n13056__, new_new_n13057__, new_new_n13058__, new_new_n13059__,
    new_new_n13060__, new_new_n13061__, new_new_n13062__, new_new_n13063__,
    new_new_n13064__, new_new_n13065__, new_new_n13066__, new_new_n13067__,
    new_new_n13068__, new_new_n13069__, new_new_n13070__, new_new_n13071__,
    new_new_n13072__, new_new_n13073__, new_new_n13074__, new_new_n13075__,
    new_new_n13076__, new_new_n13077__, new_new_n13078__, new_new_n13079__,
    new_new_n13080__, new_new_n13081__, new_new_n13082__, new_new_n13083__,
    new_new_n13084__, new_new_n13085__, new_new_n13086__, new_new_n13087__,
    new_new_n13088__, new_new_n13089__, new_new_n13090__, new_new_n13091__,
    new_new_n13092__, new_new_n13093__, new_new_n13094__, new_new_n13095__,
    new_new_n13096__, new_new_n13097__, new_new_n13098__, new_new_n13099__,
    new_new_n13100__, new_new_n13101__, new_new_n13102__, new_new_n13103__,
    new_new_n13104__, new_new_n13105__, new_new_n13106__, new_new_n13107__,
    new_new_n13108__, new_new_n13109__, new_new_n13110__, new_new_n13111__,
    new_new_n13112__, new_new_n13113__, new_new_n13114__, new_new_n13115__,
    new_new_n13116__, new_new_n13117__, new_new_n13118__, new_new_n13119__,
    new_new_n13120__, new_new_n13121__, new_new_n13122__, new_new_n13123__,
    new_new_n13124__, new_new_n13125__, new_new_n13126__, new_new_n13127__,
    new_new_n13128__, new_new_n13129__, new_new_n13130__, new_new_n13131__,
    new_new_n13132__, new_new_n13133__, new_new_n13134__, new_new_n13135__,
    new_new_n13136__, new_new_n13137__, new_new_n13138__, new_new_n13139__,
    new_new_n13140__, new_new_n13141__, new_new_n13142__, new_new_n13143__,
    new_new_n13144__, new_new_n13145__, new_new_n13146__, new_new_n13147__,
    new_new_n13148__, new_new_n13149__, new_new_n13150__, new_new_n13151__,
    new_new_n13152__, new_new_n13153__, new_new_n13154__, new_new_n13155__,
    new_new_n13156__, new_new_n13157__, new_new_n13158__, new_new_n13159__,
    new_new_n13160__, new_new_n13161__, new_new_n13162__, new_new_n13163__,
    new_new_n13164__, new_new_n13165__, new_new_n13166__, new_new_n13167__,
    new_new_n13168__, new_new_n13169__, new_new_n13170__, new_new_n13171__,
    new_new_n13172__, new_new_n13173__, new_new_n13174__, new_new_n13175__,
    new_new_n13176__, new_new_n13177__, new_new_n13178__, new_new_n13179__,
    new_new_n13180__, new_new_n13181__, new_new_n13182__, new_new_n13183__,
    new_new_n13184__, new_new_n13185__, new_new_n13186__, new_new_n13187__,
    new_new_n13188__, new_new_n13189__, new_new_n13190__, new_new_n13191__,
    new_new_n13192__, new_new_n13193__, new_new_n13194__, new_new_n13195__,
    new_new_n13196__, new_new_n13197__, new_new_n13198__, new_new_n13199__,
    new_new_n13200__, new_new_n13201__, new_new_n13202__, new_new_n13203__,
    new_new_n13204__, new_new_n13205__, new_new_n13206__, new_new_n13207__,
    new_new_n13208__, new_new_n13209__, new_new_n13210__, new_new_n13211__,
    new_new_n13212__, new_new_n13213__, new_new_n13214__, new_new_n13215__,
    new_new_n13216__, new_new_n13217__, new_new_n13218__, new_new_n13219__,
    new_new_n13220__, new_new_n13221__, new_new_n13222__, new_new_n13223__,
    new_new_n13224__, new_new_n13225__, new_new_n13226__, new_new_n13227__,
    new_new_n13228__, new_new_n13229__, new_new_n13230__, new_new_n13231__,
    new_new_n13232__, new_new_n13233__, new_new_n13234__, new_new_n13235__,
    new_new_n13236__, new_new_n13237__, new_new_n13238__, new_new_n13239__,
    new_new_n13240__, new_new_n13241__, new_new_n13242__, new_new_n13243__,
    new_new_n13244__, new_new_n13245__, new_new_n13246__, new_new_n13247__,
    new_new_n13248__, new_new_n13249__, new_new_n13250__, new_new_n13251__,
    new_new_n13252__, new_new_n13253__, new_new_n13254__, new_new_n13255__,
    new_new_n13256__, new_new_n13257__, new_new_n13258__, new_new_n13259__,
    new_new_n13260__, new_new_n13261__, new_new_n13262__, new_new_n13263__,
    new_new_n13264__, new_new_n13265__, new_new_n13266__, new_new_n13267__,
    new_new_n13268__, new_new_n13269__, new_new_n13270__, new_new_n13271__,
    new_new_n13272__, new_new_n13273__, new_new_n13274__, new_new_n13275__,
    new_new_n13276__, new_new_n13277__, new_new_n13278__, new_new_n13279__,
    new_new_n13280__, new_new_n13281__, new_new_n13282__, new_new_n13283__,
    new_new_n13284__, new_new_n13285__, new_new_n13286__, new_new_n13287__,
    new_new_n13288__, new_new_n13289__, new_new_n13290__, new_new_n13291__,
    new_new_n13292__, new_new_n13293__, new_new_n13294__, new_new_n13295__,
    new_new_n13296__, new_new_n13297__, new_new_n13298__, new_new_n13299__,
    new_new_n13300__, new_new_n13301__, new_new_n13302__, new_new_n13303__,
    new_new_n13304__, new_new_n13305__, new_new_n13306__, new_new_n13307__,
    new_new_n13308__, new_new_n13309__, new_new_n13310__, new_new_n13311__,
    new_new_n13312__, new_new_n13313__, new_new_n13314__, new_new_n13315__,
    new_new_n13316__, new_new_n13317__, new_new_n13318__, new_new_n13319__,
    new_new_n13320__, new_new_n13321__, new_new_n13322__, new_new_n13323__,
    new_new_n13324__, new_new_n13325__, new_new_n13326__, new_new_n13327__,
    new_new_n13328__, new_new_n13329__, new_new_n13330__, new_new_n13331__,
    new_new_n13332__, new_new_n13333__, new_new_n13334__, new_new_n13335__,
    new_new_n13336__, new_new_n13337__, new_new_n13338__, new_new_n13339__,
    new_new_n13340__, new_new_n13341__, new_new_n13342__, new_new_n13343__,
    new_new_n13344__, new_new_n13345__, new_new_n13346__, new_new_n13347__,
    new_new_n13348__, new_new_n13349__, new_new_n13350__, new_new_n13351__,
    new_new_n13352__, new_new_n13353__, new_new_n13354__, new_new_n13355__,
    new_new_n13356__, new_new_n13357__, new_new_n13358__, new_new_n13359__,
    new_new_n13360__, new_new_n13361__, new_new_n13362__, new_new_n13363__,
    new_new_n13364__, new_new_n13365__, new_new_n13366__, new_new_n13367__,
    new_new_n13368__, new_new_n13369__, new_new_n13370__, new_new_n13371__,
    new_new_n13372__, new_new_n13373__, new_new_n13374__, new_new_n13375__,
    new_new_n13376__, new_new_n13377__, new_new_n13378__, new_new_n13379__,
    new_new_n13380__, new_new_n13381__, new_new_n13382__, new_new_n13383__,
    new_new_n13384__, new_new_n13385__, new_new_n13386__, new_new_n13387__,
    new_new_n13388__, new_new_n13389__, new_new_n13390__, new_new_n13391__,
    new_new_n13392__, new_new_n13393__, new_new_n13394__, new_new_n13395__,
    new_new_n13396__, new_new_n13397__, new_new_n13398__, new_new_n13399__,
    new_new_n13400__, new_new_n13401__, new_new_n13402__, new_new_n13403__,
    new_new_n13404__, new_new_n13405__, new_new_n13406__, new_new_n13407__,
    new_new_n13408__, new_new_n13409__, new_new_n13410__, new_new_n13411__,
    new_new_n13412__, new_new_n13413__, new_new_n13414__, new_new_n13415__,
    new_new_n13416__, new_new_n13417__, new_new_n13418__, new_new_n13419__,
    new_new_n13420__, new_new_n13421__, new_new_n13422__, new_new_n13423__,
    new_new_n13424__, new_new_n13425__, new_new_n13426__, new_new_n13427__,
    new_new_n13428__, new_new_n13429__, new_new_n13430__, new_new_n13431__,
    new_new_n13432__, new_new_n13433__, new_new_n13434__, new_new_n13435__,
    new_new_n13436__, new_new_n13437__, new_new_n13438__, new_new_n13439__,
    new_new_n13440__, new_new_n13441__, new_new_n13442__, new_new_n13443__,
    new_new_n13444__, new_new_n13445__, new_new_n13446__, new_new_n13447__,
    new_new_n13448__, new_new_n13449__, new_new_n13450__, new_new_n13451__,
    new_new_n13452__, new_new_n13453__, new_new_n13454__, new_new_n13455__,
    new_new_n13456__, new_new_n13457__, new_new_n13458__, new_new_n13459__,
    new_new_n13460__, new_new_n13461__, new_new_n13462__, new_new_n13463__,
    new_new_n13464__, new_new_n13465__, new_new_n13466__, new_new_n13467__,
    new_new_n13468__, new_new_n13469__, new_new_n13470__, new_new_n13471__,
    new_new_n13472__, new_new_n13473__, new_new_n13474__, new_new_n13475__,
    new_new_n13476__, new_new_n13477__, new_new_n13478__, new_new_n13479__,
    new_new_n13480__, new_new_n13481__, new_new_n13482__, new_new_n13483__,
    new_new_n13484__, new_new_n13485__, new_new_n13486__, new_new_n13487__,
    new_new_n13488__, new_new_n13489__, new_new_n13490__, new_new_n13491__,
    new_new_n13492__, new_new_n13493__, new_new_n13494__, new_new_n13495__,
    new_new_n13496__, new_new_n13497__, new_new_n13498__, new_new_n13499__,
    new_new_n13500__, new_new_n13501__, new_new_n13502__, new_new_n13503__,
    new_new_n13504__, new_new_n13505__, new_new_n13506__, new_new_n13507__,
    new_new_n13508__, new_new_n13509__, new_new_n13510__, new_new_n13511__,
    new_new_n13512__, new_new_n13513__, new_new_n13514__, new_new_n13515__,
    new_new_n13516__, new_new_n13517__, new_new_n13518__, new_new_n13519__,
    new_new_n13520__, new_new_n13521__, new_new_n13522__, new_new_n13523__,
    new_new_n13524__, new_new_n13525__, new_new_n13526__, new_new_n13527__,
    new_new_n13528__, new_new_n13529__, new_new_n13530__, new_new_n13531__,
    new_new_n13532__, new_new_n13533__, new_new_n13534__, new_new_n13535__,
    new_new_n13536__, new_new_n13537__, new_new_n13538__, new_new_n13539__,
    new_new_n13540__, new_new_n13541__, new_new_n13542__, new_new_n13543__,
    new_new_n13544__, new_new_n13545__, new_new_n13546__, new_new_n13547__,
    new_new_n13548__, new_new_n13549__, new_new_n13550__, new_new_n13551__,
    new_new_n13552__, new_new_n13553__, new_new_n13554__, new_new_n13555__,
    new_new_n13556__, new_new_n13557__, new_new_n13558__, new_new_n13559__,
    new_new_n13560__, new_new_n13561__, new_new_n13562__, new_new_n13563__,
    new_new_n13564__, new_new_n13565__, new_new_n13566__, new_new_n13567__,
    new_new_n13568__, new_new_n13569__, new_new_n13570__, new_new_n13571__,
    new_new_n13572__, new_new_n13573__, new_new_n13574__, new_new_n13575__,
    new_new_n13576__, new_new_n13577__, new_new_n13578__, new_new_n13579__,
    new_new_n13580__, new_new_n13581__, new_new_n13582__, new_new_n13583__,
    new_new_n13584__, new_new_n13585__, new_new_n13586__, new_new_n13587__,
    new_new_n13588__, new_new_n13589__, new_new_n13590__, new_new_n13591__,
    new_new_n13592__, new_new_n13593__, new_new_n13594__, new_new_n13595__,
    new_new_n13596__, new_new_n13597__, new_new_n13598__, new_new_n13599__,
    new_new_n13600__, new_new_n13601__, new_new_n13602__, new_new_n13603__,
    new_new_n13604__, new_new_n13605__, new_new_n13606__, new_new_n13607__,
    new_new_n13608__, new_new_n13609__, new_new_n13610__, new_new_n13611__,
    new_new_n13612__, new_new_n13613__, new_new_n13614__, new_new_n13615__,
    new_new_n13616__, new_new_n13617__, new_new_n13618__, new_new_n13619__,
    new_new_n13620__, new_new_n13621__, new_new_n13622__, new_new_n13623__,
    new_new_n13624__, new_new_n13625__, new_new_n13626__, new_new_n13627__,
    new_new_n13628__, new_new_n13629__, new_new_n13630__, new_new_n13631__,
    new_new_n13632__, new_new_n13633__, new_new_n13634__, new_new_n13635__,
    new_new_n13636__, new_new_n13637__, new_new_n13638__, new_new_n13639__,
    new_new_n13640__, new_new_n13641__, new_new_n13642__, new_new_n13643__,
    new_new_n13644__, new_new_n13645__, new_new_n13646__, new_new_n13647__,
    new_new_n13648__, new_new_n13649__, new_new_n13650__, new_new_n13651__,
    new_new_n13652__, new_new_n13653__, new_new_n13654__, new_new_n13655__,
    new_new_n13656__, new_new_n13657__, new_new_n13658__, new_new_n13659__,
    new_new_n13660__, new_new_n13661__, new_new_n13662__, new_new_n13663__,
    new_new_n13664__, new_new_n13665__, new_new_n13666__, new_new_n13667__,
    new_new_n13668__, new_new_n13669__, new_new_n13670__, new_new_n13671__,
    new_new_n13672__, new_new_n13673__, new_new_n13674__, new_new_n13675__,
    new_new_n13676__, new_new_n13677__, new_new_n13678__, new_new_n13679__,
    new_new_n13680__, new_new_n13681__, new_new_n13682__, new_new_n13683__,
    new_new_n13684__, new_new_n13685__, new_new_n13686__, new_new_n13687__,
    new_new_n13688__, new_new_n13689__, new_new_n13690__, new_new_n13691__,
    new_new_n13692__, new_new_n13693__, new_new_n13694__, new_new_n13695__,
    new_new_n13696__, new_new_n13697__, new_new_n13698__, new_new_n13699__,
    new_new_n13700__, new_new_n13701__, new_new_n13702__, new_new_n13703__,
    new_new_n13704__, new_new_n13705__, new_new_n13706__, new_new_n13707__,
    new_new_n13708__, new_new_n13709__, new_new_n13710__, new_new_n13711__,
    new_new_n13712__, new_new_n13713__, new_new_n13714__, new_new_n13715__,
    new_new_n13716__, new_new_n13717__, new_new_n13718__, new_new_n13719__,
    new_new_n13720__, new_new_n13721__, new_new_n13722__, new_new_n13723__,
    new_new_n13724__, new_new_n13725__, new_new_n13726__, new_new_n13727__,
    new_new_n13728__, new_new_n13729__, new_new_n13730__, new_new_n13731__,
    new_new_n13732__, new_new_n13733__, new_new_n13734__, new_new_n13735__,
    new_new_n13736__, new_new_n13737__, new_new_n13738__, new_new_n13739__,
    new_new_n13740__, new_new_n13741__, new_new_n13742__, new_new_n13743__,
    new_new_n13744__, new_new_n13745__, new_new_n13746__, new_new_n13747__,
    new_new_n13748__, new_new_n13749__, new_new_n13750__, new_new_n13751__,
    new_new_n13752__, new_new_n13753__, new_new_n13754__, new_new_n13755__,
    new_new_n13756__, new_new_n13757__, new_new_n13758__, new_new_n13759__,
    new_new_n13760__, new_new_n13761__, new_new_n13762__, new_new_n13763__,
    new_new_n13764__, new_new_n13765__, new_new_n13766__, new_new_n13767__,
    new_new_n13768__, new_new_n13769__, new_new_n13770__, new_new_n13771__,
    new_new_n13772__, new_new_n13773__, new_new_n13774__, new_new_n13775__,
    new_new_n13776__, new_new_n13777__, new_new_n13778__, new_new_n13779__,
    new_new_n13780__, new_new_n13781__, new_new_n13782__, new_new_n13783__,
    new_new_n13784__, new_new_n13785__, new_new_n13786__, new_new_n13787__,
    new_new_n13788__, new_new_n13789__, new_new_n13790__, new_new_n13791__,
    new_new_n13792__, new_new_n13793__, new_new_n13794__, new_new_n13795__,
    new_new_n13796__, new_new_n13797__, new_new_n13798__, new_new_n13799__,
    new_new_n13800__, new_new_n13801__, new_new_n13802__, new_new_n13803__,
    new_new_n13804__, new_new_n13805__, new_new_n13806__, new_new_n13807__,
    new_new_n13808__, new_new_n13809__, new_new_n13810__, new_new_n13811__,
    new_new_n13812__, new_new_n13813__, new_new_n13814__, new_new_n13815__,
    new_new_n13816__, new_new_n13817__, new_new_n13818__, new_new_n13819__,
    new_new_n13820__, new_new_n13821__, new_new_n13822__, new_new_n13823__,
    new_new_n13824__, new_new_n13825__, new_new_n13826__, new_new_n13827__,
    new_new_n13828__, new_new_n13829__, new_new_n13830__, new_new_n13831__,
    new_new_n13832__, new_new_n13833__, new_new_n13834__, new_new_n13835__,
    new_new_n13836__, new_new_n13837__, new_new_n13838__, new_new_n13839__,
    new_new_n13840__, new_new_n13841__, new_new_n13842__, new_new_n13843__,
    new_new_n13844__, new_new_n13845__, new_new_n13846__, new_new_n13847__,
    new_new_n13848__, new_new_n13849__, new_new_n13850__, new_new_n13851__,
    new_new_n13852__, new_new_n13853__, new_new_n13854__, new_new_n13855__,
    new_new_n13856__, new_new_n13857__, new_new_n13858__, new_new_n13859__,
    new_new_n13860__, new_new_n13861__, new_new_n13862__, new_new_n13863__,
    new_new_n13864__, new_new_n13865__, new_new_n13866__, new_new_n13867__,
    new_new_n13868__, new_new_n13869__, new_new_n13870__, new_new_n13871__,
    new_new_n13872__, new_new_n13873__, new_new_n13874__, new_new_n13875__,
    new_new_n13876__, new_new_n13877__, new_new_n13878__, new_new_n13879__,
    new_new_n13880__, new_new_n13881__, new_new_n13882__, new_new_n13883__,
    new_new_n13884__, new_new_n13885__, new_new_n13886__, new_new_n13887__,
    new_new_n13888__, new_new_n13889__, new_new_n13890__, new_new_n13891__,
    new_new_n13893__, new_new_n13894__, new_new_n13895__, new_new_n13896__,
    new_new_n13897__, new_new_n13898__, new_new_n13899__, new_new_n13900__,
    new_new_n13901__, new_new_n13902__, new_new_n13903__, new_new_n13904__,
    new_new_n13905__, new_new_n13906__, new_new_n13907__, new_new_n13908__,
    new_new_n13909__, new_new_n13910__, new_new_n13911__, new_new_n13912__,
    new_new_n13913__, new_new_n13914__, new_new_n13915__, new_new_n13916__,
    new_new_n13917__, new_new_n13918__, new_new_n13919__, new_new_n13920__,
    new_new_n13921__, new_new_n13922__, new_new_n13923__, new_new_n13927__,
    new_new_n13928__, new_new_n13929__, new_new_n13930__, new_new_n13931__,
    new_new_n13932__, new_new_n13933__, new_new_n13934__, new_new_n13935__,
    new_new_n13936__, new_new_n13938__, new_new_n13940__, new_new_n13941__,
    new_new_n13942__, new_new_n13945__, new_new_n13947__, new_new_n13950__,
    new_new_n13951__, new_new_n13954__, new_new_n13958__, new_new_n13959__,
    new_new_n13960__, new_new_n13961__, new_new_n13962__, new_new_n13964__,
    new_new_n13966__, new_new_n13967__, new_new_n13969__, new_new_n13970__,
    new_new_n13971__, new_new_n13972__, new_new_n13974__, new_new_n13975__,
    new_new_n13976__, new_new_n13977__, new_new_n13981__, new_new_n13982__,
    new_new_n13983__, new_new_n13984__, new_new_n13985__, new_new_n13986__,
    new_new_n13987__, new_new_n13988__, new_new_n13989__, new_new_n13990__,
    new_new_n13991__, new_new_n13992__, new_new_n13999__, new_new_n14000__,
    new_new_n14001__, new_new_n14002__, new_new_n14003__, new_new_n14004__,
    new_new_n14006__, new_new_n14012__, new_new_n14013__, new_new_n14014__,
    new_new_n14015__, new_new_n14016__, new_new_n14017__, new_new_n14018__,
    new_new_n14019__, new_new_n14020__, new_new_n14021__, new_new_n14022__,
    new_new_n14024__, new_new_n14025__, new_new_n14026__, new_new_n14027__,
    new_new_n14028__, new_new_n14029__, new_new_n14030__, new_new_n14031__,
    new_new_n14032__, new_new_n14033__, new_new_n14034__, new_new_n14035__,
    new_new_n14036__, new_new_n14037__, new_new_n14038__, new_new_n14039__,
    new_new_n14040__, new_new_n14041__, new_new_n14042__, new_new_n14043__,
    new_new_n14044__, new_new_n14045__, new_new_n14046__, new_new_n14047__,
    new_new_n14048__, new_new_n14049__, new_new_n14050__, new_new_n14051__,
    new_new_n14052__, new_new_n14053__, new_new_n14054__, new_new_n14055__,
    new_new_n14056__, new_new_n14057__, new_new_n14058__, new_new_n14059__,
    new_new_n14060__, new_new_n14061__, new_new_n14062__, new_new_n14063__,
    new_new_n14064__, new_new_n14065__, new_new_n14066__, new_new_n14067__,
    new_new_n14068__, new_new_n14069__, new_new_n14070__, new_new_n14071__,
    new_new_n14072__, new_new_n14073__, new_new_n14074__, new_new_n14075__,
    new_new_n14076__, new_new_n14077__, new_new_n14078__, new_new_n14079__,
    new_new_n14080__, new_new_n14081__, new_new_n14082__, new_new_n14083__,
    new_new_n14084__, new_new_n14085__, new_new_n14086__, new_new_n14087__,
    new_new_n14088__, new_new_n14089__, new_new_n14090__, new_new_n14091__,
    new_new_n14092__, new_new_n14093__, new_new_n14094__, new_new_n14095__,
    new_new_n14096__, new_new_n14097__, new_new_n14098__, new_new_n14099__,
    new_new_n14100__, new_new_n14101__, new_new_n14102__, new_new_n14103__,
    new_new_n14104__, new_new_n14105__, new_new_n14106__, new_new_n14107__,
    new_new_n14108__, new_new_n14109__, new_new_n14110__, new_new_n14111__,
    new_new_n14112__, new_new_n14113__, new_new_n14114__, new_new_n14115__,
    new_new_n14116__, new_new_n14117__, new_new_n14118__, new_new_n14119__,
    new_new_n14120__, new_new_n14121__, new_new_n14122__, new_new_n14123__,
    new_new_n14124__, new_new_n14125__, new_new_n14126__, new_new_n14127__,
    new_new_n14128__, new_new_n14129__, new_new_n14130__, new_new_n14131__,
    new_new_n14132__, new_new_n14133__, new_new_n14134__, new_new_n14135__,
    new_new_n14136__, new_new_n14137__, new_new_n14138__, new_new_n14139__,
    new_new_n14140__, new_new_n14141__, new_new_n14142__, new_new_n14143__,
    new_new_n14144__, new_new_n14145__, new_new_n14146__, new_new_n14147__,
    new_new_n14148__, new_new_n14149__, new_new_n14150__, new_new_n14151__,
    new_new_n14152__, new_new_n14153__, new_new_n14154__, new_new_n14155__,
    new_new_n14156__, new_new_n14157__, new_new_n14158__, new_new_n14159__,
    new_new_n14160__, new_new_n14161__, new_new_n14162__, new_new_n14163__,
    new_new_n14164__, new_new_n14165__, new_new_n14166__, new_new_n14167__,
    new_new_n14168__, new_new_n14169__, new_new_n14170__, new_new_n14171__,
    new_new_n14172__, new_new_n14173__, new_new_n14174__, new_new_n14175__,
    new_new_n14176__, new_new_n14177__, new_new_n14178__, new_new_n14179__,
    new_new_n14180__, new_new_n14181__, new_new_n14182__, new_new_n14183__,
    new_new_n14184__, new_new_n14185__, new_new_n14186__, new_new_n14187__,
    new_new_n14188__, new_new_n14189__, new_new_n14190__, new_new_n14191__,
    new_new_n14192__, new_new_n14193__, new_new_n14194__, new_new_n14195__,
    new_new_n14196__, new_new_n14197__, new_new_n14198__, new_new_n14199__,
    new_new_n14200__, new_new_n14201__, new_new_n14202__, new_new_n14203__,
    new_new_n14204__, new_new_n14205__, new_new_n14206__, new_new_n14207__,
    new_new_n14208__, new_new_n14209__, new_new_n14210__, new_new_n14211__,
    new_new_n14212__, new_new_n14213__, new_new_n14214__, new_new_n14215__,
    new_new_n14216__, new_new_n14217__, new_new_n14218__, new_new_n14219__,
    new_new_n14220__, new_new_n14221__, new_new_n14222__, new_new_n14223__,
    new_new_n14224__, new_new_n14225__, new_new_n14226__, new_new_n14227__,
    new_new_n14228__, new_new_n14229__, new_new_n14230__, new_new_n14231__,
    new_new_n14232__, new_new_n14233__, new_new_n14234__, new_new_n14235__,
    new_new_n14236__, new_new_n14237__, new_new_n14238__, new_new_n14239__,
    new_new_n14240__, new_new_n14241__, new_new_n14242__, new_new_n14243__,
    new_new_n14244__, new_new_n14245__, new_new_n14246__, new_new_n14247__,
    new_new_n14248__, new_new_n14249__, new_new_n14250__, new_new_n14251__,
    new_new_n14252__, new_new_n14253__, new_new_n14254__, new_new_n14255__,
    new_new_n14256__, new_new_n14257__, new_new_n14258__, new_new_n14259__,
    new_new_n14260__, new_new_n14261__, new_new_n14262__, new_new_n14263__,
    new_new_n14264__, new_new_n14265__, new_new_n14266__, new_new_n14267__,
    new_new_n14268__, new_new_n14269__, new_new_n14270__, new_new_n14271__,
    new_new_n14272__, new_new_n14273__, new_new_n14274__, new_new_n14275__,
    new_new_n14276__, new_new_n14277__, new_new_n14278__, new_new_n14279__,
    new_new_n14280__, new_new_n14281__, new_new_n14282__, new_new_n14283__,
    new_new_n14284__, new_new_n14285__, new_new_n14286__, new_new_n14287__,
    new_new_n14288__, new_new_n14289__, new_new_n14290__, new_new_n14291__,
    new_new_n14292__, new_new_n14293__, new_new_n14294__, new_new_n14295__,
    new_new_n14296__, new_new_n14297__, new_new_n14298__, new_new_n14299__,
    new_new_n14300__, new_new_n14301__, new_new_n14302__, new_new_n14303__,
    new_new_n14304__, new_new_n14305__, new_new_n14306__, new_new_n14307__,
    new_new_n14308__, new_new_n14309__, new_new_n14310__, new_new_n14311__,
    new_new_n14312__, new_new_n14313__, new_new_n14314__, new_new_n14315__,
    new_new_n14316__, new_new_n14317__, new_new_n14318__, new_new_n14319__,
    new_new_n14320__, new_new_n14321__, new_new_n14322__, new_new_n14323__,
    new_new_n14324__, new_new_n14325__, new_new_n14326__, new_new_n14327__,
    new_new_n14328__, new_new_n14329__, new_new_n14330__, new_new_n14331__,
    new_new_n14332__, new_new_n14333__, new_new_n14334__, new_new_n14335__,
    new_new_n14336__, new_new_n14337__, new_new_n14338__, new_new_n14339__,
    new_new_n14340__, new_new_n14341__, new_new_n14342__, new_new_n14343__,
    new_new_n14344__, new_new_n14345__, new_new_n14346__, new_new_n14347__,
    new_new_n14348__, new_new_n14349__, new_new_n14350__, new_new_n14351__,
    new_new_n14352__, new_new_n14353__, new_new_n14354__, new_new_n14355__,
    new_new_n14356__, new_new_n14357__, new_new_n14358__, new_new_n14359__,
    new_new_n14360__, new_new_n14361__, new_new_n14362__, new_new_n14363__,
    new_new_n14364__, new_new_n14365__, new_new_n14366__, new_new_n14367__,
    new_new_n14368__, new_new_n14369__, new_new_n14370__, new_new_n14371__,
    new_new_n14372__, new_new_n14373__, new_new_n14374__, new_new_n14375__,
    new_new_n14376__, new_new_n14377__, new_new_n14378__, new_new_n14379__,
    new_new_n14380__, new_new_n14381__, new_new_n14382__, new_new_n14383__,
    new_new_n14384__, new_new_n14385__, new_new_n14386__, new_new_n14387__,
    new_new_n14388__, new_new_n14389__, new_new_n14390__, new_new_n14391__,
    new_new_n14392__, new_new_n14393__, new_new_n14394__, new_new_n14395__,
    new_new_n14396__, new_new_n14397__, new_new_n14398__, new_new_n14399__,
    new_new_n14400__, new_new_n14401__, new_new_n14402__, new_new_n14403__,
    new_new_n14404__, new_new_n14405__, new_new_n14406__, new_new_n14407__,
    new_new_n14408__, new_new_n14409__, new_new_n14410__, new_new_n14411__,
    new_new_n14412__, new_new_n14413__, new_new_n14414__, new_new_n14415__,
    new_new_n14416__, new_new_n14417__, new_new_n14418__, new_new_n14419__,
    new_new_n14420__, new_new_n14421__, new_new_n14422__, new_new_n14423__,
    new_new_n14424__, new_new_n14425__, new_new_n14426__, new_new_n14427__,
    new_new_n14428__, new_new_n14429__, new_new_n14430__, new_new_n14431__,
    new_new_n14432__, new_new_n14433__, new_new_n14434__, new_new_n14435__,
    new_new_n14436__, new_new_n14437__, new_new_n14438__, new_new_n14439__,
    new_new_n14440__, new_new_n14441__, new_new_n14442__, new_new_n14443__,
    new_new_n14444__, new_new_n14445__, new_new_n14446__, new_new_n14447__,
    new_new_n14448__, new_new_n14449__, new_new_n14450__, new_new_n14451__,
    new_new_n14452__, new_new_n14453__, new_new_n14454__, new_new_n14455__,
    new_new_n14456__, new_new_n14457__, new_new_n14458__, new_new_n14459__,
    new_new_n14460__, new_new_n14461__, new_new_n14462__, new_new_n14463__,
    new_new_n14464__, new_new_n14465__, new_new_n14466__, new_new_n14467__,
    new_new_n14468__, new_new_n14469__, new_new_n14470__, new_new_n14471__,
    new_new_n14472__, new_new_n14473__, new_new_n14474__, new_new_n14475__,
    new_new_n14476__, new_new_n14477__, new_new_n14478__, new_new_n14479__,
    new_new_n14480__, new_new_n14481__, new_new_n14482__, new_new_n14483__,
    new_new_n14484__, new_new_n14485__, new_new_n14486__, new_new_n14487__,
    new_new_n14488__, new_new_n14489__, new_new_n14490__, new_new_n14491__,
    new_new_n14492__, new_new_n14493__, new_new_n14494__, new_new_n14495__,
    new_new_n14496__, new_new_n14497__, new_new_n14498__, new_new_n14499__,
    new_new_n14500__, new_new_n14501__, new_new_n14502__, new_new_n14503__,
    new_new_n14504__, new_new_n14505__, new_new_n14506__, new_new_n14507__,
    new_new_n14508__, new_new_n14509__, new_new_n14510__, new_new_n14511__,
    new_new_n14512__, new_new_n14513__, new_new_n14514__, new_new_n14515__,
    new_new_n14516__, new_new_n14517__, new_new_n14518__, new_new_n14519__,
    new_new_n14520__, new_new_n14521__, new_new_n14522__, new_new_n14523__,
    new_new_n14524__, new_new_n14525__, new_new_n14526__, new_new_n14527__,
    new_new_n14528__, new_new_n14529__, new_new_n14530__, new_new_n14531__,
    new_new_n14532__, new_new_n14533__, new_new_n14534__, new_new_n14535__,
    new_new_n14536__, new_new_n14537__, new_new_n14538__, new_new_n14539__,
    new_new_n14540__, new_new_n14541__, new_new_n14542__, new_new_n14543__,
    new_new_n14544__, new_new_n14545__, new_new_n14546__, new_new_n14547__,
    new_new_n14548__, new_new_n14549__, new_new_n14550__, new_new_n14551__,
    new_new_n14552__, new_new_n14553__, new_new_n14554__, new_new_n14555__,
    new_new_n14556__, new_new_n14557__, new_new_n14558__, new_new_n14559__,
    new_new_n14560__, new_new_n14561__, new_new_n14562__, new_new_n14563__,
    new_new_n14564__, new_new_n14565__, new_new_n14566__, new_new_n14567__,
    new_new_n14568__, new_new_n14569__, new_new_n14570__, new_new_n14571__,
    new_new_n14572__, new_new_n14573__, new_new_n14574__, new_new_n14575__,
    new_new_n14576__, new_new_n14577__, new_new_n14578__, new_new_n14579__,
    new_new_n14580__, new_new_n14581__, new_new_n14582__, new_new_n14583__,
    new_new_n14584__, new_new_n14585__, new_new_n14586__, new_new_n14587__,
    new_new_n14588__, new_new_n14589__, new_new_n14590__, new_new_n14591__,
    new_new_n14592__, new_new_n14593__, new_new_n14594__, new_new_n14595__,
    new_new_n14596__, new_new_n14597__, new_new_n14598__, new_new_n14599__,
    new_new_n14600__, new_new_n14601__, new_new_n14602__, new_new_n14603__,
    new_new_n14604__, new_new_n14605__, new_new_n14606__, new_new_n14607__,
    new_new_n14608__, new_new_n14609__, new_new_n14610__, new_new_n14611__,
    new_new_n14612__, new_new_n14613__, new_new_n14614__, new_new_n14615__,
    new_new_n14616__, new_new_n14617__, new_new_n14618__, new_new_n14619__,
    new_new_n14620__, new_new_n14621__, new_new_n14622__, new_new_n14623__,
    new_new_n14624__, new_new_n14625__, new_new_n14626__, new_new_n14627__,
    new_new_n14628__, new_new_n14629__, new_new_n14630__, new_new_n14631__,
    new_new_n14632__, new_new_n14633__, new_new_n14634__, new_new_n14635__,
    new_new_n14636__, new_new_n14637__, new_new_n14638__, new_new_n14639__,
    new_new_n14640__, new_new_n14641__, new_new_n14642__, new_new_n14643__,
    new_new_n14644__, new_new_n14645__, new_new_n14646__, new_new_n14647__,
    new_new_n14648__, new_new_n14649__, new_new_n14650__, new_new_n14651__,
    new_new_n14652__, new_new_n14653__, new_new_n14654__, new_new_n14655__,
    new_new_n14656__, new_new_n14657__, new_new_n14658__, new_new_n14659__,
    new_new_n14660__, new_new_n14661__, new_new_n14662__, new_new_n14663__,
    new_new_n14664__, new_new_n14665__, new_new_n14666__, new_new_n14667__,
    new_new_n14668__, new_new_n14669__, new_new_n14670__, new_new_n14671__,
    new_new_n14672__, new_new_n14673__, new_new_n14674__, new_new_n14675__,
    new_new_n14676__, new_new_n14677__, new_new_n14678__, new_new_n14679__,
    new_new_n14680__, new_new_n14681__, new_new_n14682__, new_new_n14683__,
    new_new_n14684__, new_new_n14685__, new_new_n14686__, new_new_n14687__,
    new_new_n14688__, new_new_n14689__, new_new_n14690__, new_new_n14691__,
    new_new_n14692__, new_new_n14693__, new_new_n14694__, new_new_n14695__,
    new_new_n14696__, new_new_n14697__, new_new_n14698__, new_new_n14699__,
    new_new_n14700__, new_new_n14701__, new_new_n14702__, new_new_n14703__,
    new_new_n14704__, new_new_n14705__, new_new_n14706__, new_new_n14707__,
    new_new_n14708__, new_new_n14709__, new_new_n14710__, new_new_n14711__,
    new_new_n14712__, new_new_n14713__, new_new_n14714__, new_new_n14715__,
    new_new_n14716__, new_new_n14717__, new_new_n14718__, new_new_n14719__,
    new_new_n14720__, new_new_n14721__, new_new_n14722__, new_new_n14723__,
    new_new_n14724__, new_new_n14725__, new_new_n14726__, new_new_n14727__,
    new_new_n14728__, new_new_n14729__, new_new_n14730__, new_new_n14731__,
    new_new_n14732__, new_new_n14733__, new_new_n14734__, new_new_n14735__,
    new_new_n14736__, new_new_n14737__, new_new_n14738__, new_new_n14739__,
    new_new_n14740__, new_new_n14741__, new_new_n14742__, new_new_n14743__,
    new_new_n14744__, new_new_n14745__, new_new_n14746__, new_new_n14747__,
    new_new_n14748__, new_new_n14749__, new_new_n14750__, new_new_n14751__,
    new_new_n14752__, new_new_n14753__, new_new_n14754__, new_new_n14755__,
    new_new_n14756__, new_new_n14757__, new_new_n14758__, new_new_n14759__,
    new_new_n14760__, new_new_n14761__, new_new_n14762__, new_new_n14763__,
    new_new_n14764__, new_new_n14765__, new_new_n14766__, new_new_n14767__,
    new_new_n14768__, new_new_n14769__, new_new_n14770__, new_new_n14771__,
    new_new_n14772__, new_new_n14773__, new_new_n14774__, new_new_n14775__,
    new_new_n14776__, new_new_n14777__, new_new_n14778__, new_new_n14779__,
    new_new_n14780__, new_new_n14781__, new_new_n14782__, new_new_n14783__,
    new_new_n14784__, new_new_n14785__, new_new_n14786__, new_new_n14787__,
    new_new_n14788__, new_new_n14789__, new_new_n14790__, new_new_n14791__,
    new_new_n14792__, new_new_n14793__, new_new_n14794__, new_new_n14795__,
    new_new_n14796__, new_new_n14797__, new_new_n14798__, new_new_n14799__,
    new_new_n14800__, new_new_n14801__, new_new_n14802__, new_new_n14803__,
    new_new_n14804__, new_new_n14805__, new_new_n14806__, new_new_n14807__,
    new_new_n14808__, new_new_n14809__, new_new_n14810__, new_new_n14811__,
    new_new_n14812__, new_new_n14813__, new_new_n14814__, new_new_n14815__,
    new_new_n14816__, new_new_n14817__, new_new_n14818__, new_new_n14819__,
    new_new_n14820__, new_new_n14821__, new_new_n14822__, new_new_n14823__,
    new_new_n14824__, new_new_n14825__, new_new_n14826__, new_new_n14827__,
    new_new_n14828__, new_new_n14829__, new_new_n14830__, new_new_n14831__,
    new_new_n14832__, new_new_n14833__, new_new_n14834__, new_new_n14835__,
    new_new_n14836__, new_new_n14837__, new_new_n14838__, new_new_n14839__,
    new_new_n14840__, new_new_n14841__, new_new_n14842__, new_new_n14843__,
    new_new_n14844__, new_new_n14845__, new_new_n14846__, new_new_n14847__,
    new_new_n14848__, new_new_n14849__, new_new_n14850__, new_new_n14851__,
    new_new_n14852__, new_new_n14853__, new_new_n14854__, new_new_n14855__,
    new_new_n14856__, new_new_n14857__, new_new_n14858__, new_new_n14859__,
    new_new_n14860__, new_new_n14861__, new_new_n14862__, new_new_n14863__,
    new_new_n14864__, new_new_n14865__, new_new_n14866__, new_new_n14867__,
    new_new_n14868__, new_new_n14869__, new_new_n14870__, new_new_n14871__,
    new_new_n14872__, new_new_n14873__, new_new_n14874__, new_new_n14875__,
    new_new_n14876__, new_new_n14877__, new_new_n14878__, new_new_n14879__,
    new_new_n14880__, new_new_n14881__, new_new_n14882__, new_new_n14883__,
    new_new_n14884__, new_new_n14885__, new_new_n14886__, new_new_n14887__,
    new_new_n14888__, new_new_n14889__, new_new_n14890__, new_new_n14891__,
    new_new_n14892__, new_new_n14893__, new_new_n14894__, new_new_n14895__,
    new_new_n14896__, new_new_n14897__, new_new_n14898__, new_new_n14899__,
    new_new_n14900__, new_new_n14901__, new_new_n14902__, new_new_n14903__,
    new_new_n14904__, new_new_n14905__, new_new_n14906__, new_new_n14907__,
    new_new_n14908__, new_new_n14909__, new_new_n14910__, new_new_n14911__,
    new_new_n14912__, new_new_n14913__, new_new_n14914__, new_new_n14915__,
    new_new_n14916__, new_new_n14917__, new_new_n14918__, new_new_n14919__,
    new_new_n14920__, new_new_n14921__, new_new_n14922__, new_new_n14923__,
    new_new_n14924__, new_new_n14925__, new_new_n14926__, new_new_n14927__,
    new_new_n14928__, new_new_n14929__, new_new_n14930__, new_new_n14931__,
    new_new_n14932__, new_new_n14933__, new_new_n14934__, new_new_n14935__,
    new_new_n14936__, new_new_n14937__, new_new_n14938__, new_new_n14939__,
    new_new_n14940__, new_new_n14941__, new_new_n14942__, new_new_n14943__,
    new_new_n14944__, new_new_n14945__, new_new_n14946__, new_new_n14947__,
    new_new_n14948__, new_new_n14949__, new_new_n14950__, new_new_n14951__,
    new_new_n14952__, new_new_n14953__, new_new_n14954__, new_new_n14955__,
    new_new_n14956__, new_new_n14957__, new_new_n14958__, new_new_n14959__,
    new_new_n14960__, new_new_n14961__, new_new_n14962__, new_new_n14963__,
    new_new_n14964__, new_new_n14965__, new_new_n14966__, new_new_n14967__,
    new_new_n14968__, new_new_n14969__, new_new_n14970__, new_new_n14971__,
    new_new_n14972__, new_new_n14973__, new_new_n14974__, new_new_n14975__,
    new_new_n14976__, new_new_n14977__, new_new_n14978__, new_new_n14979__,
    new_new_n14980__, new_new_n14981__, new_new_n14982__, new_new_n14983__,
    new_new_n14984__, new_new_n14985__, new_new_n14986__, new_new_n14987__,
    new_new_n14988__, new_new_n14989__, new_new_n14990__, new_new_n14991__,
    new_new_n14992__, new_new_n14993__, new_new_n14994__, new_new_n14995__,
    new_new_n14996__, new_new_n14997__, new_new_n14998__, new_new_n14999__,
    new_new_n15000__, new_new_n15001__, new_new_n15002__, new_new_n15003__,
    new_new_n15004__, new_new_n15005__, new_new_n15006__, new_new_n15007__,
    new_new_n15008__, new_new_n15009__, new_new_n15010__, new_new_n15011__,
    new_new_n15012__, new_new_n15013__, new_new_n15014__, new_new_n15015__,
    new_new_n15016__, new_new_n15017__, new_new_n15018__, new_new_n15019__,
    new_new_n15020__, new_new_n15021__, new_new_n15022__, new_new_n15023__,
    new_new_n15024__, new_new_n15025__, new_new_n15026__, new_new_n15027__,
    new_new_n15028__, new_new_n15029__, new_new_n15030__, new_new_n15031__,
    new_new_n15032__, new_new_n15033__, new_new_n15034__, new_new_n15035__,
    new_new_n15036__, new_new_n15037__, new_new_n15038__, new_new_n15039__,
    new_new_n15040__, new_new_n15041__, new_new_n15042__, new_new_n15043__,
    new_new_n15044__, new_new_n15045__, new_new_n15046__, new_new_n15047__,
    new_new_n15048__, new_new_n15049__, new_new_n15050__, new_new_n15051__,
    new_new_n15052__, new_new_n15053__, new_new_n15054__, new_new_n15055__,
    new_new_n15056__, new_new_n15057__, new_new_n15058__, new_new_n15059__,
    new_new_n15060__, new_new_n15061__, new_new_n15062__, new_new_n15063__,
    new_new_n15064__, new_new_n15065__, new_new_n15066__, new_new_n15067__,
    new_new_n15068__, new_new_n15069__, new_new_n15070__, new_new_n15071__,
    new_new_n15072__, new_new_n15073__, new_new_n15074__, new_new_n15075__,
    new_new_n15076__, new_new_n15077__, new_new_n15078__, new_new_n15079__,
    new_new_n15080__, new_new_n15081__, new_new_n15082__, new_new_n15083__,
    new_new_n15084__, new_new_n15085__, new_new_n15086__, new_new_n15087__,
    new_new_n15088__, new_new_n15089__, new_new_n15090__, new_new_n15091__,
    new_new_n15092__, new_new_n15093__, new_new_n15094__, new_new_n15095__,
    new_new_n15096__, new_new_n15097__, new_new_n15098__, new_new_n15099__,
    new_new_n15100__, new_new_n15101__, new_new_n15102__, new_new_n15103__,
    new_new_n15104__, new_new_n15105__, new_new_n15106__, new_new_n15107__,
    new_new_n15108__, new_new_n15109__, new_new_n15110__, new_new_n15111__,
    new_new_n15112__, new_new_n15113__, new_new_n15114__, new_new_n15115__,
    new_new_n15116__, new_new_n15117__, new_new_n15118__, new_new_n15119__,
    new_new_n15120__, new_new_n15121__, new_new_n15122__, new_new_n15123__,
    new_new_n15124__, new_new_n15125__, new_new_n15126__, new_new_n15127__,
    new_new_n15128__, new_new_n15129__, new_new_n15130__, new_new_n15131__,
    new_new_n15132__, new_new_n15133__, new_new_n15134__, new_new_n15135__,
    new_new_n15136__, new_new_n15137__, new_new_n15138__, new_new_n15139__,
    new_new_n15140__, new_new_n15141__, new_new_n15142__, new_new_n15143__,
    new_new_n15144__, new_new_n15145__, new_new_n15146__, new_new_n15147__,
    new_new_n15148__, new_new_n15149__, new_new_n15150__, new_new_n15151__,
    new_new_n15152__, new_new_n15153__, new_new_n15154__, new_new_n15155__,
    new_new_n15156__, new_new_n15157__, new_new_n15158__, new_new_n15159__,
    new_new_n15160__, new_new_n15161__, new_new_n15162__, new_new_n15163__,
    new_new_n15164__, new_new_n15165__, new_new_n15166__, new_new_n15167__,
    new_new_n15168__, new_new_n15169__, new_new_n15170__, new_new_n15171__,
    new_new_n15172__, new_new_n15173__, new_new_n15174__, new_new_n15175__,
    new_new_n15176__, new_new_n15177__, new_new_n15178__, new_new_n15179__,
    new_new_n15180__, new_new_n15181__, new_new_n15182__, new_new_n15183__,
    new_new_n15184__, new_new_n15185__, new_new_n15186__, new_new_n15187__,
    new_new_n15188__, new_new_n15189__, new_new_n15190__, new_new_n15191__,
    new_new_n15192__, new_new_n15193__, new_new_n15194__, new_new_n15195__,
    new_new_n15196__, new_new_n15197__, new_new_n15198__, new_new_n15199__,
    new_new_n15200__, new_new_n15201__, new_new_n15202__, new_new_n15203__,
    new_new_n15204__, new_new_n15205__, new_new_n15206__, new_new_n15207__,
    new_new_n15208__, new_new_n15209__, new_new_n15210__, new_new_n15211__,
    new_new_n15212__, new_new_n15213__, new_new_n15214__, new_new_n15215__,
    new_new_n15216__, new_new_n15217__, new_new_n15218__, new_new_n15219__,
    new_new_n15220__, new_new_n15221__, new_new_n15222__, new_new_n15223__,
    new_new_n15224__, new_new_n15225__, new_new_n15226__, new_new_n15227__,
    new_new_n15228__, new_new_n15229__, new_new_n15230__, new_new_n15231__,
    new_new_n15232__, new_new_n15233__, new_new_n15234__, new_new_n15235__,
    new_new_n15236__, new_new_n15237__, new_new_n15238__, new_new_n15239__,
    new_new_n15240__, new_new_n15241__, new_new_n15242__, new_new_n15243__,
    new_new_n15244__, new_new_n15245__, new_new_n15246__, new_new_n15247__,
    new_new_n15248__, new_new_n15249__, new_new_n15250__, new_new_n15251__,
    new_new_n15252__, new_new_n15253__, new_new_n15254__, new_new_n15255__,
    new_new_n15256__, new_new_n15257__, new_new_n15258__, new_new_n15259__,
    new_new_n15260__, new_new_n15261__, new_new_n15262__, new_new_n15263__,
    new_new_n15264__, new_new_n15265__, new_new_n15266__, new_new_n15267__,
    new_new_n15268__, new_new_n15269__, new_new_n15270__, new_new_n15271__,
    new_new_n15272__, new_new_n15273__, new_new_n15274__, new_new_n15275__,
    new_new_n15276__, new_new_n15277__, new_new_n15278__, new_new_n15279__,
    new_new_n15280__, new_new_n15281__, new_new_n15282__, new_new_n15283__,
    new_new_n15284__, new_new_n15285__, new_new_n15286__, new_new_n15287__,
    new_new_n15288__, new_new_n15289__, new_new_n15290__, new_new_n15291__,
    new_new_n15292__, new_new_n15293__, new_new_n15294__, new_new_n15295__,
    new_new_n15296__, new_new_n15297__, new_new_n15298__, new_new_n15299__,
    new_new_n15300__, new_new_n15301__, new_new_n15302__, new_new_n15303__,
    new_new_n15304__, new_new_n15305__, new_new_n15306__, new_new_n15307__,
    new_new_n15308__, new_new_n15309__, new_new_n15310__, new_new_n15311__,
    new_new_n15312__, new_new_n15313__, new_new_n15314__, new_new_n15315__,
    new_new_n15316__, new_new_n15317__, new_new_n15318__, new_new_n15319__,
    new_new_n15320__, new_new_n15321__, new_new_n15322__, new_new_n15323__,
    new_new_n15324__, new_new_n15325__, new_new_n15326__, new_new_n15327__,
    new_new_n15328__, new_new_n15329__, new_new_n15330__, new_new_n15331__,
    new_new_n15332__, new_new_n15333__, new_new_n15334__, new_new_n15335__,
    new_new_n15336__, new_new_n15337__, new_new_n15338__, new_new_n15339__,
    new_new_n15340__, new_new_n15341__, new_new_n15342__, new_new_n15343__,
    new_new_n15344__, new_new_n15345__, new_new_n15346__, new_new_n15347__,
    new_new_n15348__, new_new_n15349__, new_new_n15350__, new_new_n15351__,
    new_new_n15352__, new_new_n15353__, new_new_n15354__, new_new_n15355__,
    new_new_n15356__, new_new_n15357__, new_new_n15358__, new_new_n15359__,
    new_new_n15360__, new_new_n15361__, new_new_n15362__, new_new_n15363__,
    new_new_n15364__, new_new_n15365__, new_new_n15366__, new_new_n15367__,
    new_new_n15368__, new_new_n15369__, new_new_n15370__, new_new_n15371__,
    new_new_n15372__, new_new_n15373__, new_new_n15374__, new_new_n15375__,
    new_new_n15376__, new_new_n15377__, new_new_n15378__, new_new_n15379__,
    new_new_n15380__, new_new_n15381__, new_new_n15382__, new_new_n15383__,
    new_new_n15384__, new_new_n15385__, new_new_n15386__, new_new_n15387__,
    new_new_n15388__, new_new_n15389__, new_new_n15390__, new_new_n15391__,
    new_new_n15392__, new_new_n15393__, new_new_n15394__, new_new_n15395__,
    new_new_n15396__, new_new_n15397__, new_new_n15398__, new_new_n15399__,
    new_new_n15400__, new_new_n15401__, new_new_n15402__, new_new_n15403__,
    new_new_n15404__, new_new_n15405__, new_new_n15406__, new_new_n15407__,
    new_new_n15408__, new_new_n15409__, new_new_n15410__, new_new_n15411__,
    new_new_n15412__, new_new_n15413__, new_new_n15414__, new_new_n15415__,
    new_new_n15416__, new_new_n15417__, new_new_n15418__, new_new_n15419__,
    new_new_n15420__, new_new_n15421__, new_new_n15422__, new_new_n15423__,
    new_new_n15424__, new_new_n15425__, new_new_n15426__, new_new_n15427__,
    new_new_n15428__, new_new_n15429__, new_new_n15430__, new_new_n15431__,
    new_new_n15432__, new_new_n15433__, new_new_n15434__, new_new_n15435__,
    new_new_n15436__, new_new_n15437__, new_new_n15438__, new_new_n15439__,
    new_new_n15440__, new_new_n15441__, new_new_n15442__, new_new_n15443__,
    new_new_n15444__, new_new_n15445__, new_new_n15446__, new_new_n15447__,
    new_new_n15448__, new_new_n15449__, new_new_n15450__, new_new_n15451__,
    new_new_n15452__, new_new_n15453__, new_new_n15454__, new_new_n15455__,
    new_new_n15456__, new_new_n15457__, new_new_n15458__, new_new_n15459__,
    new_new_n15460__, new_new_n15461__, new_new_n15462__, new_new_n15463__,
    new_new_n15464__, new_new_n15465__, new_new_n15466__, new_new_n15467__,
    new_new_n15468__, new_new_n15469__, new_new_n15470__, new_new_n15471__,
    new_new_n15472__, new_new_n15473__, new_new_n15474__, new_new_n15475__,
    new_new_n15476__, new_new_n15477__, new_new_n15478__, new_new_n15479__,
    new_new_n15480__, new_new_n15481__, new_new_n15482__, new_new_n15483__,
    new_new_n15484__, new_new_n15485__, new_new_n15486__, new_new_n15487__,
    new_new_n15488__, new_new_n15489__, new_new_n15490__, new_new_n15491__,
    new_new_n15492__, new_new_n15493__, new_new_n15494__, new_new_n15495__,
    new_new_n15496__, new_new_n15497__, new_new_n15498__, new_new_n15499__,
    new_new_n15500__, new_new_n15501__, new_new_n15502__, new_new_n15503__,
    new_new_n15504__, new_new_n15505__, new_new_n15506__, new_new_n15507__,
    new_new_n15508__, new_new_n15509__, new_new_n15510__, new_new_n15511__,
    new_new_n15512__, new_new_n15513__, new_new_n15514__, new_new_n15515__,
    new_new_n15516__, new_new_n15517__, new_new_n15518__, new_new_n15519__,
    new_new_n15520__, new_new_n15521__, new_new_n15522__, new_new_n15523__,
    new_new_n15524__, new_new_n15525__, new_new_n15526__, new_new_n15527__,
    new_new_n15528__, new_new_n15529__, new_new_n15530__, new_new_n15531__,
    new_new_n15532__, new_new_n15533__, new_new_n15534__, new_new_n15535__,
    new_new_n15536__, new_new_n15537__, new_new_n15538__, new_new_n15539__,
    new_new_n15540__, new_new_n15541__, new_new_n15542__, new_new_n15543__,
    new_new_n15544__, new_new_n15545__, new_new_n15546__, new_new_n15547__,
    new_new_n15548__, new_new_n15549__, new_new_n15550__, new_new_n15551__,
    new_new_n15552__, new_new_n15553__, new_new_n15554__, new_new_n15555__,
    new_new_n15556__, new_new_n15557__, new_new_n15558__, new_new_n15559__,
    new_new_n15560__, new_new_n15561__, new_new_n15562__, new_new_n15563__,
    new_new_n15564__, new_new_n15565__, new_new_n15566__, new_new_n15567__,
    new_new_n15568__, new_new_n15569__, new_new_n15570__, new_new_n15571__,
    new_new_n15572__, new_new_n15573__, new_new_n15574__, new_new_n15575__,
    new_new_n15576__, new_new_n15577__, new_new_n15578__, new_new_n15579__,
    new_new_n15580__, new_new_n15581__, new_new_n15582__, new_new_n15583__,
    new_new_n15584__, new_new_n15585__, new_new_n15586__, new_new_n15587__,
    new_new_n15588__, new_new_n15589__, new_new_n15590__, new_new_n15591__,
    new_new_n15592__, new_new_n15593__, new_new_n15594__, new_new_n15595__,
    new_new_n15596__, new_new_n15597__, new_new_n15598__, new_new_n15599__,
    new_new_n15600__, new_new_n15601__, new_new_n15602__, new_new_n15603__,
    new_new_n15604__, new_new_n15605__, new_new_n15606__, new_new_n15607__,
    new_new_n15608__, new_new_n15609__, new_new_n15610__, new_new_n15611__,
    new_new_n15612__, new_new_n15613__, new_new_n15614__, new_new_n15615__,
    new_new_n15616__, new_new_n15617__, new_new_n15618__, new_new_n15619__,
    new_new_n15620__, new_new_n15621__, new_new_n15622__, new_new_n15623__,
    new_new_n15624__, new_new_n15625__, new_new_n15626__, new_new_n15627__,
    new_new_n15628__, new_new_n15629__, new_new_n15630__, new_new_n15631__,
    new_new_n15632__, new_new_n15633__, new_new_n15634__, new_new_n15635__,
    new_new_n15636__, new_new_n15637__, new_new_n15638__, new_new_n15639__,
    new_new_n15640__, new_new_n15641__, new_new_n15642__, new_new_n15643__,
    new_new_n15644__, new_new_n15645__, new_new_n15646__, new_new_n15647__,
    new_new_n15648__, new_new_n15649__, new_new_n15650__, new_new_n15651__,
    new_new_n15652__, new_new_n15653__, new_new_n15654__, new_new_n15655__,
    new_new_n15656__, new_new_n15657__, new_new_n15658__, new_new_n15659__,
    new_new_n15660__, new_new_n15661__, new_new_n15662__, new_new_n15663__,
    new_new_n15664__, new_new_n15665__, new_new_n15666__, new_new_n15667__,
    new_new_n15668__, new_new_n15669__, new_new_n15670__, new_new_n15671__,
    new_new_n15672__, new_new_n15673__, new_new_n15674__, new_new_n15675__,
    new_new_n15676__, new_new_n15677__, new_new_n15678__, new_new_n15679__,
    new_new_n15680__, new_new_n15681__, new_new_n15682__, new_new_n15683__,
    new_new_n15684__, new_new_n15685__, new_new_n15686__, new_new_n15687__,
    new_new_n15688__, new_new_n15689__, new_new_n15690__, new_new_n15691__,
    new_new_n15692__, new_new_n15693__, new_new_n15694__, new_new_n15695__,
    new_new_n15696__, new_new_n15697__, new_new_n15698__, new_new_n15699__,
    new_new_n15700__, new_new_n15701__, new_new_n15702__, new_new_n15703__,
    new_new_n15704__, new_new_n15705__, new_new_n15706__, new_new_n15707__,
    new_new_n15708__, new_new_n15709__, new_new_n15710__, new_new_n15711__,
    new_new_n15712__, new_new_n15713__, new_new_n15714__, new_new_n15715__,
    new_new_n15716__, new_new_n15717__, new_new_n15718__, new_new_n15719__,
    new_new_n15720__, new_new_n15721__, new_new_n15722__, new_new_n15723__,
    new_new_n15724__, new_new_n15725__, new_new_n15726__, new_new_n15727__,
    new_new_n15728__, new_new_n15729__, new_new_n15730__, new_new_n15731__,
    new_new_n15732__, new_new_n15733__, new_new_n15734__, new_new_n15735__,
    new_new_n15736__, new_new_n15737__, new_new_n15738__, new_new_n15739__,
    new_new_n15740__, new_new_n15741__, new_new_n15742__, new_new_n15743__,
    new_new_n15744__, new_new_n15745__, new_new_n15746__, new_new_n15747__,
    new_new_n15748__, new_new_n15749__, new_new_n15750__, new_new_n15751__,
    new_new_n15752__, new_new_n15753__, new_new_n15754__, new_new_n15755__,
    new_new_n15756__, new_new_n15757__, new_new_n15758__, new_new_n15759__,
    new_new_n15760__, new_new_n15761__, new_new_n15762__, new_new_n15763__,
    new_new_n15764__, new_new_n15765__, new_new_n15766__, new_new_n15767__,
    new_new_n15768__, new_new_n15769__, new_new_n15770__, new_new_n15771__,
    new_new_n15772__, new_new_n15773__, new_new_n15774__, new_new_n15775__,
    new_new_n15776__, new_new_n15777__, new_new_n15778__, new_new_n15779__,
    new_new_n15780__, new_new_n15781__, new_new_n15782__, new_new_n15783__,
    new_new_n15784__, new_new_n15785__, new_new_n15786__, new_new_n15787__,
    new_new_n15788__, new_new_n15789__, new_new_n15790__, new_new_n15791__,
    new_new_n15792__, new_new_n15793__, new_new_n15794__, new_new_n15795__,
    new_new_n15796__, new_new_n15797__, new_new_n15798__, new_new_n15799__,
    new_new_n15800__, new_new_n15801__, new_new_n15802__, new_new_n15803__,
    new_new_n15804__, new_new_n15805__, new_new_n15806__, new_new_n15807__,
    new_new_n15808__, new_new_n15809__, new_new_n15810__, new_new_n15811__,
    new_new_n15812__, new_new_n15813__, new_new_n15814__, new_new_n15815__,
    new_new_n15816__, new_new_n15817__, new_new_n15818__, new_new_n15819__,
    new_new_n15820__, new_new_n15821__, new_new_n15822__, new_new_n15823__,
    new_new_n15824__, new_new_n15825__, new_new_n15826__, new_new_n15827__,
    new_new_n15828__, new_new_n15829__, new_new_n15830__, new_new_n15831__,
    new_new_n15832__, new_new_n15833__, new_new_n15834__, new_new_n15835__,
    new_new_n15836__, new_new_n15837__, new_new_n15838__, new_new_n15839__,
    new_new_n15840__, new_new_n15841__, new_new_n15842__, new_new_n15843__,
    new_new_n15844__, new_new_n15845__, new_new_n15847__, new_new_n15848__,
    new_new_n15849__, new_new_n15850__, new_new_n15852__, new_new_n15853__,
    new_new_n15854__, new_new_n15855__, new_new_n15856__, new_new_n15857__,
    new_new_n15859__, new_new_n15861__, new_new_n15862__, new_new_n15863__,
    new_new_n15864__, new_new_n15865__, new_new_n15867__, new_new_n15868__,
    new_new_n15869__, new_new_n15870__, new_new_n15872__, new_new_n15873__,
    new_new_n15874__, new_new_n15875__, new_new_n15877__, new_new_n15878__,
    new_new_n15879__, new_new_n15880__, new_new_n15881__, new_new_n15882__,
    new_new_n15884__, new_new_n15886__, new_new_n15887__, new_new_n15888__,
    new_new_n15889__, new_new_n15890__, new_new_n15892__, new_new_n15893__,
    new_new_n15894__, new_new_n15895__, new_new_n15897__, new_new_n15898__,
    new_new_n15900__, new_new_n15901__, new_new_n15902__, new_new_n15903__,
    new_new_n15904__, new_new_n15905__, new_new_n15906__, new_new_n15907__,
    new_new_n15908__, new_new_n15909__, new_new_n15910__, new_new_n15911__,
    new_new_n15912__, new_new_n15913__, new_new_n15914__, new_new_n15915__,
    new_new_n15916__, new_new_n15917__, new_new_n15918__, new_new_n15919__,
    new_new_n15920__, new_new_n15921__, new_new_n15922__, new_new_n15923__,
    new_new_n15924__, new_new_n15925__, new_new_n15926__, new_new_n15927__,
    new_new_n15928__, new_new_n15929__, new_new_n15930__, new_new_n15931__,
    new_new_n15932__, new_new_n15933__, new_new_n15934__, new_new_n15935__,
    new_new_n15936__, new_new_n15937__, new_new_n15938__, new_new_n15939__,
    new_new_n15940__, new_new_n15941__, new_new_n15942__, new_new_n15943__,
    new_new_n15944__, new_new_n15945__, new_new_n15946__, new_new_n15947__,
    new_new_n15948__, new_new_n15949__, new_new_n15950__, new_new_n15951__,
    new_new_n15952__, new_new_n15956__, new_new_n15957__, new_new_n15958__,
    new_new_n15959__, new_new_n15960__, new_new_n15961__, new_new_n15962__,
    new_new_n15963__, new_new_n15964__, new_new_n15965__, new_new_n15966__,
    new_new_n15967__, new_new_n15968__, new_new_n15969__, new_new_n15970__,
    new_new_n15971__, new_new_n15972__, new_new_n15973__, new_new_n15974__,
    new_new_n15975__, new_new_n15976__, new_new_n15977__, new_new_n15978__,
    new_new_n15980__, new_new_n15981__, new_new_n15982__, new_new_n15983__,
    new_new_n15984__, new_new_n15985__, new_new_n15986__, new_new_n15987__,
    new_new_n15988__, new_new_n15989__, new_new_n15990__, new_new_n15991__,
    new_new_n15992__, new_new_n15993__, new_new_n15994__, new_new_n15995__,
    new_new_n15997__, new_new_n15998__, new_new_n15999__, new_new_n16000__,
    new_new_n16001__, new_new_n16002__, new_new_n16003__, new_new_n16004__,
    new_new_n16005__, new_new_n16006__, new_new_n16007__, new_new_n16008__,
    new_new_n16009__, new_new_n16010__, new_new_n16011__, new_new_n16012__,
    new_new_n16013__, new_new_n16014__, new_new_n16015__, new_new_n16016__,
    new_new_n16017__, new_new_n16018__, new_new_n16019__, new_new_n16020__,
    new_new_n16021__, new_new_n16022__, new_new_n16023__, new_new_n16024__,
    new_new_n16025__, new_new_n16026__, new_new_n16027__, new_new_n16028__,
    new_new_n16029__, new_new_n16030__, new_new_n16032__, new_new_n16033__,
    new_new_n16034__, new_new_n16035__, new_new_n16036__, new_new_n16037__,
    new_new_n16038__, new_new_n16039__, new_new_n16040__, new_new_n16041__,
    new_new_n16042__, new_new_n16043__, new_new_n16044__, new_new_n16045__,
    new_new_n16046__, new_new_n16047__, new_new_n16048__, new_new_n16049__,
    new_new_n16050__, new_new_n16051__, new_new_n16052__, new_new_n16053__,
    new_new_n16054__, new_new_n16055__, new_new_n16056__, new_new_n16057__,
    new_new_n16058__, new_new_n16059__, new_new_n16060__, new_new_n16061__,
    new_new_n16062__, new_new_n16063__, new_new_n16064__, new_new_n16065__,
    new_new_n16066__, new_new_n16067__, new_new_n16068__, new_new_n16069__,
    new_new_n16070__, new_new_n16071__, new_new_n16072__, new_new_n16073__,
    new_new_n16074__, new_new_n16075__, new_new_n16076__, new_new_n16077__,
    new_new_n16078__, new_new_n16079__, new_new_n16080__, new_new_n16081__,
    new_new_n16082__, new_new_n16083__, new_new_n16084__, new_new_n16085__,
    new_new_n16086__, new_new_n16087__, new_new_n16088__, new_new_n16089__,
    new_new_n16090__, new_new_n16091__, new_new_n16092__, new_new_n16093__,
    new_new_n16094__, new_new_n16095__, new_new_n16096__, new_new_n16097__,
    new_new_n16098__, new_new_n16099__, new_new_n16100__, new_new_n16101__,
    new_new_n16102__, new_new_n16103__, new_new_n16104__, new_new_n16105__,
    new_new_n16106__, new_new_n16107__, new_new_n16108__, new_new_n16109__,
    new_new_n16110__, new_new_n16111__, new_new_n16112__, new_new_n16113__,
    new_new_n16114__, new_new_n16115__, new_new_n16116__, new_new_n16117__,
    new_new_n16118__, new_new_n16119__, new_new_n16120__, new_new_n16121__,
    new_new_n16122__, new_new_n16123__, new_new_n16124__, new_new_n16125__,
    new_new_n16126__, new_new_n16127__, new_new_n16128__, new_new_n16129__,
    new_new_n16130__, new_new_n16131__, new_new_n16132__, new_new_n16133__,
    new_new_n16134__, new_new_n16135__, new_new_n16136__, new_new_n16137__,
    new_new_n16138__, new_new_n16139__, new_new_n16140__, new_new_n16141__,
    new_new_n16142__, new_new_n16143__, new_new_n16144__, new_new_n16145__,
    new_new_n16146__, new_new_n16147__, new_new_n16148__, new_new_n16149__,
    new_new_n16150__, new_new_n16151__, new_new_n16152__, new_new_n16153__,
    new_new_n16154__, new_new_n16155__, new_new_n16156__, new_new_n16157__,
    new_new_n16158__, new_new_n16159__, new_new_n16160__, new_new_n16161__,
    new_new_n16162__, new_new_n16163__, new_new_n16164__, new_new_n16165__,
    new_new_n16166__, new_new_n16167__, new_new_n16168__, new_new_n16169__,
    new_new_n16170__, new_new_n16171__, new_new_n16172__, new_new_n16173__,
    new_new_n16174__, new_new_n16175__, new_new_n16176__, new_new_n16177__,
    new_new_n16178__, new_new_n16179__, new_new_n16180__, new_new_n16181__,
    new_new_n16182__, new_new_n16183__, new_new_n16184__, new_new_n16185__,
    new_new_n16186__, new_new_n16187__, new_new_n16188__, new_new_n16189__,
    new_new_n16190__, new_new_n16191__, new_new_n16192__, new_new_n16193__,
    new_new_n16194__, new_new_n16195__, new_new_n16196__, new_new_n16197__,
    new_new_n16198__, new_new_n16199__, new_new_n16200__, new_new_n16201__,
    new_new_n16202__, new_new_n16203__, new_new_n16204__, new_new_n16205__,
    new_new_n16206__, new_new_n16207__, new_new_n16208__, new_new_n16209__,
    new_new_n16210__, new_new_n16211__, new_new_n16212__, new_new_n16213__,
    new_new_n16214__, new_new_n16215__, new_new_n16216__, new_new_n16217__,
    new_new_n16218__, new_new_n16219__, new_new_n16220__, new_new_n16221__,
    new_new_n16222__, new_new_n16223__, new_new_n16225__, new_new_n16226__,
    new_new_n16227__, new_new_n16230__, new_new_n16231__, new_new_n16234__,
    new_new_n16235__, new_new_n16236__, new_new_n16238__, new_new_n16239__,
    new_new_n16240__, new_new_n16241__, new_new_n16243__, new_new_n16244__,
    new_new_n16245__, new_new_n16246__, new_new_n16247__, new_new_n16248__,
    new_new_n16250__, new_new_n16251__, new_new_n16252__, new_new_n16253__,
    new_new_n16254__, new_new_n16256__, new_new_n16257__, new_new_n16258__,
    new_new_n16259__, new_new_n16260__, new_new_n16261__, new_new_n16263__,
    new_new_n16264__, new_new_n16265__, new_new_n16267__, new_new_n16268__,
    new_new_n16271__, new_new_n16272__, new_new_n16273__, new_new_n16275__,
    new_new_n16276__, new_new_n16277__, new_new_n16278__, new_new_n16279__,
    new_new_n16281__, new_new_n16282__, new_new_n16283__, new_new_n16284__,
    new_new_n16285__, new_new_n16287__, new_new_n16288__, new_new_n16289__,
    new_new_n16290__, new_new_n16291__, new_new_n16293__, new_new_n16294__,
    new_new_n16295__, new_new_n16296__, new_new_n16297__, new_new_n16299__,
    new_new_n16300__, new_new_n16301__, new_new_n16302__, new_new_n16303__,
    new_new_n16305__, new_new_n16306__, new_new_n16307__, new_new_n16308__,
    new_new_n16309__, new_new_n16311__, new_new_n16312__, new_new_n16313__,
    new_new_n16314__, new_new_n16315__, new_new_n16317__, new_new_n16318__,
    new_new_n16319__, new_new_n16320__, new_new_n16321__, new_new_n16323__,
    new_new_n16324__, new_new_n16325__, new_new_n16326__, new_new_n16327__,
    new_new_n16329__, new_new_n16330__, new_new_n16331__, new_new_n16332__,
    new_new_n16333__, new_new_n16335__, new_new_n16336__, new_new_n16337__,
    new_new_n16338__, new_new_n16339__, new_new_n16341__, new_new_n16342__,
    new_new_n16343__, new_new_n16344__, new_new_n16345__, new_new_n16347__,
    new_new_n16348__, new_new_n16349__, new_new_n16350__, new_new_n16351__,
    new_new_n16353__, new_new_n16354__, new_new_n16355__, new_new_n16356__,
    new_new_n16357__, new_new_n16359__, new_new_n16360__, new_new_n16361__,
    new_new_n16362__, new_new_n16363__, new_new_n16365__, new_new_n16366__,
    new_new_n16367__, new_new_n16368__, new_new_n16369__, new_new_n16371__,
    new_new_n16372__, new_new_n16373__, new_new_n16374__, new_new_n16375__,
    new_new_n16377__, new_new_n16378__, new_new_n16379__, new_new_n16380__,
    new_new_n16381__, new_new_n16383__, new_new_n16384__, new_new_n16385__,
    new_new_n16386__, new_new_n16387__, new_new_n16389__, new_new_n16390__,
    new_new_n16391__, new_new_n16392__, new_new_n16393__, new_new_n16395__,
    new_new_n16396__, new_new_n16397__, new_new_n16398__, new_new_n16399__,
    new_new_n16401__, new_new_n16402__, new_new_n16403__, new_new_n16404__,
    new_new_n16405__, new_new_n16407__, new_new_n16408__, new_new_n16409__,
    new_new_n16410__, new_new_n16411__, new_new_n16413__, new_new_n16414__,
    new_new_n16415__, new_new_n16416__, new_new_n16417__, new_new_n16419__,
    new_new_n16420__, new_new_n16421__, new_new_n16422__, new_new_n16423__,
    new_new_n16425__, new_new_n16426__, new_new_n16427__, new_new_n16428__,
    new_new_n16429__, new_new_n16431__, new_new_n16432__, new_new_n16433__,
    new_new_n16434__, new_new_n16435__, new_new_n16437__, new_new_n16438__,
    new_new_n16439__, new_new_n16440__, new_new_n16441__, new_new_n16443__,
    new_new_n16444__, new_new_n16445__, new_new_n16446__, new_new_n16448__,
    new_new_n16449__, new_new_n16450__, new_new_n16451__, new_new_n16453__,
    new_new_n16454__, new_new_n16455__, new_new_n16456__, new_new_n16458__,
    new_new_n16460__, new_new_n16461__, new_new_n16463__, new_new_n16464__,
    new_new_n16466__, new_new_n16468__, new_new_n16469__, new_new_n16471__,
    new_new_n16472__, new_new_n16474__, new_new_n16476__, new_new_n16477__,
    new_new_n16479__, new_new_n16480__, new_new_n16482__, new_new_n16483__,
    new_new_n16484__, new_new_n16485__, new_new_n16486__, new_new_n16488__,
    new_new_n16490__, new_new_n16491__, new_new_n16492__, new_new_n16493__,
    new_new_n16494__, new_new_n16496__, new_new_n16497__, new_new_n16498__,
    new_new_n16499__, new_new_n16500__, new_new_n16502__, new_new_n16503__,
    new_new_n16505__, new_new_n16506__, new_new_n16507__, new_new_n16508__,
    new_new_n16509__, new_new_n16510__, new_new_n16511__, new_new_n16512__,
    new_new_n16513__, new_new_n16514__, new_new_n16516__, new_new_n16517__,
    new_new_n16518__, new_new_n16520__, new_new_n16521__, new_new_n16522__,
    new_new_n16523__, new_new_n16524__, new_new_n16525__, new_new_n16526__,
    new_new_n16527__, new_new_n16528__, new_new_n16530__, new_new_n16531__,
    new_new_n16532__, new_new_n16533__, new_new_n16534__, new_new_n16535__,
    new_new_n16538__, new_new_n16539__, new_new_n16540__, new_new_n16541__,
    new_new_n16542__, new_new_n16546__, new_new_n16547__, new_new_n16548__,
    new_new_n16550__, new_new_n16551__, new_new_n16552__, new_new_n16554__,
    new_new_n16555__, new_new_n16556__, new_new_n16557__, new_new_n16558__,
    new_new_n16559__, new_new_n16560__, new_new_n16561__, new_new_n16562__,
    new_new_n16563__, new_new_n16564__, new_new_n16565__, new_new_n16566__,
    new_new_n16568__, new_new_n16569__, new_new_n16570__, new_new_n16571__,
    new_new_n16572__, new_new_n16573__, new_new_n16574__, new_new_n16575__,
    new_new_n16576__, new_new_n16577__, new_new_n16578__, new_new_n16579__,
    new_new_n16580__, new_new_n16581__, new_new_n16582__, new_new_n16583__,
    new_new_n16584__, new_new_n16585__, new_new_n16586__, new_new_n16587__,
    new_new_n16588__, new_new_n16589__, new_new_n16590__, new_new_n16591__,
    new_new_n16592__, new_new_n16593__, new_new_n16594__, new_new_n16595__,
    new_new_n16596__, new_new_n16597__, new_new_n16598__, new_new_n16599__,
    new_new_n16601__, new_new_n16602__, new_new_n16603__, new_new_n16604__,
    new_new_n16605__, new_new_n16606__, new_new_n16608__, new_new_n16609__,
    new_new_n16610__, new_new_n16611__, new_new_n16612__, new_new_n16613__,
    new_new_n16614__, new_new_n16615__, new_new_n16616__, new_new_n16617__,
    new_new_n16618__, new_new_n16619__, new_new_n16620__, new_new_n16621__,
    new_new_n16622__, new_new_n16623__, new_new_n16624__, new_new_n16625__,
    new_new_n16626__, new_new_n16627__, new_new_n16629__, new_new_n16630__,
    new_new_n16631__, new_new_n16632__, new_new_n16633__, new_new_n16634__,
    new_new_n16637__, new_new_n16638__, new_new_n16639__, new_new_n16641__,
    new_new_n16642__, new_new_n16643__, new_new_n16644__, new_new_n16645__,
    new_new_n16646__, new_new_n16647__, new_new_n16648__, new_new_n16649__,
    new_new_n16650__, new_new_n16651__, new_new_n16652__, new_new_n16653__,
    new_new_n16654__, new_new_n16655__, new_new_n16656__, new_new_n16657__,
    new_new_n16658__, new_new_n16659__, new_new_n16660__, new_new_n16661__,
    new_new_n16662__, new_new_n16663__, new_new_n16664__, new_new_n16665__,
    new_new_n16666__, new_new_n16667__, new_new_n16668__, new_new_n16669__,
    new_new_n16670__, new_new_n16671__, new_new_n16672__, new_new_n16673__,
    new_new_n16674__, new_new_n16675__, new_new_n16676__, new_new_n16677__,
    new_new_n16678__, new_new_n16679__, new_new_n16680__, new_new_n16681__,
    new_new_n16682__, new_new_n16683__, new_new_n16684__, new_new_n16685__,
    new_new_n16686__, new_new_n16687__, new_new_n16688__, new_new_n16689__,
    new_new_n16690__, new_new_n16691__, new_new_n16692__, new_new_n16693__,
    new_new_n16694__, new_new_n16695__, new_new_n16696__, new_new_n16697__,
    new_new_n16698__, new_new_n16699__, new_new_n16700__, new_new_n16701__,
    new_new_n16702__, new_new_n16703__, new_new_n16705__, new_new_n16706__,
    new_new_n16707__, new_new_n16710__, new_new_n16711__, new_new_n16712__,
    new_new_n16713__, new_new_n16714__, new_new_n16715__, new_new_n16717__,
    new_new_n16718__, new_new_n16719__, new_new_n16721__, new_new_n16722__,
    new_new_n16723__, new_new_n16724__, new_new_n16726__, new_new_n16727__,
    new_new_n16728__, new_new_n16731__, new_new_n16732__, new_new_n16733__,
    new_new_n16734__, new_new_n16735__, new_new_n16736__, new_new_n16737__,
    new_new_n16738__, new_new_n16739__, new_new_n16740__, new_new_n16741__,
    new_new_n16742__, new_new_n16743__, new_new_n16744__, new_new_n16745__,
    new_new_n16746__, new_new_n16747__, new_new_n16748__, new_new_n16749__,
    new_new_n16750__, new_new_n16751__, new_new_n16752__, new_new_n16753__,
    new_new_n16754__, new_new_n16755__, new_new_n16756__, new_new_n16757__,
    new_new_n16758__, new_new_n16759__, new_new_n16760__, new_new_n16761__,
    new_new_n16762__, new_new_n16763__, new_new_n16764__, new_new_n16765__,
    new_new_n16766__, new_new_n16767__, new_new_n16768__, new_new_n16769__,
    new_new_n16770__, new_new_n16771__, new_new_n16772__, new_new_n16773__,
    new_new_n16774__, new_new_n16775__, new_new_n16776__, new_new_n16777__,
    new_new_n16778__, new_new_n16779__, new_new_n16780__, new_new_n16781__,
    new_new_n16782__, new_new_n16783__, new_new_n16784__, new_new_n16785__,
    new_new_n16786__, new_new_n16787__, new_new_n16788__, new_new_n16789__,
    new_new_n16790__, new_new_n16791__, new_new_n16792__, new_new_n16793__,
    new_new_n16794__, new_new_n16795__, new_new_n16796__, new_new_n16797__,
    new_new_n16798__, new_new_n16799__, new_new_n16800__, new_new_n16801__,
    new_new_n16802__, new_new_n16803__, new_new_n16804__, new_new_n16805__,
    new_new_n16806__, new_new_n16807__, new_new_n16808__, new_new_n16809__,
    new_new_n16810__, new_new_n16811__, new_new_n16812__, new_new_n16813__,
    new_new_n16814__, new_new_n16815__, new_new_n16816__, new_new_n16817__,
    new_new_n16818__, new_new_n16819__, new_new_n16820__, new_new_n16821__,
    new_new_n16822__, new_new_n16823__, new_new_n16824__, new_new_n16825__,
    new_new_n16826__, new_new_n16827__, new_new_n16828__, new_new_n16829__,
    new_new_n16830__, new_new_n16831__, new_new_n16832__, new_new_n16833__,
    new_new_n16834__, new_new_n16835__, new_new_n16836__, new_new_n16837__,
    new_new_n16838__, new_new_n16839__, new_new_n16840__, new_new_n16841__,
    new_new_n16842__, new_new_n16844__, new_new_n16845__, new_new_n16846__,
    new_new_n16847__, new_new_n16848__, new_new_n16849__, new_new_n16850__,
    new_new_n16851__, new_new_n16852__, new_new_n16853__, new_new_n16856__,
    new_new_n16857__, new_new_n16858__, new_new_n16859__, new_new_n16860__,
    new_new_n16861__, new_new_n16862__, new_new_n16865__, new_new_n16866__,
    new_new_n16867__, new_new_n16869__, new_new_n16870__, new_new_n16871__,
    new_new_n16872__, new_new_n16873__, new_new_n16874__, new_new_n16875__,
    new_new_n16876__, new_new_n16877__, new_new_n16878__, new_new_n16879__,
    new_new_n16880__, new_new_n16882__, new_new_n16883__, new_new_n16885__,
    new_new_n16886__, new_new_n16888__, new_new_n16889__, new_new_n16890__,
    new_new_n16891__, new_new_n16892__, new_new_n16893__, new_new_n16894__,
    new_new_n16895__, new_new_n16896__, new_new_n16897__, new_new_n16899__,
    new_new_n16900__, new_new_n16901__, new_new_n16903__, new_new_n16904__,
    new_new_n16905__, new_new_n16906__, new_new_n16907__, new_new_n16908__,
    new_new_n16909__, new_new_n16910__, new_new_n16911__, new_new_n16912__,
    new_new_n16914__, new_new_n16915__, new_new_n16916__, new_new_n16918__,
    new_new_n16921__, new_new_n16922__, new_new_n16923__, new_new_n16924__,
    new_new_n16925__, new_new_n16927__, new_new_n16928__, new_new_n16929__,
    new_new_n16930__, new_new_n16931__, new_new_n16932__, new_new_n16934__,
    new_new_n16935__, new_new_n16937__, new_new_n16938__, new_new_n16939__,
    new_new_n16941__, new_new_n16942__, new_new_n16943__, new_new_n16945__,
    new_new_n16946__, new_new_n16947__, new_new_n16949__, new_new_n16950__,
    new_new_n16951__, new_new_n16953__, new_new_n16954__, new_new_n16955__,
    new_new_n16957__, new_new_n16958__, new_new_n16959__, new_new_n16961__,
    new_new_n16962__, new_new_n16963__, new_new_n16965__, new_new_n16966__,
    new_new_n16967__, new_new_n16969__, new_new_n16970__, new_new_n16971__,
    new_new_n16973__, new_new_n16974__, new_new_n16975__, new_new_n16977__,
    new_new_n16978__, new_new_n16979__, new_new_n16981__, new_new_n16982__,
    new_new_n16983__, new_new_n16985__, new_new_n16986__, new_new_n16987__,
    new_new_n16989__, new_new_n16990__, new_new_n16991__, new_new_n16993__,
    new_new_n16994__, new_new_n16995__, new_new_n16996__, new_new_n16997__,
    new_new_n16998__, new_new_n16999__, new_new_n17000__, new_new_n17001__,
    new_new_n17002__, new_new_n17003__, new_new_n17004__, new_new_n17005__,
    new_new_n17006__, new_new_n17007__, new_new_n17008__, new_new_n17009__,
    new_new_n17010__, new_new_n17011__, new_new_n17013__, new_new_n17015__,
    new_new_n17016__, new_new_n17017__, new_new_n17018__, new_new_n17019__,
    new_new_n17020__, new_new_n17021__, new_new_n17022__, new_new_n17023__,
    new_new_n17024__, new_new_n17025__, new_new_n17027__, new_new_n17029__,
    new_new_n17030__, new_new_n17031__, new_new_n17033__, new_new_n17034__,
    new_new_n17035__, new_new_n17036__, new_new_n17037__, new_new_n17039__,
    new_new_n17041__, new_new_n17042__, new_new_n17043__, new_new_n17044__,
    new_new_n17045__, new_new_n17046__, new_new_n17047__, new_new_n17049__,
    new_new_n17051__, new_new_n17052__, new_new_n17053__, new_new_n17055__,
    new_new_n17056__, new_new_n17057__, new_new_n17058__, new_new_n17059__,
    new_new_n17060__, new_new_n17061__, new_new_n17063__, new_new_n17065__,
    new_new_n17066__, new_new_n17067__, new_new_n17069__, new_new_n17070__,
    new_new_n17071__, new_new_n17072__, new_new_n17073__, new_new_n17074__,
    new_new_n17075__, new_new_n17077__, new_new_n17078__, new_new_n17079__,
    new_new_n17080__, new_new_n17081__, new_new_n17082__, new_new_n17083__,
    new_new_n17084__, new_new_n17085__, new_new_n17086__, new_new_n17087__,
    new_new_n17088__, new_new_n17089__, new_new_n17090__, new_new_n17092__,
    new_new_n17093__, new_new_n17095__, new_new_n17096__, new_new_n17097__,
    new_new_n17099__, new_new_n17100__, new_new_n17101__, new_new_n17102__,
    new_new_n17104__, new_new_n17105__, new_new_n17106__, new_new_n17107__,
    new_new_n17108__, new_new_n17109__, new_new_n17110__, new_new_n17112__,
    new_new_n17114__, new_new_n17115__, new_new_n17116__, new_new_n17118__,
    new_new_n17119__, new_new_n17120__, new_new_n17121__, new_new_n17123__,
    new_new_n17124__, new_new_n17126__, new_new_n17127__, new_new_n17128__,
    new_new_n17129__, new_new_n17131__, new_new_n17132__, new_new_n17133__,
    new_new_n17134__, new_new_n17135__, new_new_n17136__, new_new_n17137__,
    new_new_n17139__, new_new_n17141__, new_new_n17142__, new_new_n17143__,
    new_new_n17145__, new_new_n17146__, new_new_n17147__, new_new_n17148__,
    new_new_n17150__, new_new_n17151__, new_new_n17153__, new_new_n17154__,
    new_new_n17155__, new_new_n17156__, new_new_n17158__, new_new_n17159__,
    new_new_n17160__, new_new_n17161__, new_new_n17162__, new_new_n17163__,
    new_new_n17164__, new_new_n17165__, new_new_n17167__, new_new_n17169__,
    new_new_n17170__, new_new_n17171__, new_new_n17172__, new_new_n17173__,
    new_new_n17174__, new_new_n17175__, new_new_n17177__, new_new_n17178__,
    new_new_n17179__, new_new_n17180__, new_new_n17182__, new_new_n17183__,
    new_new_n17185__, new_new_n17186__, new_new_n17187__, new_new_n17188__,
    new_new_n17190__, new_new_n17191__, new_new_n17192__, new_new_n17193__,
    new_new_n17194__, new_new_n17195__, new_new_n17196__, new_new_n17198__,
    new_new_n17200__, new_new_n17201__, new_new_n17202__, new_new_n17203__,
    new_new_n17204__, new_new_n17205__, new_new_n17207__, new_new_n17208__,
    new_new_n17209__, new_new_n17210__, new_new_n17212__, new_new_n17213__,
    new_new_n17215__, new_new_n17216__, new_new_n17217__, new_new_n17218__,
    new_new_n17220__, new_new_n17221__, new_new_n17222__, new_new_n17223__,
    new_new_n17224__, new_new_n17225__, new_new_n17227__, new_new_n17229__,
    new_new_n17230__, new_new_n17231__, new_new_n17232__, new_new_n17233__,
    new_new_n17235__, new_new_n17236__, new_new_n17237__, new_new_n17238__,
    new_new_n17240__, new_new_n17241__, new_new_n17243__, new_new_n17244__,
    new_new_n17245__, new_new_n17246__, new_new_n17248__, new_new_n17249__,
    new_new_n17250__, new_new_n17251__, new_new_n17252__, new_new_n17253__,
    new_new_n17255__, new_new_n17257__, new_new_n17258__, new_new_n17259__,
    new_new_n17260__, new_new_n17261__, new_new_n17263__, new_new_n17264__,
    new_new_n17265__, new_new_n17266__, new_new_n17268__, new_new_n17269__,
    new_new_n17271__, new_new_n17272__, new_new_n17273__, new_new_n17274__,
    new_new_n17276__, new_new_n17277__, new_new_n17278__, new_new_n17279__,
    new_new_n17280__, new_new_n17281__, new_new_n17283__, new_new_n17285__,
    new_new_n17286__, new_new_n17287__, new_new_n17288__, new_new_n17289__,
    new_new_n17291__, new_new_n17292__, new_new_n17293__, new_new_n17294__,
    new_new_n17296__, new_new_n17297__, new_new_n17299__, new_new_n17300__,
    new_new_n17301__, new_new_n17302__, new_new_n17304__, new_new_n17305__,
    new_new_n17306__, new_new_n17307__, new_new_n17308__, new_new_n17309__,
    new_new_n17311__, new_new_n17313__, new_new_n17314__, new_new_n17315__,
    new_new_n17316__, new_new_n17317__, new_new_n17319__, new_new_n17320__,
    new_new_n17321__, new_new_n17322__, new_new_n17324__, new_new_n17325__,
    new_new_n17327__, new_new_n17328__, new_new_n17329__, new_new_n17330__,
    new_new_n17332__, new_new_n17333__, new_new_n17334__, new_new_n17335__,
    new_new_n17336__, new_new_n17337__, new_new_n17339__, new_new_n17341__,
    new_new_n17342__, new_new_n17343__, new_new_n17344__, new_new_n17345__,
    new_new_n17347__, new_new_n17348__, new_new_n17349__, new_new_n17350__,
    new_new_n17352__, new_new_n17353__, new_new_n17355__, new_new_n17356__,
    new_new_n17357__, new_new_n17358__, new_new_n17360__, new_new_n17361__,
    new_new_n17362__, new_new_n17363__, new_new_n17364__, new_new_n17365__,
    new_new_n17367__, new_new_n17369__, new_new_n17370__, new_new_n17371__,
    new_new_n17372__, new_new_n17373__, new_new_n17375__, new_new_n17376__,
    new_new_n17377__, new_new_n17378__, new_new_n17380__, new_new_n17381__,
    new_new_n17383__, new_new_n17384__, new_new_n17385__, new_new_n17386__,
    new_new_n17388__, new_new_n17389__, new_new_n17390__, new_new_n17391__,
    new_new_n17392__, new_new_n17393__, new_new_n17395__, new_new_n17397__,
    new_new_n17398__, new_new_n17399__, new_new_n17400__, new_new_n17401__,
    new_new_n17403__, new_new_n17404__, new_new_n17405__, new_new_n17406__,
    new_new_n17408__, new_new_n17409__, new_new_n17411__, new_new_n17412__,
    new_new_n17413__, new_new_n17414__, new_new_n17416__, new_new_n17417__,
    new_new_n17418__, new_new_n17419__, new_new_n17420__, new_new_n17421__,
    new_new_n17423__, new_new_n17425__, new_new_n17426__, new_new_n17427__,
    new_new_n17428__, new_new_n17429__, new_new_n17431__, new_new_n17432__,
    new_new_n17433__, new_new_n17434__, new_new_n17436__, new_new_n17437__,
    new_new_n17439__, new_new_n17440__, new_new_n17441__, new_new_n17442__,
    new_new_n17444__, new_new_n17445__, new_new_n17446__, new_new_n17447__,
    new_new_n17448__, new_new_n17449__, new_new_n17451__, new_new_n17453__,
    new_new_n17454__, new_new_n17455__, new_new_n17456__, new_new_n17457__,
    new_new_n17459__, new_new_n17460__, new_new_n17461__, new_new_n17462__,
    new_new_n17464__, new_new_n17465__, new_new_n17467__, new_new_n17468__,
    new_new_n17469__, new_new_n17470__, new_new_n17472__, new_new_n17473__,
    new_new_n17474__, new_new_n17475__, new_new_n17476__, new_new_n17477__,
    new_new_n17479__, new_new_n17481__, new_new_n17482__, new_new_n17483__,
    new_new_n17484__, new_new_n17485__, new_new_n17487__, new_new_n17488__,
    new_new_n17489__, new_new_n17490__, new_new_n17492__, new_new_n17493__,
    new_new_n17495__, new_new_n17496__, new_new_n17497__, new_new_n17498__,
    new_new_n17500__, new_new_n17501__, new_new_n17502__, new_new_n17503__,
    new_new_n17504__, new_new_n17505__, new_new_n17507__, new_new_n17509__,
    new_new_n17510__, new_new_n17511__, new_new_n17512__, new_new_n17513__,
    new_new_n17515__, new_new_n17516__, new_new_n17517__, new_new_n17518__,
    new_new_n17520__, new_new_n17521__, new_new_n17523__, new_new_n17524__,
    new_new_n17525__, new_new_n17526__, new_new_n17528__, new_new_n17529__,
    new_new_n17530__, new_new_n17531__, new_new_n17532__, new_new_n17533__,
    new_new_n17535__, new_new_n17537__, new_new_n17538__, new_new_n17539__,
    new_new_n17540__, new_new_n17541__, new_new_n17543__, new_new_n17544__,
    new_new_n17545__, new_new_n17546__, new_new_n17548__, new_new_n17549__,
    new_new_n17551__, new_new_n17552__, new_new_n17553__, new_new_n17554__,
    new_new_n17556__, new_new_n17557__, new_new_n17558__, new_new_n17559__,
    new_new_n17560__, new_new_n17561__, new_new_n17563__, new_new_n17565__,
    new_new_n17566__, new_new_n17567__, new_new_n17568__, new_new_n17569__,
    new_new_n17571__, new_new_n17572__, new_new_n17573__, new_new_n17574__,
    new_new_n17576__, new_new_n17577__, new_new_n17579__, new_new_n17580__,
    new_new_n17581__, new_new_n17582__, new_new_n17584__, new_new_n17585__,
    new_new_n17586__, new_new_n17587__, new_new_n17588__, new_new_n17589__,
    new_new_n17591__, new_new_n17593__, new_new_n17594__, new_new_n17595__,
    new_new_n17596__, new_new_n17597__, new_new_n17599__, new_new_n17600__,
    new_new_n17601__, new_new_n17602__, new_new_n17604__, new_new_n17605__,
    new_new_n17607__, new_new_n17608__, new_new_n17609__, new_new_n17610__,
    new_new_n17612__, new_new_n17613__, new_new_n17614__, new_new_n17615__,
    new_new_n17616__, new_new_n17617__, new_new_n17619__, new_new_n17621__,
    new_new_n17622__, new_new_n17623__, new_new_n17624__, new_new_n17625__,
    new_new_n17627__, new_new_n17628__, new_new_n17629__, new_new_n17630__,
    new_new_n17632__, new_new_n17633__, new_new_n17635__, new_new_n17636__,
    new_new_n17637__, new_new_n17638__, new_new_n17640__, new_new_n17641__,
    new_new_n17642__, new_new_n17643__, new_new_n17644__, new_new_n17645__,
    new_new_n17647__, new_new_n17649__, new_new_n17650__, new_new_n17651__,
    new_new_n17652__, new_new_n17653__, new_new_n17655__, new_new_n17656__,
    new_new_n17657__, new_new_n17658__, new_new_n17660__, new_new_n17661__,
    new_new_n17663__, new_new_n17664__, new_new_n17665__, new_new_n17666__,
    new_new_n17668__, new_new_n17669__, new_new_n17670__, new_new_n17671__,
    new_new_n17672__, new_new_n17673__, new_new_n17675__, new_new_n17677__,
    new_new_n17678__, new_new_n17679__, new_new_n17680__, new_new_n17681__,
    new_new_n17683__, new_new_n17684__, new_new_n17685__, new_new_n17686__,
    new_new_n17688__, new_new_n17689__, new_new_n17691__, new_new_n17692__,
    new_new_n17694__, new_new_n17695__, new_new_n17697__, new_new_n17698__,
    new_new_n17700__, new_new_n17701__, new_new_n17703__, new_new_n17704__,
    new_new_n17706__, new_new_n17707__, new_new_n17709__, new_new_n17710__,
    new_new_n17712__, new_new_n17713__, new_new_n17715__, new_new_n17716__,
    new_new_n17718__, new_new_n17719__, new_new_n17721__, new_new_n17722__,
    new_new_n17724__, new_new_n17725__, new_new_n17726__, new_new_n17727__,
    new_new_n17728__, new_new_n17730__, new_new_n17731__, new_new_n17733__,
    new_new_n17734__, new_new_n17735__, new_new_n17736__, new_new_n17737__,
    new_new_n17739__, new_new_n17740__, new_new_n17742__, new_new_n17743__,
    new_new_n17744__, new_new_n17745__, new_new_n17746__, new_new_n17748__,
    new_new_n17749__, new_new_n17751__, new_new_n17752__, new_new_n17753__,
    new_new_n17754__, new_new_n17755__, new_new_n17757__, new_new_n17758__,
    new_new_n17760__, new_new_n17761__, new_new_n17762__, new_new_n17763__,
    new_new_n17764__, new_new_n17766__, new_new_n17767__, new_new_n17769__,
    new_new_n17770__, new_new_n17771__, new_new_n17772__, new_new_n17773__,
    new_new_n17775__, new_new_n17776__, new_new_n17778__, new_new_n17779__,
    new_new_n17780__, new_new_n17781__, new_new_n17782__, new_new_n17784__,
    new_new_n17785__, new_new_n17787__, new_new_n17788__, new_new_n17789__,
    new_new_n17790__, new_new_n17791__, new_new_n17793__, new_new_n17794__,
    new_new_n17796__, new_new_n17797__, new_new_n17798__, new_new_n17799__,
    new_new_n17800__, new_new_n17802__, new_new_n17803__, new_new_n17805__,
    new_new_n17806__, new_new_n17807__, new_new_n17808__, new_new_n17809__,
    new_new_n17811__, new_new_n17812__, new_new_n17814__, new_new_n17815__,
    new_new_n17816__, new_new_n17817__, new_new_n17818__, new_new_n17820__,
    new_new_n17821__, new_new_n17823__, new_new_n17824__, new_new_n17825__,
    new_new_n17826__, new_new_n17827__, new_new_n17829__, new_new_n17830__,
    new_new_n17832__, new_new_n17833__, new_new_n17834__, new_new_n17835__,
    new_new_n17836__, new_new_n17838__, new_new_n17839__, new_new_n17841__,
    new_new_n17842__, new_new_n17843__, new_new_n17844__, new_new_n17845__,
    new_new_n17847__, new_new_n17848__, new_new_n17850__, new_new_n17851__,
    new_new_n17852__, new_new_n17853__, new_new_n17854__, new_new_n17856__,
    new_new_n17857__, new_new_n17859__, new_new_n17860__, new_new_n17861__,
    new_new_n17862__, new_new_n17863__, new_new_n17865__, new_new_n17866__,
    new_new_n17868__, new_new_n17869__, new_new_n17870__, new_new_n17871__,
    new_new_n17872__, new_new_n17874__, new_new_n17875__, new_new_n17877__,
    new_new_n17878__, new_new_n17879__, new_new_n17880__, new_new_n17881__,
    new_new_n17883__, new_new_n17884__, new_new_n17886__, new_new_n17887__,
    new_new_n17888__, new_new_n17889__, new_new_n17890__, new_new_n17892__,
    new_new_n17893__, new_new_n17895__, new_new_n17896__, new_new_n17897__,
    new_new_n17898__, new_new_n17899__, new_new_n17901__, new_new_n17902__,
    new_new_n17904__, new_new_n17905__, new_new_n17906__, new_new_n17907__,
    new_new_n17908__, new_new_n17910__, new_new_n17911__, new_new_n17913__,
    new_new_n17914__, new_new_n17915__, new_new_n17916__, new_new_n17917__,
    new_new_n17919__, new_new_n17920__, new_new_n17922__, new_new_n17923__,
    new_new_n17924__, new_new_n17925__, new_new_n17926__, new_new_n17928__,
    new_new_n17929__, new_new_n17931__, new_new_n17932__, new_new_n17933__,
    new_new_n17934__, new_new_n17935__, new_new_n17937__, new_new_n17938__,
    new_new_n17940__, new_new_n17941__, new_new_n17942__, new_new_n17943__,
    new_new_n17944__, new_new_n17946__, new_new_n17947__, new_new_n17949__,
    new_new_n17950__, new_new_n17951__, new_new_n17952__, new_new_n17953__,
    new_new_n17955__, new_new_n17956__, new_new_n17958__, new_new_n17959__,
    new_new_n17960__, new_new_n17961__, new_new_n17962__, new_new_n17964__,
    new_new_n17965__, new_new_n17967__, new_new_n17968__, new_new_n17969__,
    new_new_n17970__, new_new_n17971__, new_new_n17973__, new_new_n17974__,
    new_new_n17976__, new_new_n17977__, new_new_n17978__, new_new_n17979__,
    new_new_n17980__, new_new_n17982__, new_new_n17983__, new_new_n17985__,
    new_new_n17986__, new_new_n17987__, new_new_n17988__, new_new_n17989__,
    new_new_n17991__, new_new_n17992__, new_new_n17994__, new_new_n17995__,
    new_new_n17996__, new_new_n17997__, new_new_n17998__, new_new_n18000__,
    new_new_n18001__, new_new_n18003__, new_new_n18004__, new_new_n18005__,
    new_new_n18006__, new_new_n18007__, new_new_n18009__, new_new_n18010__,
    new_new_n18012__, new_new_n18014__, new_new_n18015__, new_new_n18017__,
    new_new_n18018__, new_new_n18019__, new_new_n18020__, new_new_n18022__,
    new_new_n18023__, new_new_n18024__, new_new_n18025__, new_new_n18026__,
    new_new_n18028__, new_new_n18029__, new_new_n18032__, new_new_n18033__,
    new_new_n18034__, new_new_n18035__, new_new_n18036__, new_new_n18037__,
    new_new_n18038__, new_new_n18039__, new_new_n18040__, new_new_n18041__,
    new_new_n18042__, new_new_n18043__, new_new_n18044__, new_new_n18046__,
    new_new_n18047__, new_new_n18049__, new_new_n18050__, new_new_n18052__,
    new_new_n18053__, new_new_n18055__, new_new_n18056__, new_new_n18057__,
    new_new_n18059__, new_new_n18060__, new_new_n18061__, new_new_n18062__,
    new_new_n18063__, new_new_n18064__, new_new_n18065__, new_new_n18066__,
    new_new_n18067__, new_new_n18068__, new_new_n18069__, new_new_n18071__,
    new_new_n18072__, new_new_n18074__, new_new_n18075__, new_new_n18076__,
    new_new_n18078__, new_new_n18079__, new_new_n18080__, new_new_n18082__,
    new_new_n18083__, new_new_n18084__, new_new_n18086__, new_new_n18087__,
    new_new_n18088__, new_new_n18090__, new_new_n18091__, new_new_n18092__,
    new_new_n18094__, new_new_n18095__, new_new_n18096__, new_new_n18097__,
    new_new_n18098__, new_new_n18100__, new_new_n18101__, new_new_n18102__,
    new_new_n18104__, new_new_n18106__, new_new_n18107__, new_new_n18108__,
    new_new_n18109__, new_new_n18110__, new_new_n18112__, new_new_n18113__,
    new_new_n18114__, new_new_n18116__, new_new_n18117__, new_new_n18118__,
    new_new_n18119__, new_new_n18120__, new_new_n18121__, new_new_n18122__,
    new_new_n18123__, new_new_n18124__, new_new_n18125__, new_new_n18126__,
    new_new_n18127__, new_new_n18128__, new_new_n18129__, new_new_n18130__,
    new_new_n18131__, new_new_n18132__, new_new_n18133__, new_new_n18134__,
    new_new_n18135__, new_new_n18136__, new_new_n18137__, new_new_n18138__,
    new_new_n18139__, new_new_n18140__, new_new_n18141__, new_new_n18142__,
    new_new_n18143__, new_new_n18144__, new_new_n18145__, new_new_n18146__,
    new_new_n18147__, new_new_n18148__, new_new_n18149__, new_new_n18150__,
    new_new_n18151__, new_new_n18152__, new_new_n18153__, new_new_n18154__,
    new_new_n18155__, new_new_n18156__, new_new_n18157__, new_new_n18158__,
    new_new_n18159__, new_new_n18160__, new_new_n18161__, new_new_n18162__,
    new_new_n18163__, new_new_n18164__, new_new_n18165__, new_new_n18166__,
    new_new_n18167__, new_new_n18168__, new_new_n18169__, new_new_n18170__,
    new_new_n18171__, new_new_n18172__, new_new_n18173__, new_new_n18174__,
    new_new_n18175__, new_new_n18176__, new_new_n18177__, new_new_n18178__,
    new_new_n18179__, new_new_n18180__, new_new_n18181__, new_new_n18182__,
    new_new_n18183__, new_new_n18184__, new_new_n18185__, new_new_n18186__,
    new_new_n18187__, new_new_n18188__, new_new_n18189__, new_new_n18190__,
    new_new_n18191__, new_new_n18192__, new_new_n18193__, new_new_n18194__,
    new_new_n18195__, new_new_n18196__, new_new_n18197__, new_new_n18198__,
    new_new_n18199__, new_new_n18200__, new_new_n18201__, new_new_n18202__,
    new_new_n18203__, new_new_n18204__, new_new_n18205__, new_new_n18206__,
    new_new_n18207__, new_new_n18208__, new_new_n18209__, new_new_n18210__,
    new_new_n18211__, new_new_n18212__, new_new_n18213__, new_new_n18214__,
    new_new_n18215__, new_new_n18216__, new_new_n18217__, new_new_n18218__,
    new_new_n18219__, new_new_n18220__, new_new_n18221__, new_new_n18222__,
    new_new_n18223__, new_new_n18224__, new_new_n18225__, new_new_n18226__,
    new_new_n18227__, new_new_n18228__, new_new_n18229__, new_new_n18230__,
    new_new_n18231__, new_new_n18232__, new_new_n18233__, new_new_n18234__,
    new_new_n18235__, new_new_n18236__, new_new_n18237__, new_new_n18238__,
    new_new_n18239__, new_new_n18240__, new_new_n18241__, new_new_n18242__,
    new_new_n18243__, new_new_n18244__, new_new_n18245__, new_new_n18246__,
    new_new_n18247__, new_new_n18248__, new_new_n18249__, new_new_n18250__,
    new_new_n18251__, new_new_n18252__, new_new_n18253__, new_new_n18254__,
    new_new_n18255__, new_new_n18256__, new_new_n18257__, new_new_n18258__,
    new_new_n18259__, new_new_n18260__, new_new_n18261__, new_new_n18262__,
    new_new_n18263__, new_new_n18264__, new_new_n18265__, new_new_n18266__,
    new_new_n18267__, new_new_n18268__, new_new_n18269__, new_new_n18270__,
    new_new_n18271__, new_new_n18272__, new_new_n18273__, new_new_n18274__,
    new_new_n18275__, new_new_n18276__, new_new_n18277__, new_new_n18278__,
    new_new_n18279__, new_new_n18280__, new_new_n18281__, new_new_n18282__,
    new_new_n18283__, new_new_n18284__, new_new_n18285__, new_new_n18286__,
    new_new_n18287__, new_new_n18288__, new_new_n18289__, new_new_n18290__,
    new_new_n18291__, new_new_n18292__, new_new_n18293__, new_new_n18294__,
    new_new_n18295__, new_new_n18296__, new_new_n18297__, new_new_n18298__,
    new_new_n18299__, new_new_n18300__, new_new_n18301__, new_new_n18302__,
    new_new_n18303__, new_new_n18304__, new_new_n18305__, new_new_n18306__,
    new_new_n18307__, new_new_n18308__, new_new_n18309__, new_new_n18310__,
    new_new_n18311__, new_new_n18312__, new_new_n18313__, new_new_n18314__,
    new_new_n18315__, new_new_n18316__, new_new_n18317__, new_new_n18318__,
    new_new_n18319__, new_new_n18320__, new_new_n18321__, new_new_n18322__,
    new_new_n18323__, new_new_n18324__, new_new_n18325__, new_new_n18326__,
    new_new_n18327__, new_new_n18328__, new_new_n18329__, new_new_n18330__,
    new_new_n18331__, new_new_n18332__, new_new_n18333__, new_new_n18334__,
    new_new_n18335__, new_new_n18336__, new_new_n18337__, new_new_n18338__,
    new_new_n18339__, new_new_n18340__, new_new_n18341__, new_new_n18342__,
    new_new_n18343__, new_new_n18344__, new_new_n18345__, new_new_n18346__,
    new_new_n18347__, new_new_n18348__, new_new_n18349__, new_new_n18350__,
    new_new_n18351__, new_new_n18352__, new_new_n18353__, new_new_n18354__,
    new_new_n18355__, new_new_n18356__, new_new_n18357__, new_new_n18358__,
    new_new_n18359__, new_new_n18360__, new_new_n18361__, new_new_n18362__,
    new_new_n18363__, new_new_n18364__, new_new_n18365__, new_new_n18366__,
    new_new_n18367__, new_new_n18368__, new_new_n18369__, new_new_n18370__,
    new_new_n18371__, new_new_n18372__, new_new_n18373__, new_new_n18374__,
    new_new_n18375__, new_new_n18376__, new_new_n18377__, new_new_n18378__,
    new_new_n18379__, new_new_n18380__, new_new_n18381__, new_new_n18382__,
    new_new_n18383__, new_new_n18384__, new_new_n18385__, new_new_n18386__,
    new_new_n18387__, new_new_n18388__, new_new_n18389__, new_new_n18390__,
    new_new_n18391__, new_new_n18392__, new_new_n18393__, new_new_n18394__,
    new_new_n18395__, new_new_n18396__, new_new_n18397__, new_new_n18398__,
    new_new_n18399__, new_new_n18400__, new_new_n18401__, new_new_n18402__,
    new_new_n18403__, new_new_n18404__, new_new_n18405__, new_new_n18406__,
    new_new_n18407__, new_new_n18408__, new_new_n18409__, new_new_n18410__,
    new_new_n18411__, new_new_n18412__, new_new_n18413__, new_new_n18414__,
    new_new_n18415__, new_new_n18416__, new_new_n18417__, new_new_n18418__,
    new_new_n18419__, new_new_n18420__, new_new_n18421__, new_new_n18422__,
    new_new_n18423__, new_new_n18424__, new_new_n18425__, new_new_n18426__,
    new_new_n18427__, new_new_n18428__, new_new_n18429__, new_new_n18430__,
    new_new_n18431__, new_new_n18432__, new_new_n18433__, new_new_n18434__,
    new_new_n18435__, new_new_n18436__, new_new_n18437__, new_new_n18438__,
    new_new_n18439__, new_new_n18440__, new_new_n18441__, new_new_n18442__,
    new_new_n18443__, new_new_n18444__, new_new_n18445__, new_new_n18446__,
    new_new_n18447__, new_new_n18448__, new_new_n18449__, new_new_n18450__,
    new_new_n18451__, new_new_n18452__, new_new_n18453__, new_new_n18454__,
    new_new_n18456__, new_new_n18457__, new_new_n18458__, new_new_n18459__,
    new_new_n18460__, new_new_n18461__, new_new_n18462__, new_new_n18463__,
    new_new_n18464__, new_new_n18465__, new_new_n18466__, new_new_n18467__,
    new_new_n18468__, new_new_n18469__, new_new_n18470__, new_new_n18471__,
    new_new_n18472__, new_new_n18473__, new_new_n18474__, new_new_n18475__,
    new_new_n18476__, new_new_n18477__, new_new_n18478__, new_new_n18479__,
    new_new_n18480__, new_new_n18481__, new_new_n18482__, new_new_n18483__,
    new_new_n18484__, new_new_n18485__, new_new_n18486__, new_new_n18487__,
    new_new_n18488__, new_new_n18489__, new_new_n18490__, new_new_n18491__,
    new_new_n18492__, new_new_n18493__, new_new_n18494__, new_new_n18495__,
    new_new_n18496__, new_new_n18497__, new_new_n18498__, new_new_n18499__,
    new_new_n18500__, new_new_n18501__, new_new_n18502__, new_new_n18503__,
    new_new_n18504__, new_new_n18505__, new_new_n18506__, new_new_n18507__,
    new_new_n18508__, new_new_n18509__, new_new_n18510__, new_new_n18511__,
    new_new_n18512__, new_new_n18513__, new_new_n18514__, new_new_n18515__,
    new_new_n18516__, new_new_n18517__, new_new_n18518__, new_new_n18519__,
    new_new_n18520__, new_new_n18521__, new_new_n18522__, new_new_n18523__,
    new_new_n18524__, new_new_n18525__, new_new_n18526__, new_new_n18527__,
    new_new_n18528__, new_new_n18529__, new_new_n18530__, new_new_n18531__,
    new_new_n18532__, new_new_n18533__, new_new_n18534__, new_new_n18535__,
    new_new_n18536__, new_new_n18537__, new_new_n18538__, new_new_n18539__,
    new_new_n18540__, new_new_n18541__, new_new_n18542__, new_new_n18543__,
    new_new_n18544__, new_new_n18545__, new_new_n18546__, new_new_n18547__,
    new_new_n18548__, new_new_n18549__, new_new_n18550__, new_new_n18551__,
    new_new_n18552__, new_new_n18553__, new_new_n18554__, new_new_n18555__,
    new_new_n18556__, new_new_n18557__, new_new_n18558__, new_new_n18559__,
    new_new_n18560__, new_new_n18561__, new_new_n18562__, new_new_n18563__,
    new_new_n18564__, new_new_n18565__, new_new_n18566__, new_new_n18567__,
    new_new_n18568__, new_new_n18569__, new_new_n18570__, new_new_n18571__,
    new_new_n18572__, new_new_n18573__, new_new_n18574__, new_new_n18575__,
    new_new_n18576__, new_new_n18577__, new_new_n18578__, new_new_n18579__,
    new_new_n18580__, new_new_n18581__, new_new_n18582__, new_new_n18583__,
    new_new_n18584__, new_new_n18585__, new_new_n18586__, new_new_n18587__,
    new_new_n18588__, new_new_n18589__, new_new_n18590__, new_new_n18591__,
    new_new_n18592__, new_new_n18593__, new_new_n18594__, new_new_n18595__,
    new_new_n18596__, new_new_n18597__, new_new_n18598__, new_new_n18599__,
    new_new_n18600__, new_new_n18601__, new_new_n18602__, new_new_n18603__,
    new_new_n18605__, new_new_n18606__, new_new_n18607__, new_new_n18608__,
    new_new_n18609__, new_new_n18610__, new_new_n18611__, new_new_n18612__,
    new_new_n18613__, new_new_n18614__, new_new_n18615__, new_new_n18616__,
    new_new_n18617__, new_new_n18618__, new_new_n18619__, new_new_n18620__,
    new_new_n18621__, new_new_n18622__, new_new_n18623__, new_new_n18624__,
    new_new_n18625__, new_new_n18626__, new_new_n18627__, new_new_n18628__,
    new_new_n18629__, new_new_n18630__, new_new_n18631__, new_new_n18632__,
    new_new_n18633__, new_new_n18634__, new_new_n18635__, new_new_n18636__,
    new_new_n18637__, new_new_n18638__, new_new_n18639__, new_new_n18640__,
    new_new_n18641__, new_new_n18642__, new_new_n18643__, new_new_n18644__,
    new_new_n18645__, new_new_n18646__, new_new_n18647__, new_new_n18648__,
    new_new_n18649__, new_new_n18650__, new_new_n18651__, new_new_n18652__,
    new_new_n18653__, new_new_n18654__, new_new_n18655__, new_new_n18656__,
    new_new_n18657__, new_new_n18658__, new_new_n18659__, new_new_n18660__,
    new_new_n18661__, new_new_n18662__, new_new_n18663__, new_new_n18664__,
    new_new_n18665__, new_new_n18666__, new_new_n18667__, new_new_n18668__,
    new_new_n18669__, new_new_n18670__, new_new_n18671__, new_new_n18672__,
    new_new_n18673__, new_new_n18674__, new_new_n18675__, new_new_n18676__,
    new_new_n18677__, new_new_n18678__, new_new_n18679__, new_new_n18680__,
    new_new_n18681__, new_new_n18682__, new_new_n18683__, new_new_n18684__,
    new_new_n18685__, new_new_n18686__, new_new_n18687__, new_new_n18688__,
    new_new_n18689__, new_new_n18690__, new_new_n18691__, new_new_n18692__,
    new_new_n18693__, new_new_n18694__, new_new_n18695__, new_new_n18696__,
    new_new_n18697__, new_new_n18698__, new_new_n18699__, new_new_n18700__,
    new_new_n18701__, new_new_n18702__, new_new_n18703__, new_new_n18704__,
    new_new_n18705__, new_new_n18706__, new_new_n18707__, new_new_n18709__,
    new_new_n18710__, new_new_n18711__, new_new_n18712__, new_new_n18713__,
    new_new_n18714__, new_new_n18715__, new_new_n18716__, new_new_n18717__,
    new_new_n18718__, new_new_n18719__, new_new_n18720__, new_new_n18721__,
    new_new_n18722__, new_new_n18723__, new_new_n18724__, new_new_n18725__,
    new_new_n18726__, new_new_n18727__, new_new_n18728__, new_new_n18729__,
    new_new_n18730__, new_new_n18731__, new_new_n18732__, new_new_n18733__,
    new_new_n18734__, new_new_n18735__, new_new_n18736__, new_new_n18737__,
    new_new_n18738__, new_new_n18739__, new_new_n18740__, new_new_n18741__,
    new_new_n18742__, new_new_n18743__, new_new_n18744__, new_new_n18745__,
    new_new_n18746__, new_new_n18747__, new_new_n18748__, new_new_n18749__,
    new_new_n18750__, new_new_n18751__, new_new_n18752__, new_new_n18753__,
    new_new_n18754__, new_new_n18755__, new_new_n18756__, new_new_n18757__,
    new_new_n18758__, new_new_n18759__, new_new_n18760__, new_new_n18761__,
    new_new_n18762__, new_new_n18763__, new_new_n18764__, new_new_n18765__,
    new_new_n18766__, new_new_n18767__, new_new_n18768__, new_new_n18769__,
    new_new_n18770__, new_new_n18771__, new_new_n18772__, new_new_n18773__,
    new_new_n18774__, new_new_n18775__, new_new_n18776__, new_new_n18777__,
    new_new_n18778__, new_new_n18779__, new_new_n18780__, new_new_n18781__,
    new_new_n18782__, new_new_n18783__, new_new_n18784__, new_new_n18785__,
    new_new_n18786__, new_new_n18787__, new_new_n18788__, new_new_n18789__,
    new_new_n18790__, new_new_n18791__, new_new_n18792__, new_new_n18793__,
    new_new_n18794__, new_new_n18795__, new_new_n18796__, new_new_n18797__,
    new_new_n18798__, new_new_n18799__, new_new_n18800__, new_new_n18801__,
    new_new_n18802__, new_new_n18803__, new_new_n18804__, new_new_n18805__,
    new_new_n18806__, new_new_n18807__, new_new_n18808__, new_new_n18809__,
    new_new_n18810__, new_new_n18811__, new_new_n18812__, new_new_n18813__,
    new_new_n18814__, new_new_n18816__, new_new_n18817__, new_new_n18818__,
    new_new_n18819__, new_new_n18820__, new_new_n18821__, new_new_n18822__,
    new_new_n18823__, new_new_n18824__, new_new_n18825__, new_new_n18826__,
    new_new_n18827__, new_new_n18828__, new_new_n18829__, new_new_n18830__,
    new_new_n18831__, new_new_n18832__, new_new_n18833__, new_new_n18834__,
    new_new_n18835__, new_new_n18836__, new_new_n18837__, new_new_n18838__,
    new_new_n18839__, new_new_n18840__, new_new_n18841__, new_new_n18842__,
    new_new_n18843__, new_new_n18844__, new_new_n18845__, new_new_n18846__,
    new_new_n18847__, new_new_n18848__, new_new_n18849__, new_new_n18850__,
    new_new_n18851__, new_new_n18852__, new_new_n18853__, new_new_n18854__,
    new_new_n18855__, new_new_n18856__, new_new_n18857__, new_new_n18858__,
    new_new_n18859__, new_new_n18860__, new_new_n18861__, new_new_n18862__,
    new_new_n18863__, new_new_n18864__, new_new_n18865__, new_new_n18866__,
    new_new_n18867__, new_new_n18868__, new_new_n18869__, new_new_n18870__,
    new_new_n18871__, new_new_n18872__, new_new_n18873__, new_new_n18874__,
    new_new_n18875__, new_new_n18876__, new_new_n18877__, new_new_n18878__,
    new_new_n18879__, new_new_n18880__, new_new_n18881__, new_new_n18882__,
    new_new_n18883__, new_new_n18884__, new_new_n18885__, new_new_n18886__,
    new_new_n18887__, new_new_n18888__, new_new_n18889__, new_new_n18890__,
    new_new_n18891__, new_new_n18892__, new_new_n18893__, new_new_n18894__,
    new_new_n18896__, new_new_n18897__, new_new_n18898__, new_new_n18899__,
    new_new_n18900__, new_new_n18901__, new_new_n18902__, new_new_n18903__,
    new_new_n18904__, new_new_n18905__, new_new_n18906__, new_new_n18907__,
    new_new_n18908__, new_new_n18909__, new_new_n18910__, new_new_n18911__,
    new_new_n18912__, new_new_n18913__, new_new_n18914__, new_new_n18915__,
    new_new_n18916__, new_new_n18917__, new_new_n18918__, new_new_n18919__,
    new_new_n18920__, new_new_n18921__, new_new_n18922__, new_new_n18923__,
    new_new_n18924__, new_new_n18925__, new_new_n18926__, new_new_n18927__,
    new_new_n18928__, new_new_n18929__, new_new_n18930__, new_new_n18931__,
    new_new_n18932__, new_new_n18933__, new_new_n18934__, new_new_n18935__,
    new_new_n18936__, new_new_n18937__, new_new_n18938__, new_new_n18939__,
    new_new_n18940__, new_new_n18941__, new_new_n18942__, new_new_n18943__,
    new_new_n18944__, new_new_n18945__, new_new_n18946__, new_new_n18947__,
    new_new_n18948__, new_new_n18949__, new_new_n18950__, new_new_n18951__,
    new_new_n18952__, new_new_n18953__, new_new_n18954__, new_new_n18955__,
    new_new_n18956__, new_new_n18957__, new_new_n18958__, new_new_n18959__,
    new_new_n18960__, new_new_n18961__, new_new_n18962__, new_new_n18963__,
    new_new_n18964__, new_new_n18965__, new_new_n18966__, new_new_n18967__,
    new_new_n18968__, new_new_n18969__, new_new_n18970__, new_new_n18971__,
    new_new_n18972__, new_new_n18973__, new_new_n18974__, new_new_n18975__,
    new_new_n18976__, new_new_n18977__, new_new_n18978__, new_new_n18979__,
    new_new_n18981__, new_new_n18982__, new_new_n18983__, new_new_n18984__,
    new_new_n18985__, new_new_n18986__, new_new_n18987__, new_new_n18988__,
    new_new_n18989__, new_new_n18990__, new_new_n18991__, new_new_n18992__,
    new_new_n18993__, new_new_n18994__, new_new_n18995__, new_new_n18996__,
    new_new_n18997__, new_new_n18998__, new_new_n18999__, new_new_n19000__,
    new_new_n19001__, new_new_n19002__, new_new_n19003__, new_new_n19004__,
    new_new_n19005__, new_new_n19006__, new_new_n19007__, new_new_n19008__,
    new_new_n19009__, new_new_n19010__, new_new_n19011__, new_new_n19012__,
    new_new_n19013__, new_new_n19014__, new_new_n19015__, new_new_n19016__,
    new_new_n19017__, new_new_n19018__, new_new_n19019__, new_new_n19020__,
    new_new_n19021__, new_new_n19022__, new_new_n19023__, new_new_n19024__,
    new_new_n19025__, new_new_n19026__, new_new_n19027__, new_new_n19028__,
    new_new_n19029__, new_new_n19030__, new_new_n19031__, new_new_n19032__,
    new_new_n19033__, new_new_n19034__, new_new_n19035__, new_new_n19036__,
    new_new_n19037__, new_new_n19038__, new_new_n19039__, new_new_n19040__,
    new_new_n19041__, new_new_n19042__, new_new_n19043__, new_new_n19044__,
    new_new_n19045__, new_new_n19046__, new_new_n19047__, new_new_n19048__,
    new_new_n19049__, new_new_n19050__, new_new_n19051__, new_new_n19052__,
    new_new_n19053__, new_new_n19054__, new_new_n19055__, new_new_n19056__,
    new_new_n19057__, new_new_n19058__, new_new_n19059__, new_new_n19060__,
    new_new_n19061__, new_new_n19062__, new_new_n19063__, new_new_n19064__,
    new_new_n19066__, new_new_n19067__, new_new_n19068__, new_new_n19069__,
    new_new_n19070__, new_new_n19071__, new_new_n19072__, new_new_n19073__,
    new_new_n19074__, new_new_n19075__, new_new_n19076__, new_new_n19077__,
    new_new_n19078__, new_new_n19079__, new_new_n19080__, new_new_n19081__,
    new_new_n19082__, new_new_n19083__, new_new_n19084__, new_new_n19085__,
    new_new_n19086__, new_new_n19087__, new_new_n19088__, new_new_n19089__,
    new_new_n19090__, new_new_n19091__, new_new_n19092__, new_new_n19093__,
    new_new_n19094__, new_new_n19095__, new_new_n19096__, new_new_n19097__,
    new_new_n19098__, new_new_n19099__, new_new_n19100__, new_new_n19101__,
    new_new_n19102__, new_new_n19103__, new_new_n19104__, new_new_n19105__,
    new_new_n19106__, new_new_n19107__, new_new_n19108__, new_new_n19109__,
    new_new_n19110__, new_new_n19111__, new_new_n19112__, new_new_n19113__,
    new_new_n19114__, new_new_n19115__, new_new_n19116__, new_new_n19117__,
    new_new_n19118__, new_new_n19119__, new_new_n19120__, new_new_n19121__,
    new_new_n19122__, new_new_n19123__, new_new_n19124__, new_new_n19125__,
    new_new_n19126__, new_new_n19127__, new_new_n19128__, new_new_n19129__,
    new_new_n19130__, new_new_n19131__, new_new_n19132__, new_new_n19133__,
    new_new_n19134__, new_new_n19135__, new_new_n19136__, new_new_n19137__,
    new_new_n19138__, new_new_n19139__, new_new_n19140__, new_new_n19141__,
    new_new_n19142__, new_new_n19143__, new_new_n19144__, new_new_n19145__,
    new_new_n19146__, new_new_n19147__, new_new_n19149__, new_new_n19150__,
    new_new_n19151__, new_new_n19152__, new_new_n19153__, new_new_n19154__,
    new_new_n19155__, new_new_n19156__, new_new_n19157__, new_new_n19158__,
    new_new_n19159__, new_new_n19160__, new_new_n19161__, new_new_n19162__,
    new_new_n19163__, new_new_n19164__, new_new_n19165__, new_new_n19166__,
    new_new_n19167__, new_new_n19168__, new_new_n19169__, new_new_n19170__,
    new_new_n19171__, new_new_n19172__, new_new_n19173__, new_new_n19174__,
    new_new_n19175__, new_new_n19176__, new_new_n19177__, new_new_n19178__,
    new_new_n19179__, new_new_n19180__, new_new_n19181__, new_new_n19182__,
    new_new_n19183__, new_new_n19184__, new_new_n19185__, new_new_n19186__,
    new_new_n19187__, new_new_n19188__, new_new_n19189__, new_new_n19190__,
    new_new_n19191__, new_new_n19192__, new_new_n19193__, new_new_n19194__,
    new_new_n19195__, new_new_n19196__, new_new_n19197__, new_new_n19198__,
    new_new_n19199__, new_new_n19200__, new_new_n19201__, new_new_n19202__,
    new_new_n19203__, new_new_n19204__, new_new_n19205__, new_new_n19206__,
    new_new_n19207__, new_new_n19208__, new_new_n19209__, new_new_n19210__,
    new_new_n19211__, new_new_n19212__, new_new_n19213__, new_new_n19214__,
    new_new_n19215__, new_new_n19217__, new_new_n19218__, new_new_n19219__,
    new_new_n19220__, new_new_n19221__, new_new_n19222__, new_new_n19223__,
    new_new_n19224__, new_new_n19225__, new_new_n19226__, new_new_n19227__,
    new_new_n19228__, new_new_n19229__, new_new_n19230__, new_new_n19231__,
    new_new_n19232__, new_new_n19233__, new_new_n19234__, new_new_n19235__,
    new_new_n19236__, new_new_n19237__, new_new_n19238__, new_new_n19239__,
    new_new_n19240__, new_new_n19241__, new_new_n19242__, new_new_n19243__,
    new_new_n19244__, new_new_n19245__, new_new_n19246__, new_new_n19247__,
    new_new_n19248__, new_new_n19249__, new_new_n19250__, new_new_n19251__,
    new_new_n19252__, new_new_n19253__, new_new_n19254__, new_new_n19255__,
    new_new_n19256__, new_new_n19257__, new_new_n19258__, new_new_n19259__,
    new_new_n19260__, new_new_n19261__, new_new_n19262__, new_new_n19263__,
    new_new_n19264__, new_new_n19265__, new_new_n19266__, new_new_n19267__,
    new_new_n19268__, new_new_n19269__, new_new_n19270__, new_new_n19271__,
    new_new_n19272__, new_new_n19273__, new_new_n19274__, new_new_n19275__,
    new_new_n19276__, new_new_n19277__, new_new_n19278__, new_new_n19279__,
    new_new_n19280__, new_new_n19281__, new_new_n19282__, new_new_n19283__,
    new_new_n19284__, new_new_n19285__, new_new_n19286__, new_new_n19287__,
    new_new_n19288__, new_new_n19290__, new_new_n19291__, new_new_n19292__,
    new_new_n19293__, new_new_n19294__, new_new_n19295__, new_new_n19296__,
    new_new_n19297__, new_new_n19298__, new_new_n19299__, new_new_n19300__,
    new_new_n19301__, new_new_n19302__, new_new_n19303__, new_new_n19304__,
    new_new_n19305__, new_new_n19306__, new_new_n19307__, new_new_n19308__,
    new_new_n19309__, new_new_n19310__, new_new_n19311__, new_new_n19312__,
    new_new_n19313__, new_new_n19314__, new_new_n19315__, new_new_n19316__,
    new_new_n19317__, new_new_n19318__, new_new_n19319__, new_new_n19320__,
    new_new_n19321__, new_new_n19322__, new_new_n19323__, new_new_n19324__,
    new_new_n19325__, new_new_n19326__, new_new_n19327__, new_new_n19328__,
    new_new_n19329__, new_new_n19330__, new_new_n19331__, new_new_n19332__,
    new_new_n19333__, new_new_n19334__, new_new_n19335__, new_new_n19336__,
    new_new_n19337__, new_new_n19338__, new_new_n19339__, new_new_n19340__,
    new_new_n19341__, new_new_n19342__, new_new_n19343__, new_new_n19344__,
    new_new_n19345__, new_new_n19346__, new_new_n19347__, new_new_n19348__,
    new_new_n19349__, new_new_n19350__, new_new_n19351__, new_new_n19352__,
    new_new_n19353__, new_new_n19354__, new_new_n19355__, new_new_n19356__,
    new_new_n19357__, new_new_n19358__, new_new_n19359__, new_new_n19360__,
    new_new_n19361__, new_new_n19363__, new_new_n19364__, new_new_n19365__,
    new_new_n19366__, new_new_n19367__, new_new_n19368__, new_new_n19369__,
    new_new_n19370__, new_new_n19371__, new_new_n19372__, new_new_n19373__,
    new_new_n19374__, new_new_n19375__, new_new_n19376__, new_new_n19377__,
    new_new_n19378__, new_new_n19379__, new_new_n19380__, new_new_n19381__,
    new_new_n19382__, new_new_n19383__, new_new_n19384__, new_new_n19385__,
    new_new_n19386__, new_new_n19387__, new_new_n19388__, new_new_n19389__,
    new_new_n19390__, new_new_n19391__, new_new_n19392__, new_new_n19393__,
    new_new_n19394__, new_new_n19395__, new_new_n19396__, new_new_n19397__,
    new_new_n19398__, new_new_n19399__, new_new_n19400__, new_new_n19401__,
    new_new_n19402__, new_new_n19403__, new_new_n19404__, new_new_n19405__,
    new_new_n19406__, new_new_n19407__, new_new_n19408__, new_new_n19409__,
    new_new_n19410__, new_new_n19411__, new_new_n19412__, new_new_n19413__,
    new_new_n19414__, new_new_n19415__, new_new_n19416__, new_new_n19417__,
    new_new_n19418__, new_new_n19419__, new_new_n19420__, new_new_n19421__,
    new_new_n19422__, new_new_n19423__, new_new_n19424__, new_new_n19425__,
    new_new_n19426__, new_new_n19427__, new_new_n19428__, new_new_n19429__,
    new_new_n19430__, new_new_n19431__, new_new_n19432__, new_new_n19433__,
    new_new_n19434__, new_new_n19436__, new_new_n19437__, new_new_n19438__,
    new_new_n19439__, new_new_n19440__, new_new_n19441__, new_new_n19442__,
    new_new_n19443__, new_new_n19444__, new_new_n19445__, new_new_n19446__,
    new_new_n19447__, new_new_n19448__, new_new_n19449__, new_new_n19450__,
    new_new_n19451__, new_new_n19452__, new_new_n19453__, new_new_n19454__,
    new_new_n19455__, new_new_n19456__, new_new_n19457__, new_new_n19458__,
    new_new_n19459__, new_new_n19460__, new_new_n19461__, new_new_n19462__,
    new_new_n19463__, new_new_n19464__, new_new_n19465__, new_new_n19466__,
    new_new_n19467__, new_new_n19468__, new_new_n19469__, new_new_n19470__,
    new_new_n19471__, new_new_n19472__, new_new_n19473__, new_new_n19474__,
    new_new_n19475__, new_new_n19476__, new_new_n19477__, new_new_n19478__,
    new_new_n19479__, new_new_n19480__, new_new_n19481__, new_new_n19482__,
    new_new_n19483__, new_new_n19484__, new_new_n19485__, new_new_n19486__,
    new_new_n19487__, new_new_n19488__, new_new_n19489__, new_new_n19490__,
    new_new_n19491__, new_new_n19492__, new_new_n19493__, new_new_n19494__,
    new_new_n19495__, new_new_n19496__, new_new_n19497__, new_new_n19498__,
    new_new_n19499__, new_new_n19500__, new_new_n19501__, new_new_n19502__,
    new_new_n19503__, new_new_n19504__, new_new_n19505__, new_new_n19506__,
    new_new_n19507__, new_new_n19509__, new_new_n19510__, new_new_n19511__,
    new_new_n19512__, new_new_n19513__, new_new_n19514__, new_new_n19515__,
    new_new_n19516__, new_new_n19517__, new_new_n19518__, new_new_n19519__,
    new_new_n19520__, new_new_n19521__, new_new_n19522__, new_new_n19523__,
    new_new_n19524__, new_new_n19525__, new_new_n19526__, new_new_n19527__,
    new_new_n19528__, new_new_n19529__, new_new_n19530__, new_new_n19531__,
    new_new_n19532__, new_new_n19533__, new_new_n19534__, new_new_n19535__,
    new_new_n19536__, new_new_n19537__, new_new_n19538__, new_new_n19539__,
    new_new_n19540__, new_new_n19541__, new_new_n19542__, new_new_n19543__,
    new_new_n19544__, new_new_n19545__, new_new_n19546__, new_new_n19547__,
    new_new_n19548__, new_new_n19549__, new_new_n19550__, new_new_n19551__,
    new_new_n19552__, new_new_n19553__, new_new_n19554__, new_new_n19555__,
    new_new_n19556__, new_new_n19557__, new_new_n19558__, new_new_n19559__,
    new_new_n19560__, new_new_n19561__, new_new_n19562__, new_new_n19563__,
    new_new_n19564__, new_new_n19565__, new_new_n19566__, new_new_n19567__,
    new_new_n19568__, new_new_n19569__, new_new_n19570__, new_new_n19571__,
    new_new_n19572__, new_new_n19573__, new_new_n19574__, new_new_n19575__,
    new_new_n19576__, new_new_n19577__, new_new_n19578__, new_new_n19579__,
    new_new_n19580__, new_new_n19582__, new_new_n19583__, new_new_n19584__,
    new_new_n19585__, new_new_n19586__, new_new_n19587__, new_new_n19588__,
    new_new_n19589__, new_new_n19590__, new_new_n19591__, new_new_n19592__,
    new_new_n19593__, new_new_n19594__, new_new_n19595__, new_new_n19596__,
    new_new_n19597__, new_new_n19598__, new_new_n19599__, new_new_n19600__,
    new_new_n19601__, new_new_n19602__, new_new_n19603__, new_new_n19604__,
    new_new_n19605__, new_new_n19606__, new_new_n19607__, new_new_n19608__,
    new_new_n19609__, new_new_n19610__, new_new_n19611__, new_new_n19612__,
    new_new_n19613__, new_new_n19614__, new_new_n19615__, new_new_n19616__,
    new_new_n19617__, new_new_n19618__, new_new_n19619__, new_new_n19620__,
    new_new_n19621__, new_new_n19622__, new_new_n19623__, new_new_n19624__,
    new_new_n19625__, new_new_n19626__, new_new_n19627__, new_new_n19628__,
    new_new_n19629__, new_new_n19630__, new_new_n19631__, new_new_n19632__,
    new_new_n19633__, new_new_n19634__, new_new_n19635__, new_new_n19636__,
    new_new_n19637__, new_new_n19638__, new_new_n19639__, new_new_n19640__,
    new_new_n19641__, new_new_n19642__, new_new_n19643__, new_new_n19644__,
    new_new_n19645__, new_new_n19646__, new_new_n19647__, new_new_n19648__,
    new_new_n19649__, new_new_n19650__, new_new_n19651__, new_new_n19652__,
    new_new_n19653__, new_new_n19655__, new_new_n19656__, new_new_n19657__,
    new_new_n19658__, new_new_n19659__, new_new_n19660__, new_new_n19661__,
    new_new_n19662__, new_new_n19663__, new_new_n19664__, new_new_n19665__,
    new_new_n19666__, new_new_n19667__, new_new_n19668__, new_new_n19669__,
    new_new_n19670__, new_new_n19671__, new_new_n19672__, new_new_n19673__,
    new_new_n19674__, new_new_n19675__, new_new_n19676__, new_new_n19677__,
    new_new_n19678__, new_new_n19679__, new_new_n19680__, new_new_n19681__,
    new_new_n19682__, new_new_n19683__, new_new_n19684__, new_new_n19685__,
    new_new_n19686__, new_new_n19687__, new_new_n19688__, new_new_n19689__,
    new_new_n19690__, new_new_n19691__, new_new_n19692__, new_new_n19693__,
    new_new_n19694__, new_new_n19695__, new_new_n19696__, new_new_n19697__,
    new_new_n19698__, new_new_n19699__, new_new_n19700__, new_new_n19701__,
    new_new_n19702__, new_new_n19703__, new_new_n19704__, new_new_n19705__,
    new_new_n19706__, new_new_n19707__, new_new_n19708__, new_new_n19709__,
    new_new_n19710__, new_new_n19711__, new_new_n19712__, new_new_n19713__,
    new_new_n19714__, new_new_n19715__, new_new_n19716__, new_new_n19717__,
    new_new_n19718__, new_new_n19719__, new_new_n19720__, new_new_n19721__,
    new_new_n19722__, new_new_n19723__, new_new_n19724__, new_new_n19726__,
    new_new_n19727__, new_new_n19728__, new_new_n19729__, new_new_n19730__,
    new_new_n19731__, new_new_n19732__, new_new_n19733__, new_new_n19734__,
    new_new_n19735__, new_new_n19736__, new_new_n19737__, new_new_n19738__,
    new_new_n19739__, new_new_n19740__, new_new_n19741__, new_new_n19742__,
    new_new_n19743__, new_new_n19744__, new_new_n19745__, new_new_n19746__,
    new_new_n19747__, new_new_n19748__, new_new_n19749__, new_new_n19750__,
    new_new_n19751__, new_new_n19752__, new_new_n19753__, new_new_n19754__,
    new_new_n19755__, new_new_n19756__, new_new_n19757__, new_new_n19758__,
    new_new_n19759__, new_new_n19760__, new_new_n19761__, new_new_n19762__,
    new_new_n19763__, new_new_n19764__, new_new_n19765__, new_new_n19766__,
    new_new_n19767__, new_new_n19768__, new_new_n19769__, new_new_n19770__,
    new_new_n19771__, new_new_n19772__, new_new_n19773__, new_new_n19774__,
    new_new_n19775__, new_new_n19776__, new_new_n19777__, new_new_n19778__,
    new_new_n19779__, new_new_n19780__, new_new_n19781__, new_new_n19782__,
    new_new_n19783__, new_new_n19784__, new_new_n19785__, new_new_n19786__,
    new_new_n19787__, new_new_n19788__, new_new_n19790__, new_new_n19791__,
    new_new_n19792__, new_new_n19793__, new_new_n19794__, new_new_n19795__,
    new_new_n19796__, new_new_n19797__, new_new_n19798__, new_new_n19799__,
    new_new_n19800__, new_new_n19801__, new_new_n19802__, new_new_n19803__,
    new_new_n19804__, new_new_n19805__, new_new_n19806__, new_new_n19807__,
    new_new_n19808__, new_new_n19809__, new_new_n19810__, new_new_n19811__,
    new_new_n19812__, new_new_n19813__, new_new_n19814__, new_new_n19815__,
    new_new_n19816__, new_new_n19817__, new_new_n19818__, new_new_n19819__,
    new_new_n19820__, new_new_n19821__, new_new_n19822__, new_new_n19823__,
    new_new_n19824__, new_new_n19825__, new_new_n19826__, new_new_n19827__,
    new_new_n19828__, new_new_n19829__, new_new_n19830__, new_new_n19831__,
    new_new_n19832__, new_new_n19833__, new_new_n19834__, new_new_n19835__,
    new_new_n19836__, new_new_n19837__, new_new_n19838__, new_new_n19839__,
    new_new_n19840__, new_new_n19841__, new_new_n19842__, new_new_n19843__,
    new_new_n19844__, new_new_n19845__, new_new_n19846__, new_new_n19847__,
    new_new_n19848__, new_new_n19849__, new_new_n19850__, new_new_n19851__,
    new_new_n19852__, new_new_n19853__, new_new_n19854__, new_new_n19855__,
    new_new_n19856__, new_new_n19857__, new_new_n19859__, new_new_n19860__,
    new_new_n19861__, new_new_n19862__, new_new_n19863__, new_new_n19864__,
    new_new_n19865__, new_new_n19866__, new_new_n19867__, new_new_n19868__,
    new_new_n19869__, new_new_n19870__, new_new_n19871__, new_new_n19872__,
    new_new_n19873__, new_new_n19874__, new_new_n19875__, new_new_n19876__,
    new_new_n19877__, new_new_n19878__, new_new_n19879__, new_new_n19880__,
    new_new_n19881__, new_new_n19882__, new_new_n19883__, new_new_n19884__,
    new_new_n19885__, new_new_n19886__, new_new_n19887__, new_new_n19888__,
    new_new_n19889__, new_new_n19890__, new_new_n19891__, new_new_n19892__,
    new_new_n19893__, new_new_n19894__, new_new_n19895__, new_new_n19896__,
    new_new_n19897__, new_new_n19898__, new_new_n19899__, new_new_n19900__,
    new_new_n19901__, new_new_n19902__, new_new_n19903__, new_new_n19904__,
    new_new_n19905__, new_new_n19906__, new_new_n19907__, new_new_n19908__,
    new_new_n19909__, new_new_n19910__, new_new_n19911__, new_new_n19912__,
    new_new_n19913__, new_new_n19914__, new_new_n19915__, new_new_n19916__,
    new_new_n19917__, new_new_n19918__, new_new_n19919__, new_new_n19920__,
    new_new_n19921__, new_new_n19922__, new_new_n19923__, new_new_n19924__,
    new_new_n19925__, new_new_n19927__, new_new_n19928__, new_new_n19929__,
    new_new_n19930__, new_new_n19931__, new_new_n19932__, new_new_n19933__,
    new_new_n19934__, new_new_n19935__, new_new_n19936__, new_new_n19937__,
    new_new_n19938__, new_new_n19939__, new_new_n19940__, new_new_n19941__,
    new_new_n19942__, new_new_n19943__, new_new_n19944__, new_new_n19945__,
    new_new_n19946__, new_new_n19947__, new_new_n19948__, new_new_n19949__,
    new_new_n19950__, new_new_n19951__, new_new_n19952__, new_new_n19953__,
    new_new_n19954__, new_new_n19955__, new_new_n19956__, new_new_n19957__,
    new_new_n19958__, new_new_n19959__, new_new_n19960__, new_new_n19961__,
    new_new_n19962__, new_new_n19963__, new_new_n19964__, new_new_n19965__,
    new_new_n19966__, new_new_n19967__, new_new_n19968__, new_new_n19969__,
    new_new_n19970__, new_new_n19971__, new_new_n19972__, new_new_n19973__,
    new_new_n19974__, new_new_n19975__, new_new_n19976__, new_new_n19977__,
    new_new_n19978__, new_new_n19979__, new_new_n19980__, new_new_n19981__,
    new_new_n19982__, new_new_n19983__, new_new_n19984__, new_new_n19985__,
    new_new_n19986__, new_new_n19987__, new_new_n19988__, new_new_n19989__,
    new_new_n19990__, new_new_n19991__, new_new_n19992__, new_new_n19993__,
    new_new_n19995__, new_new_n19996__, new_new_n19997__, new_new_n19998__,
    new_new_n19999__, new_new_n20000__, new_new_n20001__, new_new_n20002__,
    new_new_n20003__, new_new_n20004__, new_new_n20005__, new_new_n20006__,
    new_new_n20007__, new_new_n20008__, new_new_n20009__, new_new_n20010__,
    new_new_n20011__, new_new_n20012__, new_new_n20013__, new_new_n20014__,
    new_new_n20015__, new_new_n20016__, new_new_n20017__, new_new_n20018__,
    new_new_n20019__, new_new_n20020__, new_new_n20021__, new_new_n20022__,
    new_new_n20023__, new_new_n20024__, new_new_n20025__, new_new_n20026__,
    new_new_n20027__, new_new_n20028__, new_new_n20029__, new_new_n20030__,
    new_new_n20031__, new_new_n20032__, new_new_n20033__, new_new_n20034__,
    new_new_n20035__, new_new_n20036__, new_new_n20037__, new_new_n20038__,
    new_new_n20039__, new_new_n20040__, new_new_n20041__, new_new_n20042__,
    new_new_n20043__, new_new_n20044__, new_new_n20045__, new_new_n20046__,
    new_new_n20047__, new_new_n20048__, new_new_n20049__, new_new_n20050__,
    new_new_n20051__, new_new_n20052__, new_new_n20053__, new_new_n20054__,
    new_new_n20055__, new_new_n20056__, new_new_n20057__, new_new_n20058__,
    new_new_n20059__, new_new_n20060__, new_new_n20061__, new_new_n20063__,
    new_new_n20064__, new_new_n20065__, new_new_n20066__, new_new_n20067__,
    new_new_n20068__, new_new_n20069__, new_new_n20070__, new_new_n20071__,
    new_new_n20072__, new_new_n20073__, new_new_n20074__, new_new_n20075__,
    new_new_n20076__, new_new_n20077__, new_new_n20078__, new_new_n20079__,
    new_new_n20080__, new_new_n20081__, new_new_n20082__, new_new_n20083__,
    new_new_n20084__, new_new_n20085__, new_new_n20086__, new_new_n20087__,
    new_new_n20088__, new_new_n20089__, new_new_n20090__, new_new_n20091__,
    new_new_n20092__, new_new_n20093__, new_new_n20094__, new_new_n20095__,
    new_new_n20096__, new_new_n20097__, new_new_n20098__, new_new_n20099__,
    new_new_n20100__, new_new_n20101__, new_new_n20102__, new_new_n20103__,
    new_new_n20104__, new_new_n20105__, new_new_n20106__, new_new_n20107__,
    new_new_n20108__, new_new_n20109__, new_new_n20110__, new_new_n20111__,
    new_new_n20112__, new_new_n20113__, new_new_n20114__, new_new_n20115__,
    new_new_n20116__, new_new_n20117__, new_new_n20118__, new_new_n20119__,
    new_new_n20120__, new_new_n20121__, new_new_n20122__, new_new_n20123__,
    new_new_n20124__, new_new_n20125__, new_new_n20126__, new_new_n20127__,
    new_new_n20128__, new_new_n20129__, new_new_n20131__, new_new_n20132__,
    new_new_n20133__, new_new_n20134__, new_new_n20135__, new_new_n20136__,
    new_new_n20137__, new_new_n20138__, new_new_n20139__, new_new_n20140__,
    new_new_n20141__, new_new_n20142__, new_new_n20143__, new_new_n20144__,
    new_new_n20145__, new_new_n20146__, new_new_n20147__, new_new_n20148__,
    new_new_n20149__, new_new_n20150__, new_new_n20151__, new_new_n20152__,
    new_new_n20153__, new_new_n20154__, new_new_n20155__, new_new_n20156__,
    new_new_n20157__, new_new_n20158__, new_new_n20159__, new_new_n20160__,
    new_new_n20161__, new_new_n20162__, new_new_n20163__, new_new_n20164__,
    new_new_n20165__, new_new_n20166__, new_new_n20167__, new_new_n20168__,
    new_new_n20169__, new_new_n20170__, new_new_n20171__, new_new_n20172__,
    new_new_n20173__, new_new_n20174__, new_new_n20175__, new_new_n20176__,
    new_new_n20177__, new_new_n20178__, new_new_n20179__, new_new_n20180__,
    new_new_n20181__, new_new_n20182__, new_new_n20183__, new_new_n20184__,
    new_new_n20185__, new_new_n20186__, new_new_n20187__, new_new_n20188__,
    new_new_n20189__, new_new_n20190__, new_new_n20191__, new_new_n20192__,
    new_new_n20193__, new_new_n20194__, new_new_n20195__, new_new_n20196__,
    new_new_n20197__, new_new_n20199__, new_new_n20200__, new_new_n20201__,
    new_new_n20202__, new_new_n20203__, new_new_n20204__, new_new_n20205__,
    new_new_n20206__, new_new_n20207__, new_new_n20208__, new_new_n20209__,
    new_new_n20210__, new_new_n20211__, new_new_n20212__, new_new_n20213__,
    new_new_n20214__, new_new_n20215__, new_new_n20216__, new_new_n20217__,
    new_new_n20218__, new_new_n20219__, new_new_n20220__, new_new_n20221__,
    new_new_n20222__, new_new_n20223__, new_new_n20224__, new_new_n20225__,
    new_new_n20226__, new_new_n20227__, new_new_n20228__, new_new_n20229__,
    new_new_n20230__, new_new_n20231__, new_new_n20232__, new_new_n20233__,
    new_new_n20234__, new_new_n20235__, new_new_n20236__, new_new_n20237__,
    new_new_n20238__, new_new_n20239__, new_new_n20240__, new_new_n20241__,
    new_new_n20242__, new_new_n20243__, new_new_n20244__, new_new_n20245__,
    new_new_n20246__, new_new_n20247__, new_new_n20248__, new_new_n20249__,
    new_new_n20250__, new_new_n20251__, new_new_n20252__, new_new_n20253__,
    new_new_n20254__, new_new_n20255__, new_new_n20256__, new_new_n20257__,
    new_new_n20258__, new_new_n20259__, new_new_n20260__, new_new_n20261__,
    new_new_n20262__, new_new_n20263__, new_new_n20264__, new_new_n20265__,
    new_new_n20267__, new_new_n20268__, new_new_n20269__, new_new_n20270__,
    new_new_n20271__, new_new_n20272__, new_new_n20273__, new_new_n20274__,
    new_new_n20275__, new_new_n20276__, new_new_n20277__, new_new_n20278__,
    new_new_n20279__, new_new_n20280__, new_new_n20281__, new_new_n20282__,
    new_new_n20283__, new_new_n20284__, new_new_n20285__, new_new_n20286__,
    new_new_n20287__, new_new_n20288__, new_new_n20289__, new_new_n20290__,
    new_new_n20291__, new_new_n20292__, new_new_n20293__, new_new_n20294__,
    new_new_n20295__, new_new_n20296__, new_new_n20297__, new_new_n20298__,
    new_new_n20299__, new_new_n20300__, new_new_n20301__, new_new_n20302__,
    new_new_n20303__, new_new_n20304__, new_new_n20305__, new_new_n20306__,
    new_new_n20307__, new_new_n20308__, new_new_n20309__, new_new_n20310__,
    new_new_n20311__, new_new_n20312__, new_new_n20313__, new_new_n20314__,
    new_new_n20315__, new_new_n20316__, new_new_n20317__, new_new_n20318__,
    new_new_n20319__, new_new_n20320__, new_new_n20321__, new_new_n20322__,
    new_new_n20323__, new_new_n20324__, new_new_n20325__, new_new_n20326__,
    new_new_n20327__, new_new_n20328__, new_new_n20329__, new_new_n20330__,
    new_new_n20331__, new_new_n20333__, new_new_n20334__, new_new_n20335__,
    new_new_n20336__, new_new_n20337__, new_new_n20338__, new_new_n20339__,
    new_new_n20340__, new_new_n20341__, new_new_n20342__, new_new_n20343__,
    new_new_n20344__, new_new_n20345__, new_new_n20346__, new_new_n20347__,
    new_new_n20348__, new_new_n20349__, new_new_n20350__, new_new_n20351__,
    new_new_n20352__, new_new_n20353__, new_new_n20354__, new_new_n20355__,
    new_new_n20356__, new_new_n20357__, new_new_n20358__, new_new_n20359__,
    new_new_n20360__, new_new_n20361__, new_new_n20362__, new_new_n20363__,
    new_new_n20364__, new_new_n20365__, new_new_n20366__, new_new_n20367__,
    new_new_n20368__, new_new_n20369__, new_new_n20370__, new_new_n20371__,
    new_new_n20372__, new_new_n20373__, new_new_n20374__, new_new_n20375__,
    new_new_n20376__, new_new_n20377__, new_new_n20378__, new_new_n20379__,
    new_new_n20380__, new_new_n20381__, new_new_n20382__, new_new_n20383__,
    new_new_n20384__, new_new_n20385__, new_new_n20386__, new_new_n20387__,
    new_new_n20388__, new_new_n20389__, new_new_n20390__, new_new_n20391__,
    new_new_n20392__, new_new_n20393__, new_new_n20394__, new_new_n20395__,
    new_new_n20396__, new_new_n20397__, new_new_n20398__, new_new_n20399__,
    new_new_n20401__, new_new_n20402__, new_new_n20403__, new_new_n20404__,
    new_new_n20405__, new_new_n20406__, new_new_n20407__, new_new_n20408__,
    new_new_n20409__, new_new_n20410__, new_new_n20411__, new_new_n20412__,
    new_new_n20413__, new_new_n20414__, new_new_n20415__, new_new_n20416__,
    new_new_n20417__, new_new_n20418__, new_new_n20419__, new_new_n20420__,
    new_new_n20421__, new_new_n20422__, new_new_n20423__, new_new_n20424__,
    new_new_n20425__, new_new_n20426__, new_new_n20427__, new_new_n20428__,
    new_new_n20429__, new_new_n20430__, new_new_n20431__, new_new_n20432__,
    new_new_n20433__, new_new_n20434__, new_new_n20435__, new_new_n20436__,
    new_new_n20437__, new_new_n20438__, new_new_n20439__, new_new_n20440__,
    new_new_n20441__, new_new_n20442__, new_new_n20443__, new_new_n20444__,
    new_new_n20445__, new_new_n20446__, new_new_n20447__, new_new_n20448__,
    new_new_n20449__, new_new_n20450__, new_new_n20451__, new_new_n20452__,
    new_new_n20453__, new_new_n20454__, new_new_n20455__, new_new_n20456__,
    new_new_n20457__, new_new_n20458__, new_new_n20459__, new_new_n20460__,
    new_new_n20461__, new_new_n20462__, new_new_n20463__, new_new_n20464__,
    new_new_n20465__, new_new_n20466__, new_new_n20467__, new_new_n20469__,
    new_new_n20470__, new_new_n20471__, new_new_n20472__, new_new_n20473__,
    new_new_n20474__, new_new_n20475__, new_new_n20476__, new_new_n20477__,
    new_new_n20478__, new_new_n20479__, new_new_n20480__, new_new_n20481__,
    new_new_n20482__, new_new_n20483__, new_new_n20484__, new_new_n20485__,
    new_new_n20486__, new_new_n20487__, new_new_n20488__, new_new_n20489__,
    new_new_n20490__, new_new_n20491__, new_new_n20492__, new_new_n20493__,
    new_new_n20494__, new_new_n20495__, new_new_n20496__, new_new_n20497__,
    new_new_n20498__, new_new_n20499__, new_new_n20500__, new_new_n20501__,
    new_new_n20502__, new_new_n20503__, new_new_n20504__, new_new_n20505__,
    new_new_n20506__, new_new_n20507__, new_new_n20508__, new_new_n20509__,
    new_new_n20510__, new_new_n20511__, new_new_n20512__, new_new_n20513__,
    new_new_n20514__, new_new_n20515__, new_new_n20516__, new_new_n20517__,
    new_new_n20518__, new_new_n20519__, new_new_n20520__, new_new_n20521__,
    new_new_n20522__, new_new_n20523__, new_new_n20524__, new_new_n20525__,
    new_new_n20526__, new_new_n20527__, new_new_n20528__, new_new_n20529__,
    new_new_n20530__, new_new_n20531__, new_new_n20532__, new_new_n20533__,
    new_new_n20534__, new_new_n20535__, new_new_n20537__, new_new_n20538__,
    new_new_n20539__, new_new_n20540__, new_new_n20541__, new_new_n20542__,
    new_new_n20543__, new_new_n20544__, new_new_n20545__, new_new_n20546__,
    new_new_n20547__, new_new_n20548__, new_new_n20549__, new_new_n20550__,
    new_new_n20551__, new_new_n20552__, new_new_n20553__, new_new_n20554__,
    new_new_n20555__, new_new_n20556__, new_new_n20557__, new_new_n20558__,
    new_new_n20559__, new_new_n20560__, new_new_n20561__, new_new_n20562__,
    new_new_n20563__, new_new_n20564__, new_new_n20565__, new_new_n20566__,
    new_new_n20567__, new_new_n20568__, new_new_n20569__, new_new_n20570__,
    new_new_n20571__, new_new_n20572__, new_new_n20573__, new_new_n20574__,
    new_new_n20575__, new_new_n20576__, new_new_n20577__, new_new_n20578__,
    new_new_n20579__, new_new_n20580__, new_new_n20581__, new_new_n20582__,
    new_new_n20583__, new_new_n20584__, new_new_n20585__, new_new_n20586__,
    new_new_n20587__, new_new_n20588__, new_new_n20589__, new_new_n20590__,
    new_new_n20591__, new_new_n20592__, new_new_n20593__, new_new_n20594__,
    new_new_n20595__, new_new_n20596__, new_new_n20597__, new_new_n20598__,
    new_new_n20599__, new_new_n20600__, new_new_n20601__, new_new_n20603__,
    new_new_n20604__, new_new_n20605__, new_new_n20606__, new_new_n20607__,
    new_new_n20608__, new_new_n20609__, new_new_n20610__, new_new_n20611__,
    new_new_n20612__, new_new_n20613__, new_new_n20614__, new_new_n20615__,
    new_new_n20616__, new_new_n20617__, new_new_n20618__, new_new_n20619__,
    new_new_n20620__, new_new_n20621__, new_new_n20622__, new_new_n20623__,
    new_new_n20624__, new_new_n20625__, new_new_n20626__, new_new_n20627__,
    new_new_n20628__, new_new_n20629__, new_new_n20630__, new_new_n20631__,
    new_new_n20632__, new_new_n20633__, new_new_n20634__, new_new_n20635__,
    new_new_n20636__, new_new_n20637__, new_new_n20638__, new_new_n20639__,
    new_new_n20640__, new_new_n20641__, new_new_n20642__, new_new_n20643__,
    new_new_n20644__, new_new_n20645__, new_new_n20646__, new_new_n20647__,
    new_new_n20648__, new_new_n20649__, new_new_n20650__, new_new_n20651__,
    new_new_n20652__, new_new_n20653__, new_new_n20654__, new_new_n20655__,
    new_new_n20656__, new_new_n20657__, new_new_n20658__, new_new_n20659__,
    new_new_n20660__, new_new_n20661__, new_new_n20662__, new_new_n20663__,
    new_new_n20664__, new_new_n20666__, new_new_n20667__, new_new_n20668__,
    new_new_n20669__, new_new_n20670__, new_new_n20671__, new_new_n20672__,
    new_new_n20673__, new_new_n20674__, new_new_n20675__, new_new_n20676__,
    new_new_n20677__, new_new_n20678__, new_new_n20679__, new_new_n20680__,
    new_new_n20681__, new_new_n20682__, new_new_n20683__, new_new_n20684__,
    new_new_n20685__, new_new_n20686__, new_new_n20687__, new_new_n20688__,
    new_new_n20689__, new_new_n20690__, new_new_n20691__, new_new_n20692__,
    new_new_n20693__, new_new_n20694__, new_new_n20695__, new_new_n20696__,
    new_new_n20697__, new_new_n20698__, new_new_n20699__, new_new_n20700__,
    new_new_n20701__, new_new_n20702__, new_new_n20703__, new_new_n20704__,
    new_new_n20705__, new_new_n20706__, new_new_n20707__, new_new_n20708__,
    new_new_n20709__, new_new_n20710__, new_new_n20711__, new_new_n20712__,
    new_new_n20713__, new_new_n20714__, new_new_n20715__, new_new_n20716__,
    new_new_n20717__, new_new_n20718__, new_new_n20719__, new_new_n20720__,
    new_new_n20721__, new_new_n20722__, new_new_n20723__, new_new_n20724__,
    new_new_n20725__, new_new_n20726__, new_new_n20727__, new_new_n20729__,
    new_new_n20730__, new_new_n20731__, new_new_n20732__, new_new_n20733__,
    new_new_n20734__, new_new_n20735__, new_new_n20736__, new_new_n20737__,
    new_new_n20738__, new_new_n20739__, new_new_n20740__, new_new_n20741__,
    new_new_n20742__, new_new_n20743__, new_new_n20744__, new_new_n20745__,
    new_new_n20746__, new_new_n20747__, new_new_n20748__, new_new_n20749__,
    new_new_n20750__, new_new_n20751__, new_new_n20752__, new_new_n20753__,
    new_new_n20754__, new_new_n20755__, new_new_n20756__, new_new_n20757__,
    new_new_n20758__, new_new_n20759__, new_new_n20760__, new_new_n20761__,
    new_new_n20762__, new_new_n20763__, new_new_n20764__, new_new_n20765__,
    new_new_n20766__, new_new_n20767__, new_new_n20768__, new_new_n20769__,
    new_new_n20770__, new_new_n20771__, new_new_n20772__, new_new_n20773__,
    new_new_n20774__, new_new_n20775__, new_new_n20776__, new_new_n20777__,
    new_new_n20778__, new_new_n20779__, new_new_n20780__, new_new_n20781__,
    new_new_n20782__, new_new_n20783__, new_new_n20784__, new_new_n20785__,
    new_new_n20786__, new_new_n20787__, new_new_n20788__, new_new_n20790__,
    new_new_n20792__, new_new_n20794__, new_new_n20796__, new_new_n20798__,
    new_new_n20800__, new_new_n20802__, new_new_n20804__, new_new_n20806__,
    new_new_n20808__, new_new_n20810__, new_new_n20812__, new_new_n20814__,
    new_new_n20816__, new_new_n20818__, new_new_n20820__, new_new_n20822__,
    new_new_n20824__, new_new_n20826__, new_new_n20828__, new_new_n20830__,
    new_new_n20832__, new_new_n20834__, new_new_n20836__, new_new_n20838__,
    new_new_n20840__, new_new_n20842__, new_new_n20844__, new_new_n20846__,
    new_new_n20848__, new_new_n20849__, new_new_n20851__, new_new_n20852__,
    new_new_n20854__, new_new_n20855__, new_new_n20856__, new_new_n20857__,
    new_new_n20858__, new_new_n20859__, new_new_n20860__, new_new_n20861__,
    new_new_n20862__, new_new_n20863__, new_new_n20865__, new_new_n20866__,
    new_new_n20867__, new_new_n20868__, new_new_n20869__, new_new_n20870__,
    new_new_n20871__, new_new_n20872__, new_new_n20873__, new_new_n20875__,
    new_new_n20876__, new_new_n20877__, new_new_n20878__, new_new_n20879__,
    new_new_n20880__, new_new_n20881__, new_new_n20882__, new_new_n20884__,
    new_new_n20885__, new_new_n20886__, new_new_n20887__, new_new_n20888__,
    new_new_n20889__, new_new_n20890__, new_new_n20891__, new_new_n20893__,
    new_new_n20894__, new_new_n20895__, new_new_n20896__, new_new_n20897__,
    new_new_n20898__, new_new_n20899__, new_new_n20900__, new_new_n20902__,
    new_new_n20903__, new_new_n20904__, new_new_n20905__, new_new_n20906__,
    new_new_n20907__, new_new_n20908__, new_new_n20909__, new_new_n20911__,
    new_new_n20912__, new_new_n20913__, new_new_n20914__, new_new_n20915__,
    new_new_n20916__, new_new_n20917__, new_new_n20918__, new_new_n20920__,
    new_new_n20921__, new_new_n20922__, new_new_n20923__, new_new_n20924__,
    new_new_n20925__, new_new_n20926__, new_new_n20927__, new_new_n20929__,
    new_new_n20930__, new_new_n20931__, new_new_n20932__, new_new_n20933__,
    new_new_n20934__, new_new_n20935__, new_new_n20936__, new_new_n20938__,
    new_new_n20939__, new_new_n20940__, new_new_n20941__, new_new_n20942__,
    new_new_n20943__, new_new_n20944__, new_new_n20946__, new_new_n20947__,
    new_new_n20948__, new_new_n20949__, new_new_n20950__, new_new_n20951__,
    new_new_n20952__, new_new_n20954__, new_new_n20955__, new_new_n20956__,
    new_new_n20957__, new_new_n20958__, new_new_n20959__, new_new_n20960__,
    new_new_n20962__, new_new_n20963__, new_new_n20964__, new_new_n20965__,
    new_new_n20966__, new_new_n20967__, new_new_n20968__, new_new_n20970__,
    new_new_n20971__, new_new_n20972__, new_new_n20973__, new_new_n20974__,
    new_new_n20975__, new_new_n20976__, new_new_n20978__, new_new_n20979__,
    new_new_n20980__, new_new_n20981__, new_new_n20982__, new_new_n20983__,
    new_new_n20984__, new_new_n20986__, new_new_n20987__, new_new_n20988__,
    new_new_n20989__, new_new_n20990__, new_new_n20991__, new_new_n20992__,
    new_new_n20994__, new_new_n20995__, new_new_n20996__, new_new_n20997__,
    new_new_n20998__, new_new_n20999__, new_new_n21000__, new_new_n21002__,
    new_new_n21003__, new_new_n21004__, new_new_n21005__, new_new_n21006__,
    new_new_n21007__, new_new_n21009__, new_new_n21010__, new_new_n21011__,
    new_new_n21012__, new_new_n21013__, new_new_n21014__, new_new_n21016__,
    new_new_n21017__, new_new_n21018__, new_new_n21019__, new_new_n21020__,
    new_new_n21021__, new_new_n21023__, new_new_n21024__, new_new_n21025__,
    new_new_n21026__, new_new_n21027__, new_new_n21028__, new_new_n21030__,
    new_new_n21031__, new_new_n21032__, new_new_n21033__, new_new_n21034__,
    new_new_n21035__, new_new_n21037__, new_new_n21038__, new_new_n21039__,
    new_new_n21040__, new_new_n21041__, new_new_n21042__, new_new_n21044__,
    new_new_n21045__, new_new_n21046__, new_new_n21047__, new_new_n21048__,
    new_new_n21049__, new_new_n21051__, new_new_n21052__, new_new_n21053__,
    new_new_n21054__, new_new_n21055__, new_new_n21056__, new_new_n21058__,
    new_new_n21059__, new_new_n21060__, new_new_n21061__, new_new_n21062__,
    new_new_n21063__, new_new_n21065__, new_new_n21066__, new_new_n21067__,
    new_new_n21068__, new_new_n21069__, new_new_n21070__, new_new_n21072__,
    new_new_n21073__, new_new_n21074__, new_new_n21075__, new_new_n21076__,
    new_new_n21077__, new_new_n21079__, new_new_n21080__, new_new_n21081__,
    new_new_n21082__, new_new_n21083__, new_new_n21084__, new_new_n21086__,
    new_new_n21087__, new_new_n21088__, new_new_n21089__, new_new_n21090__,
    new_new_n21091__, new_new_n21093__, new_new_n21094__, new_new_n21095__,
    new_new_n21096__, new_new_n21097__, new_new_n21098__, new_new_n21100__,
    new_new_n21101__, new_new_n21102__, new_new_n21103__, new_new_n21104__,
    new_new_n21105__, new_new_n21107__, new_new_n21108__, new_new_n21109__,
    new_new_n21110__, new_new_n21111__, new_new_n21112__, new_new_n21114__,
    new_new_n21115__, new_new_n21116__, new_new_n21117__, new_new_n21118__,
    new_new_n21119__, new_new_n21121__, new_new_n21122__, new_new_n21123__,
    new_new_n21124__, new_new_n21125__, new_new_n21126__, new_new_n21128__,
    new_new_n21129__, new_new_n21130__, new_new_n21131__, new_new_n21132__,
    new_new_n21133__, new_new_n21135__, new_new_n21136__, new_new_n21137__,
    new_new_n21138__, new_new_n21139__, new_new_n21140__, new_new_n21142__,
    new_new_n21143__, new_new_n21144__, new_new_n21145__, new_new_n21146__,
    new_new_n21147__, new_new_n21149__, new_new_n21150__, new_new_n21151__,
    new_new_n21152__, new_new_n21153__, new_new_n21154__, new_new_n21156__,
    new_new_n21157__, new_new_n21158__, new_new_n21159__, new_new_n21160__,
    new_new_n21161__, new_new_n21163__, new_new_n21164__, new_new_n21165__,
    new_new_n21166__, new_new_n21167__, new_new_n21168__, new_new_n21170__,
    new_new_n21171__, new_new_n21172__, new_new_n21173__, new_new_n21174__,
    new_new_n21175__, new_new_n21177__, new_new_n21178__, new_new_n21179__,
    new_new_n21180__, new_new_n21181__, new_new_n21182__, new_new_n21184__,
    new_new_n21185__, new_new_n21186__, new_new_n21187__, new_new_n21188__,
    new_new_n21189__, new_new_n21191__, new_new_n21192__, new_new_n21193__,
    new_new_n21194__, new_new_n21195__, new_new_n21196__, new_new_n21198__,
    new_new_n21199__, new_new_n21200__, new_new_n21201__, new_new_n21202__,
    new_new_n21203__, new_new_n21205__, new_new_n21206__, new_new_n21207__,
    new_new_n21208__, new_new_n21209__, new_new_n21210__, new_new_n21212__,
    new_new_n21213__, new_new_n21214__, new_new_n21215__, new_new_n21216__,
    new_new_n21217__, new_new_n21219__, new_new_n21220__, new_new_n21221__,
    new_new_n21222__, new_new_n21223__, new_new_n21224__, new_new_n21226__,
    new_new_n21227__, new_new_n21228__, new_new_n21229__, new_new_n21230__,
    new_new_n21231__, new_new_n21233__, new_new_n21234__, new_new_n21235__,
    new_new_n21236__, new_new_n21237__, new_new_n21238__, new_new_n21240__,
    new_new_n21241__, new_new_n21242__, new_new_n21243__, new_new_n21244__,
    new_new_n21245__, new_new_n21247__, new_new_n21248__, new_new_n21249__,
    new_new_n21250__, new_new_n21251__, new_new_n21252__, new_new_n21254__,
    new_new_n21255__, new_new_n21256__, new_new_n21257__, new_new_n21258__,
    new_new_n21259__, new_new_n21261__, new_new_n21262__, new_new_n21263__,
    new_new_n21264__, new_new_n21265__, new_new_n21266__, new_new_n21268__,
    new_new_n21269__, new_new_n21270__, new_new_n21271__, new_new_n21272__,
    new_new_n21273__, new_new_n21275__, new_new_n21276__, new_new_n21277__,
    new_new_n21278__, new_new_n21279__, new_new_n21280__, new_new_n21282__,
    new_new_n21283__, new_new_n21284__, new_new_n21285__, new_new_n21286__,
    new_new_n21287__, new_new_n21289__, new_new_n21290__, new_new_n21291__,
    new_new_n21292__, new_new_n21293__, new_new_n21294__, new_new_n21296__,
    new_new_n21297__, new_new_n21298__, new_new_n21299__, new_new_n21300__,
    new_new_n21301__, new_new_n21303__, new_new_n21304__, new_new_n21305__,
    new_new_n21306__, new_new_n21307__, new_new_n21308__, new_new_n21310__,
    new_new_n21311__, new_new_n21312__, new_new_n21313__, new_new_n21314__,
    new_new_n21315__, new_new_n21317__, new_new_n21318__, new_new_n21319__,
    new_new_n21320__, new_new_n21321__, new_new_n21322__, new_new_n21324__,
    new_new_n21325__, new_new_n21326__, new_new_n21327__, new_new_n21328__,
    new_new_n21329__, new_new_n21331__, new_new_n21332__, new_new_n21333__,
    new_new_n21334__, new_new_n21335__, new_new_n21336__, new_new_n21338__,
    new_new_n21339__, new_new_n21340__, new_new_n21341__, new_new_n21342__,
    new_new_n21343__, new_new_n21344__, new_new_n21345__, new_new_n21346__,
    new_new_n21347__, new_new_n21348__, new_new_n21350__, new_new_n21351__,
    new_new_n21353__, new_new_n21354__, new_new_n21356__, new_new_n21357__,
    new_new_n21359__, new_new_n21360__, new_new_n21361__, new_new_n21362__,
    new_new_n21364__, new_new_n21365__, new_new_n21367__, new_new_n21368__,
    new_new_n21369__, new_new_n21371__, new_new_n21372__, new_new_n21373__,
    new_new_n21375__, new_new_n21376__, new_new_n21377__, new_new_n21379__,
    new_new_n21380__, new_new_n21382__, new_new_n21383__, new_new_n21384__,
    new_new_n21386__, new_new_n21387__, new_new_n21388__, new_new_n21390__,
    new_new_n21391__, new_new_n21392__, new_new_n21394__, new_new_n21395__,
    new_new_n21396__, new_new_n21398__, new_new_n21399__, new_new_n21400__,
    new_new_n21402__, new_new_n21403__, new_new_n21404__, new_new_n21406__,
    new_new_n21407__, new_new_n21408__, new_new_n21410__, new_new_n21411__,
    new_new_n21413__, new_new_n21414__, new_new_n21415__, new_new_n21416__,
    new_new_n21417__, new_new_n21419__, new_new_n21420__, new_new_n21421__,
    new_new_n21422__, new_new_n21423__, new_new_n21425__, new_new_n21426__,
    new_new_n21427__, new_new_n21428__, new_new_n21429__, new_new_n21430__,
    new_new_n21432__, new_new_n21433__, new_new_n21434__, new_new_n21435__,
    new_new_n21436__, new_new_n21438__, new_new_n21439__, new_new_n21440__,
    new_new_n21441__, new_new_n21442__, new_new_n21443__, new_new_n21445__,
    new_new_n21446__, new_new_n21447__, new_new_n21448__, new_new_n21449__,
    new_new_n21450__, new_new_n21452__, new_new_n21453__, new_new_n21454__,
    new_new_n21455__, new_new_n21456__, new_new_n21457__, new_new_n21459__,
    new_new_n21460__, new_new_n21461__, new_new_n21462__, new_new_n21463__,
    new_new_n21465__, new_new_n21466__, new_new_n21467__, new_new_n21468__,
    new_new_n21469__, new_new_n21470__, new_new_n21472__, new_new_n21473__,
    new_new_n21474__, new_new_n21475__, new_new_n21476__, new_new_n21477__,
    new_new_n21479__, new_new_n21480__, new_new_n21481__, new_new_n21482__,
    new_new_n21483__, new_new_n21484__, new_new_n21486__, new_new_n21487__,
    new_new_n21488__, new_new_n21489__, new_new_n21490__, new_new_n21492__,
    new_new_n21493__, new_new_n21494__, new_new_n21495__, new_new_n21496__,
    new_new_n21497__, new_new_n21498__, new_new_n21499__, new_new_n21500__,
    new_new_n21501__, new_new_n21502__, new_new_n21503__, new_new_n21504__,
    new_new_n21505__, new_new_n21506__, new_new_n21507__, new_new_n21509__,
    new_new_n21510__, new_new_n21511__, new_new_n21512__, new_new_n21513__,
    new_new_n21515__, new_new_n21516__, new_new_n21517__, new_new_n21518__,
    new_new_n21519__, new_new_n21520__, new_new_n21521__, new_new_n21522__,
    new_new_n21523__, new_new_n21524__, new_new_n21525__, new_new_n21526__,
    new_new_n21527__, new_new_n21528__, new_new_n21529__, new_new_n21530__,
    new_new_n21531__, new_new_n21532__, new_new_n21533__, new_new_n21534__,
    new_new_n21535__, new_new_n21536__, new_new_n21537__, new_new_n21538__,
    new_new_n21539__, new_new_n21540__, new_new_n21541__, new_new_n21542__,
    new_new_n21543__, new_new_n21544__, new_new_n21545__, new_new_n21546__,
    new_new_n21547__, new_new_n21548__, new_new_n21549__, new_new_n21550__,
    new_new_n21551__, new_new_n21552__, new_new_n21553__, new_new_n21554__,
    new_new_n21555__, new_new_n21556__, new_new_n21557__, new_new_n21558__,
    new_new_n21559__, new_new_n21560__, new_new_n21561__, new_new_n21562__,
    new_new_n21563__, new_new_n21564__, new_new_n21565__, new_new_n21566__,
    new_new_n21567__, new_new_n21568__, new_new_n21569__, new_new_n21570__,
    new_new_n21571__, new_new_n21572__, new_new_n21573__, new_new_n21574__,
    new_new_n21575__, new_new_n21576__, new_new_n21577__, new_new_n21578__,
    new_new_n21579__, new_new_n21580__, new_new_n21581__, new_new_n21582__,
    new_new_n21583__, new_new_n21584__, new_new_n21585__, new_new_n21586__,
    new_new_n21587__, new_new_n21588__, new_new_n21589__, new_new_n21590__,
    new_new_n21591__, new_new_n21592__, new_new_n21593__, new_new_n21594__,
    new_new_n21596__, new_new_n21597__, new_new_n21598__, new_new_n21599__,
    new_new_n21600__, new_new_n21601__, new_new_n21602__, new_new_n21603__,
    new_new_n21604__, new_new_n21605__, new_new_n21606__, new_new_n21607__,
    new_new_n21608__, new_new_n21609__, new_new_n21611__, new_new_n21612__,
    new_new_n21613__, new_new_n21614__, new_new_n21615__, new_new_n21616__,
    new_new_n21617__, new_new_n21618__, new_new_n21619__, new_new_n21620__,
    new_new_n21621__, new_new_n21622__, new_new_n21623__, new_new_n21624__,
    new_new_n21626__, new_new_n21627__, new_new_n21628__, new_new_n21629__,
    new_new_n21630__, new_new_n21631__, new_new_n21632__, new_new_n21633__,
    new_new_n21634__, new_new_n21635__, new_new_n21636__, new_new_n21637__,
    new_new_n21638__, new_new_n21639__, new_new_n21641__, new_new_n21642__,
    new_new_n21643__, new_new_n21644__, new_new_n21645__, new_new_n21646__,
    new_new_n21647__, new_new_n21648__, new_new_n21649__, new_new_n21650__,
    new_new_n21651__, new_new_n21652__, new_new_n21653__, new_new_n21654__,
    new_new_n21656__, new_new_n21657__, new_new_n21658__, new_new_n21659__,
    new_new_n21660__, new_new_n21662__, new_new_n21663__, new_new_n21664__,
    new_new_n21665__, new_new_n21666__, new_new_n21667__, new_new_n21668__,
    new_new_n21669__, new_new_n21670__, new_new_n21671__, new_new_n21672__,
    new_new_n21673__, new_new_n21674__, new_new_n21675__, new_new_n21676__,
    new_new_n21677__, new_new_n21678__, new_new_n21679__, new_new_n21680__,
    new_new_n21681__, new_new_n21682__, new_new_n21683__, new_new_n21684__,
    new_new_n21685__, new_new_n21686__, new_new_n21687__, new_new_n21688__,
    new_new_n21689__, new_new_n21690__, new_new_n21691__, new_new_n21692__,
    new_new_n21693__, new_new_n21694__, new_new_n21695__, new_new_n21696__,
    new_new_n21697__, new_new_n21698__, new_new_n21699__, new_new_n21700__,
    new_new_n21701__, new_new_n21702__, new_new_n21703__, new_new_n21704__,
    new_new_n21705__, new_new_n21706__, new_new_n21707__, new_new_n21708__,
    new_new_n21709__, new_new_n21710__, new_new_n21711__, new_new_n21712__,
    new_new_n21713__, new_new_n21714__, new_new_n21715__, new_new_n21716__,
    new_new_n21717__, new_new_n21718__, new_new_n21719__, new_new_n21720__,
    new_new_n21721__, new_new_n21722__, new_new_n21723__, new_new_n21724__,
    new_new_n21725__, new_new_n21726__, new_new_n21727__, new_new_n21728__,
    new_new_n21729__, new_new_n21730__, new_new_n21731__, new_new_n21732__,
    new_new_n21733__, new_new_n21734__, new_new_n21735__, new_new_n21736__,
    new_new_n21737__, new_new_n21738__, new_new_n21739__, new_new_n21740__,
    new_new_n21741__, new_new_n21743__, new_new_n21744__, new_new_n21745__,
    new_new_n21746__, new_new_n21747__, new_new_n21748__, new_new_n21749__,
    new_new_n21750__, new_new_n21751__, new_new_n21752__, new_new_n21753__,
    new_new_n21754__, new_new_n21755__, new_new_n21756__, new_new_n21758__,
    new_new_n21759__, new_new_n21760__, new_new_n21761__, new_new_n21762__,
    new_new_n21763__, new_new_n21764__, new_new_n21765__, new_new_n21766__,
    new_new_n21767__, new_new_n21768__, new_new_n21769__, new_new_n21770__,
    new_new_n21771__, new_new_n21773__, new_new_n21774__, new_new_n21775__,
    new_new_n21776__, new_new_n21777__, new_new_n21778__, new_new_n21779__,
    new_new_n21780__, new_new_n21781__, new_new_n21782__, new_new_n21783__,
    new_new_n21784__, new_new_n21785__, new_new_n21786__, new_new_n21788__,
    new_new_n21789__, new_new_n21790__, new_new_n21791__, new_new_n21792__,
    new_new_n21793__, new_new_n21794__, new_new_n21795__, new_new_n21796__,
    new_new_n21797__, new_new_n21798__, new_new_n21799__, new_new_n21800__,
    new_new_n21801__, new_new_n21803__, new_new_n21804__, new_new_n21805__,
    new_new_n21806__, new_new_n21807__, new_new_n21809__, new_new_n21810__,
    new_new_n21811__, new_new_n21812__, new_new_n21813__, new_new_n21814__,
    new_new_n21815__, new_new_n21816__, new_new_n21817__, new_new_n21818__,
    new_new_n21819__, new_new_n21820__, new_new_n21821__, new_new_n21822__,
    new_new_n21823__, new_new_n21824__, new_new_n21825__, new_new_n21826__,
    new_new_n21827__, new_new_n21828__, new_new_n21829__, new_new_n21830__,
    new_new_n21831__, new_new_n21832__, new_new_n21833__, new_new_n21834__,
    new_new_n21835__, new_new_n21836__, new_new_n21837__, new_new_n21838__,
    new_new_n21839__, new_new_n21840__, new_new_n21841__, new_new_n21842__,
    new_new_n21843__, new_new_n21844__, new_new_n21845__, new_new_n21846__,
    new_new_n21847__, new_new_n21848__, new_new_n21849__, new_new_n21850__,
    new_new_n21851__, new_new_n21852__, new_new_n21853__, new_new_n21854__,
    new_new_n21855__, new_new_n21856__, new_new_n21857__, new_new_n21858__,
    new_new_n21859__, new_new_n21860__, new_new_n21861__, new_new_n21862__,
    new_new_n21863__, new_new_n21864__, new_new_n21865__, new_new_n21866__,
    new_new_n21867__, new_new_n21868__, new_new_n21869__, new_new_n21870__,
    new_new_n21871__, new_new_n21872__, new_new_n21873__, new_new_n21874__,
    new_new_n21875__, new_new_n21876__, new_new_n21877__, new_new_n21878__,
    new_new_n21879__, new_new_n21880__, new_new_n21881__, new_new_n21882__,
    new_new_n21883__, new_new_n21884__, new_new_n21885__, new_new_n21886__,
    new_new_n21887__, new_new_n21888__, new_new_n21890__, new_new_n21891__,
    new_new_n21892__, new_new_n21893__, new_new_n21894__, new_new_n21895__,
    new_new_n21896__, new_new_n21897__, new_new_n21898__, new_new_n21899__,
    new_new_n21900__, new_new_n21901__, new_new_n21902__, new_new_n21903__,
    new_new_n21905__, new_new_n21906__, new_new_n21907__, new_new_n21908__,
    new_new_n21909__, new_new_n21910__, new_new_n21911__, new_new_n21912__,
    new_new_n21913__, new_new_n21914__, new_new_n21915__, new_new_n21916__,
    new_new_n21917__, new_new_n21918__, new_new_n21920__, new_new_n21921__,
    new_new_n21922__, new_new_n21923__, new_new_n21924__, new_new_n21925__,
    new_new_n21926__, new_new_n21927__, new_new_n21928__, new_new_n21929__,
    new_new_n21930__, new_new_n21931__, new_new_n21932__, new_new_n21933__,
    new_new_n21935__, new_new_n21936__, new_new_n21937__, new_new_n21938__,
    new_new_n21939__, new_new_n21940__, new_new_n21941__, new_new_n21942__,
    new_new_n21943__, new_new_n21944__, new_new_n21945__, new_new_n21946__,
    new_new_n21947__, new_new_n21948__, new_new_n21950__, new_new_n21951__,
    new_new_n21952__, new_new_n21953__, new_new_n21954__, new_new_n21957__,
    new_new_n21958__, new_new_n21959__, new_new_n21960__, new_new_n21961__,
    new_new_n21962__, new_new_n21963__, new_new_n21964__, new_new_n21965__,
    new_new_n21968__, new_new_n21969__, new_new_n21971__, new_new_n21972__,
    new_new_n21973__, new_new_n21974__, new_new_n21975__, new_new_n21976__,
    new_new_n21977__, new_new_n21978__, new_new_n21979__, new_new_n21980__,
    new_new_n21981__, new_new_n21983__, new_new_n21984__, new_new_n21985__,
    new_new_n21986__, new_new_n21987__, new_new_n21988__, new_new_n21989__,
    new_new_n21990__, new_new_n21991__, new_new_n21992__, new_new_n21993__,
    new_new_n21994__, new_new_n21995__, new_new_n21996__, new_new_n21997__,
    new_new_n21998__, new_new_n21999__, new_new_n22000__, new_new_n22001__,
    new_new_n22002__, new_new_n22003__, new_new_n22004__, new_new_n22005__,
    new_new_n22006__, new_new_n22007__, new_new_n22008__, new_new_n22010__,
    new_new_n22011__, new_new_n22012__, new_new_n22013__, new_new_n22014__,
    new_new_n22015__, new_new_n22016__, new_new_n22017__, new_new_n22019__,
    new_new_n22020__, new_new_n22021__, new_new_n22022__, new_new_n22023__,
    new_new_n22024__, new_new_n22026__, new_new_n22027__, new_new_n22029__,
    new_new_n22030__, new_new_n22031__, new_new_n22033__, new_new_n22034__,
    new_new_n22035__, new_new_n22036__, new_new_n22037__, new_new_n22038__,
    new_new_n22039__, new_new_n22040__, new_new_n22041__, new_new_n22042__,
    new_new_n22043__, new_new_n22044__, new_new_n22045__, new_new_n22046__,
    new_new_n22047__, new_new_n22048__, new_new_n22050__, new_new_n22051__,
    new_new_n22052__, new_new_n22053__, new_new_n22054__, new_new_n22055__,
    new_new_n22056__, new_new_n22058__, new_new_n22059__, new_new_n22060__,
    new_new_n22061__, new_new_n22062__, new_new_n22063__, new_new_n22064__,
    new_new_n22065__, new_new_n22066__, new_new_n22067__, new_new_n22068__,
    new_new_n22069__, new_new_n22070__, new_new_n22072__, new_new_n22073__,
    new_new_n22074__, new_new_n22075__, new_new_n22076__, new_new_n22077__,
    new_new_n22080__, new_new_n22081__, new_new_n22082__, new_new_n22083__,
    new_new_n22085__, new_new_n22086__, new_new_n22087__, new_new_n22088__,
    new_new_n22089__, new_new_n22090__, new_new_n22091__, new_new_n22092__,
    new_new_n22093__, new_new_n22094__, new_new_n22095__, new_new_n22096__,
    new_new_n22097__, new_new_n22098__, new_new_n22099__, new_new_n22100__,
    new_new_n22101__, new_new_n22102__, new_new_n22103__, new_new_n22104__,
    new_new_n22105__, new_new_n22106__, new_new_n22107__, new_new_n22110__,
    new_new_n22111__, new_new_n22112__, new_new_n22113__, new_new_n22114__,
    new_new_n22115__, new_new_n22116__, new_new_n22117__, new_new_n22118__,
    new_new_n22121__, new_new_n22122__, new_new_n22124__, new_new_n22125__,
    new_new_n22126__, new_new_n22127__, new_new_n22128__, new_new_n22129__,
    new_new_n22130__, new_new_n22131__, new_new_n22132__, new_new_n22133__,
    new_new_n22134__, new_new_n22136__, new_new_n22137__, new_new_n22138__,
    new_new_n22139__, new_new_n22140__, new_new_n22141__, new_new_n22143__,
    new_new_n22144__, new_new_n22145__, new_new_n22146__, new_new_n22147__,
    new_new_n22148__, new_new_n22149__, new_new_n22150__, new_new_n22151__,
    new_new_n22152__, new_new_n22153__, new_new_n22154__, new_new_n22155__,
    new_new_n22156__, new_new_n22157__, new_new_n22158__, new_new_n22159__,
    new_new_n22160__, new_new_n22161__, new_new_n22162__, new_new_n22163__,
    new_new_n22164__, new_new_n22165__, new_new_n22166__, new_new_n22167__,
    new_new_n22168__, new_new_n22170__, new_new_n22171__, new_new_n22172__,
    new_new_n22173__, new_new_n22174__, new_new_n22175__, new_new_n22176__,
    new_new_n22177__, new_new_n22178__, new_new_n22180__, new_new_n22181__,
    new_new_n22182__, new_new_n22183__, new_new_n22184__, new_new_n22185__,
    new_new_n22186__, new_new_n22187__, new_new_n22188__, new_new_n22189__,
    new_new_n22190__, new_new_n22191__, new_new_n22192__, new_new_n22193__,
    new_new_n22194__, new_new_n22195__, new_new_n22196__, new_new_n22197__,
    new_new_n22198__, new_new_n22199__, new_new_n22200__, new_new_n22201__,
    new_new_n22202__, new_new_n22203__, new_new_n22204__, new_new_n22205__,
    new_new_n22206__, new_new_n22207__, new_new_n22209__, new_new_n22210__,
    new_new_n22211__, new_new_n22212__, new_new_n22213__, new_new_n22214__,
    new_new_n22215__, new_new_n22216__, new_new_n22218__, new_new_n22219__,
    new_new_n22220__, new_new_n22221__, new_new_n22222__, new_new_n22223__,
    new_new_n22224__, new_new_n22225__, new_new_n22226__, new_new_n22227__,
    new_new_n22228__, new_new_n22229__, new_new_n22230__, new_new_n22231__,
    new_new_n22232__, new_new_n22233__, new_new_n22234__, new_new_n22235__,
    new_new_n22236__, new_new_n22237__, new_new_n22238__, new_new_n22239__,
    new_new_n22240__, new_new_n22241__, new_new_n22242__, new_new_n22243__,
    new_new_n22244__, new_new_n22245__, new_new_n22247__, new_new_n22248__,
    new_new_n22249__, new_new_n22250__, new_new_n22251__, new_new_n22252__,
    new_new_n22253__, new_new_n22254__, new_new_n22256__, new_new_n22257__,
    new_new_n22258__, new_new_n22259__, new_new_n22260__, new_new_n22261__,
    new_new_n22262__, new_new_n22263__, new_new_n22264__, new_new_n22265__,
    new_new_n22266__, new_new_n22267__, new_new_n22268__, new_new_n22269__,
    new_new_n22270__, new_new_n22271__, new_new_n22272__, new_new_n22273__,
    new_new_n22274__, new_new_n22275__, new_new_n22276__, new_new_n22277__,
    new_new_n22278__, new_new_n22279__, new_new_n22280__, new_new_n22281__,
    new_new_n22282__, new_new_n22283__, new_new_n22284__, new_new_n22285__,
    new_new_n22286__, new_new_n22288__, new_new_n22289__, new_new_n22290__,
    new_new_n22291__, new_new_n22292__, new_new_n22293__, new_new_n22294__,
    new_new_n22295__, new_new_n22297__, new_new_n22298__, new_new_n22299__,
    new_new_n22300__, new_new_n22301__, new_new_n22302__, new_new_n22303__,
    new_new_n22304__, new_new_n22305__, new_new_n22306__, new_new_n22307__,
    new_new_n22308__, new_new_n22309__, new_new_n22310__, new_new_n22311__,
    new_new_n22312__, new_new_n22313__, new_new_n22314__, new_new_n22315__,
    new_new_n22316__, new_new_n22317__, new_new_n22318__, new_new_n22319__,
    new_new_n22320__, new_new_n22321__, new_new_n22322__, new_new_n22323__,
    new_new_n22324__, new_new_n22325__, new_new_n22327__, new_new_n22328__,
    new_new_n22329__, new_new_n22330__, new_new_n22331__, new_new_n22332__,
    new_new_n22333__, new_new_n22334__, new_new_n22336__, new_new_n22337__,
    new_new_n22338__, new_new_n22339__, new_new_n22340__, new_new_n22341__,
    new_new_n22342__, new_new_n22343__, new_new_n22344__, new_new_n22345__,
    new_new_n22346__, new_new_n22347__, new_new_n22348__, new_new_n22349__,
    new_new_n22350__, new_new_n22351__, new_new_n22352__, new_new_n22353__,
    new_new_n22354__, new_new_n22355__, new_new_n22356__, new_new_n22357__,
    new_new_n22358__, new_new_n22359__, new_new_n22360__, new_new_n22361__,
    new_new_n22362__, new_new_n22363__, new_new_n22364__, new_new_n22365__,
    new_new_n22366__, new_new_n22368__, new_new_n22369__, new_new_n22370__,
    new_new_n22371__, new_new_n22372__, new_new_n22373__, new_new_n22374__,
    new_new_n22375__, new_new_n22376__, new_new_n22377__, new_new_n22378__,
    new_new_n22380__, new_new_n22381__, new_new_n22382__, new_new_n22383__,
    new_new_n22384__, new_new_n22385__, new_new_n22386__, new_new_n22387__,
    new_new_n22388__, new_new_n22389__, new_new_n22390__, new_new_n22391__,
    new_new_n22392__, new_new_n22394__, new_new_n22395__, new_new_n22396__,
    new_new_n22398__, new_new_n22399__, new_new_n22400__, new_new_n22402__,
    new_new_n22403__, new_new_n22404__, new_new_n22405__, new_new_n22406__,
    new_new_n22407__, new_new_n22408__, new_new_n22409__, new_new_n22410__,
    new_new_n22411__, new_new_n22414__, new_new_n22415__, new_new_n22416__,
    new_new_n22417__, new_new_n22419__, new_new_n22420__, new_new_n22421__,
    new_new_n22422__, new_new_n22423__, new_new_n22425__, new_new_n22426__,
    new_new_n22428__, new_new_n22429__, new_new_n22430__, new_new_n22431__,
    new_new_n22432__, new_new_n22433__, new_new_n22434__, new_new_n22435__,
    new_new_n22436__, new_new_n22437__, new_new_n22438__, new_new_n22439__,
    new_new_n22440__, new_new_n22441__, new_new_n22442__, new_new_n22443__,
    new_new_n22444__, new_new_n22445__, new_new_n22446__, new_new_n22447__,
    new_new_n22448__, new_new_n22449__, new_new_n22450__, new_new_n22451__,
    new_new_n22452__, new_new_n22453__, new_new_n22454__, new_new_n22455__,
    new_new_n22456__, new_new_n22457__, new_new_n22458__, new_new_n22459__,
    new_new_n22460__, new_new_n22461__, new_new_n22462__, new_new_n22463__,
    new_new_n22464__, new_new_n22465__, new_new_n22466__, new_new_n22467__,
    new_new_n22468__, new_new_n22469__, new_new_n22470__, new_new_n22471__,
    new_new_n22472__, new_new_n22473__, new_new_n22474__, new_new_n22475__,
    new_new_n22476__, new_new_n22477__, new_new_n22478__, new_new_n22480__,
    new_new_n22481__, new_new_n22482__, new_new_n22483__, new_new_n22484__,
    new_new_n22485__, new_new_n22486__, new_new_n22487__, new_new_n22488__,
    new_new_n22489__, new_new_n22491__, new_new_n22492__, new_new_n22493__,
    new_new_n22494__, new_new_n22496__, new_new_n22498__, new_new_n22501__,
    new_new_n22502__, new_new_n22503__, new_new_n22505__, new_new_n22506__,
    new_new_n22507__, new_new_n22508__, new_new_n22509__, new_new_n22511__,
    new_new_n22512__, new_new_n22513__, new_new_n22514__, new_new_n22515__,
    new_new_n22516__, new_new_n22517__, new_new_n22518__, new_new_n22519__,
    new_new_n22520__, new_new_n22522__, new_new_n22523__, new_new_n22524__,
    new_new_n22525__, new_new_n22527__, new_new_n22528__, new_new_n22529__,
    new_new_n22530__, new_new_n22531__, new_new_n22534__, new_new_n22535__,
    new_new_n22536__, new_new_n22538__, new_new_n22539__, new_new_n22540__,
    new_new_n22541__, new_new_n22542__, new_new_n22545__, new_new_n22546__,
    new_new_n22547__, new_new_n22548__, new_new_n22549__, new_new_n22550__,
    new_new_n22551__, new_new_n22552__, new_new_n22553__, new_new_n22556__,
    new_new_n22557__, new_new_n22559__, new_new_n22560__, new_new_n22561__,
    new_new_n22562__, new_new_n22563__, new_new_n22564__, new_new_n22565__,
    new_new_n22566__, new_new_n22567__, new_new_n22568__, new_new_n22569__,
    new_new_n22571__, new_new_n22572__, new_new_n22573__, new_new_n22574__,
    new_new_n22575__, new_new_n22576__, new_new_n22577__, new_new_n22578__,
    new_new_n22579__, new_new_n22580__, new_new_n22581__, new_new_n22582__,
    new_new_n22583__, new_new_n22584__, new_new_n22585__, new_new_n22586__,
    new_new_n22587__, new_new_n22588__, new_new_n22589__, new_new_n22590__,
    new_new_n22591__, new_new_n22592__, new_new_n22593__, new_new_n22594__,
    new_new_n22595__, new_new_n22596__, new_new_n22597__, new_new_n22598__,
    new_new_n22599__, new_new_n22600__, new_new_n22601__, new_new_n22602__,
    new_new_n22603__, new_new_n22604__, new_new_n22605__, new_new_n22606__,
    new_new_n22607__, new_new_n22608__, new_new_n22609__, new_new_n22610__,
    new_new_n22611__, new_new_n22612__, new_new_n22613__, new_new_n22614__,
    new_new_n22615__, new_new_n22616__, new_new_n22617__, new_new_n22618__,
    new_new_n22619__, new_new_n22620__, new_new_n22621__, new_new_n22622__,
    new_new_n22623__, new_new_n22624__, new_new_n22625__, new_new_n22626__,
    new_new_n22627__, new_new_n22628__, new_new_n22629__, new_new_n22630__,
    new_new_n22631__, new_new_n22633__, new_new_n22634__, new_new_n22635__,
    new_new_n22636__, new_new_n22637__, new_new_n22638__, new_new_n22639__,
    new_new_n22640__, new_new_n22641__, new_new_n22642__, new_new_n22643__,
    new_new_n22644__, new_new_n22645__, new_new_n22646__, new_new_n22648__,
    new_new_n22649__, new_new_n22650__, new_new_n22651__, new_new_n22652__,
    new_new_n22653__, new_new_n22654__, new_new_n22655__, new_new_n22656__,
    new_new_n22657__, new_new_n22658__, new_new_n22659__, new_new_n22660__,
    new_new_n22661__, new_new_n22663__, new_new_n22664__, new_new_n22665__,
    new_new_n22666__, new_new_n22667__, new_new_n22668__, new_new_n22669__,
    new_new_n22670__, new_new_n22671__, new_new_n22672__, new_new_n22673__,
    new_new_n22674__, new_new_n22675__, new_new_n22676__, new_new_n22678__,
    new_new_n22679__, new_new_n22680__, new_new_n22681__, new_new_n22682__,
    new_new_n22683__, new_new_n22684__, new_new_n22685__, new_new_n22686__,
    new_new_n22687__, new_new_n22688__, new_new_n22689__, new_new_n22690__,
    new_new_n22691__, new_new_n22693__, new_new_n22694__, new_new_n22695__,
    new_new_n22696__, new_new_n22697__, new_new_n22698__, new_new_n22699__,
    new_new_n22700__, new_new_n22701__, new_new_n22702__, new_new_n22703__,
    new_new_n22704__, new_new_n22705__, new_new_n22706__, new_new_n22708__,
    new_new_n22709__, new_new_n22710__, new_new_n22711__, new_new_n22712__,
    new_new_n22713__, new_new_n22714__, new_new_n22715__, new_new_n22716__,
    new_new_n22717__, new_new_n22718__, new_new_n22719__, new_new_n22720__,
    new_new_n22721__, new_new_n22723__, new_new_n22724__, new_new_n22725__,
    new_new_n22726__, new_new_n22727__, new_new_n22728__, new_new_n22729__,
    new_new_n22730__, new_new_n22731__, new_new_n22732__, new_new_n22733__,
    new_new_n22734__, new_new_n22735__, new_new_n22736__, new_new_n22738__,
    new_new_n22739__, new_new_n22740__, new_new_n22741__, new_new_n22742__,
    new_new_n22743__, new_new_n22745__, new_new_n22746__, new_new_n22748__,
    new_new_n22749__, new_new_n22751__, new_new_n22752__, new_new_n22754__,
    new_new_n22755__, new_new_n22757__, new_new_n22758__, new_new_n22760__,
    new_new_n22761__, new_new_n22763__, new_new_n22764__, new_new_n22766__,
    new_new_n22767__, new_new_n22768__, new_new_n22769__, new_new_n22770__,
    new_new_n22771__, new_new_n22772__, new_new_n22773__, new_new_n22774__,
    new_new_n22775__, new_new_n22776__, new_new_n22777__, new_new_n22778__,
    new_new_n22779__, new_new_n22781__, new_new_n22782__, new_new_n22783__,
    new_new_n22784__, new_new_n22785__, new_new_n22786__, new_new_n22787__,
    new_new_n22788__, new_new_n22789__, new_new_n22790__, new_new_n22791__,
    new_new_n22792__, new_new_n22793__, new_new_n22794__, new_new_n22796__,
    new_new_n22797__, new_new_n22798__, new_new_n22799__, new_new_n22800__,
    new_new_n22801__, new_new_n22802__, new_new_n22803__, new_new_n22804__,
    new_new_n22805__, new_new_n22806__, new_new_n22807__, new_new_n22808__,
    new_new_n22809__, new_new_n22811__, new_new_n22812__, new_new_n22813__,
    new_new_n22814__, new_new_n22815__, new_new_n22816__, new_new_n22817__,
    new_new_n22818__, new_new_n22819__, new_new_n22820__, new_new_n22821__,
    new_new_n22822__, new_new_n22823__, new_new_n22824__, new_new_n22826__,
    new_new_n22827__, new_new_n22828__, new_new_n22829__, new_new_n22830__,
    new_new_n22831__, new_new_n22832__, new_new_n22833__, new_new_n22834__,
    new_new_n22835__, new_new_n22836__, new_new_n22837__, new_new_n22838__,
    new_new_n22839__, new_new_n22841__, new_new_n22842__, new_new_n22843__,
    new_new_n22844__, new_new_n22845__, new_new_n22846__, new_new_n22847__,
    new_new_n22848__, new_new_n22849__, new_new_n22850__, new_new_n22851__,
    new_new_n22852__, new_new_n22853__, new_new_n22854__, new_new_n22856__,
    new_new_n22857__, new_new_n22858__, new_new_n22859__, new_new_n22860__,
    new_new_n22861__, new_new_n22862__, new_new_n22863__, new_new_n22864__,
    new_new_n22865__, new_new_n22866__, new_new_n22867__, new_new_n22868__,
    new_new_n22869__, new_new_n22871__, new_new_n22872__, new_new_n22873__,
    new_new_n22874__, new_new_n22875__, new_new_n22876__, new_new_n22877__,
    new_new_n22878__, new_new_n22879__, new_new_n22880__, new_new_n22881__,
    new_new_n22882__, new_new_n22883__, new_new_n22884__, new_new_n22886__,
    new_new_n22887__, new_new_n22888__, new_new_n22889__, new_new_n22890__,
    new_new_n22891__, new_new_n22893__, new_new_n22894__, new_new_n22896__,
    new_new_n22897__, new_new_n22899__, new_new_n22900__, new_new_n22902__,
    new_new_n22903__, new_new_n22905__, new_new_n22906__, new_new_n22908__,
    new_new_n22909__, new_new_n22911__, new_new_n22912__, new_new_n22914__,
    new_new_n22915__, new_new_n22916__, new_new_n22917__, new_new_n22918__,
    new_new_n22919__, new_new_n22920__, new_new_n22921__, new_new_n22922__,
    new_new_n22923__, new_new_n22924__, new_new_n22925__, new_new_n22926__,
    new_new_n22927__, new_new_n22928__, new_new_n22929__, new_new_n22930__,
    new_new_n22931__, new_new_n22932__, new_new_n22933__, new_new_n22934__,
    new_new_n22935__, new_new_n22936__, new_new_n22937__, new_new_n22938__,
    new_new_n22939__, new_new_n22941__, new_new_n22942__, new_new_n22943__,
    new_new_n22944__, new_new_n22945__, new_new_n22946__, new_new_n22947__,
    new_new_n22948__, new_new_n22949__, new_new_n22950__, new_new_n22951__,
    new_new_n22952__, new_new_n22953__, new_new_n22954__, new_new_n22955__,
    new_new_n22956__, new_new_n22957__, new_new_n22959__, new_new_n22960__,
    new_new_n22961__, new_new_n22962__, new_new_n22963__, new_new_n22964__,
    new_new_n22965__, new_new_n22966__, new_new_n22967__, new_new_n22968__,
    new_new_n22969__, new_new_n22970__, new_new_n22971__, new_new_n22972__,
    new_new_n22973__, new_new_n22974__, new_new_n22975__, new_new_n22977__,
    new_new_n22978__, new_new_n22979__, new_new_n22980__, new_new_n22981__,
    new_new_n22982__, new_new_n22983__, new_new_n22984__, new_new_n22985__,
    new_new_n22986__, new_new_n22987__, new_new_n22988__, new_new_n22989__,
    new_new_n22990__, new_new_n22991__, new_new_n22992__, new_new_n22993__,
    new_new_n22995__, new_new_n22996__, new_new_n22997__, new_new_n22998__,
    new_new_n22999__, new_new_n23000__, new_new_n23001__, new_new_n23002__,
    new_new_n23003__, new_new_n23004__, new_new_n23005__, new_new_n23006__,
    new_new_n23007__, new_new_n23008__, new_new_n23009__, new_new_n23010__,
    new_new_n23011__, new_new_n23013__, new_new_n23014__, new_new_n23015__,
    new_new_n23016__, new_new_n23017__, new_new_n23018__, new_new_n23019__,
    new_new_n23020__, new_new_n23021__, new_new_n23022__, new_new_n23023__,
    new_new_n23024__, new_new_n23025__, new_new_n23026__, new_new_n23027__,
    new_new_n23028__, new_new_n23029__, new_new_n23031__, new_new_n23032__,
    new_new_n23033__, new_new_n23034__, new_new_n23035__, new_new_n23036__,
    new_new_n23037__, new_new_n23038__, new_new_n23039__, new_new_n23040__,
    new_new_n23041__, new_new_n23042__, new_new_n23043__, new_new_n23044__,
    new_new_n23045__, new_new_n23046__, new_new_n23047__, new_new_n23049__,
    new_new_n23050__, new_new_n23051__, new_new_n23052__, new_new_n23053__,
    new_new_n23054__, new_new_n23055__, new_new_n23056__, new_new_n23057__,
    new_new_n23058__, new_new_n23059__, new_new_n23060__, new_new_n23061__,
    new_new_n23062__, new_new_n23063__, new_new_n23064__, new_new_n23065__,
    new_new_n23067__, new_new_n23068__, new_new_n23069__, new_new_n23070__,
    new_new_n23071__, new_new_n23072__, new_new_n23074__, new_new_n23075__,
    new_new_n23077__, new_new_n23078__, new_new_n23080__, new_new_n23081__,
    new_new_n23083__, new_new_n23084__, new_new_n23086__, new_new_n23087__,
    new_new_n23089__, new_new_n23090__, new_new_n23092__, new_new_n23093__,
    new_new_n23095__, new_new_n23096__, new_new_n23097__, new_new_n23098__,
    new_new_n23099__, new_new_n23100__, new_new_n23101__, new_new_n23102__,
    new_new_n23103__, new_new_n23104__, new_new_n23105__, new_new_n23106__,
    new_new_n23107__, new_new_n23108__, new_new_n23109__, new_new_n23110__,
    new_new_n23111__, new_new_n23112__, new_new_n23113__, new_new_n23114__,
    new_new_n23115__, new_new_n23116__, new_new_n23117__, new_new_n23118__,
    new_new_n23119__, new_new_n23120__, new_new_n23121__, new_new_n23122__,
    new_new_n23123__, new_new_n23124__, new_new_n23125__, new_new_n23127__,
    new_new_n23128__, new_new_n23129__, new_new_n23130__, new_new_n23131__,
    new_new_n23132__, new_new_n23133__, new_new_n23134__, new_new_n23135__,
    new_new_n23136__, new_new_n23137__, new_new_n23138__, new_new_n23139__,
    new_new_n23140__, new_new_n23141__, new_new_n23142__, new_new_n23143__,
    new_new_n23144__, new_new_n23146__, new_new_n23147__, new_new_n23148__,
    new_new_n23149__, new_new_n23150__, new_new_n23151__, new_new_n23152__,
    new_new_n23153__, new_new_n23154__, new_new_n23155__, new_new_n23156__,
    new_new_n23157__, new_new_n23158__, new_new_n23159__, new_new_n23160__,
    new_new_n23161__, new_new_n23162__, new_new_n23163__, new_new_n23165__,
    new_new_n23166__, new_new_n23167__, new_new_n23168__, new_new_n23169__,
    new_new_n23170__, new_new_n23171__, new_new_n23172__, new_new_n23173__,
    new_new_n23174__, new_new_n23175__, new_new_n23176__, new_new_n23177__,
    new_new_n23178__, new_new_n23179__, new_new_n23180__, new_new_n23181__,
    new_new_n23182__, new_new_n23184__, new_new_n23185__, new_new_n23186__,
    new_new_n23187__, new_new_n23188__, new_new_n23189__, new_new_n23190__,
    new_new_n23191__, new_new_n23192__, new_new_n23193__, new_new_n23194__,
    new_new_n23195__, new_new_n23196__, new_new_n23197__, new_new_n23198__,
    new_new_n23199__, new_new_n23200__, new_new_n23201__, new_new_n23203__,
    new_new_n23204__, new_new_n23205__, new_new_n23206__, new_new_n23207__,
    new_new_n23208__, new_new_n23209__, new_new_n23210__, new_new_n23211__,
    new_new_n23212__, new_new_n23213__, new_new_n23214__, new_new_n23215__,
    new_new_n23216__, new_new_n23217__, new_new_n23218__, new_new_n23219__,
    new_new_n23220__, new_new_n23222__, new_new_n23223__, new_new_n23224__,
    new_new_n23225__, new_new_n23226__, new_new_n23227__, new_new_n23228__,
    new_new_n23229__, new_new_n23230__, new_new_n23231__, new_new_n23232__,
    new_new_n23233__, new_new_n23234__, new_new_n23235__, new_new_n23236__,
    new_new_n23237__, new_new_n23238__, new_new_n23239__, new_new_n23241__,
    new_new_n23242__, new_new_n23243__, new_new_n23244__, new_new_n23245__,
    new_new_n23246__, new_new_n23247__, new_new_n23248__, new_new_n23249__,
    new_new_n23250__, new_new_n23251__, new_new_n23252__, new_new_n23253__,
    new_new_n23254__, new_new_n23255__, new_new_n23256__, new_new_n23257__,
    new_new_n23258__, new_new_n23260__, new_new_n23261__, new_new_n23262__,
    new_new_n23263__, new_new_n23264__, new_new_n23265__, new_new_n23266__,
    new_new_n23267__, new_new_n23269__, new_new_n23270__, new_new_n23271__,
    new_new_n23273__, new_new_n23274__, new_new_n23276__, new_new_n23277__,
    new_new_n23279__, new_new_n23280__, new_new_n23282__, new_new_n23283__,
    new_new_n23285__, new_new_n23286__, new_new_n23288__, new_new_n23289__,
    new_new_n23291__, new_new_n23292__, new_new_n23293__, new_new_n23294__,
    new_new_n23295__, new_new_n23296__, new_new_n23297__, new_new_n23298__,
    new_new_n23299__, new_new_n23300__, new_new_n23301__, new_new_n23302__,
    new_new_n23303__, new_new_n23304__, new_new_n23306__, new_new_n23307__,
    new_new_n23308__, new_new_n23309__, new_new_n23310__, new_new_n23311__,
    new_new_n23313__, new_new_n23314__, new_new_n23316__, new_new_n23318__,
    new_new_n23319__, new_new_n23320__, new_new_n23321__, new_new_n23322__,
    new_new_n23324__, new_new_n23325__, new_new_n23326__, new_new_n23328__,
    new_new_n23329__, new_new_n23330__, new_new_n23331__, new_new_n23332__,
    new_new_n23333__, new_new_n23334__, new_new_n23335__, new_new_n23336__,
    new_new_n23337__, new_new_n23338__, new_new_n23339__, new_new_n23340__,
    new_new_n23341__, new_new_n23342__, new_new_n23344__, new_new_n23345__,
    new_new_n23346__, new_new_n23347__, new_new_n23348__, new_new_n23349__,
    new_new_n23350__, new_new_n23351__, new_new_n23352__, new_new_n23353__,
    new_new_n23354__, new_new_n23355__, new_new_n23356__, new_new_n23358__,
    new_new_n23359__, new_new_n23360__, new_new_n23361__, new_new_n23362__,
    new_new_n23363__, new_new_n23364__, new_new_n23365__, new_new_n23366__,
    new_new_n23367__, new_new_n23368__, new_new_n23369__, new_new_n23371__,
    new_new_n23372__, new_new_n23373__, new_new_n23374__, new_new_n23375__,
    new_new_n23376__, new_new_n23378__, new_new_n23379__, new_new_n23380__,
    new_new_n23381__, new_new_n23383__, new_new_n23384__, new_new_n23386__,
    new_new_n23387__, new_new_n23388__, new_new_n23389__, new_new_n23390__,
    new_new_n23393__, new_new_n23394__, new_new_n23395__, new_new_n23396__,
    new_new_n23397__, new_new_n23398__, new_new_n23399__, new_new_n23400__,
    new_new_n23401__, new_new_n23402__, new_new_n23403__, new_new_n23404__,
    new_new_n23405__, new_new_n23407__, new_new_n23408__, new_new_n23409__,
    new_new_n23411__, new_new_n23412__, new_new_n23413__, new_new_n23415__,
    new_new_n23416__, new_new_n23417__, new_new_n23418__, new_new_n23419__,
    new_new_n23420__, new_new_n23421__, new_new_n23422__, new_new_n23423__,
    new_new_n23424__, new_new_n23425__, new_new_n23426__, new_new_n23427__,
    new_new_n23428__, new_new_n23429__, new_new_n23430__, new_new_n23431__,
    new_new_n23432__, new_new_n23433__, new_new_n23434__, new_new_n23435__,
    new_new_n23436__, new_new_n23437__, new_new_n23438__, new_new_n23439__,
    new_new_n23440__, new_new_n23441__, new_new_n23442__, new_new_n23443__,
    new_new_n23444__, new_new_n23445__, new_new_n23446__, new_new_n23447__,
    new_new_n23448__, new_new_n23449__, new_new_n23451__, new_new_n23452__,
    new_new_n23453__, new_new_n23454__, new_new_n23455__, new_new_n23456__,
    new_new_n23457__, new_new_n23458__, new_new_n23459__, new_new_n23461__,
    new_new_n23463__, new_new_n23465__, new_new_n23466__, new_new_n23467__,
    new_new_n23469__, new_new_n23470__, new_new_n23471__, new_new_n23472__,
    new_new_n23476__, new_new_n23477__, new_new_n23478__, new_new_n23479__,
    new_new_n23480__, new_new_n23481__, new_new_n23482__, new_new_n23483__,
    new_new_n23484__, new_new_n23485__, new_new_n23486__, new_new_n23487__,
    new_new_n23488__, new_new_n23489__, new_new_n23490__, new_new_n23491__,
    new_new_n23492__, new_new_n23493__, new_new_n23494__, new_new_n23495__,
    new_new_n23496__, new_new_n23497__, new_new_n23498__, new_new_n23499__,
    new_new_n23500__, new_new_n23501__, new_new_n23502__, new_new_n23503__,
    new_new_n23504__, new_new_n23505__, new_new_n23506__, new_new_n23507__,
    new_new_n23508__, new_new_n23509__, new_new_n23510__, new_new_n23511__,
    new_new_n23512__, new_new_n23513__, new_new_n23514__, new_new_n23515__,
    new_new_n23516__, new_new_n23517__, new_new_n23518__, new_new_n23519__,
    new_new_n23520__, new_new_n23521__, new_new_n23522__, new_new_n23523__,
    new_new_n23524__, new_new_n23525__, new_new_n23526__, new_new_n23527__,
    new_new_n23528__, new_new_n23529__, new_new_n23530__, new_new_n23531__,
    new_new_n23532__, new_new_n23533__, new_new_n23534__, new_new_n23535__,
    new_new_n23536__, new_new_n23537__, new_new_n23538__, new_new_n23539__,
    new_new_n23540__, new_new_n23541__, new_new_n23542__, new_new_n23543__,
    new_new_n23544__, new_new_n23545__, new_new_n23546__, new_new_n23547__,
    new_new_n23548__, new_new_n23549__, new_new_n23550__, new_new_n23551__,
    new_new_n23552__, new_new_n23553__, new_new_n23554__, new_new_n23555__,
    new_new_n23556__, new_new_n23557__, new_new_n23558__, new_new_n23559__,
    new_new_n23560__, new_new_n23561__, new_new_n23562__, new_new_n23563__,
    new_new_n23564__, new_new_n23565__, new_new_n23566__, new_new_n23567__,
    new_new_n23568__, new_new_n23569__, new_new_n23570__, new_new_n23571__,
    new_new_n23572__, new_new_n23573__, new_new_n23574__, new_new_n23575__,
    new_new_n23576__, new_new_n23577__, new_new_n23578__, new_new_n23579__,
    new_new_n23580__, new_new_n23581__, new_new_n23582__, new_new_n23583__,
    new_new_n23584__, new_new_n23585__, new_new_n23586__, new_new_n23587__,
    new_new_n23588__, new_new_n23589__, new_new_n23590__, new_new_n23591__,
    new_new_n23592__, new_new_n23593__, new_new_n23594__, new_new_n23595__,
    new_new_n23596__, new_new_n23597__, new_new_n23598__, new_new_n23599__,
    new_new_n23600__, new_new_n23601__, new_new_n23602__, new_new_n23603__,
    new_new_n23604__, new_new_n23605__, new_new_n23606__, new_new_n23607__,
    new_new_n23608__, new_new_n23609__, new_new_n23610__, new_new_n23611__,
    new_new_n23612__, new_new_n23613__, new_new_n23614__, new_new_n23615__,
    new_new_n23616__, new_new_n23617__, new_new_n23618__, new_new_n23619__,
    new_new_n23620__, new_new_n23621__, new_new_n23622__, new_new_n23623__,
    new_new_n23624__, new_new_n23625__, new_new_n23626__, new_new_n23627__,
    new_new_n23628__, new_new_n23629__, new_new_n23630__, new_new_n23631__,
    new_new_n23632__, new_new_n23633__, new_new_n23634__, new_new_n23635__,
    new_new_n23636__, new_new_n23637__, new_new_n23638__, new_new_n23639__,
    new_new_n23640__, new_new_n23641__, new_new_n23642__, new_new_n23643__,
    new_new_n23644__, new_new_n23645__, new_new_n23646__, new_new_n23647__,
    new_new_n23648__, new_new_n23649__, new_new_n23650__, new_new_n23651__,
    new_new_n23652__, new_new_n23653__, new_new_n23654__, new_new_n23655__,
    new_new_n23656__, new_new_n23657__, new_new_n23658__, new_new_n23659__,
    new_new_n23660__, new_new_n23661__, new_new_n23662__, new_new_n23663__,
    new_new_n23664__, new_new_n23665__, new_new_n23666__, new_new_n23667__,
    new_new_n23668__, new_new_n23669__, new_new_n23670__, new_new_n23671__,
    new_new_n23672__, new_new_n23673__, new_new_n23674__, new_new_n23675__,
    new_new_n23676__, new_new_n23677__, new_new_n23678__, new_new_n23679__,
    new_new_n23680__, new_new_n23681__, new_new_n23682__, new_new_n23683__,
    new_new_n23684__, new_new_n23685__, new_new_n23686__, new_new_n23687__,
    new_new_n23688__, new_new_n23689__, new_new_n23690__, new_new_n23691__,
    new_new_n23692__, new_new_n23693__, new_new_n23694__, new_new_n23695__,
    new_new_n23696__, new_new_n23697__, new_new_n23698__, new_new_n23699__,
    new_new_n23700__, new_new_n23701__, new_new_n23702__, new_new_n23703__,
    new_new_n23704__, new_new_n23705__, new_new_n23706__, new_new_n23707__,
    new_new_n23708__, new_new_n23709__, new_new_n23710__, new_new_n23711__,
    new_new_n23712__, new_new_n23713__, new_new_n23714__, new_new_n23715__,
    new_new_n23716__, new_new_n23717__, new_new_n23718__, new_new_n23719__,
    new_new_n23720__, new_new_n23721__, new_new_n23722__, new_new_n23723__,
    new_new_n23724__, new_new_n23725__, new_new_n23726__, new_new_n23727__,
    new_new_n23728__, new_new_n23729__, new_new_n23730__, new_new_n23731__,
    new_new_n23732__, new_new_n23733__, new_new_n23734__, new_new_n23735__,
    new_new_n23736__, new_new_n23737__, new_new_n23738__, new_new_n23739__,
    new_new_n23740__, new_new_n23741__, new_new_n23742__, new_new_n23743__,
    new_new_n23744__, new_new_n23745__, new_new_n23746__, new_new_n23747__,
    new_new_n23748__, new_new_n23749__, new_new_n23750__, new_new_n23751__,
    new_new_n23752__, new_new_n23753__, new_new_n23754__, new_new_n23755__,
    new_new_n23756__, new_new_n23757__, new_new_n23758__, new_new_n23759__,
    new_new_n23760__, new_new_n23761__, new_new_n23762__, new_new_n23763__,
    new_new_n23764__, new_new_n23765__, new_new_n23766__, new_new_n23767__,
    new_new_n23768__, new_new_n23769__, new_new_n23770__, new_new_n23771__,
    new_new_n23772__, new_new_n23773__, new_new_n23774__, new_new_n23775__,
    new_new_n23776__, new_new_n23777__, new_new_n23778__, new_new_n23779__,
    new_new_n23780__, new_new_n23781__, new_new_n23782__, new_new_n23783__,
    new_new_n23784__, new_new_n23785__, new_new_n23786__, new_new_n23787__,
    new_new_n23788__, new_new_n23789__, new_new_n23790__, new_new_n23791__,
    new_new_n23792__, new_new_n23793__, new_new_n23794__, new_new_n23795__,
    new_new_n23796__, new_new_n23797__, new_new_n23798__, new_new_n23799__,
    new_new_n23800__, new_new_n23801__, new_new_n23802__, new_new_n23803__,
    new_new_n23804__, new_new_n23805__, new_new_n23806__, new_new_n23807__,
    new_new_n23808__, new_new_n23809__, new_new_n23810__, new_new_n23811__,
    new_new_n23812__, new_new_n23813__, new_new_n23814__, new_new_n23815__,
    new_new_n23816__, new_new_n23817__, new_new_n23818__, new_new_n23819__,
    new_new_n23820__, new_new_n23821__, new_new_n23822__, new_new_n23823__,
    new_new_n23824__, new_new_n23825__, new_new_n23826__, new_new_n23827__,
    new_new_n23828__, new_new_n23829__, new_new_n23830__, new_new_n23831__,
    new_new_n23832__, new_new_n23833__, new_new_n23834__, new_new_n23835__,
    new_new_n23836__, new_new_n23837__, new_new_n23838__, new_new_n23839__,
    new_new_n23840__, new_new_n23841__, new_new_n23842__, new_new_n23843__,
    new_new_n23844__, new_new_n23845__, new_new_n23846__, new_new_n23847__,
    new_new_n23848__, new_new_n23849__, new_new_n23850__, new_new_n23851__,
    new_new_n23852__, new_new_n23853__, new_new_n23854__, new_new_n23855__,
    new_new_n23856__, new_new_n23857__, new_new_n23858__, new_new_n23859__,
    new_new_n23860__, new_new_n23861__, new_new_n23862__, new_new_n23863__,
    new_new_n23864__, new_new_n23865__, new_new_n23866__, new_new_n23867__,
    new_new_n23868__, new_new_n23869__, new_new_n23870__, new_new_n23871__,
    new_new_n23872__, new_new_n23873__, new_new_n23874__, new_new_n23875__,
    new_new_n23876__, new_new_n23877__, new_new_n23878__, new_new_n23879__,
    new_new_n23880__, new_new_n23881__, new_new_n23882__, new_new_n23883__,
    new_new_n23884__, new_new_n23885__, new_new_n23886__, new_new_n23887__,
    new_new_n23888__, new_new_n23889__, new_new_n23890__, new_new_n23891__,
    new_new_n23892__, new_new_n23893__, new_new_n23894__, new_new_n23895__,
    new_new_n23896__, new_new_n23897__, new_new_n23898__, new_new_n23899__,
    new_new_n23900__, new_new_n23901__, new_new_n23902__, new_new_n23903__,
    new_new_n23904__, new_new_n23905__, new_new_n23906__, new_new_n23907__,
    new_new_n23908__, new_new_n23909__, new_new_n23910__, new_new_n23911__,
    new_new_n23912__, new_new_n23913__, new_new_n23914__, new_new_n23915__,
    new_new_n23916__, new_new_n23917__, new_new_n23918__, new_new_n23919__,
    new_new_n23920__, new_new_n23921__, new_new_n23922__, new_new_n23923__,
    new_new_n23924__, new_new_n23925__, new_new_n23926__, new_new_n23927__,
    new_new_n23928__, new_new_n23929__, new_new_n23930__, new_new_n23931__,
    new_new_n23932__, new_new_n23933__, new_new_n23934__, new_new_n23935__,
    new_new_n23936__, new_new_n23937__, new_new_n23938__, new_new_n23939__,
    new_new_n23940__, new_new_n23941__, new_new_n23942__, new_new_n23943__,
    new_new_n23944__, new_new_n23945__, new_new_n23946__, new_new_n23947__,
    new_new_n23948__, new_new_n23949__, new_new_n23950__, new_new_n23951__,
    new_new_n23952__, new_new_n23953__, new_new_n23954__, new_new_n23955__,
    new_new_n23956__, new_new_n23957__, new_new_n23958__, new_new_n23959__,
    new_new_n23960__, new_new_n23961__, new_new_n23962__, new_new_n23963__,
    new_new_n23964__, new_new_n23965__, new_new_n23966__, new_new_n23967__,
    new_new_n23968__, new_new_n23969__, new_new_n23970__, new_new_n23971__,
    new_new_n23972__, new_new_n23973__, new_new_n23974__, new_new_n23975__,
    new_new_n23976__, new_new_n23977__, new_new_n23978__, new_new_n23979__,
    new_new_n23980__, new_new_n23981__, new_new_n23982__, new_new_n23983__,
    new_new_n23984__, new_new_n23985__, new_new_n23986__, new_new_n23987__,
    new_new_n23988__, new_new_n23989__, new_new_n23990__, new_new_n23991__,
    new_new_n23992__, new_new_n23993__, new_new_n23994__, new_new_n23995__,
    new_new_n23996__, new_new_n23997__, new_new_n23998__, new_new_n23999__,
    new_new_n24000__, new_new_n24001__, new_new_n24002__, new_new_n24003__,
    new_new_n24004__, new_new_n24005__, new_new_n24006__, new_new_n24007__,
    new_new_n24008__, new_new_n24009__, new_new_n24010__, new_new_n24011__,
    new_new_n24012__, new_new_n24013__, new_new_n24014__, new_new_n24015__,
    new_new_n24016__, new_new_n24017__, new_new_n24018__, new_new_n24019__,
    new_new_n24020__, new_new_n24021__, new_new_n24022__, new_new_n24023__,
    new_new_n24024__, new_new_n24025__, new_new_n24026__, new_new_n24027__,
    new_new_n24028__, new_new_n24029__, new_new_n24030__, new_new_n24031__,
    new_new_n24032__, new_new_n24033__, new_new_n24034__, new_new_n24035__,
    new_new_n24036__, new_new_n24037__, new_new_n24038__, new_new_n24039__,
    new_new_n24040__, new_new_n24041__, new_new_n24042__, new_new_n24043__,
    new_new_n24044__, new_new_n24045__, new_new_n24046__, new_new_n24047__,
    new_new_n24048__, new_new_n24049__, new_new_n24050__, new_new_n24051__,
    new_new_n24052__, new_new_n24053__, new_new_n24054__, new_new_n24055__,
    new_new_n24056__, new_new_n24057__, new_new_n24058__, new_new_n24059__,
    new_new_n24060__, new_new_n24061__, new_new_n24062__, new_new_n24063__,
    new_new_n24064__, new_new_n24065__, new_new_n24066__, new_new_n24067__,
    new_new_n24068__, new_new_n24069__, new_new_n24070__, new_new_n24071__,
    new_new_n24072__, new_new_n24073__, new_new_n24074__, new_new_n24075__,
    new_new_n24076__, new_new_n24077__, new_new_n24078__, new_new_n24079__,
    new_new_n24080__, new_new_n24081__, new_new_n24082__, new_new_n24083__,
    new_new_n24084__, new_new_n24085__, new_new_n24086__, new_new_n24087__,
    new_new_n24088__, new_new_n24089__, new_new_n24090__, new_new_n24091__,
    new_new_n24092__, new_new_n24093__, new_new_n24094__, new_new_n24095__,
    new_new_n24096__, new_new_n24097__, new_new_n24098__, new_new_n24099__,
    new_new_n24100__, new_new_n24101__, new_new_n24102__, new_new_n24103__,
    new_new_n24104__, new_new_n24105__, new_new_n24106__, new_new_n24107__,
    new_new_n24108__, new_new_n24109__, new_new_n24110__, new_new_n24111__,
    new_new_n24112__, new_new_n24113__, new_new_n24114__, new_new_n24115__,
    new_new_n24116__, new_new_n24117__, new_new_n24118__, new_new_n24119__,
    new_new_n24120__, new_new_n24121__, new_new_n24122__, new_new_n24123__,
    new_new_n24124__, new_new_n24125__, new_new_n24126__, new_new_n24127__,
    new_new_n24128__, new_new_n24129__, new_new_n24130__, new_new_n24131__,
    new_new_n24132__, new_new_n24133__, new_new_n24134__, new_new_n24135__,
    new_new_n24136__, new_new_n24137__, new_new_n24138__, new_new_n24139__,
    new_new_n24140__, new_new_n24141__, new_new_n24142__, new_new_n24143__,
    new_new_n24144__, new_new_n24145__, new_new_n24146__, new_new_n24147__,
    new_new_n24148__, new_new_n24149__, new_new_n24150__, new_new_n24151__,
    new_new_n24152__, new_new_n24153__, new_new_n24154__, new_new_n24155__,
    new_new_n24156__, new_new_n24157__, new_new_n24158__, new_new_n24159__,
    new_new_n24160__, new_new_n24161__, new_new_n24162__, new_new_n24163__,
    new_new_n24164__, new_new_n24165__, new_new_n24166__, new_new_n24167__,
    new_new_n24168__, new_new_n24169__, new_new_n24170__, new_new_n24171__,
    new_new_n24172__, new_new_n24173__, new_new_n24174__, new_new_n24175__,
    new_new_n24176__, new_new_n24177__, new_new_n24178__, new_new_n24179__,
    new_new_n24180__, new_new_n24181__, new_new_n24182__, new_new_n24183__,
    new_new_n24184__, new_new_n24185__, new_new_n24186__, new_new_n24187__,
    new_new_n24188__, new_new_n24189__, new_new_n24190__, new_new_n24191__,
    new_new_n24192__, new_new_n24193__, new_new_n24194__, new_new_n24195__,
    new_new_n24196__, new_new_n24197__, new_new_n24198__, new_new_n24199__,
    new_new_n24200__, new_new_n24201__, new_new_n24202__, new_new_n24203__,
    new_new_n24204__, new_new_n24205__, new_new_n24206__, new_new_n24207__,
    new_new_n24208__, new_new_n24209__, new_new_n24210__, new_new_n24211__,
    new_new_n24212__, new_new_n24213__, new_new_n24214__, new_new_n24215__,
    new_new_n24216__, new_new_n24217__, new_new_n24218__, new_new_n24219__,
    new_new_n24220__, new_new_n24221__, new_new_n24222__, new_new_n24223__,
    new_new_n24224__, new_new_n24225__, new_new_n24226__, new_new_n24227__,
    new_new_n24228__, new_new_n24229__, new_new_n24230__, new_new_n24231__,
    new_new_n24232__, new_new_n24233__, new_new_n24234__, new_new_n24235__,
    new_new_n24236__, new_new_n24237__, new_new_n24238__, new_new_n24239__,
    new_new_n24240__, new_new_n24241__, new_new_n24242__, new_new_n24243__,
    new_new_n24244__, new_new_n24245__, new_new_n24246__, new_new_n24247__,
    new_new_n24248__, new_new_n24249__, new_new_n24250__, new_new_n24251__,
    new_new_n24252__, new_new_n24253__, new_new_n24254__, new_new_n24255__,
    new_new_n24256__, new_new_n24257__, new_new_n24258__, new_new_n24259__,
    new_new_n24260__, new_new_n24261__, new_new_n24262__, new_new_n24263__,
    new_new_n24264__, new_new_n24265__, new_new_n24266__, new_new_n24267__,
    new_new_n24268__, new_new_n24269__, new_new_n24270__, new_new_n24271__,
    new_new_n24272__, new_new_n24274__, new_new_n24275__, new_new_n24276__,
    new_new_n24277__, new_new_n24278__, new_new_n24279__, new_new_n24280__,
    new_new_n24281__, new_new_n24282__, new_new_n24283__, new_new_n24284__,
    new_new_n24285__, new_new_n24286__, new_new_n24287__, new_new_n24288__,
    new_new_n24289__, new_new_n24290__, new_new_n24291__, new_new_n24292__,
    new_new_n24293__, new_new_n24294__, new_new_n24295__, new_new_n24296__,
    new_new_n24297__, new_new_n24298__, new_new_n24299__, new_new_n24300__,
    new_new_n24301__, new_new_n24302__, new_new_n24303__, new_new_n24304__,
    new_new_n24305__, new_new_n24306__, new_new_n24307__, new_new_n24308__,
    new_new_n24309__, new_new_n24310__, new_new_n24311__, new_new_n24312__,
    new_new_n24313__, new_new_n24314__, new_new_n24315__, new_new_n24316__,
    new_new_n24317__, new_new_n24318__, new_new_n24319__, new_new_n24320__,
    new_new_n24321__, new_new_n24322__, new_new_n24323__, new_new_n24324__,
    new_new_n24325__, new_new_n24326__, new_new_n24327__, new_new_n24328__,
    new_new_n24329__, new_new_n24330__, new_new_n24331__, new_new_n24332__,
    new_new_n24333__, new_new_n24334__, new_new_n24335__, new_new_n24336__,
    new_new_n24337__, new_new_n24338__, new_new_n24340__, new_new_n24341__,
    new_new_n24342__, new_new_n24343__, new_new_n24344__, new_new_n24345__,
    new_new_n24346__, new_new_n24347__, new_new_n24348__, new_new_n24349__,
    new_new_n24350__, new_new_n24351__, new_new_n24352__, new_new_n24353__,
    new_new_n24354__, new_new_n24355__, new_new_n24356__, new_new_n24357__,
    new_new_n24358__, new_new_n24359__, new_new_n24360__, new_new_n24361__,
    new_new_n24362__, new_new_n24363__, new_new_n24364__, new_new_n24365__,
    new_new_n24366__, new_new_n24367__, new_new_n24368__, new_new_n24369__,
    new_new_n24370__, new_new_n24371__, new_new_n24372__, new_new_n24373__,
    new_new_n24374__, new_new_n24375__, new_new_n24376__, new_new_n24377__,
    new_new_n24378__, new_new_n24379__, new_new_n24380__, new_new_n24381__,
    new_new_n24382__, new_new_n24383__, new_new_n24384__, new_new_n24385__,
    new_new_n24386__, new_new_n24387__, new_new_n24388__, new_new_n24389__,
    new_new_n24390__, new_new_n24391__, new_new_n24392__, new_new_n24393__,
    new_new_n24394__, new_new_n24395__, new_new_n24396__, new_new_n24397__,
    new_new_n24398__, new_new_n24399__, new_new_n24400__, new_new_n24401__,
    new_new_n24402__, new_new_n24403__, new_new_n24404__, new_new_n24405__,
    new_new_n24406__, new_new_n24407__, new_new_n24408__, new_new_n24409__,
    new_new_n24410__, new_new_n24412__, new_new_n24413__, new_new_n24414__,
    new_new_n24415__, new_new_n24416__, new_new_n24417__, new_new_n24418__,
    new_new_n24419__, new_new_n24420__, new_new_n24421__, new_new_n24422__,
    new_new_n24423__, new_new_n24424__, new_new_n24425__, new_new_n24426__,
    new_new_n24427__, new_new_n24428__, new_new_n24429__, new_new_n24430__,
    new_new_n24431__, new_new_n24432__, new_new_n24433__, new_new_n24434__,
    new_new_n24435__, new_new_n24436__, new_new_n24437__, new_new_n24438__,
    new_new_n24439__, new_new_n24440__, new_new_n24441__, new_new_n24442__,
    new_new_n24443__, new_new_n24444__, new_new_n24445__, new_new_n24446__,
    new_new_n24447__, new_new_n24448__, new_new_n24449__, new_new_n24450__,
    new_new_n24451__, new_new_n24452__, new_new_n24453__, new_new_n24454__,
    new_new_n24455__, new_new_n24456__, new_new_n24457__, new_new_n24458__,
    new_new_n24459__, new_new_n24460__, new_new_n24461__, new_new_n24462__,
    new_new_n24463__, new_new_n24464__, new_new_n24465__, new_new_n24466__,
    new_new_n24467__, new_new_n24468__, new_new_n24469__, new_new_n24470__,
    new_new_n24471__, new_new_n24472__, new_new_n24473__, new_new_n24474__,
    new_new_n24475__, new_new_n24476__, new_new_n24477__, new_new_n24478__,
    new_new_n24479__, new_new_n24480__, new_new_n24481__, new_new_n24482__,
    new_new_n24483__, new_new_n24484__, new_new_n24485__, new_new_n24487__,
    new_new_n24488__, new_new_n24489__, new_new_n24490__, new_new_n24491__,
    new_new_n24492__, new_new_n24493__, new_new_n24494__, new_new_n24495__,
    new_new_n24496__, new_new_n24497__, new_new_n24498__, new_new_n24499__,
    new_new_n24500__, new_new_n24501__, new_new_n24502__, new_new_n24503__,
    new_new_n24504__, new_new_n24505__, new_new_n24506__, new_new_n24507__,
    new_new_n24508__, new_new_n24509__, new_new_n24510__, new_new_n24511__,
    new_new_n24512__, new_new_n24513__, new_new_n24514__, new_new_n24515__,
    new_new_n24516__, new_new_n24517__, new_new_n24518__, new_new_n24519__,
    new_new_n24520__, new_new_n24521__, new_new_n24522__, new_new_n24523__,
    new_new_n24524__, new_new_n24525__, new_new_n24526__, new_new_n24527__,
    new_new_n24528__, new_new_n24529__, new_new_n24530__, new_new_n24531__,
    new_new_n24532__, new_new_n24533__, new_new_n24534__, new_new_n24535__,
    new_new_n24536__, new_new_n24537__, new_new_n24538__, new_new_n24539__,
    new_new_n24540__, new_new_n24541__, new_new_n24542__, new_new_n24543__,
    new_new_n24544__, new_new_n24545__, new_new_n24546__, new_new_n24547__,
    new_new_n24548__, new_new_n24549__, new_new_n24550__, new_new_n24551__,
    new_new_n24552__, new_new_n24553__, new_new_n24554__, new_new_n24555__,
    new_new_n24556__, new_new_n24557__, new_new_n24558__, new_new_n24559__,
    new_new_n24560__, new_new_n24561__, new_new_n24562__, new_new_n24564__,
    new_new_n24565__, new_new_n24566__, new_new_n24567__, new_new_n24568__,
    new_new_n24569__, new_new_n24570__, new_new_n24571__, new_new_n24572__,
    new_new_n24573__, new_new_n24574__, new_new_n24575__, new_new_n24576__,
    new_new_n24577__, new_new_n24578__, new_new_n24579__, new_new_n24580__,
    new_new_n24581__, new_new_n24582__, new_new_n24583__, new_new_n24584__,
    new_new_n24585__, new_new_n24586__, new_new_n24587__, new_new_n24588__,
    new_new_n24589__, new_new_n24590__, new_new_n24591__, new_new_n24592__,
    new_new_n24593__, new_new_n24594__, new_new_n24595__, new_new_n24596__,
    new_new_n24597__, new_new_n24598__, new_new_n24599__, new_new_n24600__,
    new_new_n24601__, new_new_n24602__, new_new_n24603__, new_new_n24604__,
    new_new_n24605__, new_new_n24606__, new_new_n24607__, new_new_n24608__,
    new_new_n24609__, new_new_n24610__, new_new_n24611__, new_new_n24612__,
    new_new_n24613__, new_new_n24614__, new_new_n24615__, new_new_n24616__,
    new_new_n24617__, new_new_n24618__, new_new_n24619__, new_new_n24620__,
    new_new_n24621__, new_new_n24622__, new_new_n24623__, new_new_n24624__,
    new_new_n24625__, new_new_n24626__, new_new_n24627__, new_new_n24628__,
    new_new_n24629__, new_new_n24630__, new_new_n24631__, new_new_n24632__,
    new_new_n24633__, new_new_n24634__, new_new_n24635__, new_new_n24636__,
    new_new_n24637__, new_new_n24638__, new_new_n24640__, new_new_n24641__,
    new_new_n24642__, new_new_n24643__, new_new_n24644__, new_new_n24645__,
    new_new_n24646__, new_new_n24647__, new_new_n24648__, new_new_n24649__,
    new_new_n24650__, new_new_n24651__, new_new_n24652__, new_new_n24653__,
    new_new_n24654__, new_new_n24655__, new_new_n24656__, new_new_n24657__,
    new_new_n24658__, new_new_n24659__, new_new_n24660__, new_new_n24661__,
    new_new_n24662__, new_new_n24663__, new_new_n24664__, new_new_n24665__,
    new_new_n24666__, new_new_n24667__, new_new_n24668__, new_new_n24669__,
    new_new_n24670__, new_new_n24671__, new_new_n24672__, new_new_n24673__,
    new_new_n24674__, new_new_n24675__, new_new_n24676__, new_new_n24677__,
    new_new_n24678__, new_new_n24679__, new_new_n24680__, new_new_n24681__,
    new_new_n24682__, new_new_n24683__, new_new_n24684__, new_new_n24685__,
    new_new_n24686__, new_new_n24687__, new_new_n24688__, new_new_n24689__,
    new_new_n24690__, new_new_n24691__, new_new_n24692__, new_new_n24693__,
    new_new_n24694__, new_new_n24695__, new_new_n24696__, new_new_n24697__,
    new_new_n24698__, new_new_n24699__, new_new_n24700__, new_new_n24701__,
    new_new_n24702__, new_new_n24703__, new_new_n24704__, new_new_n24705__,
    new_new_n24706__, new_new_n24707__, new_new_n24708__, new_new_n24709__,
    new_new_n24710__, new_new_n24711__, new_new_n24712__, new_new_n24713__,
    new_new_n24714__, new_new_n24715__, new_new_n24716__, new_new_n24717__,
    new_new_n24718__, new_new_n24720__, new_new_n24721__, new_new_n24722__,
    new_new_n24723__, new_new_n24724__, new_new_n24725__, new_new_n24726__,
    new_new_n24727__, new_new_n24728__, new_new_n24729__, new_new_n24730__,
    new_new_n24731__, new_new_n24732__, new_new_n24733__, new_new_n24734__,
    new_new_n24735__, new_new_n24736__, new_new_n24737__, new_new_n24738__,
    new_new_n24739__, new_new_n24740__, new_new_n24741__, new_new_n24742__,
    new_new_n24743__, new_new_n24744__, new_new_n24745__, new_new_n24746__,
    new_new_n24747__, new_new_n24748__, new_new_n24749__, new_new_n24750__,
    new_new_n24751__, new_new_n24752__, new_new_n24753__, new_new_n24754__,
    new_new_n24755__, new_new_n24756__, new_new_n24757__, new_new_n24758__,
    new_new_n24759__, new_new_n24760__, new_new_n24761__, new_new_n24762__,
    new_new_n24763__, new_new_n24764__, new_new_n24765__, new_new_n24766__,
    new_new_n24767__, new_new_n24768__, new_new_n24769__, new_new_n24770__,
    new_new_n24771__, new_new_n24772__, new_new_n24773__, new_new_n24774__,
    new_new_n24775__, new_new_n24776__, new_new_n24777__, new_new_n24778__,
    new_new_n24779__, new_new_n24780__, new_new_n24781__, new_new_n24782__,
    new_new_n24783__, new_new_n24784__, new_new_n24785__, new_new_n24786__,
    new_new_n24787__, new_new_n24788__, new_new_n24789__, new_new_n24790__,
    new_new_n24791__, new_new_n24792__, new_new_n24793__, new_new_n24794__,
    new_new_n24796__, new_new_n24797__, new_new_n24798__, new_new_n24799__,
    new_new_n24800__, new_new_n24801__, new_new_n24802__, new_new_n24803__,
    new_new_n24804__, new_new_n24805__, new_new_n24806__, new_new_n24807__,
    new_new_n24808__, new_new_n24809__, new_new_n24810__, new_new_n24811__,
    new_new_n24812__, new_new_n24813__, new_new_n24814__, new_new_n24815__,
    new_new_n24816__, new_new_n24817__, new_new_n24818__, new_new_n24819__,
    new_new_n24820__, new_new_n24821__, new_new_n24822__, new_new_n24823__,
    new_new_n24824__, new_new_n24825__, new_new_n24826__, new_new_n24827__,
    new_new_n24828__, new_new_n24829__, new_new_n24830__, new_new_n24831__,
    new_new_n24832__, new_new_n24833__, new_new_n24834__, new_new_n24835__,
    new_new_n24836__, new_new_n24837__, new_new_n24838__, new_new_n24839__,
    new_new_n24840__, new_new_n24841__, new_new_n24842__, new_new_n24843__,
    new_new_n24844__, new_new_n24845__, new_new_n24846__, new_new_n24847__,
    new_new_n24848__, new_new_n24849__, new_new_n24850__, new_new_n24851__,
    new_new_n24852__, new_new_n24853__, new_new_n24854__, new_new_n24855__,
    new_new_n24856__, new_new_n24857__, new_new_n24858__, new_new_n24859__,
    new_new_n24860__, new_new_n24861__, new_new_n24862__, new_new_n24863__,
    new_new_n24864__, new_new_n24865__, new_new_n24866__, new_new_n24867__,
    new_new_n24868__, new_new_n24869__, new_new_n24870__, new_new_n24871__,
    new_new_n24872__, new_new_n24873__, new_new_n24874__, new_new_n24875__,
    new_new_n24877__, new_new_n24878__, new_new_n24879__, new_new_n24880__,
    new_new_n24881__, new_new_n24882__, new_new_n24883__, new_new_n24884__,
    new_new_n24885__, new_new_n24886__, new_new_n24887__, new_new_n24888__,
    new_new_n24889__, new_new_n24890__, new_new_n24891__, new_new_n24892__,
    new_new_n24893__, new_new_n24894__, new_new_n24895__, new_new_n24896__,
    new_new_n24897__, new_new_n24898__, new_new_n24899__, new_new_n24900__,
    new_new_n24901__, new_new_n24902__, new_new_n24903__, new_new_n24904__,
    new_new_n24905__, new_new_n24906__, new_new_n24907__, new_new_n24908__,
    new_new_n24909__, new_new_n24910__, new_new_n24911__, new_new_n24912__,
    new_new_n24913__, new_new_n24914__, new_new_n24915__, new_new_n24916__,
    new_new_n24917__, new_new_n24918__, new_new_n24919__, new_new_n24920__,
    new_new_n24921__, new_new_n24922__, new_new_n24923__, new_new_n24924__,
    new_new_n24925__, new_new_n24926__, new_new_n24927__, new_new_n24928__,
    new_new_n24929__, new_new_n24930__, new_new_n24931__, new_new_n24932__,
    new_new_n24933__, new_new_n24934__, new_new_n24935__, new_new_n24936__,
    new_new_n24937__, new_new_n24938__, new_new_n24939__, new_new_n24940__,
    new_new_n24941__, new_new_n24942__, new_new_n24943__, new_new_n24944__,
    new_new_n24945__, new_new_n24946__, new_new_n24947__, new_new_n24948__,
    new_new_n24949__, new_new_n24950__, new_new_n24951__, new_new_n24953__,
    new_new_n24954__, new_new_n24955__, new_new_n24956__, new_new_n24957__,
    new_new_n24958__, new_new_n24959__, new_new_n24960__, new_new_n24961__,
    new_new_n24962__, new_new_n24963__, new_new_n24964__, new_new_n24965__,
    new_new_n24966__, new_new_n24967__, new_new_n24968__, new_new_n24969__,
    new_new_n24970__, new_new_n24971__, new_new_n24972__, new_new_n24973__,
    new_new_n24974__, new_new_n24975__, new_new_n24976__, new_new_n24977__,
    new_new_n24978__, new_new_n24979__, new_new_n24980__, new_new_n24981__,
    new_new_n24982__, new_new_n24983__, new_new_n24984__, new_new_n24985__,
    new_new_n24986__, new_new_n24987__, new_new_n24988__, new_new_n24989__,
    new_new_n24990__, new_new_n24991__, new_new_n24992__, new_new_n24993__,
    new_new_n24994__, new_new_n24995__, new_new_n24996__, new_new_n24997__,
    new_new_n24998__, new_new_n24999__, new_new_n25000__, new_new_n25001__,
    new_new_n25002__, new_new_n25003__, new_new_n25004__, new_new_n25005__,
    new_new_n25006__, new_new_n25007__, new_new_n25008__, new_new_n25009__,
    new_new_n25010__, new_new_n25011__, new_new_n25012__, new_new_n25013__,
    new_new_n25014__, new_new_n25015__, new_new_n25016__, new_new_n25017__,
    new_new_n25018__, new_new_n25019__, new_new_n25020__, new_new_n25021__,
    new_new_n25022__, new_new_n25023__, new_new_n25024__, new_new_n25025__,
    new_new_n25026__, new_new_n25027__, new_new_n25028__, new_new_n25029__,
    new_new_n25030__, new_new_n25031__, new_new_n25033__, new_new_n25034__,
    new_new_n25035__, new_new_n25036__, new_new_n25037__, new_new_n25038__,
    new_new_n25039__, new_new_n25040__, new_new_n25041__, new_new_n25042__,
    new_new_n25043__, new_new_n25044__, new_new_n25045__, new_new_n25046__,
    new_new_n25047__, new_new_n25048__, new_new_n25049__, new_new_n25050__,
    new_new_n25051__, new_new_n25052__, new_new_n25053__, new_new_n25054__,
    new_new_n25055__, new_new_n25056__, new_new_n25057__, new_new_n25058__,
    new_new_n25059__, new_new_n25060__, new_new_n25061__, new_new_n25062__,
    new_new_n25063__, new_new_n25064__, new_new_n25065__, new_new_n25066__,
    new_new_n25067__, new_new_n25068__, new_new_n25069__, new_new_n25070__,
    new_new_n25071__, new_new_n25072__, new_new_n25073__, new_new_n25074__,
    new_new_n25075__, new_new_n25076__, new_new_n25077__, new_new_n25078__,
    new_new_n25079__, new_new_n25080__, new_new_n25081__, new_new_n25082__,
    new_new_n25083__, new_new_n25084__, new_new_n25085__, new_new_n25086__,
    new_new_n25087__, new_new_n25088__, new_new_n25089__, new_new_n25090__,
    new_new_n25091__, new_new_n25092__, new_new_n25093__, new_new_n25094__,
    new_new_n25095__, new_new_n25096__, new_new_n25097__, new_new_n25098__,
    new_new_n25099__, new_new_n25100__, new_new_n25101__, new_new_n25102__,
    new_new_n25103__, new_new_n25104__, new_new_n25105__, new_new_n25106__,
    new_new_n25107__, new_new_n25109__, new_new_n25110__, new_new_n25111__,
    new_new_n25112__, new_new_n25113__, new_new_n25114__, new_new_n25115__,
    new_new_n25116__, new_new_n25117__, new_new_n25118__, new_new_n25119__,
    new_new_n25120__, new_new_n25121__, new_new_n25122__, new_new_n25123__,
    new_new_n25124__, new_new_n25125__, new_new_n25126__, new_new_n25127__,
    new_new_n25128__, new_new_n25129__, new_new_n25130__, new_new_n25131__,
    new_new_n25132__, new_new_n25133__, new_new_n25134__, new_new_n25135__,
    new_new_n25136__, new_new_n25137__, new_new_n25138__, new_new_n25139__,
    new_new_n25140__, new_new_n25141__, new_new_n25142__, new_new_n25143__,
    new_new_n25144__, new_new_n25145__, new_new_n25146__, new_new_n25147__,
    new_new_n25148__, new_new_n25149__, new_new_n25150__, new_new_n25151__,
    new_new_n25152__, new_new_n25153__, new_new_n25154__, new_new_n25155__,
    new_new_n25156__, new_new_n25157__, new_new_n25158__, new_new_n25159__,
    new_new_n25160__, new_new_n25161__, new_new_n25162__, new_new_n25163__,
    new_new_n25164__, new_new_n25165__, new_new_n25166__, new_new_n25167__,
    new_new_n25168__, new_new_n25169__, new_new_n25170__, new_new_n25171__,
    new_new_n25172__, new_new_n25173__, new_new_n25174__, new_new_n25175__,
    new_new_n25176__, new_new_n25177__, new_new_n25178__, new_new_n25179__,
    new_new_n25180__, new_new_n25181__, new_new_n25182__, new_new_n25183__,
    new_new_n25184__, new_new_n25185__, new_new_n25186__, new_new_n25187__,
    new_new_n25188__, new_new_n25189__, new_new_n25190__, new_new_n25191__,
    new_new_n25193__, new_new_n25194__, new_new_n25195__, new_new_n25196__,
    new_new_n25197__, new_new_n25198__, new_new_n25199__, new_new_n25200__,
    new_new_n25201__, new_new_n25202__, new_new_n25203__, new_new_n25204__,
    new_new_n25205__, new_new_n25206__, new_new_n25207__, new_new_n25208__,
    new_new_n25209__, new_new_n25210__, new_new_n25211__, new_new_n25212__,
    new_new_n25213__, new_new_n25214__, new_new_n25215__, new_new_n25216__,
    new_new_n25217__, new_new_n25218__, new_new_n25219__, new_new_n25220__,
    new_new_n25221__, new_new_n25222__, new_new_n25223__, new_new_n25224__,
    new_new_n25225__, new_new_n25226__, new_new_n25227__, new_new_n25228__,
    new_new_n25229__, new_new_n25230__, new_new_n25231__, new_new_n25232__,
    new_new_n25233__, new_new_n25234__, new_new_n25235__, new_new_n25236__,
    new_new_n25237__, new_new_n25238__, new_new_n25239__, new_new_n25240__,
    new_new_n25241__, new_new_n25242__, new_new_n25243__, new_new_n25244__,
    new_new_n25245__, new_new_n25246__, new_new_n25247__, new_new_n25248__,
    new_new_n25249__, new_new_n25250__, new_new_n25251__, new_new_n25252__,
    new_new_n25253__, new_new_n25254__, new_new_n25255__, new_new_n25256__,
    new_new_n25257__, new_new_n25258__, new_new_n25259__, new_new_n25260__,
    new_new_n25261__, new_new_n25262__, new_new_n25263__, new_new_n25264__,
    new_new_n25265__, new_new_n25266__, new_new_n25267__, new_new_n25269__,
    new_new_n25270__, new_new_n25271__, new_new_n25272__, new_new_n25273__,
    new_new_n25274__, new_new_n25275__, new_new_n25276__, new_new_n25277__,
    new_new_n25278__, new_new_n25279__, new_new_n25280__, new_new_n25281__,
    new_new_n25282__, new_new_n25283__, new_new_n25284__, new_new_n25285__,
    new_new_n25286__, new_new_n25287__, new_new_n25288__, new_new_n25289__,
    new_new_n25290__, new_new_n25291__, new_new_n25292__, new_new_n25293__,
    new_new_n25294__, new_new_n25295__, new_new_n25296__, new_new_n25297__,
    new_new_n25298__, new_new_n25299__, new_new_n25300__, new_new_n25301__,
    new_new_n25302__, new_new_n25303__, new_new_n25304__, new_new_n25305__,
    new_new_n25306__, new_new_n25307__, new_new_n25308__, new_new_n25309__,
    new_new_n25310__, new_new_n25311__, new_new_n25312__, new_new_n25313__,
    new_new_n25314__, new_new_n25315__, new_new_n25316__, new_new_n25317__,
    new_new_n25318__, new_new_n25319__, new_new_n25320__, new_new_n25321__,
    new_new_n25322__, new_new_n25323__, new_new_n25324__, new_new_n25325__,
    new_new_n25326__, new_new_n25327__, new_new_n25328__, new_new_n25329__,
    new_new_n25330__, new_new_n25331__, new_new_n25332__, new_new_n25333__,
    new_new_n25334__, new_new_n25335__, new_new_n25336__, new_new_n25337__,
    new_new_n25338__, new_new_n25339__, new_new_n25340__, new_new_n25341__,
    new_new_n25342__, new_new_n25343__, new_new_n25344__, new_new_n25345__,
    new_new_n25346__, new_new_n25347__, new_new_n25349__, new_new_n25350__,
    new_new_n25351__, new_new_n25352__, new_new_n25353__, new_new_n25354__,
    new_new_n25355__, new_new_n25356__, new_new_n25357__, new_new_n25358__,
    new_new_n25359__, new_new_n25360__, new_new_n25361__, new_new_n25362__,
    new_new_n25363__, new_new_n25364__, new_new_n25365__, new_new_n25366__,
    new_new_n25367__, new_new_n25368__, new_new_n25369__, new_new_n25370__,
    new_new_n25371__, new_new_n25372__, new_new_n25373__, new_new_n25374__,
    new_new_n25375__, new_new_n25376__, new_new_n25377__, new_new_n25378__,
    new_new_n25379__, new_new_n25380__, new_new_n25381__, new_new_n25382__,
    new_new_n25383__, new_new_n25384__, new_new_n25385__, new_new_n25386__,
    new_new_n25387__, new_new_n25388__, new_new_n25389__, new_new_n25390__,
    new_new_n25391__, new_new_n25392__, new_new_n25393__, new_new_n25394__,
    new_new_n25395__, new_new_n25396__, new_new_n25397__, new_new_n25398__,
    new_new_n25399__, new_new_n25400__, new_new_n25401__, new_new_n25402__,
    new_new_n25403__, new_new_n25404__, new_new_n25405__, new_new_n25406__,
    new_new_n25407__, new_new_n25408__, new_new_n25409__, new_new_n25410__,
    new_new_n25411__, new_new_n25412__, new_new_n25413__, new_new_n25414__,
    new_new_n25415__, new_new_n25416__, new_new_n25417__, new_new_n25418__,
    new_new_n25419__, new_new_n25420__, new_new_n25421__, new_new_n25423__,
    new_new_n25424__, new_new_n25425__, new_new_n25426__, new_new_n25427__,
    new_new_n25428__, new_new_n25429__, new_new_n25430__, new_new_n25431__,
    new_new_n25432__, new_new_n25433__, new_new_n25434__, new_new_n25435__,
    new_new_n25436__, new_new_n25437__, new_new_n25438__, new_new_n25439__,
    new_new_n25440__, new_new_n25441__, new_new_n25442__, new_new_n25443__,
    new_new_n25444__, new_new_n25445__, new_new_n25446__, new_new_n25447__,
    new_new_n25448__, new_new_n25449__, new_new_n25450__, new_new_n25451__,
    new_new_n25452__, new_new_n25453__, new_new_n25454__, new_new_n25455__,
    new_new_n25456__, new_new_n25457__, new_new_n25458__, new_new_n25459__,
    new_new_n25460__, new_new_n25461__, new_new_n25462__, new_new_n25463__,
    new_new_n25464__, new_new_n25465__, new_new_n25466__, new_new_n25467__,
    new_new_n25468__, new_new_n25469__, new_new_n25470__, new_new_n25471__,
    new_new_n25472__, new_new_n25473__, new_new_n25474__, new_new_n25475__,
    new_new_n25476__, new_new_n25477__, new_new_n25478__, new_new_n25479__,
    new_new_n25480__, new_new_n25481__, new_new_n25482__, new_new_n25483__,
    new_new_n25484__, new_new_n25485__, new_new_n25486__, new_new_n25487__,
    new_new_n25488__, new_new_n25489__, new_new_n25490__, new_new_n25491__,
    new_new_n25492__, new_new_n25493__, new_new_n25494__, new_new_n25495__,
    new_new_n25496__, new_new_n25497__, new_new_n25498__, new_new_n25499__,
    new_new_n25500__, new_new_n25501__, new_new_n25502__, new_new_n25503__,
    new_new_n25504__, new_new_n25505__, new_new_n25506__, new_new_n25507__,
    new_new_n25508__, new_new_n25509__, new_new_n25510__, new_new_n25511__,
    new_new_n25512__, new_new_n25514__, new_new_n25515__, new_new_n25516__,
    new_new_n25517__, new_new_n25518__, new_new_n25519__, new_new_n25520__,
    new_new_n25521__, new_new_n25522__, new_new_n25523__, new_new_n25524__,
    new_new_n25525__, new_new_n25526__, new_new_n25527__, new_new_n25528__,
    new_new_n25529__, new_new_n25530__, new_new_n25531__, new_new_n25532__,
    new_new_n25533__, new_new_n25534__, new_new_n25535__, new_new_n25536__,
    new_new_n25537__, new_new_n25539__, new_new_n25540__, new_new_n25541__,
    new_new_n25542__, new_new_n25543__, new_new_n25544__, new_new_n25545__,
    new_new_n25546__, new_new_n25547__, new_new_n25548__, new_new_n25549__,
    new_new_n25550__, new_new_n25551__, new_new_n25552__, new_new_n25553__,
    new_new_n25554__, new_new_n25555__, new_new_n25556__, new_new_n25557__,
    new_new_n25558__, new_new_n25559__, new_new_n25560__, new_new_n25561__,
    new_new_n25562__, new_new_n25563__, new_new_n25564__, new_new_n25566__,
    new_new_n25567__, new_new_n25568__, new_new_n25569__, new_new_n25570__,
    new_new_n25571__, new_new_n25572__, new_new_n25573__, new_new_n25574__,
    new_new_n25575__, new_new_n25576__, new_new_n25577__, new_new_n25578__,
    new_new_n25579__, new_new_n25580__, new_new_n25581__, new_new_n25582__,
    new_new_n25583__, new_new_n25584__, new_new_n25585__, new_new_n25586__,
    new_new_n25587__, new_new_n25588__, new_new_n25589__, new_new_n25590__,
    new_new_n25591__, new_new_n25593__, new_new_n25594__, new_new_n25595__,
    new_new_n25596__, new_new_n25597__, new_new_n25598__, new_new_n25599__,
    new_new_n25600__, new_new_n25601__, new_new_n25602__, new_new_n25603__,
    new_new_n25604__, new_new_n25605__, new_new_n25606__, new_new_n25607__,
    new_new_n25608__, new_new_n25609__, new_new_n25610__, new_new_n25611__,
    new_new_n25612__, new_new_n25613__, new_new_n25614__, new_new_n25615__,
    new_new_n25616__, new_new_n25617__, new_new_n25618__, new_new_n25619__,
    new_new_n25620__, new_new_n25621__, new_new_n25623__, new_new_n25624__,
    new_new_n25625__, new_new_n25626__, new_new_n25627__, new_new_n25628__,
    new_new_n25629__, new_new_n25630__, new_new_n25631__, new_new_n25632__,
    new_new_n25633__, new_new_n25634__, new_new_n25635__, new_new_n25636__,
    new_new_n25637__, new_new_n25638__, new_new_n25639__, new_new_n25640__,
    new_new_n25641__, new_new_n25642__, new_new_n25643__, new_new_n25644__,
    new_new_n25645__, new_new_n25646__, new_new_n25647__, new_new_n25648__,
    new_new_n25650__, new_new_n25651__, new_new_n25652__, new_new_n25653__,
    new_new_n25654__, new_new_n25655__, new_new_n25656__, new_new_n25657__,
    new_new_n25658__, new_new_n25659__, new_new_n25660__, new_new_n25661__,
    new_new_n25662__, new_new_n25663__, new_new_n25664__, new_new_n25665__,
    new_new_n25666__, new_new_n25667__, new_new_n25668__, new_new_n25669__,
    new_new_n25670__, new_new_n25671__, new_new_n25672__, new_new_n25673__,
    new_new_n25674__, new_new_n25675__, new_new_n25676__, new_new_n25677__,
    new_new_n25678__, new_new_n25680__, new_new_n25681__, new_new_n25682__,
    new_new_n25683__, new_new_n25684__, new_new_n25685__, new_new_n25686__,
    new_new_n25687__, new_new_n25688__, new_new_n25689__, new_new_n25690__,
    new_new_n25691__, new_new_n25692__, new_new_n25693__, new_new_n25694__,
    new_new_n25695__, new_new_n25696__, new_new_n25697__, new_new_n25698__,
    new_new_n25699__, new_new_n25700__, new_new_n25701__, new_new_n25702__,
    new_new_n25703__, new_new_n25704__, new_new_n25705__, new_new_n25707__,
    new_new_n25708__, new_new_n25709__, new_new_n25710__, new_new_n25711__,
    new_new_n25712__, new_new_n25713__, new_new_n25714__, new_new_n25715__,
    new_new_n25716__, new_new_n25717__, new_new_n25718__, new_new_n25719__,
    new_new_n25720__, new_new_n25721__, new_new_n25722__, new_new_n25723__,
    new_new_n25724__, new_new_n25725__, new_new_n25726__, new_new_n25727__,
    new_new_n25728__, new_new_n25729__, new_new_n25730__, new_new_n25731__,
    new_new_n25732__, new_new_n25733__, new_new_n25734__, new_new_n25735__,
    new_new_n25736__, new_new_n25737__, new_new_n25738__, new_new_n25740__,
    new_new_n25741__, new_new_n25742__, new_new_n25743__, new_new_n25744__,
    new_new_n25745__, new_new_n25746__, new_new_n25747__, new_new_n25748__,
    new_new_n25749__, new_new_n25750__, new_new_n25751__, new_new_n25752__,
    new_new_n25753__, new_new_n25754__, new_new_n25755__, new_new_n25756__,
    new_new_n25757__, new_new_n25758__, new_new_n25759__, new_new_n25760__,
    new_new_n25761__, new_new_n25762__, new_new_n25763__, new_new_n25764__,
    new_new_n25765__, new_new_n25767__, new_new_n25768__, new_new_n25769__,
    new_new_n25770__, new_new_n25771__, new_new_n25772__, new_new_n25773__,
    new_new_n25774__, new_new_n25775__, new_new_n25776__, new_new_n25777__,
    new_new_n25778__, new_new_n25779__, new_new_n25780__, new_new_n25781__,
    new_new_n25782__, new_new_n25783__, new_new_n25784__, new_new_n25785__,
    new_new_n25786__, new_new_n25787__, new_new_n25788__, new_new_n25789__,
    new_new_n25790__, new_new_n25791__, new_new_n25792__, new_new_n25793__,
    new_new_n25794__, new_new_n25795__, new_new_n25797__, new_new_n25798__,
    new_new_n25799__, new_new_n25800__, new_new_n25801__, new_new_n25802__,
    new_new_n25803__, new_new_n25804__, new_new_n25805__, new_new_n25806__,
    new_new_n25807__, new_new_n25808__, new_new_n25809__, new_new_n25810__,
    new_new_n25811__, new_new_n25812__, new_new_n25813__, new_new_n25814__,
    new_new_n25815__, new_new_n25816__, new_new_n25817__, new_new_n25818__,
    new_new_n25819__, new_new_n25820__, new_new_n25821__, new_new_n25822__,
    new_new_n25824__, new_new_n25825__, new_new_n25826__, new_new_n25827__,
    new_new_n25828__, new_new_n25829__, new_new_n25830__, new_new_n25831__,
    new_new_n25832__, new_new_n25833__, new_new_n25834__, new_new_n25835__,
    new_new_n25836__, new_new_n25837__, new_new_n25838__, new_new_n25839__,
    new_new_n25840__, new_new_n25841__, new_new_n25842__, new_new_n25843__,
    new_new_n25844__, new_new_n25845__, new_new_n25846__, new_new_n25847__,
    new_new_n25848__, new_new_n25849__, new_new_n25850__, new_new_n25851__,
    new_new_n25852__, new_new_n25853__, new_new_n25854__, new_new_n25855__,
    new_new_n25857__, new_new_n25858__, new_new_n25859__, new_new_n25860__,
    new_new_n25861__, new_new_n25862__, new_new_n25863__, new_new_n25864__,
    new_new_n25865__, new_new_n25866__, new_new_n25867__, new_new_n25868__,
    new_new_n25869__, new_new_n25870__, new_new_n25871__, new_new_n25872__,
    new_new_n25873__, new_new_n25874__, new_new_n25875__, new_new_n25876__,
    new_new_n25877__, new_new_n25878__, new_new_n25879__, new_new_n25880__,
    new_new_n25881__, new_new_n25882__, new_new_n25884__, new_new_n25885__,
    new_new_n25886__, new_new_n25887__, new_new_n25888__, new_new_n25889__,
    new_new_n25890__, new_new_n25891__, new_new_n25892__, new_new_n25893__,
    new_new_n25894__, new_new_n25895__, new_new_n25896__, new_new_n25897__,
    new_new_n25898__, new_new_n25899__, new_new_n25900__, new_new_n25901__,
    new_new_n25902__, new_new_n25903__, new_new_n25904__, new_new_n25905__,
    new_new_n25906__, new_new_n25907__, new_new_n25908__, new_new_n25909__,
    new_new_n25910__, new_new_n25911__, new_new_n25912__, new_new_n25914__,
    new_new_n25915__, new_new_n25916__, new_new_n25917__, new_new_n25918__,
    new_new_n25919__, new_new_n25920__, new_new_n25921__, new_new_n25922__,
    new_new_n25923__, new_new_n25924__, new_new_n25925__, new_new_n25926__,
    new_new_n25927__, new_new_n25928__, new_new_n25929__, new_new_n25930__,
    new_new_n25931__, new_new_n25932__, new_new_n25933__, new_new_n25934__,
    new_new_n25935__, new_new_n25936__, new_new_n25937__, new_new_n25938__,
    new_new_n25939__, new_new_n25941__, new_new_n25942__, new_new_n25943__,
    new_new_n25944__, new_new_n25945__, new_new_n25946__, new_new_n25947__,
    new_new_n25948__, new_new_n25949__, new_new_n25950__, new_new_n25951__,
    new_new_n25952__, new_new_n25953__, new_new_n25954__, new_new_n25955__,
    new_new_n25956__, new_new_n25957__, new_new_n25958__, new_new_n25959__,
    new_new_n25960__, new_new_n25961__, new_new_n25962__, new_new_n25963__,
    new_new_n25964__, new_new_n25966__, new_new_n25967__, new_new_n25968__,
    new_new_n25969__, new_new_n25970__, new_new_n25971__, new_new_n25972__,
    new_new_n25973__, new_new_n25974__, new_new_n25976__, new_new_n25977__,
    new_new_n25978__, new_new_n25980__, new_new_n25981__, new_new_n25982__,
    new_new_n25983__, new_new_n25984__, new_new_n25985__, new_new_n25986__,
    new_new_n25987__, new_new_n25988__, new_new_n25990__, new_new_n25991__,
    new_new_n25992__, new_new_n25993__, new_new_n25994__, new_new_n25995__,
    new_new_n25996__, new_new_n25997__, new_new_n25998__, new_new_n26000__,
    new_new_n26001__, new_new_n26002__, new_new_n26003__, new_new_n26004__,
    new_new_n26005__, new_new_n26006__, new_new_n26007__, new_new_n26008__,
    new_new_n26010__, new_new_n26011__, new_new_n26012__, new_new_n26013__,
    new_new_n26014__, new_new_n26015__, new_new_n26016__, new_new_n26017__,
    new_new_n26018__, new_new_n26020__, new_new_n26021__, new_new_n26022__,
    new_new_n26023__, new_new_n26024__, new_new_n26025__, new_new_n26026__,
    new_new_n26027__, new_new_n26028__, new_new_n26030__, new_new_n26031__,
    new_new_n26032__, new_new_n26033__, new_new_n26034__, new_new_n26035__,
    new_new_n26036__, new_new_n26037__, new_new_n26038__, new_new_n26040__,
    new_new_n26041__, new_new_n26042__, new_new_n26043__, new_new_n26044__,
    new_new_n26045__, new_new_n26046__, new_new_n26047__, new_new_n26048__,
    new_new_n26050__, new_new_n26051__, new_new_n26052__, new_new_n26053__,
    new_new_n26054__, new_new_n26055__, new_new_n26056__, new_new_n26057__,
    new_new_n26058__, new_new_n26060__, new_new_n26061__, new_new_n26062__,
    new_new_n26063__, new_new_n26064__, new_new_n26065__, new_new_n26066__,
    new_new_n26067__, new_new_n26068__, new_new_n26070__, new_new_n26071__,
    new_new_n26072__, new_new_n26073__, new_new_n26074__, new_new_n26075__,
    new_new_n26076__, new_new_n26077__, new_new_n26078__, new_new_n26080__,
    new_new_n26081__, new_new_n26082__, new_new_n26083__, new_new_n26084__,
    new_new_n26085__, new_new_n26086__, new_new_n26087__, new_new_n26088__,
    new_new_n26090__, new_new_n26091__, new_new_n26092__, new_new_n26093__,
    new_new_n26094__, new_new_n26095__, new_new_n26096__, new_new_n26097__,
    new_new_n26098__, new_new_n26100__, new_new_n26101__, new_new_n26102__,
    new_new_n26103__, new_new_n26104__, new_new_n26105__, new_new_n26106__,
    new_new_n26107__, new_new_n26108__, new_new_n26110__, new_new_n26111__,
    new_new_n26112__, new_new_n26113__, new_new_n26114__, new_new_n26115__,
    new_new_n26116__, new_new_n26117__, new_new_n26118__, new_new_n26120__,
    new_new_n26121__, new_new_n26122__, new_new_n26123__, new_new_n26124__,
    new_new_n26125__, new_new_n26126__, new_new_n26127__, new_new_n26128__,
    new_new_n26130__, new_new_n26131__, new_new_n26132__, new_new_n26133__,
    new_new_n26134__, new_new_n26135__, new_new_n26136__, new_new_n26137__,
    new_new_n26138__, new_new_n26140__, new_new_n26141__, new_new_n26142__,
    new_new_n26144__, new_new_n26145__, new_new_n26146__, new_new_n26147__,
    new_new_n26148__, new_new_n26149__, new_new_n26150__, new_new_n26151__,
    new_new_n26152__, new_new_n26154__, new_new_n26155__, new_new_n26157__,
    new_new_n26158__, new_new_n26160__, new_new_n26161__, new_new_n26163__,
    new_new_n26164__, new_new_n26166__, new_new_n26167__, new_new_n26168__,
    new_new_n26169__, new_new_n26170__, new_new_n26171__, new_new_n26172__,
    new_new_n26173__, new_new_n26174__, new_new_n26175__, new_new_n26177__,
    new_new_n26178__, new_new_n26179__, new_new_n26180__, new_new_n26181__,
    new_new_n26182__, new_new_n26183__, new_new_n26184__, new_new_n26185__,
    new_new_n26186__, new_new_n26188__, new_new_n26189__, new_new_n26190__,
    new_new_n26191__, new_new_n26192__, new_new_n26193__, new_new_n26194__,
    new_new_n26195__, new_new_n26196__, new_new_n26197__, new_new_n26199__,
    new_new_n26200__, new_new_n26201__, new_new_n26202__, new_new_n26203__,
    new_new_n26204__, new_new_n26205__, new_new_n26206__, new_new_n26207__,
    new_new_n26208__, new_new_n26209__, new_new_n26211__, new_new_n26212__,
    new_new_n26213__, new_new_n26214__, new_new_n26216__, new_new_n26217__,
    new_new_n26218__, new_new_n26219__, new_new_n26220__, new_new_n26222__,
    new_new_n26223__, new_new_n26225__, new_new_n26226__, new_new_n26227__,
    new_new_n26228__, new_new_n26229__, new_new_n26230__, new_new_n26231__,
    new_new_n26232__, new_new_n26233__, new_new_n26234__, new_new_n26235__,
    new_new_n26236__, new_new_n26237__, new_new_n26239__, new_new_n26240__,
    new_new_n26242__, new_new_n26243__, new_new_n26244__, new_new_n26245__,
    new_new_n26246__, new_new_n26247__, new_new_n26248__, new_new_n26249__,
    new_new_n26250__, new_new_n26252__, new_new_n26253__, new_new_n26254__,
    new_new_n26255__, new_new_n26256__, new_new_n26257__, new_new_n26258__,
    new_new_n26260__, new_new_n26261__, new_new_n26262__, new_new_n26263__,
    new_new_n26265__, new_new_n26271__, new_new_n26272__, new_new_n26273__,
    new_new_n26274__, new_new_n26275__, new_new_n26276__, new_new_n26277__,
    new_new_n26278__, new_new_n26280__, new_new_n26281__, new_new_n26282__,
    new_new_n26283__, new_new_n26285__, new_new_n26286__, new_new_n26287__,
    new_new_n26288__, new_new_n26289__, new_new_n26291__, new_new_n26292__,
    new_new_n26293__, new_new_n26294__, new_new_n26295__, new_new_n26296__,
    new_new_n26297__, new_new_n26298__, new_new_n26299__, new_new_n26300__,
    new_new_n26301__, new_new_n26302__, new_new_n26304__, new_new_n26306__,
    new_new_n26307__, new_new_n26308__, new_new_n26310__, new_new_n26311__,
    new_new_n26312__, new_new_n26313__, new_new_n26314__, new_new_n26315__,
    new_new_n26316__, new_new_n26317__, new_new_n26318__, new_new_n26319__,
    new_new_n26320__, new_new_n26321__, new_new_n26323__, new_new_n26324__,
    new_new_n26325__, new_new_n26326__, new_new_n26328__, new_new_n26329__,
    new_new_n26330__, new_new_n26331__, new_new_n26332__, new_new_n26333__,
    new_new_n26334__, new_new_n26335__, new_new_n26336__, new_new_n26337__,
    new_new_n26338__, new_new_n26339__, new_new_n26340__, new_new_n26342__,
    new_new_n26343__, new_new_n26344__, new_new_n26345__, new_new_n26346__,
    new_new_n26347__, new_new_n26348__, new_new_n26349__, new_new_n26350__,
    new_new_n26352__, new_new_n26353__, new_new_n26354__, new_new_n26355__,
    new_new_n26356__, new_new_n26357__, new_new_n26358__, new_new_n26359__,
    new_new_n26360__, new_new_n26361__, new_new_n26363__, new_new_n26364__,
    new_new_n26365__, new_new_n26366__, new_new_n26367__, new_new_n26368__,
    new_new_n26369__, new_new_n26370__, new_new_n26371__, new_new_n26372__,
    new_new_n26374__, new_new_n26375__, new_new_n26376__, new_new_n26377__,
    new_new_n26378__, new_new_n26379__, new_new_n26380__, new_new_n26381__,
    new_new_n26382__, new_new_n26384__, new_new_n26385__, new_new_n26386__,
    new_new_n26387__, new_new_n26388__, new_new_n26389__, new_new_n26390__,
    new_new_n26391__, new_new_n26392__, new_new_n26394__, new_new_n26395__,
    new_new_n26396__, new_new_n26397__, new_new_n26398__, new_new_n26399__,
    new_new_n26400__, new_new_n26401__, new_new_n26402__, new_new_n26404__,
    new_new_n26405__, new_new_n26406__, new_new_n26407__, new_new_n26408__,
    new_new_n26409__, new_new_n26410__, new_new_n26411__, new_new_n26412__,
    new_new_n26414__, new_new_n26415__, new_new_n26416__, new_new_n26417__,
    new_new_n26418__, new_new_n26419__, new_new_n26420__, new_new_n26421__,
    new_new_n26422__, new_new_n26424__, new_new_n26425__, new_new_n26426__,
    new_new_n26427__, new_new_n26428__, new_new_n26429__, new_new_n26430__,
    new_new_n26431__, new_new_n26432__, new_new_n26434__, new_new_n26435__,
    new_new_n26436__, new_new_n26437__, new_new_n26438__, new_new_n26439__,
    new_new_n26440__, new_new_n26441__, new_new_n26442__, new_new_n26444__,
    new_new_n26445__, new_new_n26446__, new_new_n26447__, new_new_n26448__,
    new_new_n26449__, new_new_n26450__, new_new_n26451__, new_new_n26452__,
    new_new_n26454__, new_new_n26455__, new_new_n26456__, new_new_n26457__,
    new_new_n26458__, new_new_n26459__, new_new_n26460__, new_new_n26461__,
    new_new_n26462__, new_new_n26464__, new_new_n26465__, new_new_n26466__,
    new_new_n26467__, new_new_n26468__, new_new_n26469__, new_new_n26470__,
    new_new_n26471__, new_new_n26472__, new_new_n26474__, new_new_n26475__,
    new_new_n26476__, new_new_n26477__, new_new_n26478__, new_new_n26479__,
    new_new_n26480__, new_new_n26481__, new_new_n26482__, new_new_n26484__,
    new_new_n26485__, new_new_n26486__, new_new_n26487__, new_new_n26488__,
    new_new_n26489__, new_new_n26490__, new_new_n26491__, new_new_n26492__,
    new_new_n26494__, new_new_n26495__, new_new_n26496__, new_new_n26497__,
    new_new_n26498__, new_new_n26499__, new_new_n26500__, new_new_n26501__,
    new_new_n26502__, new_new_n26504__, new_new_n26505__, new_new_n26506__,
    new_new_n26507__, new_new_n26508__, new_new_n26509__, new_new_n26510__,
    new_new_n26511__, new_new_n26512__, new_new_n26514__, new_new_n26515__,
    new_new_n26516__, new_new_n26517__, new_new_n26518__, new_new_n26519__,
    new_new_n26520__, new_new_n26521__, new_new_n26522__, new_new_n26524__,
    new_new_n26525__, new_new_n26526__, new_new_n26527__, new_new_n26528__,
    new_new_n26529__, new_new_n26530__, new_new_n26531__, new_new_n26532__,
    new_new_n26533__, new_new_n26535__, new_new_n26536__, new_new_n26537__,
    new_new_n26538__, new_new_n26539__, new_new_n26540__, new_new_n26541__,
    new_new_n26542__, new_new_n26543__, new_new_n26544__, new_new_n26546__,
    new_new_n26547__, new_new_n26548__, new_new_n26549__, new_new_n26550__,
    new_new_n26551__, new_new_n26552__, new_new_n26553__, new_new_n26554__,
    new_new_n26556__, new_new_n26557__, new_new_n26558__, new_new_n26559__,
    new_new_n26560__, new_new_n26561__, new_new_n26562__, new_new_n26563__,
    new_new_n26564__, new_new_n26566__, new_new_n26567__, new_new_n26568__,
    new_new_n26569__, new_new_n26570__, new_new_n26571__, new_new_n26572__,
    new_new_n26573__, new_new_n26574__, new_new_n26576__, new_new_n26577__,
    new_new_n26578__, new_new_n26579__, new_new_n26580__, new_new_n26581__,
    new_new_n26582__, new_new_n26583__, new_new_n26584__, new_new_n26586__,
    new_new_n26587__, new_new_n26588__, new_new_n26589__, new_new_n26590__,
    new_new_n26591__, new_new_n26592__, new_new_n26593__, new_new_n26594__,
    new_new_n26596__, new_new_n26597__, new_new_n26598__, new_new_n26599__,
    new_new_n26600__, new_new_n26601__, new_new_n26602__, new_new_n26603__,
    new_new_n26604__, new_new_n26605__, new_new_n26607__, new_new_n26608__,
    new_new_n26609__, new_new_n26610__, new_new_n26611__, new_new_n26612__,
    new_new_n26613__, new_new_n26614__, new_new_n26615__, new_new_n26617__,
    new_new_n26618__, new_new_n26619__, new_new_n26620__, new_new_n26621__,
    new_new_n26622__, new_new_n26623__, new_new_n26624__, new_new_n26625__,
    new_new_n26627__, new_new_n26628__, new_new_n26629__, new_new_n26630__,
    new_new_n26631__, new_new_n26632__, new_new_n26633__, new_new_n26634__,
    new_new_n26635__, new_new_n26636__, new_new_n26638__, new_new_n26639__,
    new_new_n26640__, new_new_n26641__, new_new_n26642__, new_new_n26643__,
    new_new_n26644__, new_new_n26645__, new_new_n26646__, new_new_n26648__,
    new_new_n26649__, new_new_n26650__, new_new_n26651__, new_new_n26652__,
    new_new_n26653__, new_new_n26654__, new_new_n26655__, new_new_n26656__,
    new_new_n26658__, new_new_n26659__, new_new_n26660__, new_new_n26661__,
    new_new_n26662__, new_new_n26663__, new_new_n26664__, new_new_n26665__,
    new_new_n26666__, new_new_n26667__, new_new_n26668__, new_new_n26669__,
    new_new_n26670__, new_new_n26671__, new_new_n26672__, new_new_n26673__,
    new_new_n26674__, new_new_n26675__, new_new_n26676__, new_new_n26677__,
    new_new_n26678__, new_new_n26679__, new_new_n26680__, new_new_n26681__,
    new_new_n26682__, new_new_n26683__, new_new_n26684__, new_new_n26685__,
    new_new_n26686__, new_new_n26687__, new_new_n26688__, new_new_n26689__,
    new_new_n26690__, new_new_n26691__, new_new_n26692__, new_new_n26693__,
    new_new_n26694__, new_new_n26696__, new_new_n26697__, new_new_n26698__,
    new_new_n26699__, new_new_n26700__, new_new_n26701__, new_new_n26702__,
    new_new_n26703__, new_new_n26704__, new_new_n26705__, new_new_n26706__,
    new_new_n26707__, new_new_n26709__, new_new_n26710__, new_new_n26711__,
    new_new_n26712__, new_new_n26713__, new_new_n26714__, new_new_n26716__,
    new_new_n26717__, new_new_n26718__, new_new_n26719__, new_new_n26720__,
    new_new_n26721__, new_new_n26723__, new_new_n26724__, new_new_n26725__,
    new_new_n26726__, new_new_n26727__, new_new_n26728__, new_new_n26734__,
    new_new_n26735__, new_new_n26736__, new_new_n26737__, new_new_n26738__,
    new_new_n26739__, new_new_n26740__, new_new_n26741__, new_new_n26742__,
    new_new_n26743__, new_new_n26745__, new_new_n26746__, new_new_n26747__,
    new_new_n26748__, new_new_n26749__, new_new_n26751__, new_new_n26752__,
    new_new_n26753__, new_new_n26754__, new_new_n26755__, new_new_n26757__,
    new_new_n26758__, new_new_n26759__, new_new_n26760__, new_new_n26761__,
    new_new_n26763__, new_new_n26764__, new_new_n26765__, new_new_n26766__,
    new_new_n26767__, new_new_n26768__, new_new_n26769__, new_new_n26770__,
    new_new_n26771__, new_new_n26772__, new_new_n26773__, new_new_n26774__,
    new_new_n26775__, new_new_n26776__, new_new_n26777__, new_new_n26778__,
    new_new_n26779__, new_new_n26780__, new_new_n26781__, new_new_n26782__,
    new_new_n26783__, new_new_n26784__, new_new_n26785__, new_new_n26786__,
    new_new_n26787__, new_new_n26788__, new_new_n26789__, new_new_n26790__,
    new_new_n26791__, new_new_n26792__, new_new_n26793__, new_new_n26794__,
    new_new_n26795__, new_new_n26796__, new_new_n26797__, new_new_n26798__,
    new_new_n26799__, new_new_n26800__, new_new_n26801__, new_new_n26802__,
    new_new_n26803__, new_new_n26804__, new_new_n26805__, new_new_n26806__,
    new_new_n26807__, new_new_n26808__, new_new_n26809__, new_new_n26810__,
    new_new_n26811__, new_new_n26812__, new_new_n26813__, new_new_n26814__,
    new_new_n26815__, new_new_n26816__, new_new_n26817__, new_new_n26818__,
    new_new_n26819__, new_new_n26820__, new_new_n26821__, new_new_n26822__,
    new_new_n26823__, new_new_n26824__, new_new_n26825__, new_new_n26826__,
    new_new_n26827__, new_new_n26828__, new_new_n26829__, new_new_n26830__,
    new_new_n26831__, new_new_n26832__, new_new_n26833__, new_new_n26834__,
    new_new_n26835__, new_new_n26836__, new_new_n26837__, new_new_n26838__,
    new_new_n26839__, new_new_n26840__, new_new_n26841__, new_new_n26842__,
    new_new_n26843__, new_new_n26844__, new_new_n26845__, new_new_n26846__,
    new_new_n26847__, new_new_n26848__, new_new_n26849__, new_new_n26850__,
    new_new_n26851__, new_new_n26852__, new_new_n26853__, new_new_n26854__,
    new_new_n26855__, new_new_n26856__, new_new_n26857__, new_new_n26858__,
    new_new_n26859__, new_new_n26860__, new_new_n26861__, new_new_n26862__,
    new_new_n26863__, new_new_n26864__, new_new_n26865__, new_new_n26866__,
    new_new_n26867__, new_new_n26868__, new_new_n26869__, new_new_n26870__,
    new_new_n26871__, new_new_n26872__, new_new_n26873__, new_new_n26874__,
    new_new_n26875__, new_new_n26876__, new_new_n26877__, new_new_n26878__,
    new_new_n26879__, new_new_n26880__, new_new_n26881__, new_new_n26882__,
    new_new_n26883__, new_new_n26884__, new_new_n26886__, new_new_n26887__,
    new_new_n26888__, new_new_n26889__, new_new_n26890__, new_new_n26891__,
    new_new_n26892__, new_new_n26893__, new_new_n26894__, new_new_n26895__,
    new_new_n26896__, new_new_n26897__, new_new_n26898__, new_new_n26899__,
    new_new_n26900__, new_new_n26901__, new_new_n26902__, new_new_n26903__,
    new_new_n26904__, new_new_n26905__, new_new_n26906__, new_new_n26907__,
    new_new_n26908__, new_new_n26909__, new_new_n26910__, new_new_n26911__,
    new_new_n26912__, new_new_n26913__, new_new_n26914__, new_new_n26915__,
    new_new_n26916__, new_new_n26917__, new_new_n26918__, new_new_n26919__,
    new_new_n26920__, new_new_n26921__, new_new_n26922__, new_new_n26923__,
    new_new_n26924__, new_new_n26925__, new_new_n26926__, new_new_n26927__,
    new_new_n26928__, new_new_n26929__, new_new_n26930__, new_new_n26931__,
    new_new_n26932__, new_new_n26933__, new_new_n26934__, new_new_n26935__,
    new_new_n26936__, new_new_n26937__, new_new_n26938__, new_new_n26939__,
    new_new_n26940__, new_new_n26941__, new_new_n26942__, new_new_n26943__,
    new_new_n26944__, new_new_n26945__, new_new_n26946__, new_new_n26947__,
    new_new_n26948__, new_new_n26949__, new_new_n26950__, new_new_n26951__,
    new_new_n26952__, new_new_n26953__, new_new_n26954__, new_new_n26955__,
    new_new_n26956__, new_new_n26957__, new_new_n26958__, new_new_n26959__,
    new_new_n26960__, new_new_n26961__, new_new_n26962__, new_new_n26963__,
    new_new_n26964__, new_new_n26965__, new_new_n26966__, new_new_n26967__,
    new_new_n26968__, new_new_n26969__, new_new_n26970__, new_new_n26971__,
    new_new_n26972__, new_new_n26974__, new_new_n26975__, new_new_n26976__,
    new_new_n26977__, new_new_n26978__, new_new_n26979__, new_new_n26980__,
    new_new_n26981__, new_new_n26982__, new_new_n26983__, new_new_n26984__,
    new_new_n26985__, new_new_n26986__, new_new_n26987__, new_new_n26988__,
    new_new_n26989__, new_new_n26990__, new_new_n26991__, new_new_n26992__,
    new_new_n26993__, new_new_n26994__, new_new_n26995__, new_new_n26996__,
    new_new_n26997__, new_new_n26998__, new_new_n26999__, new_new_n27000__,
    new_new_n27001__, new_new_n27002__, new_new_n27003__, new_new_n27004__,
    new_new_n27005__, new_new_n27006__, new_new_n27007__, new_new_n27008__,
    new_new_n27009__, new_new_n27010__, new_new_n27011__, new_new_n27012__,
    new_new_n27013__, new_new_n27014__, new_new_n27015__, new_new_n27016__,
    new_new_n27017__, new_new_n27018__, new_new_n27019__, new_new_n27020__,
    new_new_n27021__, new_new_n27022__, new_new_n27023__, new_new_n27024__,
    new_new_n27025__, new_new_n27026__, new_new_n27027__, new_new_n27028__,
    new_new_n27029__, new_new_n27030__, new_new_n27031__, new_new_n27032__,
    new_new_n27033__, new_new_n27034__, new_new_n27035__, new_new_n27036__,
    new_new_n27037__, new_new_n27038__, new_new_n27039__, new_new_n27040__,
    new_new_n27041__, new_new_n27042__, new_new_n27043__, new_new_n27044__,
    new_new_n27045__, new_new_n27046__, new_new_n27047__, new_new_n27048__,
    new_new_n27049__, new_new_n27050__, new_new_n27051__, new_new_n27052__,
    new_new_n27053__, new_new_n27054__, new_new_n27055__, new_new_n27056__,
    new_new_n27057__, new_new_n27058__, new_new_n27059__, new_new_n27060__,
    new_new_n27062__, new_new_n27063__, new_new_n27064__, new_new_n27065__,
    new_new_n27066__, new_new_n27067__, new_new_n27068__, new_new_n27069__,
    new_new_n27070__, new_new_n27071__, new_new_n27072__, new_new_n27073__,
    new_new_n27074__, new_new_n27075__, new_new_n27076__, new_new_n27077__,
    new_new_n27078__, new_new_n27079__, new_new_n27080__, new_new_n27081__,
    new_new_n27082__, new_new_n27083__, new_new_n27084__, new_new_n27085__,
    new_new_n27086__, new_new_n27087__, new_new_n27088__, new_new_n27089__,
    new_new_n27090__, new_new_n27091__, new_new_n27092__, new_new_n27093__,
    new_new_n27094__, new_new_n27095__, new_new_n27096__, new_new_n27097__,
    new_new_n27098__, new_new_n27099__, new_new_n27100__, new_new_n27101__,
    new_new_n27102__, new_new_n27103__, new_new_n27104__, new_new_n27105__,
    new_new_n27106__, new_new_n27107__, new_new_n27108__, new_new_n27109__,
    new_new_n27110__, new_new_n27111__, new_new_n27112__, new_new_n27113__,
    new_new_n27114__, new_new_n27115__, new_new_n27116__, new_new_n27117__,
    new_new_n27118__, new_new_n27119__, new_new_n27120__, new_new_n27121__,
    new_new_n27122__, new_new_n27123__, new_new_n27124__, new_new_n27125__,
    new_new_n27126__, new_new_n27127__, new_new_n27128__, new_new_n27129__,
    new_new_n27130__, new_new_n27131__, new_new_n27132__, new_new_n27133__,
    new_new_n27134__, new_new_n27135__, new_new_n27136__, new_new_n27137__,
    new_new_n27138__, new_new_n27139__, new_new_n27140__, new_new_n27141__,
    new_new_n27142__, new_new_n27143__, new_new_n27144__, new_new_n27145__,
    new_new_n27146__, new_new_n27147__, new_new_n27148__, new_new_n27150__,
    new_new_n27151__, new_new_n27152__, new_new_n27153__, new_new_n27154__,
    new_new_n27155__, new_new_n27156__, new_new_n27157__, new_new_n27158__,
    new_new_n27159__, new_new_n27160__, new_new_n27161__, new_new_n27162__,
    new_new_n27163__, new_new_n27164__, new_new_n27165__, new_new_n27166__,
    new_new_n27167__, new_new_n27168__, new_new_n27169__, new_new_n27170__,
    new_new_n27171__, new_new_n27172__, new_new_n27173__, new_new_n27174__,
    new_new_n27175__, new_new_n27176__, new_new_n27177__, new_new_n27178__,
    new_new_n27179__, new_new_n27180__, new_new_n27181__, new_new_n27182__,
    new_new_n27183__, new_new_n27184__, new_new_n27185__, new_new_n27186__,
    new_new_n27187__, new_new_n27188__, new_new_n27189__, new_new_n27190__,
    new_new_n27191__, new_new_n27192__, new_new_n27193__, new_new_n27194__,
    new_new_n27195__, new_new_n27196__, new_new_n27197__, new_new_n27198__,
    new_new_n27199__, new_new_n27200__, new_new_n27201__, new_new_n27202__,
    new_new_n27203__, new_new_n27204__, new_new_n27205__, new_new_n27206__,
    new_new_n27207__, new_new_n27208__, new_new_n27209__, new_new_n27210__,
    new_new_n27211__, new_new_n27212__, new_new_n27213__, new_new_n27214__,
    new_new_n27215__, new_new_n27216__, new_new_n27217__, new_new_n27218__,
    new_new_n27219__, new_new_n27220__, new_new_n27221__, new_new_n27222__,
    new_new_n27223__, new_new_n27224__, new_new_n27225__, new_new_n27226__,
    new_new_n27227__, new_new_n27228__, new_new_n27229__, new_new_n27230__,
    new_new_n27231__, new_new_n27232__, new_new_n27233__, new_new_n27234__,
    new_new_n27235__, new_new_n27236__, new_new_n27238__, new_new_n27239__,
    new_new_n27240__, new_new_n27241__, new_new_n27242__, new_new_n27243__,
    new_new_n27244__, new_new_n27245__, new_new_n27246__, new_new_n27247__,
    new_new_n27248__, new_new_n27249__, new_new_n27250__, new_new_n27251__,
    new_new_n27252__, new_new_n27253__, new_new_n27254__, new_new_n27255__,
    new_new_n27256__, new_new_n27257__, new_new_n27258__, new_new_n27259__,
    new_new_n27260__, new_new_n27261__, new_new_n27262__, new_new_n27263__,
    new_new_n27264__, new_new_n27265__, new_new_n27266__, new_new_n27267__,
    new_new_n27268__, new_new_n27269__, new_new_n27270__, new_new_n27271__,
    new_new_n27272__, new_new_n27273__, new_new_n27274__, new_new_n27275__,
    new_new_n27276__, new_new_n27277__, new_new_n27278__, new_new_n27279__,
    new_new_n27280__, new_new_n27281__, new_new_n27282__, new_new_n27283__,
    new_new_n27284__, new_new_n27285__, new_new_n27286__, new_new_n27287__,
    new_new_n27288__, new_new_n27289__, new_new_n27290__, new_new_n27291__,
    new_new_n27292__, new_new_n27293__, new_new_n27294__, new_new_n27295__,
    new_new_n27296__, new_new_n27297__, new_new_n27298__, new_new_n27299__,
    new_new_n27300__, new_new_n27301__, new_new_n27302__, new_new_n27303__,
    new_new_n27304__, new_new_n27305__, new_new_n27306__, new_new_n27307__,
    new_new_n27308__, new_new_n27309__, new_new_n27310__, new_new_n27311__,
    new_new_n27312__, new_new_n27313__, new_new_n27314__, new_new_n27315__,
    new_new_n27316__, new_new_n27317__, new_new_n27318__, new_new_n27319__,
    new_new_n27320__, new_new_n27321__, new_new_n27322__, new_new_n27323__,
    new_new_n27324__, new_new_n27326__, new_new_n27327__, new_new_n27328__,
    new_new_n27329__, new_new_n27330__, new_new_n27331__, new_new_n27332__,
    new_new_n27333__, new_new_n27334__, new_new_n27335__, new_new_n27336__,
    new_new_n27337__, new_new_n27338__, new_new_n27339__, new_new_n27340__,
    new_new_n27341__, new_new_n27342__, new_new_n27343__, new_new_n27344__,
    new_new_n27345__, new_new_n27346__, new_new_n27347__, new_new_n27348__,
    new_new_n27349__, new_new_n27350__, new_new_n27351__, new_new_n27352__,
    new_new_n27353__, new_new_n27354__, new_new_n27355__, new_new_n27356__,
    new_new_n27357__, new_new_n27358__, new_new_n27359__, new_new_n27360__,
    new_new_n27361__, new_new_n27362__, new_new_n27363__, new_new_n27364__,
    new_new_n27365__, new_new_n27366__, new_new_n27367__, new_new_n27368__,
    new_new_n27369__, new_new_n27370__, new_new_n27371__, new_new_n27372__,
    new_new_n27373__, new_new_n27374__, new_new_n27375__, new_new_n27376__,
    new_new_n27377__, new_new_n27378__, new_new_n27379__, new_new_n27380__,
    new_new_n27381__, new_new_n27382__, new_new_n27383__, new_new_n27384__,
    new_new_n27385__, new_new_n27386__, new_new_n27387__, new_new_n27388__,
    new_new_n27389__, new_new_n27390__, new_new_n27391__, new_new_n27392__,
    new_new_n27393__, new_new_n27394__, new_new_n27395__, new_new_n27396__,
    new_new_n27397__, new_new_n27398__, new_new_n27399__, new_new_n27400__,
    new_new_n27401__, new_new_n27402__, new_new_n27403__, new_new_n27404__,
    new_new_n27405__, new_new_n27406__, new_new_n27407__, new_new_n27408__,
    new_new_n27409__, new_new_n27410__, new_new_n27411__, new_new_n27412__,
    new_new_n27414__, new_new_n27415__, new_new_n27416__, new_new_n27417__,
    new_new_n27418__, new_new_n27419__, new_new_n27420__, new_new_n27421__,
    new_new_n27422__, new_new_n27423__, new_new_n27424__, new_new_n27425__,
    new_new_n27426__, new_new_n27427__, new_new_n27428__, new_new_n27429__,
    new_new_n27430__, new_new_n27431__, new_new_n27432__, new_new_n27433__,
    new_new_n27434__, new_new_n27435__, new_new_n27436__, new_new_n27437__,
    new_new_n27438__, new_new_n27439__, new_new_n27440__, new_new_n27441__,
    new_new_n27442__, new_new_n27443__, new_new_n27444__, new_new_n27445__,
    new_new_n27446__, new_new_n27447__, new_new_n27448__, new_new_n27449__,
    new_new_n27450__, new_new_n27451__, new_new_n27452__, new_new_n27453__,
    new_new_n27454__, new_new_n27455__, new_new_n27456__, new_new_n27457__,
    new_new_n27458__, new_new_n27459__, new_new_n27460__, new_new_n27461__,
    new_new_n27462__, new_new_n27463__, new_new_n27464__, new_new_n27465__,
    new_new_n27466__, new_new_n27467__, new_new_n27468__, new_new_n27469__,
    new_new_n27470__, new_new_n27471__, new_new_n27472__, new_new_n27473__,
    new_new_n27474__, new_new_n27475__, new_new_n27476__, new_new_n27477__,
    new_new_n27478__, new_new_n27479__, new_new_n27480__, new_new_n27481__,
    new_new_n27482__, new_new_n27483__, new_new_n27484__, new_new_n27485__,
    new_new_n27486__, new_new_n27487__, new_new_n27488__, new_new_n27489__,
    new_new_n27490__, new_new_n27491__, new_new_n27492__, new_new_n27493__,
    new_new_n27494__, new_new_n27495__, new_new_n27496__, new_new_n27497__,
    new_new_n27498__, new_new_n27499__, new_new_n27500__, new_new_n27502__,
    new_new_n27503__, new_new_n27504__, new_new_n27505__, new_new_n27506__,
    new_new_n27507__, new_new_n27508__, new_new_n27509__, new_new_n27510__,
    new_new_n27511__, new_new_n27512__, new_new_n27513__, new_new_n27514__,
    new_new_n27515__, new_new_n27516__, new_new_n27517__, new_new_n27518__,
    new_new_n27519__, new_new_n27520__, new_new_n27521__, new_new_n27522__,
    new_new_n27523__, new_new_n27524__, new_new_n27525__, new_new_n27526__,
    new_new_n27527__, new_new_n27528__, new_new_n27529__, new_new_n27530__,
    new_new_n27531__, new_new_n27532__, new_new_n27533__, new_new_n27534__,
    new_new_n27535__, new_new_n27536__, new_new_n27537__, new_new_n27538__,
    new_new_n27539__, new_new_n27540__, new_new_n27541__, new_new_n27542__,
    new_new_n27543__, new_new_n27544__, new_new_n27545__, new_new_n27546__,
    new_new_n27547__, new_new_n27548__, new_new_n27549__, new_new_n27550__,
    new_new_n27551__, new_new_n27552__, new_new_n27553__, new_new_n27554__,
    new_new_n27555__, new_new_n27556__, new_new_n27557__, new_new_n27558__,
    new_new_n27559__, new_new_n27560__, new_new_n27561__, new_new_n27562__,
    new_new_n27563__, new_new_n27564__, new_new_n27565__, new_new_n27566__,
    new_new_n27567__, new_new_n27568__, new_new_n27569__, new_new_n27570__,
    new_new_n27571__, new_new_n27572__, new_new_n27573__, new_new_n27574__,
    new_new_n27575__, new_new_n27576__, new_new_n27577__, new_new_n27578__,
    new_new_n27579__, new_new_n27580__, new_new_n27581__, new_new_n27582__,
    new_new_n27583__, new_new_n27584__, new_new_n27585__, new_new_n27586__,
    new_new_n27587__, new_new_n27588__, new_new_n27590__, new_new_n27591__,
    new_new_n27592__, new_new_n27593__, new_new_n27594__, new_new_n27595__,
    new_new_n27596__, new_new_n27597__, new_new_n27598__, new_new_n27599__,
    new_new_n27600__, new_new_n27601__, new_new_n27602__, new_new_n27603__,
    new_new_n27604__, new_new_n27605__, new_new_n27606__, new_new_n27607__,
    new_new_n27608__, new_new_n27609__, new_new_n27610__, new_new_n27611__,
    new_new_n27612__, new_new_n27613__, new_new_n27614__, new_new_n27615__,
    new_new_n27616__, new_new_n27617__, new_new_n27618__, new_new_n27619__,
    new_new_n27620__, new_new_n27621__, new_new_n27622__, new_new_n27623__,
    new_new_n27624__, new_new_n27625__, new_new_n27626__, new_new_n27627__,
    new_new_n27628__, new_new_n27629__, new_new_n27630__, new_new_n27631__,
    new_new_n27632__, new_new_n27633__, new_new_n27634__, new_new_n27635__,
    new_new_n27636__, new_new_n27637__, new_new_n27638__, new_new_n27639__,
    new_new_n27640__, new_new_n27641__, new_new_n27642__, new_new_n27643__,
    new_new_n27644__, new_new_n27645__, new_new_n27646__, new_new_n27647__,
    new_new_n27648__, new_new_n27649__, new_new_n27650__, new_new_n27651__,
    new_new_n27652__, new_new_n27653__, new_new_n27654__, new_new_n27655__,
    new_new_n27656__, new_new_n27657__, new_new_n27658__, new_new_n27659__,
    new_new_n27660__, new_new_n27661__, new_new_n27662__, new_new_n27663__,
    new_new_n27664__, new_new_n27665__, new_new_n27666__, new_new_n27667__,
    new_new_n27668__, new_new_n27669__, new_new_n27670__, new_new_n27671__,
    new_new_n27672__, new_new_n27673__, new_new_n27674__, new_new_n27675__,
    new_new_n27676__, new_new_n27678__, new_new_n27679__, new_new_n27680__,
    new_new_n27681__, new_new_n27682__, new_new_n27683__, new_new_n27684__,
    new_new_n27685__, new_new_n27686__, new_new_n27687__, new_new_n27688__,
    new_new_n27689__, new_new_n27690__, new_new_n27691__, new_new_n27692__,
    new_new_n27693__, new_new_n27694__, new_new_n27695__, new_new_n27696__,
    new_new_n27697__, new_new_n27698__, new_new_n27699__, new_new_n27700__,
    new_new_n27701__, new_new_n27702__, new_new_n27703__, new_new_n27704__,
    new_new_n27705__, new_new_n27706__, new_new_n27707__, new_new_n27708__,
    new_new_n27709__, new_new_n27710__, new_new_n27711__, new_new_n27712__,
    new_new_n27713__, new_new_n27714__, new_new_n27715__, new_new_n27716__,
    new_new_n27717__, new_new_n27718__, new_new_n27719__, new_new_n27720__,
    new_new_n27721__, new_new_n27722__, new_new_n27723__, new_new_n27724__,
    new_new_n27725__, new_new_n27726__, new_new_n27727__, new_new_n27728__,
    new_new_n27729__, new_new_n27730__, new_new_n27731__, new_new_n27732__,
    new_new_n27733__, new_new_n27734__, new_new_n27735__, new_new_n27736__,
    new_new_n27737__, new_new_n27738__, new_new_n27739__, new_new_n27740__,
    new_new_n27741__, new_new_n27742__, new_new_n27743__, new_new_n27744__,
    new_new_n27745__, new_new_n27746__, new_new_n27747__, new_new_n27748__,
    new_new_n27749__, new_new_n27750__, new_new_n27751__, new_new_n27752__,
    new_new_n27753__, new_new_n27754__, new_new_n27755__, new_new_n27756__,
    new_new_n27757__, new_new_n27758__, new_new_n27759__, new_new_n27760__,
    new_new_n27761__, new_new_n27762__, new_new_n27763__, new_new_n27764__,
    new_new_n27766__, new_new_n27767__, new_new_n27768__, new_new_n27769__,
    new_new_n27770__, new_new_n27771__, new_new_n27772__, new_new_n27773__,
    new_new_n27774__, new_new_n27775__, new_new_n27776__, new_new_n27777__,
    new_new_n27778__, new_new_n27779__, new_new_n27780__, new_new_n27781__,
    new_new_n27782__, new_new_n27783__, new_new_n27784__, new_new_n27785__,
    new_new_n27786__, new_new_n27787__, new_new_n27788__, new_new_n27789__,
    new_new_n27790__, new_new_n27791__, new_new_n27792__, new_new_n27793__,
    new_new_n27794__, new_new_n27795__, new_new_n27796__, new_new_n27797__,
    new_new_n27798__, new_new_n27799__, new_new_n27800__, new_new_n27801__,
    new_new_n27802__, new_new_n27803__, new_new_n27804__, new_new_n27805__,
    new_new_n27806__, new_new_n27807__, new_new_n27808__, new_new_n27809__,
    new_new_n27810__, new_new_n27811__, new_new_n27812__, new_new_n27813__,
    new_new_n27814__, new_new_n27815__, new_new_n27816__, new_new_n27817__,
    new_new_n27818__, new_new_n27819__, new_new_n27820__, new_new_n27821__,
    new_new_n27822__, new_new_n27823__, new_new_n27824__, new_new_n27825__,
    new_new_n27826__, new_new_n27827__, new_new_n27828__, new_new_n27829__,
    new_new_n27830__, new_new_n27831__, new_new_n27832__, new_new_n27833__,
    new_new_n27834__, new_new_n27835__, new_new_n27836__, new_new_n27837__,
    new_new_n27838__, new_new_n27839__, new_new_n27840__, new_new_n27841__,
    new_new_n27842__, new_new_n27843__, new_new_n27844__, new_new_n27845__,
    new_new_n27846__, new_new_n27847__, new_new_n27848__, new_new_n27849__,
    new_new_n27850__, new_new_n27851__, new_new_n27852__, new_new_n27854__,
    new_new_n27855__, new_new_n27856__, new_new_n27857__, new_new_n27858__,
    new_new_n27859__, new_new_n27860__, new_new_n27861__, new_new_n27862__,
    new_new_n27863__, new_new_n27864__, new_new_n27865__, new_new_n27866__,
    new_new_n27867__, new_new_n27868__, new_new_n27869__, new_new_n27870__,
    new_new_n27871__, new_new_n27872__, new_new_n27873__, new_new_n27874__,
    new_new_n27875__, new_new_n27876__, new_new_n27877__, new_new_n27878__,
    new_new_n27879__, new_new_n27880__, new_new_n27881__, new_new_n27882__,
    new_new_n27883__, new_new_n27884__, new_new_n27885__, new_new_n27886__,
    new_new_n27887__, new_new_n27888__, new_new_n27889__, new_new_n27890__,
    new_new_n27891__, new_new_n27892__, new_new_n27893__, new_new_n27894__,
    new_new_n27895__, new_new_n27896__, new_new_n27897__, new_new_n27898__,
    new_new_n27899__, new_new_n27900__, new_new_n27901__, new_new_n27902__,
    new_new_n27903__, new_new_n27904__, new_new_n27905__, new_new_n27906__,
    new_new_n27907__, new_new_n27908__, new_new_n27909__, new_new_n27910__,
    new_new_n27911__, new_new_n27912__, new_new_n27913__, new_new_n27914__,
    new_new_n27915__, new_new_n27916__, new_new_n27917__, new_new_n27918__,
    new_new_n27919__, new_new_n27920__, new_new_n27921__, new_new_n27922__,
    new_new_n27923__, new_new_n27924__, new_new_n27925__, new_new_n27926__,
    new_new_n27927__, new_new_n27928__, new_new_n27929__, new_new_n27930__,
    new_new_n27931__, new_new_n27932__, new_new_n27933__, new_new_n27934__,
    new_new_n27935__, new_new_n27936__, new_new_n27937__, new_new_n27938__,
    new_new_n27939__, new_new_n27940__, new_new_n27942__, new_new_n27943__,
    new_new_n27944__, new_new_n27945__, new_new_n27946__, new_new_n27947__,
    new_new_n27948__, new_new_n27949__, new_new_n27950__, new_new_n27951__,
    new_new_n27952__, new_new_n27953__, new_new_n27954__, new_new_n27955__,
    new_new_n27956__, new_new_n27957__, new_new_n27958__, new_new_n27959__,
    new_new_n27960__, new_new_n27961__, new_new_n27962__, new_new_n27963__,
    new_new_n27964__, new_new_n27965__, new_new_n27966__, new_new_n27967__,
    new_new_n27968__, new_new_n27969__, new_new_n27970__, new_new_n27971__,
    new_new_n27972__, new_new_n27973__, new_new_n27974__, new_new_n27975__,
    new_new_n27976__, new_new_n27977__, new_new_n27978__, new_new_n27979__,
    new_new_n27980__, new_new_n27981__, new_new_n27982__, new_new_n27983__,
    new_new_n27984__, new_new_n27985__, new_new_n27986__, new_new_n27987__,
    new_new_n27988__, new_new_n27989__, new_new_n27990__, new_new_n27991__,
    new_new_n27992__, new_new_n27993__, new_new_n27994__, new_new_n27995__,
    new_new_n27996__, new_new_n27997__, new_new_n27998__, new_new_n27999__,
    new_new_n28000__, new_new_n28001__, new_new_n28002__, new_new_n28003__,
    new_new_n28004__, new_new_n28005__, new_new_n28006__, new_new_n28007__,
    new_new_n28008__, new_new_n28009__, new_new_n28010__, new_new_n28011__,
    new_new_n28012__, new_new_n28013__, new_new_n28014__, new_new_n28015__,
    new_new_n28016__, new_new_n28017__, new_new_n28018__, new_new_n28019__,
    new_new_n28020__, new_new_n28021__, new_new_n28022__, new_new_n28023__,
    new_new_n28024__, new_new_n28025__, new_new_n28026__, new_new_n28027__,
    new_new_n28028__, new_new_n28030__, new_new_n28031__, new_new_n28032__,
    new_new_n28033__, new_new_n28034__, new_new_n28035__, new_new_n28036__,
    new_new_n28037__, new_new_n28038__, new_new_n28039__, new_new_n28040__,
    new_new_n28041__, new_new_n28042__, new_new_n28043__, new_new_n28044__,
    new_new_n28045__, new_new_n28046__, new_new_n28047__, new_new_n28048__,
    new_new_n28049__, new_new_n28050__, new_new_n28051__, new_new_n28052__,
    new_new_n28053__, new_new_n28054__, new_new_n28055__, new_new_n28056__,
    new_new_n28057__, new_new_n28058__, new_new_n28059__, new_new_n28060__,
    new_new_n28061__, new_new_n28062__, new_new_n28063__, new_new_n28064__,
    new_new_n28065__, new_new_n28066__, new_new_n28067__, new_new_n28068__,
    new_new_n28069__, new_new_n28070__, new_new_n28071__, new_new_n28072__,
    new_new_n28073__, new_new_n28074__, new_new_n28075__, new_new_n28076__,
    new_new_n28077__, new_new_n28078__, new_new_n28079__, new_new_n28080__,
    new_new_n28081__, new_new_n28082__, new_new_n28083__, new_new_n28084__,
    new_new_n28085__, new_new_n28086__, new_new_n28087__, new_new_n28088__,
    new_new_n28089__, new_new_n28090__, new_new_n28091__, new_new_n28092__,
    new_new_n28093__, new_new_n28094__, new_new_n28095__, new_new_n28096__,
    new_new_n28097__, new_new_n28098__, new_new_n28099__, new_new_n28100__,
    new_new_n28101__, new_new_n28102__, new_new_n28103__, new_new_n28104__,
    new_new_n28105__, new_new_n28106__, new_new_n28107__, new_new_n28108__,
    new_new_n28109__, new_new_n28110__, new_new_n28111__, new_new_n28112__,
    new_new_n28113__, new_new_n28114__, new_new_n28115__, new_new_n28116__,
    new_new_n28118__, new_new_n28119__, new_new_n28120__, new_new_n28121__,
    new_new_n28122__, new_new_n28123__, new_new_n28124__, new_new_n28125__,
    new_new_n28126__, new_new_n28127__, new_new_n28128__, new_new_n28129__,
    new_new_n28130__, new_new_n28131__, new_new_n28132__, new_new_n28133__,
    new_new_n28134__, new_new_n28135__, new_new_n28136__, new_new_n28137__,
    new_new_n28138__, new_new_n28139__, new_new_n28140__, new_new_n28141__,
    new_new_n28142__, new_new_n28143__, new_new_n28144__, new_new_n28145__,
    new_new_n28146__, new_new_n28147__, new_new_n28148__, new_new_n28149__,
    new_new_n28150__, new_new_n28151__, new_new_n28152__, new_new_n28153__,
    new_new_n28154__, new_new_n28155__, new_new_n28156__, new_new_n28157__,
    new_new_n28158__, new_new_n28159__, new_new_n28160__, new_new_n28161__,
    new_new_n28162__, new_new_n28163__, new_new_n28164__, new_new_n28165__,
    new_new_n28166__, new_new_n28167__, new_new_n28168__, new_new_n28169__,
    new_new_n28170__, new_new_n28171__, new_new_n28172__, new_new_n28173__,
    new_new_n28174__, new_new_n28175__, new_new_n28176__, new_new_n28177__,
    new_new_n28178__, new_new_n28179__, new_new_n28180__, new_new_n28181__,
    new_new_n28182__, new_new_n28183__, new_new_n28184__, new_new_n28185__,
    new_new_n28186__, new_new_n28187__, new_new_n28188__, new_new_n28189__,
    new_new_n28190__, new_new_n28191__, new_new_n28192__, new_new_n28193__,
    new_new_n28194__, new_new_n28195__, new_new_n28196__, new_new_n28197__,
    new_new_n28198__, new_new_n28199__, new_new_n28200__, new_new_n28201__,
    new_new_n28202__, new_new_n28203__, new_new_n28204__, new_new_n28206__,
    new_new_n28207__, new_new_n28208__, new_new_n28209__, new_new_n28210__,
    new_new_n28211__, new_new_n28212__, new_new_n28213__, new_new_n28214__,
    new_new_n28215__, new_new_n28216__, new_new_n28217__, new_new_n28218__,
    new_new_n28219__, new_new_n28220__, new_new_n28221__, new_new_n28222__,
    new_new_n28223__, new_new_n28224__, new_new_n28225__, new_new_n28226__,
    new_new_n28227__, new_new_n28228__, new_new_n28229__, new_new_n28230__,
    new_new_n28231__, new_new_n28232__, new_new_n28233__, new_new_n28234__,
    new_new_n28235__, new_new_n28236__, new_new_n28237__, new_new_n28238__,
    new_new_n28239__, new_new_n28240__, new_new_n28241__, new_new_n28242__,
    new_new_n28243__, new_new_n28244__, new_new_n28245__, new_new_n28246__,
    new_new_n28247__, new_new_n28248__, new_new_n28249__, new_new_n28250__,
    new_new_n28251__, new_new_n28252__, new_new_n28253__, new_new_n28254__,
    new_new_n28255__, new_new_n28256__, new_new_n28257__, new_new_n28258__,
    new_new_n28259__, new_new_n28260__, new_new_n28261__, new_new_n28262__,
    new_new_n28263__, new_new_n28264__, new_new_n28265__, new_new_n28266__,
    new_new_n28267__, new_new_n28268__, new_new_n28269__, new_new_n28270__,
    new_new_n28271__, new_new_n28272__, new_new_n28273__, new_new_n28274__,
    new_new_n28275__, new_new_n28276__, new_new_n28277__, new_new_n28278__,
    new_new_n28279__, new_new_n28280__, new_new_n28281__, new_new_n28282__,
    new_new_n28283__, new_new_n28284__, new_new_n28285__, new_new_n28286__,
    new_new_n28287__, new_new_n28288__, new_new_n28289__, new_new_n28290__,
    new_new_n28291__, new_new_n28292__, new_new_n28294__, new_new_n28295__,
    new_new_n28296__, new_new_n28297__, new_new_n28298__, new_new_n28299__,
    new_new_n28300__, new_new_n28301__, new_new_n28302__, new_new_n28303__,
    new_new_n28304__, new_new_n28305__, new_new_n28306__, new_new_n28307__,
    new_new_n28308__, new_new_n28309__, new_new_n28310__, new_new_n28311__,
    new_new_n28312__, new_new_n28313__, new_new_n28314__, new_new_n28315__,
    new_new_n28316__, new_new_n28317__, new_new_n28318__, new_new_n28319__,
    new_new_n28320__, new_new_n28321__, new_new_n28322__, new_new_n28323__,
    new_new_n28324__, new_new_n28325__, new_new_n28326__, new_new_n28327__,
    new_new_n28328__, new_new_n28329__, new_new_n28330__, new_new_n28331__,
    new_new_n28332__, new_new_n28333__, new_new_n28334__, new_new_n28335__,
    new_new_n28336__, new_new_n28337__, new_new_n28338__, new_new_n28339__,
    new_new_n28340__, new_new_n28341__, new_new_n28342__, new_new_n28343__,
    new_new_n28344__, new_new_n28345__, new_new_n28346__, new_new_n28347__,
    new_new_n28348__, new_new_n28349__, new_new_n28350__, new_new_n28351__,
    new_new_n28352__, new_new_n28353__, new_new_n28354__, new_new_n28355__,
    new_new_n28356__, new_new_n28357__, new_new_n28358__, new_new_n28359__,
    new_new_n28360__, new_new_n28361__, new_new_n28362__, new_new_n28363__,
    new_new_n28364__, new_new_n28365__, new_new_n28366__, new_new_n28367__,
    new_new_n28368__, new_new_n28369__, new_new_n28370__, new_new_n28371__,
    new_new_n28372__, new_new_n28373__, new_new_n28374__, new_new_n28375__,
    new_new_n28376__, new_new_n28377__, new_new_n28378__, new_new_n28379__,
    new_new_n28380__, new_new_n28382__, new_new_n28383__, new_new_n28384__,
    new_new_n28385__, new_new_n28386__, new_new_n28387__, new_new_n28388__,
    new_new_n28389__, new_new_n28390__, new_new_n28391__, new_new_n28392__,
    new_new_n28393__, new_new_n28394__, new_new_n28395__, new_new_n28396__,
    new_new_n28397__, new_new_n28398__, new_new_n28399__, new_new_n28400__,
    new_new_n28401__, new_new_n28402__, new_new_n28403__, new_new_n28404__,
    new_new_n28405__, new_new_n28406__, new_new_n28407__, new_new_n28408__,
    new_new_n28409__, new_new_n28410__, new_new_n28411__, new_new_n28412__,
    new_new_n28413__, new_new_n28414__, new_new_n28415__, new_new_n28416__,
    new_new_n28417__, new_new_n28418__, new_new_n28419__, new_new_n28420__,
    new_new_n28421__, new_new_n28422__, new_new_n28423__, new_new_n28424__,
    new_new_n28425__, new_new_n28426__, new_new_n28427__, new_new_n28428__,
    new_new_n28429__, new_new_n28430__, new_new_n28431__, new_new_n28432__,
    new_new_n28433__, new_new_n28434__, new_new_n28435__, new_new_n28436__,
    new_new_n28437__, new_new_n28438__, new_new_n28439__, new_new_n28440__,
    new_new_n28441__, new_new_n28442__, new_new_n28443__, new_new_n28444__,
    new_new_n28445__, new_new_n28446__, new_new_n28447__, new_new_n28448__,
    new_new_n28449__, new_new_n28450__, new_new_n28451__, new_new_n28452__,
    new_new_n28453__, new_new_n28454__, new_new_n28455__, new_new_n28456__,
    new_new_n28457__, new_new_n28458__, new_new_n28459__, new_new_n28460__,
    new_new_n28461__, new_new_n28462__, new_new_n28463__, new_new_n28464__,
    new_new_n28465__, new_new_n28466__, new_new_n28467__, new_new_n28468__,
    new_new_n28470__, new_new_n28471__, new_new_n28472__, new_new_n28473__,
    new_new_n28474__, new_new_n28475__, new_new_n28476__, new_new_n28477__,
    new_new_n28478__, new_new_n28479__, new_new_n28480__, new_new_n28481__,
    new_new_n28482__, new_new_n28483__, new_new_n28484__, new_new_n28485__,
    new_new_n28486__, new_new_n28487__, new_new_n28488__, new_new_n28489__,
    new_new_n28490__, new_new_n28491__, new_new_n28492__, new_new_n28493__,
    new_new_n28494__, new_new_n28495__, new_new_n28496__, new_new_n28497__,
    new_new_n28498__, new_new_n28499__, new_new_n28500__, new_new_n28501__,
    new_new_n28502__, new_new_n28503__, new_new_n28504__, new_new_n28505__,
    new_new_n28506__, new_new_n28507__, new_new_n28508__, new_new_n28509__,
    new_new_n28510__, new_new_n28511__, new_new_n28512__, new_new_n28513__,
    new_new_n28514__, new_new_n28515__, new_new_n28516__, new_new_n28517__,
    new_new_n28518__, new_new_n28519__, new_new_n28520__, new_new_n28521__,
    new_new_n28522__, new_new_n28523__, new_new_n28524__, new_new_n28525__,
    new_new_n28526__, new_new_n28527__, new_new_n28528__, new_new_n28529__,
    new_new_n28530__, new_new_n28531__, new_new_n28532__, new_new_n28533__,
    new_new_n28534__, new_new_n28535__, new_new_n28536__, new_new_n28537__,
    new_new_n28538__, new_new_n28539__, new_new_n28540__, new_new_n28541__,
    new_new_n28542__, new_new_n28543__, new_new_n28544__, new_new_n28545__,
    new_new_n28546__, new_new_n28547__, new_new_n28548__, new_new_n28549__,
    new_new_n28550__, new_new_n28551__, new_new_n28552__, new_new_n28553__,
    new_new_n28554__, new_new_n28555__, new_new_n28556__, new_new_n28557__,
    new_new_n28558__, new_new_n28559__, new_new_n28560__, new_new_n28561__,
    new_new_n28563__, new_new_n28564__, new_new_n28565__, new_new_n28566__,
    new_new_n28567__, new_new_n28568__, new_new_n28569__, new_new_n28570__,
    new_new_n28571__, new_new_n28572__, new_new_n28573__, new_new_n28574__,
    new_new_n28575__, new_new_n28576__, new_new_n28577__, new_new_n28578__,
    new_new_n28579__, new_new_n28580__, new_new_n28581__, new_new_n28582__,
    new_new_n28583__, new_new_n28584__, new_new_n28585__, new_new_n28586__,
    new_new_n28587__, new_new_n28588__, new_new_n28589__, new_new_n28590__,
    new_new_n28591__, new_new_n28592__, new_new_n28593__, new_new_n28594__,
    new_new_n28595__, new_new_n28596__, new_new_n28597__, new_new_n28598__,
    new_new_n28599__, new_new_n28600__, new_new_n28601__, new_new_n28602__,
    new_new_n28603__, new_new_n28604__, new_new_n28605__, new_new_n28606__,
    new_new_n28607__, new_new_n28608__, new_new_n28609__, new_new_n28610__,
    new_new_n28611__, new_new_n28612__, new_new_n28613__, new_new_n28614__,
    new_new_n28615__, new_new_n28616__, new_new_n28617__, new_new_n28618__,
    new_new_n28619__, new_new_n28620__, new_new_n28621__, new_new_n28622__,
    new_new_n28623__, new_new_n28624__, new_new_n28625__, new_new_n28626__,
    new_new_n28627__, new_new_n28628__, new_new_n28629__, new_new_n28630__,
    new_new_n28631__, new_new_n28632__, new_new_n28633__, new_new_n28634__,
    new_new_n28635__, new_new_n28636__, new_new_n28637__, new_new_n28638__,
    new_new_n28639__, new_new_n28640__, new_new_n28641__, new_new_n28642__,
    new_new_n28643__, new_new_n28644__, new_new_n28645__, new_new_n28646__,
    new_new_n28647__, new_new_n28648__, new_new_n28649__, new_new_n28651__,
    new_new_n28652__, new_new_n28653__, new_new_n28654__, new_new_n28655__,
    new_new_n28656__, new_new_n28657__, new_new_n28658__, new_new_n28659__,
    new_new_n28660__, new_new_n28661__, new_new_n28662__, new_new_n28663__,
    new_new_n28664__, new_new_n28665__, new_new_n28666__, new_new_n28667__,
    new_new_n28668__, new_new_n28669__, new_new_n28670__, new_new_n28671__,
    new_new_n28672__, new_new_n28673__, new_new_n28674__, new_new_n28675__,
    new_new_n28676__, new_new_n28677__, new_new_n28678__, new_new_n28679__,
    new_new_n28680__, new_new_n28681__, new_new_n28682__, new_new_n28683__,
    new_new_n28684__, new_new_n28685__, new_new_n28686__, new_new_n28687__,
    new_new_n28688__, new_new_n28689__, new_new_n28690__, new_new_n28691__,
    new_new_n28692__, new_new_n28693__, new_new_n28694__, new_new_n28695__,
    new_new_n28696__, new_new_n28697__, new_new_n28698__, new_new_n28699__,
    new_new_n28700__, new_new_n28701__, new_new_n28702__, new_new_n28703__,
    new_new_n28704__, new_new_n28705__, new_new_n28706__, new_new_n28707__,
    new_new_n28708__, new_new_n28709__, new_new_n28710__, new_new_n28711__,
    new_new_n28712__, new_new_n28713__, new_new_n28714__, new_new_n28715__,
    new_new_n28716__, new_new_n28717__, new_new_n28718__, new_new_n28719__,
    new_new_n28720__, new_new_n28721__, new_new_n28722__, new_new_n28723__,
    new_new_n28724__, new_new_n28725__, new_new_n28726__, new_new_n28727__,
    new_new_n28728__, new_new_n28729__, new_new_n28730__, new_new_n28731__,
    new_new_n28732__, new_new_n28733__, new_new_n28734__, new_new_n28735__,
    new_new_n28736__, new_new_n28737__, new_new_n28739__, new_new_n28740__,
    new_new_n28741__, new_new_n28742__, new_new_n28743__, new_new_n28744__,
    new_new_n28745__, new_new_n28746__, new_new_n28747__, new_new_n28748__,
    new_new_n28749__, new_new_n28750__, new_new_n28751__, new_new_n28752__,
    new_new_n28753__, new_new_n28754__, new_new_n28755__, new_new_n28756__,
    new_new_n28757__, new_new_n28758__, new_new_n28759__, new_new_n28760__,
    new_new_n28761__, new_new_n28762__, new_new_n28763__, new_new_n28764__,
    new_new_n28765__, new_new_n28766__, new_new_n28767__, new_new_n28768__,
    new_new_n28769__, new_new_n28770__, new_new_n28771__, new_new_n28772__,
    new_new_n28773__, new_new_n28774__, new_new_n28775__, new_new_n28776__,
    new_new_n28777__, new_new_n28778__, new_new_n28779__, new_new_n28780__,
    new_new_n28781__, new_new_n28782__, new_new_n28783__, new_new_n28784__,
    new_new_n28785__, new_new_n28786__, new_new_n28787__, new_new_n28788__,
    new_new_n28789__, new_new_n28790__, new_new_n28791__, new_new_n28792__,
    new_new_n28793__, new_new_n28794__, new_new_n28795__, new_new_n28796__,
    new_new_n28797__, new_new_n28798__, new_new_n28799__, new_new_n28800__,
    new_new_n28801__, new_new_n28802__, new_new_n28803__, new_new_n28804__,
    new_new_n28805__, new_new_n28806__, new_new_n28807__, new_new_n28808__,
    new_new_n28809__, new_new_n28810__, new_new_n28811__, new_new_n28812__,
    new_new_n28813__, new_new_n28814__, new_new_n28815__, new_new_n28816__,
    new_new_n28817__, new_new_n28818__, new_new_n28819__, new_new_n28820__,
    new_new_n28821__, new_new_n28822__, new_new_n28823__, new_new_n28824__,
    new_new_n28825__, new_new_n28827__, new_new_n28828__, new_new_n28829__,
    new_new_n28830__, new_new_n28831__, new_new_n28832__, new_new_n28833__,
    new_new_n28834__, new_new_n28835__, new_new_n28836__, new_new_n28837__,
    new_new_n28838__, new_new_n28839__, new_new_n28840__, new_new_n28841__,
    new_new_n28842__, new_new_n28843__, new_new_n28844__, new_new_n28845__,
    new_new_n28846__, new_new_n28847__, new_new_n28848__, new_new_n28849__,
    new_new_n28850__, new_new_n28851__, new_new_n28852__, new_new_n28853__,
    new_new_n28854__, new_new_n28855__, new_new_n28856__, new_new_n28857__,
    new_new_n28858__, new_new_n28859__, new_new_n28860__, new_new_n28861__,
    new_new_n28862__, new_new_n28863__, new_new_n28864__, new_new_n28865__,
    new_new_n28866__, new_new_n28867__, new_new_n28868__, new_new_n28869__,
    new_new_n28870__, new_new_n28871__, new_new_n28872__, new_new_n28873__,
    new_new_n28874__, new_new_n28875__, new_new_n28876__, new_new_n28877__,
    new_new_n28878__, new_new_n28879__, new_new_n28880__, new_new_n28881__,
    new_new_n28882__, new_new_n28883__, new_new_n28884__, new_new_n28885__,
    new_new_n28886__, new_new_n28887__, new_new_n28888__, new_new_n28889__,
    new_new_n28890__, new_new_n28891__, new_new_n28892__, new_new_n28893__,
    new_new_n28894__, new_new_n28895__, new_new_n28896__, new_new_n28897__,
    new_new_n28898__, new_new_n28899__, new_new_n28900__, new_new_n28901__,
    new_new_n28903__, new_new_n28904__, new_new_n28905__, new_new_n28906__,
    new_new_n28907__, new_new_n28908__, new_new_n28909__, new_new_n28910__,
    new_new_n28911__, new_new_n28912__, new_new_n28913__, new_new_n28914__,
    new_new_n28915__, new_new_n28916__, new_new_n28917__, new_new_n28918__,
    new_new_n28919__, new_new_n28920__, new_new_n28921__, new_new_n28922__,
    new_new_n28923__, new_new_n28924__, new_new_n28925__, new_new_n28926__,
    new_new_n28927__, new_new_n28928__, new_new_n28929__, new_new_n28930__,
    new_new_n28931__, new_new_n28932__, new_new_n28933__, new_new_n28934__,
    new_new_n28935__, new_new_n28936__, new_new_n28937__, new_new_n28938__,
    new_new_n28939__, new_new_n28940__, new_new_n28941__, new_new_n28942__,
    new_new_n28943__, new_new_n28944__, new_new_n28945__, new_new_n28946__,
    new_new_n28947__, new_new_n28948__, new_new_n28949__, new_new_n28950__,
    new_new_n28951__, new_new_n28952__, new_new_n28953__, new_new_n28954__,
    new_new_n28955__, new_new_n28956__, new_new_n28957__, new_new_n28958__,
    new_new_n28959__, new_new_n28960__, new_new_n28961__, new_new_n28962__,
    new_new_n28963__, new_new_n28964__, new_new_n28965__, new_new_n28966__,
    new_new_n28967__, new_new_n28968__, new_new_n28969__, new_new_n28970__,
    new_new_n28971__, new_new_n28972__, new_new_n28973__, new_new_n28974__,
    new_new_n28975__, new_new_n28976__, new_new_n28977__, new_new_n28978__,
    new_new_n28979__, new_new_n28980__, new_new_n28981__, new_new_n28982__,
    new_new_n28983__, new_new_n28984__, new_new_n28985__, new_new_n28987__,
    new_new_n28988__, new_new_n28989__, new_new_n28990__, new_new_n28991__,
    new_new_n28992__, new_new_n28993__, new_new_n28994__, new_new_n28995__,
    new_new_n28996__, new_new_n28997__, new_new_n28998__, new_new_n28999__,
    new_new_n29000__, new_new_n29001__, new_new_n29002__, new_new_n29003__,
    new_new_n29004__, new_new_n29005__, new_new_n29006__, new_new_n29007__,
    new_new_n29008__, new_new_n29009__, new_new_n29010__, new_new_n29011__,
    new_new_n29012__, new_new_n29013__, new_new_n29014__, new_new_n29015__,
    new_new_n29016__, new_new_n29017__, new_new_n29018__, new_new_n29019__,
    new_new_n29020__, new_new_n29021__, new_new_n29022__, new_new_n29023__,
    new_new_n29024__, new_new_n29025__, new_new_n29026__, new_new_n29027__,
    new_new_n29028__, new_new_n29029__, new_new_n29030__, new_new_n29031__,
    new_new_n29032__, new_new_n29033__, new_new_n29034__, new_new_n29035__,
    new_new_n29036__, new_new_n29037__, new_new_n29038__, new_new_n29039__,
    new_new_n29040__, new_new_n29041__, new_new_n29042__, new_new_n29043__,
    new_new_n29044__, new_new_n29045__, new_new_n29046__, new_new_n29047__,
    new_new_n29048__, new_new_n29049__, new_new_n29050__, new_new_n29051__,
    new_new_n29052__, new_new_n29053__, new_new_n29054__, new_new_n29055__,
    new_new_n29056__, new_new_n29057__, new_new_n29058__, new_new_n29059__,
    new_new_n29060__, new_new_n29061__, new_new_n29062__, new_new_n29063__,
    new_new_n29064__, new_new_n29065__, new_new_n29066__, new_new_n29067__,
    new_new_n29068__, new_new_n29069__, new_new_n29070__, new_new_n29071__,
    new_new_n29072__, new_new_n29073__, new_new_n29074__, new_new_n29075__,
    new_new_n29076__, new_new_n29077__, new_new_n29078__, new_new_n29079__,
    new_new_n29080__, new_new_n29081__, new_new_n29082__, new_new_n29083__,
    new_new_n29084__, new_new_n29085__, new_new_n29086__, new_new_n29087__,
    new_new_n29088__, new_new_n29089__, new_new_n29090__, new_new_n29091__,
    new_new_n29092__, new_new_n29093__, new_new_n29094__, new_new_n29095__,
    new_new_n29096__, new_new_n29097__, new_new_n29098__, new_new_n29099__,
    new_new_n29100__, new_new_n29101__, new_new_n29102__, new_new_n29103__,
    new_new_n29104__, new_new_n29105__, new_new_n29107__, new_new_n29108__,
    new_new_n29109__, new_new_n29110__, new_new_n29111__, new_new_n29112__,
    new_new_n29113__, new_new_n29114__, new_new_n29115__, new_new_n29116__,
    new_new_n29117__, new_new_n29118__, new_new_n29119__, new_new_n29120__,
    new_new_n29121__, new_new_n29122__, new_new_n29123__, new_new_n29124__,
    new_new_n29125__, new_new_n29126__, new_new_n29127__, new_new_n29128__,
    new_new_n29129__, new_new_n29130__, new_new_n29131__, new_new_n29132__,
    new_new_n29133__, new_new_n29134__, new_new_n29135__, new_new_n29136__,
    new_new_n29137__, new_new_n29138__, new_new_n29139__, new_new_n29140__,
    new_new_n29141__, new_new_n29142__, new_new_n29143__, new_new_n29144__,
    new_new_n29145__, new_new_n29146__, new_new_n29147__, new_new_n29148__,
    new_new_n29149__, new_new_n29150__, new_new_n29151__, new_new_n29152__,
    new_new_n29153__, new_new_n29154__, new_new_n29155__, new_new_n29156__,
    new_new_n29157__, new_new_n29158__, new_new_n29159__, new_new_n29160__,
    new_new_n29161__, new_new_n29162__, new_new_n29163__, new_new_n29164__,
    new_new_n29165__, new_new_n29166__, new_new_n29167__, new_new_n29168__,
    new_new_n29169__, new_new_n29170__, new_new_n29171__, new_new_n29172__,
    new_new_n29173__, new_new_n29174__, new_new_n29175__, new_new_n29176__,
    new_new_n29177__, new_new_n29178__, new_new_n29179__, new_new_n29180__,
    new_new_n29181__, new_new_n29182__, new_new_n29183__, new_new_n29184__,
    new_new_n29185__, new_new_n29186__, new_new_n29187__, new_new_n29188__,
    new_new_n29189__, new_new_n29190__, new_new_n29191__, new_new_n29192__,
    new_new_n29193__, new_new_n29194__, new_new_n29195__, new_new_n29196__,
    new_new_n29197__, new_new_n29198__, new_new_n29199__, new_new_n29200__,
    new_new_n29201__, new_new_n29202__, new_new_n29203__, new_new_n29204__,
    new_new_n29206__, new_new_n29207__, new_new_n29208__, new_new_n29209__,
    new_new_n29210__, new_new_n29211__, new_new_n29212__, new_new_n29213__,
    new_new_n29214__, new_new_n29215__, new_new_n29216__, new_new_n29217__,
    new_new_n29218__, new_new_n29219__, new_new_n29220__, new_new_n29221__,
    new_new_n29222__, new_new_n29223__, new_new_n29224__, new_new_n29225__,
    new_new_n29226__, new_new_n29227__, new_new_n29228__, new_new_n29229__,
    new_new_n29230__, new_new_n29231__, new_new_n29232__, new_new_n29233__,
    new_new_n29234__, new_new_n29235__, new_new_n29236__, new_new_n29237__,
    new_new_n29238__, new_new_n29239__, new_new_n29240__, new_new_n29241__,
    new_new_n29242__, new_new_n29243__, new_new_n29244__, new_new_n29245__,
    new_new_n29246__, new_new_n29247__, new_new_n29248__, new_new_n29249__,
    new_new_n29250__, new_new_n29251__, new_new_n29252__, new_new_n29253__,
    new_new_n29254__, new_new_n29255__, new_new_n29256__, new_new_n29257__,
    new_new_n29258__, new_new_n29259__, new_new_n29260__, new_new_n29261__,
    new_new_n29262__, new_new_n29263__, new_new_n29264__, new_new_n29265__,
    new_new_n29266__, new_new_n29267__, new_new_n29268__, new_new_n29269__,
    new_new_n29270__, new_new_n29271__, new_new_n29272__, new_new_n29273__,
    new_new_n29274__, new_new_n29275__, new_new_n29276__, new_new_n29277__,
    new_new_n29278__, new_new_n29279__, new_new_n29280__, new_new_n29281__,
    new_new_n29282__, new_new_n29283__, new_new_n29284__, new_new_n29285__,
    new_new_n29286__, new_new_n29287__, new_new_n29288__, new_new_n29289__,
    new_new_n29290__, new_new_n29291__, new_new_n29292__, new_new_n29293__,
    new_new_n29294__, new_new_n29295__, new_new_n29296__, new_new_n29297__,
    new_new_n29298__, new_new_n29299__, new_new_n29300__, new_new_n29301__,
    new_new_n29302__, new_new_n29303__, new_new_n29304__, new_new_n29306__,
    new_new_n29307__, new_new_n29308__, new_new_n29309__, new_new_n29310__,
    new_new_n29311__, new_new_n29312__, new_new_n29313__, new_new_n29314__,
    new_new_n29315__, new_new_n29316__, new_new_n29317__, new_new_n29318__,
    new_new_n29319__, new_new_n29320__, new_new_n29321__, new_new_n29322__,
    new_new_n29323__, new_new_n29324__, new_new_n29325__, new_new_n29326__,
    new_new_n29327__, new_new_n29328__, new_new_n29329__, new_new_n29330__,
    new_new_n29331__, new_new_n29332__, new_new_n29333__, new_new_n29334__,
    new_new_n29335__, new_new_n29336__, new_new_n29337__, new_new_n29338__,
    new_new_n29339__, new_new_n29340__, new_new_n29341__, new_new_n29342__,
    new_new_n29343__, new_new_n29344__, new_new_n29345__, new_new_n29346__,
    new_new_n29347__, new_new_n29348__, new_new_n29349__, new_new_n29350__,
    new_new_n29351__, new_new_n29352__, new_new_n29353__, new_new_n29354__,
    new_new_n29355__, new_new_n29356__, new_new_n29357__, new_new_n29358__,
    new_new_n29359__, new_new_n29360__, new_new_n29361__, new_new_n29362__,
    new_new_n29363__, new_new_n29364__, new_new_n29365__, new_new_n29366__,
    new_new_n29367__, new_new_n29368__, new_new_n29369__, new_new_n29370__,
    new_new_n29371__, new_new_n29372__, new_new_n29373__, new_new_n29374__,
    new_new_n29375__, new_new_n29376__, new_new_n29377__, new_new_n29378__,
    new_new_n29379__, new_new_n29380__, new_new_n29381__, new_new_n29382__,
    new_new_n29383__, new_new_n29384__, new_new_n29385__, new_new_n29386__,
    new_new_n29387__, new_new_n29388__, new_new_n29389__, new_new_n29390__,
    new_new_n29391__, new_new_n29392__, new_new_n29393__, new_new_n29394__,
    new_new_n29395__, new_new_n29396__, new_new_n29397__, new_new_n29398__,
    new_new_n29399__, new_new_n29400__, new_new_n29401__, new_new_n29402__,
    new_new_n29403__, new_new_n29404__, new_new_n29406__, new_new_n29407__,
    new_new_n29408__, new_new_n29409__, new_new_n29410__, new_new_n29411__,
    new_new_n29412__, new_new_n29413__, new_new_n29414__, new_new_n29415__,
    new_new_n29416__, new_new_n29417__, new_new_n29418__, new_new_n29419__,
    new_new_n29420__, new_new_n29421__, new_new_n29422__, new_new_n29423__,
    new_new_n29424__, new_new_n29425__, new_new_n29426__, new_new_n29427__,
    new_new_n29428__, new_new_n29429__, new_new_n29430__, new_new_n29431__,
    new_new_n29432__, new_new_n29433__, new_new_n29434__, new_new_n29435__,
    new_new_n29436__, new_new_n29437__, new_new_n29438__, new_new_n29439__,
    new_new_n29440__, new_new_n29441__, new_new_n29442__, new_new_n29443__,
    new_new_n29444__, new_new_n29445__, new_new_n29446__, new_new_n29447__,
    new_new_n29448__, new_new_n29449__, new_new_n29450__, new_new_n29451__,
    new_new_n29452__, new_new_n29453__, new_new_n29454__, new_new_n29455__,
    new_new_n29456__, new_new_n29457__, new_new_n29458__, new_new_n29459__,
    new_new_n29460__, new_new_n29461__, new_new_n29462__, new_new_n29463__,
    new_new_n29464__, new_new_n29465__, new_new_n29466__, new_new_n29467__,
    new_new_n29468__, new_new_n29469__, new_new_n29470__, new_new_n29471__,
    new_new_n29472__, new_new_n29473__, new_new_n29474__, new_new_n29475__,
    new_new_n29476__, new_new_n29477__, new_new_n29478__, new_new_n29479__,
    new_new_n29480__, new_new_n29481__, new_new_n29482__, new_new_n29483__,
    new_new_n29484__, new_new_n29485__, new_new_n29486__, new_new_n29487__,
    new_new_n29488__, new_new_n29489__, new_new_n29490__, new_new_n29491__,
    new_new_n29492__, new_new_n29493__, new_new_n29494__, new_new_n29495__,
    new_new_n29496__, new_new_n29497__, new_new_n29498__, new_new_n29499__,
    new_new_n29500__, new_new_n29501__, new_new_n29502__, new_new_n29503__,
    new_new_n29504__, new_new_n29506__, new_new_n29507__, new_new_n29508__,
    new_new_n29509__, new_new_n29510__, new_new_n29511__, new_new_n29512__,
    new_new_n29513__, new_new_n29514__, new_new_n29515__, new_new_n29516__,
    new_new_n29517__, new_new_n29518__, new_new_n29519__, new_new_n29520__,
    new_new_n29521__, new_new_n29522__, new_new_n29523__, new_new_n29524__,
    new_new_n29525__, new_new_n29526__, new_new_n29527__, new_new_n29528__,
    new_new_n29529__, new_new_n29530__, new_new_n29531__, new_new_n29532__,
    new_new_n29533__, new_new_n29534__, new_new_n29535__, new_new_n29536__,
    new_new_n29537__, new_new_n29538__, new_new_n29539__, new_new_n29540__,
    new_new_n29541__, new_new_n29542__, new_new_n29543__, new_new_n29544__,
    new_new_n29545__, new_new_n29546__, new_new_n29547__, new_new_n29548__,
    new_new_n29549__, new_new_n29550__, new_new_n29551__, new_new_n29552__,
    new_new_n29553__, new_new_n29554__, new_new_n29555__, new_new_n29556__,
    new_new_n29557__, new_new_n29558__, new_new_n29559__, new_new_n29560__,
    new_new_n29561__, new_new_n29562__, new_new_n29563__, new_new_n29564__,
    new_new_n29565__, new_new_n29566__, new_new_n29567__, new_new_n29568__,
    new_new_n29569__, new_new_n29570__, new_new_n29571__, new_new_n29572__,
    new_new_n29573__, new_new_n29574__, new_new_n29575__, new_new_n29576__,
    new_new_n29577__, new_new_n29578__, new_new_n29579__, new_new_n29580__,
    new_new_n29581__, new_new_n29582__, new_new_n29583__, new_new_n29584__,
    new_new_n29585__, new_new_n29586__, new_new_n29587__, new_new_n29588__,
    new_new_n29589__, new_new_n29590__, new_new_n29591__, new_new_n29592__,
    new_new_n29593__, new_new_n29594__, new_new_n29595__, new_new_n29597__,
    new_new_n29598__, new_new_n29599__, new_new_n29600__, new_new_n29601__,
    new_new_n29602__, new_new_n29603__, new_new_n29604__, new_new_n29605__,
    new_new_n29606__, new_new_n29607__, new_new_n29608__, new_new_n29609__,
    new_new_n29610__, new_new_n29611__, new_new_n29612__, new_new_n29613__,
    new_new_n29614__, new_new_n29615__, new_new_n29616__, new_new_n29617__,
    new_new_n29618__, new_new_n29619__, new_new_n29620__, new_new_n29621__,
    new_new_n29622__, new_new_n29623__, new_new_n29624__, new_new_n29625__,
    new_new_n29626__, new_new_n29627__, new_new_n29628__, new_new_n29629__,
    new_new_n29630__, new_new_n29631__, new_new_n29632__, new_new_n29633__,
    new_new_n29634__, new_new_n29635__, new_new_n29636__, new_new_n29637__,
    new_new_n29638__, new_new_n29639__, new_new_n29640__, new_new_n29641__,
    new_new_n29642__, new_new_n29643__, new_new_n29644__, new_new_n29645__,
    new_new_n29646__, new_new_n29647__, new_new_n29648__, new_new_n29649__,
    new_new_n29650__, new_new_n29651__, new_new_n29652__, new_new_n29653__,
    new_new_n29654__, new_new_n29655__, new_new_n29656__, new_new_n29657__,
    new_new_n29658__, new_new_n29659__, new_new_n29660__, new_new_n29661__,
    new_new_n29662__, new_new_n29663__, new_new_n29664__, new_new_n29665__,
    new_new_n29666__, new_new_n29667__, new_new_n29668__, new_new_n29669__,
    new_new_n29670__, new_new_n29671__, new_new_n29672__, new_new_n29673__,
    new_new_n29674__, new_new_n29675__, new_new_n29676__, new_new_n29677__,
    new_new_n29678__, new_new_n29679__, new_new_n29680__, new_new_n29681__,
    new_new_n29682__, new_new_n29683__, new_new_n29684__, new_new_n29685__,
    new_new_n29686__, new_new_n29688__, new_new_n29689__, new_new_n29690__,
    new_new_n29691__, new_new_n29692__, new_new_n29693__, new_new_n29695__,
    new_new_n29696__, new_new_n29697__, new_new_n29698__, new_new_n29699__,
    new_new_n29700__, new_new_n29701__, new_new_n29702__, new_new_n29704__,
    new_new_n29705__, new_new_n29706__, new_new_n29707__, new_new_n29708__,
    new_new_n29709__, new_new_n29710__, new_new_n29711__, new_new_n29712__,
    new_new_n29714__, new_new_n29715__, new_new_n29716__, new_new_n29717__,
    new_new_n29718__, new_new_n29719__, new_new_n29720__, new_new_n29721__,
    new_new_n29722__, new_new_n29724__, new_new_n29725__, new_new_n29726__,
    new_new_n29727__, new_new_n29728__, new_new_n29729__, new_new_n29730__,
    new_new_n29731__, new_new_n29732__, new_new_n29733__, new_new_n29735__,
    new_new_n29736__, new_new_n29737__, new_new_n29738__, new_new_n29739__,
    new_new_n29740__, new_new_n29741__, new_new_n29742__, new_new_n29743__,
    new_new_n29745__, new_new_n29746__, new_new_n29747__, new_new_n29748__,
    new_new_n29749__, new_new_n29750__, new_new_n29751__, new_new_n29752__,
    new_new_n29753__, new_new_n29754__, new_new_n29755__, new_new_n29757__,
    new_new_n29758__, new_new_n29759__, new_new_n29760__, new_new_n29761__,
    new_new_n29762__, new_new_n29763__, new_new_n29764__, new_new_n29765__,
    new_new_n29767__, new_new_n29768__, new_new_n29769__, new_new_n29770__,
    new_new_n29771__, new_new_n29772__, new_new_n29773__, new_new_n29774__,
    new_new_n29775__, new_new_n29776__, new_new_n29778__, new_new_n29779__,
    new_new_n29780__, new_new_n29781__, new_new_n29782__, new_new_n29783__,
    new_new_n29784__, new_new_n29785__, new_new_n29786__, new_new_n29788__,
    new_new_n29789__, new_new_n29790__, new_new_n29791__, new_new_n29792__,
    new_new_n29793__, new_new_n29794__, new_new_n29795__, new_new_n29796__,
    new_new_n29797__, new_new_n29798__, new_new_n29800__, new_new_n29801__,
    new_new_n29802__, new_new_n29803__, new_new_n29804__, new_new_n29805__,
    new_new_n29806__, new_new_n29807__, new_new_n29808__, new_new_n29810__,
    new_new_n29811__, new_new_n29812__, new_new_n29813__, new_new_n29814__,
    new_new_n29815__, new_new_n29816__, new_new_n29817__, new_new_n29818__,
    new_new_n29819__, new_new_n29821__, new_new_n29822__, new_new_n29823__,
    new_new_n29824__, new_new_n29825__, new_new_n29826__, new_new_n29827__,
    new_new_n29828__, new_new_n29829__, new_new_n29831__, new_new_n29832__,
    new_new_n29833__, new_new_n29834__, new_new_n29835__, new_new_n29836__,
    new_new_n29837__, new_new_n29838__, new_new_n29839__, new_new_n29840__,
    new_new_n29841__, new_new_n29842__, new_new_n29844__, new_new_n29845__,
    new_new_n29846__, new_new_n29847__, new_new_n29848__, new_new_n29849__,
    new_new_n29850__, new_new_n29851__, new_new_n29852__, new_new_n29854__,
    new_new_n29855__, new_new_n29856__, new_new_n29857__, new_new_n29858__,
    new_new_n29859__, new_new_n29860__, new_new_n29861__, new_new_n29862__,
    new_new_n29863__, new_new_n29865__, new_new_n29866__, new_new_n29867__,
    new_new_n29868__, new_new_n29869__, new_new_n29870__, new_new_n29871__,
    new_new_n29872__, new_new_n29873__, new_new_n29875__, new_new_n29876__,
    new_new_n29877__, new_new_n29878__, new_new_n29879__, new_new_n29880__,
    new_new_n29881__, new_new_n29882__, new_new_n29883__, new_new_n29884__,
    new_new_n29885__, new_new_n29887__, new_new_n29888__, new_new_n29889__,
    new_new_n29890__, new_new_n29891__, new_new_n29892__, new_new_n29893__,
    new_new_n29894__, new_new_n29895__, new_new_n29897__, new_new_n29898__,
    new_new_n29899__, new_new_n29900__, new_new_n29901__, new_new_n29902__,
    new_new_n29903__, new_new_n29904__, new_new_n29905__, new_new_n29906__,
    new_new_n29908__, new_new_n29909__, new_new_n29910__, new_new_n29911__,
    new_new_n29912__, new_new_n29913__, new_new_n29914__, new_new_n29915__,
    new_new_n29916__, new_new_n29918__, new_new_n29919__, new_new_n29920__,
    new_new_n29921__, new_new_n29922__, new_new_n29923__, new_new_n29924__,
    new_new_n29925__, new_new_n29926__, new_new_n29927__, new_new_n29928__,
    new_new_n29929__, new_new_n29931__, new_new_n29932__, new_new_n29933__,
    new_new_n29934__, new_new_n29935__, new_new_n29936__, new_new_n29937__,
    new_new_n29938__, new_new_n29939__, new_new_n29941__, new_new_n29942__,
    new_new_n29943__, new_new_n29944__, new_new_n29945__, new_new_n29946__,
    new_new_n29947__, new_new_n29948__, new_new_n29949__, new_new_n29950__,
    new_new_n29952__, new_new_n29953__, new_new_n29954__, new_new_n29955__,
    new_new_n29956__, new_new_n29957__, new_new_n29958__, new_new_n29959__,
    new_new_n29960__, new_new_n29962__, new_new_n29963__, new_new_n29964__,
    new_new_n29965__, new_new_n29966__, new_new_n29967__, new_new_n29968__,
    new_new_n29969__, new_new_n29970__, new_new_n29971__, new_new_n29972__,
    new_new_n29974__, new_new_n29975__, new_new_n29976__, new_new_n29977__,
    new_new_n29978__, new_new_n29979__, new_new_n29980__, new_new_n29981__,
    new_new_n29982__, new_new_n29984__, new_new_n29985__, new_new_n29986__,
    new_new_n29987__, new_new_n29988__, new_new_n29989__, new_new_n29990__,
    new_new_n29991__, new_new_n29992__, new_new_n29993__, new_new_n29995__,
    new_new_n29996__, new_new_n29997__, new_new_n29998__, new_new_n29999__,
    new_new_n30000__, new_new_n30001__, new_new_n30002__, new_new_n30003__,
    new_new_n30005__, new_new_n30007__, new_new_n30010__, new_new_n30012__,
    new_new_n30014__, new_new_n30015__, new_new_n30016__, new_new_n30017__,
    new_new_n30018__, new_new_n30022__, new_new_n30023__, new_new_n30025__,
    new_new_n30026__, new_new_n30027__, new_new_n30028__, new_new_n30029__,
    new_new_n30030__, new_new_n30031__, new_new_n30032__, new_new_n30033__,
    new_new_n30034__, new_new_n30035__, new_new_n30036__, new_new_n30037__,
    new_new_n30038__, new_new_n30039__, new_new_n30040__, new_new_n30041__,
    new_new_n30042__, new_new_n30043__, new_new_n30044__, new_new_n30046__,
    new_new_n30047__, new_new_n30048__, new_new_n30049__, new_new_n30050__,
    new_new_n30051__, new_new_n30052__, new_new_n30053__, new_new_n30054__,
    new_new_n30055__, new_new_n30056__, new_new_n30057__, new_new_n30058__,
    new_new_n30059__, new_new_n30060__, new_new_n30061__, new_new_n30062__,
    new_new_n30063__, new_new_n30065__, new_new_n30066__, new_new_n30067__,
    new_new_n30068__, new_new_n30069__, new_new_n30070__, new_new_n30071__,
    new_new_n30072__, new_new_n30073__, new_new_n30074__, new_new_n30075__,
    new_new_n30076__, new_new_n30077__, new_new_n30078__, new_new_n30079__,
    new_new_n30080__, new_new_n30081__, new_new_n30082__, new_new_n30084__,
    new_new_n30085__, new_new_n30086__, new_new_n30087__, new_new_n30088__,
    new_new_n30089__, new_new_n30090__, new_new_n30091__, new_new_n30092__,
    new_new_n30093__, new_new_n30094__, new_new_n30095__, new_new_n30096__,
    new_new_n30097__, new_new_n30098__, new_new_n30099__, new_new_n30100__,
    new_new_n30101__, new_new_n30103__, new_new_n30104__, new_new_n30105__,
    new_new_n30106__, new_new_n30107__, new_new_n30108__, new_new_n30109__,
    new_new_n30110__, new_new_n30111__, new_new_n30112__, new_new_n30113__,
    new_new_n30114__, new_new_n30115__, new_new_n30116__, new_new_n30117__,
    new_new_n30118__, new_new_n30119__, new_new_n30120__, new_new_n30122__,
    new_new_n30123__, new_new_n30124__, new_new_n30125__, new_new_n30126__,
    new_new_n30127__, new_new_n30128__, new_new_n30129__, new_new_n30130__,
    new_new_n30131__, new_new_n30132__, new_new_n30133__, new_new_n30134__,
    new_new_n30135__, new_new_n30136__, new_new_n30137__, new_new_n30138__,
    new_new_n30139__, new_new_n30141__, new_new_n30142__, new_new_n30143__,
    new_new_n30144__, new_new_n30145__, new_new_n30146__, new_new_n30147__,
    new_new_n30148__, new_new_n30149__, new_new_n30150__, new_new_n30151__,
    new_new_n30152__, new_new_n30153__, new_new_n30154__, new_new_n30155__,
    new_new_n30156__, new_new_n30157__, new_new_n30158__, new_new_n30160__,
    new_new_n30161__, new_new_n30162__, new_new_n30163__, new_new_n30164__,
    new_new_n30165__, new_new_n30166__, new_new_n30167__, new_new_n30168__,
    new_new_n30169__, new_new_n30170__, new_new_n30171__, new_new_n30172__,
    new_new_n30173__, new_new_n30174__, new_new_n30175__, new_new_n30176__,
    new_new_n30177__, new_new_n30179__, new_new_n30180__, new_new_n30181__,
    new_new_n30182__, new_new_n30183__, new_new_n30184__, new_new_n30185__,
    new_new_n30186__, new_new_n30187__, new_new_n30188__, new_new_n30189__,
    new_new_n30190__, new_new_n30191__, new_new_n30192__, new_new_n30193__,
    new_new_n30194__, new_new_n30195__, new_new_n30196__, new_new_n30197__,
    new_new_n30198__, new_new_n30200__, new_new_n30201__, new_new_n30202__,
    new_new_n30203__, new_new_n30204__, new_new_n30205__, new_new_n30206__,
    new_new_n30207__, new_new_n30208__, new_new_n30209__, new_new_n30210__,
    new_new_n30211__, new_new_n30212__, new_new_n30213__, new_new_n30214__,
    new_new_n30215__, new_new_n30216__, new_new_n30217__, new_new_n30218__,
    new_new_n30219__, new_new_n30221__, new_new_n30222__, new_new_n30223__,
    new_new_n30224__, new_new_n30225__, new_new_n30226__, new_new_n30227__,
    new_new_n30228__, new_new_n30229__, new_new_n30230__, new_new_n30231__,
    new_new_n30232__, new_new_n30233__, new_new_n30234__, new_new_n30235__,
    new_new_n30236__, new_new_n30237__, new_new_n30238__, new_new_n30240__,
    new_new_n30241__, new_new_n30242__, new_new_n30243__, new_new_n30244__,
    new_new_n30245__, new_new_n30246__, new_new_n30247__, new_new_n30248__,
    new_new_n30249__, new_new_n30250__, new_new_n30251__, new_new_n30252__,
    new_new_n30253__, new_new_n30254__, new_new_n30255__, new_new_n30256__,
    new_new_n30257__, new_new_n30258__, new_new_n30259__, new_new_n30261__,
    new_new_n30262__, new_new_n30263__, new_new_n30264__, new_new_n30265__,
    new_new_n30266__, new_new_n30267__, new_new_n30268__, new_new_n30269__,
    new_new_n30270__, new_new_n30271__, new_new_n30272__, new_new_n30273__,
    new_new_n30274__, new_new_n30275__, new_new_n30276__, new_new_n30277__,
    new_new_n30278__, new_new_n30279__, new_new_n30280__, new_new_n30282__,
    new_new_n30283__, new_new_n30284__, new_new_n30285__, new_new_n30286__,
    new_new_n30287__, new_new_n30288__, new_new_n30289__, new_new_n30290__,
    new_new_n30291__, new_new_n30292__, new_new_n30293__, new_new_n30294__,
    new_new_n30295__, new_new_n30296__, new_new_n30297__, new_new_n30298__,
    new_new_n30299__, new_new_n30301__, new_new_n30302__, new_new_n30303__,
    new_new_n30304__, new_new_n30305__, new_new_n30306__, new_new_n30307__,
    new_new_n30308__, new_new_n30309__, new_new_n30310__, new_new_n30311__,
    new_new_n30312__, new_new_n30313__, new_new_n30314__, new_new_n30315__,
    new_new_n30316__, new_new_n30317__, new_new_n30318__, new_new_n30320__,
    new_new_n30321__, new_new_n30322__, new_new_n30323__, new_new_n30324__,
    new_new_n30325__, new_new_n30326__, new_new_n30327__, new_new_n30328__,
    new_new_n30329__, new_new_n30330__, new_new_n30331__, new_new_n30332__,
    new_new_n30333__, new_new_n30334__, new_new_n30335__, new_new_n30336__,
    new_new_n30337__, new_new_n30339__, new_new_n30340__, new_new_n30341__,
    new_new_n30342__, new_new_n30343__, new_new_n30344__, new_new_n30345__,
    new_new_n30346__, new_new_n30347__, new_new_n30348__, new_new_n30349__,
    new_new_n30350__, new_new_n30351__, new_new_n30352__, new_new_n30353__,
    new_new_n30354__, new_new_n30355__, new_new_n30356__, new_new_n30357__,
    new_new_n30359__, new_new_n30360__, new_new_n30361__, new_new_n30362__,
    new_new_n30363__, new_new_n30364__, new_new_n30365__, new_new_n30366__,
    new_new_n30367__, new_new_n30368__, new_new_n30369__, new_new_n30370__,
    new_new_n30371__, new_new_n30372__, new_new_n30373__, new_new_n30374__,
    new_new_n30375__, new_new_n30376__, new_new_n30378__, new_new_n30379__,
    new_new_n30380__, new_new_n30381__, new_new_n30382__, new_new_n30383__,
    new_new_n30384__, new_new_n30385__, new_new_n30386__, new_new_n30387__,
    new_new_n30388__, new_new_n30389__, new_new_n30390__, new_new_n30391__,
    new_new_n30392__, new_new_n30393__, new_new_n30394__, new_new_n30395__,
    new_new_n30397__, new_new_n30398__, new_new_n30399__, new_new_n30400__,
    new_new_n30401__, new_new_n30402__, new_new_n30403__, new_new_n30404__,
    new_new_n30405__, new_new_n30406__, new_new_n30407__, new_new_n30408__,
    new_new_n30409__, new_new_n30410__, new_new_n30411__, new_new_n30412__,
    new_new_n30413__, new_new_n30414__, new_new_n30416__, new_new_n30417__,
    new_new_n30418__, new_new_n30419__, new_new_n30420__, new_new_n30421__,
    new_new_n30422__, new_new_n30423__, new_new_n30424__, new_new_n30425__,
    new_new_n30426__, new_new_n30427__, new_new_n30428__, new_new_n30429__,
    new_new_n30430__, new_new_n30431__, new_new_n30432__, new_new_n30433__,
    new_new_n30435__, new_new_n30436__, new_new_n30437__, new_new_n30438__,
    new_new_n30439__, new_new_n30440__, new_new_n30441__, new_new_n30442__,
    new_new_n30443__, new_new_n30444__, new_new_n30445__, new_new_n30446__,
    new_new_n30447__, new_new_n30448__, new_new_n30449__, new_new_n30450__,
    new_new_n30451__, new_new_n30452__, new_new_n30454__, new_new_n30455__,
    new_new_n30456__, new_new_n30457__, new_new_n30458__, new_new_n30459__,
    new_new_n30460__, new_new_n30461__, new_new_n30462__, new_new_n30463__,
    new_new_n30464__, new_new_n30465__, new_new_n30466__, new_new_n30467__,
    new_new_n30468__, new_new_n30469__, new_new_n30470__, new_new_n30471__,
    new_new_n30473__, new_new_n30474__, new_new_n30475__, new_new_n30476__,
    new_new_n30477__, new_new_n30478__, new_new_n30479__, new_new_n30480__,
    new_new_n30481__, new_new_n30482__, new_new_n30483__, new_new_n30484__,
    new_new_n30485__, new_new_n30486__, new_new_n30487__, new_new_n30488__,
    new_new_n30489__, new_new_n30490__, new_new_n30491__, new_new_n30493__,
    new_new_n30494__, new_new_n30495__, new_new_n30496__, new_new_n30497__,
    new_new_n30498__, new_new_n30499__, new_new_n30500__, new_new_n30501__,
    new_new_n30502__, new_new_n30503__, new_new_n30504__, new_new_n30505__,
    new_new_n30506__, new_new_n30507__, new_new_n30508__, new_new_n30509__,
    new_new_n30510__, new_new_n30512__, new_new_n30513__, new_new_n30514__,
    new_new_n30515__, new_new_n30516__, new_new_n30517__, new_new_n30518__,
    new_new_n30519__, new_new_n30520__, new_new_n30521__, new_new_n30522__,
    new_new_n30523__, new_new_n30524__, new_new_n30525__, new_new_n30526__,
    new_new_n30527__, new_new_n30528__, new_new_n30529__, new_new_n30531__,
    new_new_n30532__, new_new_n30533__, new_new_n30534__, new_new_n30535__,
    new_new_n30536__, new_new_n30537__, new_new_n30538__, new_new_n30539__,
    new_new_n30540__, new_new_n30541__, new_new_n30542__, new_new_n30543__,
    new_new_n30544__, new_new_n30545__, new_new_n30546__, new_new_n30547__,
    new_new_n30548__, new_new_n30549__, new_new_n30550__, new_new_n30552__,
    new_new_n30553__, new_new_n30554__, new_new_n30555__, new_new_n30556__,
    new_new_n30557__, new_new_n30558__, new_new_n30559__, new_new_n30560__,
    new_new_n30561__, new_new_n30562__, new_new_n30563__, new_new_n30564__,
    new_new_n30565__, new_new_n30566__, new_new_n30567__, new_new_n30568__,
    new_new_n30569__, new_new_n30570__, new_new_n30571__, new_new_n30573__,
    new_new_n30574__, new_new_n30575__, new_new_n30576__, new_new_n30577__,
    new_new_n30578__, new_new_n30579__, new_new_n30580__, new_new_n30581__,
    new_new_n30582__, new_new_n30583__, new_new_n30584__, new_new_n30585__,
    new_new_n30586__, new_new_n30587__, new_new_n30588__, new_new_n30589__,
    new_new_n30590__, new_new_n30592__, new_new_n30593__, new_new_n30594__,
    new_new_n30595__, new_new_n30596__, new_new_n30597__, new_new_n30598__,
    new_new_n30599__, new_new_n30600__, new_new_n30601__, new_new_n30602__,
    new_new_n30603__, new_new_n30604__, new_new_n30605__, new_new_n30606__,
    new_new_n30607__, new_new_n30608__, new_new_n30609__, new_new_n30611__,
    new_new_n30612__, new_new_n30613__, new_new_n30614__, new_new_n30615__,
    new_new_n30616__, new_new_n30617__, new_new_n30618__, new_new_n30619__,
    new_new_n30620__, new_new_n30621__, new_new_n30622__, new_new_n30623__,
    new_new_n30624__, new_new_n30625__, new_new_n30626__, new_new_n30627__,
    new_new_n30628__, new_new_n30630__, new_new_n30631__, new_new_n30632__,
    new_new_n30633__, new_new_n30634__, new_new_n30635__, new_new_n30636__,
    new_new_n30637__, new_new_n30638__, new_new_n30639__, new_new_n30640__,
    new_new_n30641__, new_new_n30642__, new_new_n30643__, new_new_n30644__,
    new_new_n30645__, new_new_n30646__, new_new_n30647__, new_new_n30648__,
    new_new_n30649__, new_new_n30650__, new_new_n30651__, new_new_n30653__,
    new_new_n30654__, new_new_n30655__, new_new_n30656__, new_new_n30657__,
    new_new_n30658__, new_new_n30659__, new_new_n30660__, new_new_n30661__,
    new_new_n30662__, new_new_n30663__, new_new_n30664__, new_new_n30665__,
    new_new_n30666__, new_new_n30668__, new_new_n30669__, new_new_n30670__,
    new_new_n30671__, new_new_n30672__, new_new_n30673__, new_new_n30674__,
    new_new_n30675__, new_new_n30676__, new_new_n30677__, new_new_n30678__,
    new_new_n30679__, new_new_n30680__, new_new_n30681__, new_new_n30683__,
    new_new_n30684__, new_new_n30685__, new_new_n30686__, new_new_n30687__,
    new_new_n30688__, new_new_n30689__, new_new_n30690__, new_new_n30691__,
    new_new_n30692__, new_new_n30693__, new_new_n30694__, new_new_n30695__,
    new_new_n30696__, new_new_n30698__, new_new_n30699__, new_new_n30700__,
    new_new_n30701__, new_new_n30702__, new_new_n30703__, new_new_n30704__,
    new_new_n30705__, new_new_n30706__, new_new_n30707__, new_new_n30708__,
    new_new_n30709__, new_new_n30710__, new_new_n30711__, new_new_n30713__,
    new_new_n30714__, new_new_n30715__, new_new_n30716__, new_new_n30717__,
    new_new_n30718__, new_new_n30719__, new_new_n30720__, new_new_n30721__,
    new_new_n30722__, new_new_n30723__, new_new_n30724__, new_new_n30725__,
    new_new_n30726__, new_new_n30728__, new_new_n30729__, new_new_n30730__,
    new_new_n30731__, new_new_n30732__, new_new_n30733__, new_new_n30734__,
    new_new_n30735__, new_new_n30736__, new_new_n30737__, new_new_n30738__,
    new_new_n30739__, new_new_n30740__, new_new_n30741__, new_new_n30743__,
    new_new_n30744__, new_new_n30745__, new_new_n30746__, new_new_n30747__,
    new_new_n30748__, new_new_n30749__, new_new_n30750__, new_new_n30751__,
    new_new_n30752__, new_new_n30753__, new_new_n30754__, new_new_n30756__,
    new_new_n30757__, new_new_n30758__, new_new_n30759__, new_new_n30760__,
    new_new_n30761__, new_new_n30762__, new_new_n30763__, new_new_n30764__,
    new_new_n30765__, new_new_n30766__, new_new_n30767__, new_new_n30768__,
    new_new_n30769__, new_new_n30771__, new_new_n30772__, new_new_n30773__,
    new_new_n30774__, new_new_n30775__, new_new_n30776__, new_new_n30777__,
    new_new_n30778__, new_new_n30779__, new_new_n30780__, new_new_n30781__,
    new_new_n30782__, new_new_n30783__, new_new_n30784__, new_new_n30786__,
    new_new_n30787__, new_new_n30788__, new_new_n30789__, new_new_n30790__,
    new_new_n30791__, new_new_n30792__, new_new_n30793__, new_new_n30794__,
    new_new_n30795__, new_new_n30796__, new_new_n30797__, new_new_n30798__,
    new_new_n30799__, new_new_n30801__, new_new_n30802__, new_new_n30803__,
    new_new_n30804__, new_new_n30805__, new_new_n30806__, new_new_n30807__,
    new_new_n30808__, new_new_n30809__, new_new_n30810__, new_new_n30811__,
    new_new_n30812__, new_new_n30814__, new_new_n30815__, new_new_n30816__,
    new_new_n30817__, new_new_n30818__, new_new_n30819__, new_new_n30820__,
    new_new_n30821__, new_new_n30822__, new_new_n30823__, new_new_n30824__,
    new_new_n30825__, new_new_n30826__, new_new_n30827__, new_new_n30829__,
    new_new_n30830__, new_new_n30831__, new_new_n30832__, new_new_n30833__,
    new_new_n30834__, new_new_n30835__, new_new_n30836__, new_new_n30837__,
    new_new_n30838__, new_new_n30839__, new_new_n30840__, new_new_n30841__,
    new_new_n30842__, new_new_n30844__, new_new_n30845__, new_new_n30846__,
    new_new_n30847__, new_new_n30848__, new_new_n30849__, new_new_n30850__,
    new_new_n30851__, new_new_n30852__, new_new_n30853__, new_new_n30854__,
    new_new_n30855__, new_new_n30857__, new_new_n30858__, new_new_n30859__,
    new_new_n30860__, new_new_n30861__, new_new_n30862__, new_new_n30863__,
    new_new_n30864__, new_new_n30865__, new_new_n30866__, new_new_n30867__,
    new_new_n30868__, new_new_n30869__, new_new_n30870__, new_new_n30872__,
    new_new_n30873__, new_new_n30874__, new_new_n30875__, new_new_n30876__,
    new_new_n30877__, new_new_n30878__, new_new_n30879__, new_new_n30880__,
    new_new_n30881__, new_new_n30882__, new_new_n30883__, new_new_n30884__,
    new_new_n30885__, new_new_n30887__, new_new_n30888__, new_new_n30889__,
    new_new_n30890__, new_new_n30891__, new_new_n30892__, new_new_n30893__,
    new_new_n30894__, new_new_n30895__, new_new_n30896__, new_new_n30897__,
    new_new_n30898__, new_new_n30899__, new_new_n30900__, new_new_n30902__,
    new_new_n30903__, new_new_n30904__, new_new_n30905__, new_new_n30906__,
    new_new_n30907__, new_new_n30908__, new_new_n30909__, new_new_n30910__,
    new_new_n30911__, new_new_n30912__, new_new_n30913__, new_new_n30914__,
    new_new_n30915__, new_new_n30917__, new_new_n30918__, new_new_n30919__,
    new_new_n30920__, new_new_n30921__, new_new_n30922__, new_new_n30923__,
    new_new_n30924__, new_new_n30925__, new_new_n30926__, new_new_n30927__,
    new_new_n30928__, new_new_n30929__, new_new_n30930__, new_new_n30932__,
    new_new_n30933__, new_new_n30934__, new_new_n30935__, new_new_n30936__,
    new_new_n30937__, new_new_n30938__, new_new_n30939__, new_new_n30940__,
    new_new_n30941__, new_new_n30942__, new_new_n30943__, new_new_n30944__,
    new_new_n30945__, new_new_n30947__, new_new_n30948__, new_new_n30949__,
    new_new_n30950__, new_new_n30951__, new_new_n30952__, new_new_n30953__,
    new_new_n30954__, new_new_n30955__, new_new_n30956__, new_new_n30957__,
    new_new_n30958__, new_new_n30959__, new_new_n30960__, new_new_n30962__,
    new_new_n30963__, new_new_n30964__, new_new_n30965__, new_new_n30966__,
    new_new_n30967__, new_new_n30968__, new_new_n30969__, new_new_n30970__,
    new_new_n30971__, new_new_n30972__, new_new_n30973__, new_new_n30974__,
    new_new_n30976__, new_new_n30977__, new_new_n30978__, new_new_n30979__,
    new_new_n30980__, new_new_n30981__, new_new_n30982__, new_new_n30983__,
    new_new_n30984__, new_new_n30985__, new_new_n30986__, new_new_n30987__,
    new_new_n30988__, new_new_n30989__, new_new_n30991__, new_new_n30992__,
    new_new_n30993__, new_new_n30994__, new_new_n30995__, new_new_n30996__,
    new_new_n30997__, new_new_n30998__, new_new_n30999__, new_new_n31000__,
    new_new_n31001__, new_new_n31002__, new_new_n31003__, new_new_n31004__,
    new_new_n31006__, new_new_n31007__, new_new_n31008__, new_new_n31009__,
    new_new_n31010__, new_new_n31011__, new_new_n31012__, new_new_n31013__,
    new_new_n31014__, new_new_n31015__, new_new_n31016__, new_new_n31017__,
    new_new_n31018__, new_new_n31019__, new_new_n31021__, new_new_n31022__,
    new_new_n31023__, new_new_n31024__, new_new_n31025__, new_new_n31026__,
    new_new_n31027__, new_new_n31028__, new_new_n31029__, new_new_n31030__,
    new_new_n31031__, new_new_n31032__, new_new_n31033__, new_new_n31034__,
    new_new_n31036__, new_new_n31037__, new_new_n31038__, new_new_n31039__,
    new_new_n31040__, new_new_n31041__, new_new_n31042__, new_new_n31043__,
    new_new_n31044__, new_new_n31045__, new_new_n31046__, new_new_n31047__,
    new_new_n31049__, new_new_n31050__, new_new_n31051__, new_new_n31052__,
    new_new_n31053__, new_new_n31054__, new_new_n31055__, new_new_n31056__,
    new_new_n31057__, new_new_n31058__, new_new_n31059__, new_new_n31060__,
    new_new_n31062__, new_new_n31063__, new_new_n31064__, new_new_n31065__,
    new_new_n31066__, new_new_n31067__, new_new_n31068__, new_new_n31069__,
    new_new_n31070__, new_new_n31071__, new_new_n31072__, new_new_n31073__,
    new_new_n31075__, new_new_n31076__, new_new_n31077__, new_new_n31078__,
    new_new_n31079__, new_new_n31080__, new_new_n31081__, new_new_n31082__,
    new_new_n31083__, new_new_n31084__, new_new_n31085__, new_new_n31086__,
    new_new_n31088__, new_new_n31089__, new_new_n31090__, new_new_n31091__,
    new_new_n31092__, new_new_n31093__, new_new_n31094__, new_new_n31095__,
    new_new_n31096__, new_new_n31097__, new_new_n31098__, new_new_n31099__,
    new_new_n31101__, new_new_n31102__, new_new_n31103__, new_new_n31104__,
    new_new_n31105__, new_new_n31106__, new_new_n31107__, new_new_n31108__,
    new_new_n31109__, new_new_n31110__, new_new_n31111__, new_new_n31112__,
    new_new_n31113__, new_new_n31114__, new_new_n31116__, new_new_n31117__,
    new_new_n31118__, new_new_n31119__, new_new_n31120__, new_new_n31121__,
    new_new_n31122__, new_new_n31123__, new_new_n31124__, new_new_n31125__,
    new_new_n31126__, new_new_n31127__, new_new_n31128__, new_new_n31129__,
    new_new_n31131__, new_new_n31132__, new_new_n31133__, new_new_n31134__,
    new_new_n31135__, new_new_n31136__, new_new_n31137__, new_new_n31138__,
    new_new_n31139__, new_new_n31140__, new_new_n31141__, new_new_n31142__,
    new_new_n31143__, new_new_n31144__, new_new_n31146__, new_new_n31147__,
    new_new_n31148__, new_new_n31149__, new_new_n31150__, new_new_n31151__,
    new_new_n31152__, new_new_n31153__, new_new_n31154__, new_new_n31155__,
    new_new_n31156__, new_new_n31157__, new_new_n31158__, new_new_n31159__,
    new_new_n31161__, new_new_n31162__, new_new_n31163__, new_new_n31164__,
    new_new_n31165__, new_new_n31166__, new_new_n31167__, new_new_n31168__,
    new_new_n31169__, new_new_n31170__, new_new_n31171__, new_new_n31172__,
    new_new_n31173__, new_new_n31174__, new_new_n31176__, new_new_n31177__,
    new_new_n31178__, new_new_n31179__, new_new_n31180__, new_new_n31181__,
    new_new_n31182__, new_new_n31183__, new_new_n31184__, new_new_n31185__,
    new_new_n31186__, new_new_n31187__, new_new_n31188__, new_new_n31189__,
    new_new_n31191__, new_new_n31192__, new_new_n31193__, new_new_n31194__,
    new_new_n31195__, new_new_n31196__, new_new_n31197__, new_new_n31198__,
    new_new_n31199__, new_new_n31200__, new_new_n31201__, new_new_n31202__,
    new_new_n31203__, new_new_n31204__, new_new_n31206__, new_new_n31207__,
    new_new_n31208__, new_new_n31209__, new_new_n31210__, new_new_n31211__,
    new_new_n31212__, new_new_n31213__, new_new_n31214__, new_new_n31215__,
    new_new_n31216__, new_new_n31217__, new_new_n31218__, new_new_n31219__,
    new_new_n31221__, new_new_n31222__, new_new_n31223__, new_new_n31224__,
    new_new_n31225__, new_new_n31226__, new_new_n31227__, new_new_n31228__,
    new_new_n31229__, new_new_n31230__, new_new_n31231__, new_new_n31232__,
    new_new_n31233__, new_new_n31234__, new_new_n31236__, new_new_n31237__,
    new_new_n31238__, new_new_n31239__, new_new_n31240__, new_new_n31241__,
    new_new_n31242__, new_new_n31243__, new_new_n31244__, new_new_n31245__,
    new_new_n31246__, new_new_n31247__, new_new_n31248__, new_new_n31249__,
    new_new_n31251__, new_new_n31252__, new_new_n31253__, new_new_n31254__,
    new_new_n31255__, new_new_n31256__, new_new_n31257__, new_new_n31258__,
    new_new_n31259__, new_new_n31260__, new_new_n31261__, new_new_n31262__,
    new_new_n31263__, new_new_n31264__, new_new_n31266__, new_new_n31267__,
    new_new_n31268__, new_new_n31269__, new_new_n31270__, new_new_n31271__,
    new_new_n31272__, new_new_n31273__, new_new_n31274__, new_new_n31275__,
    new_new_n31276__, new_new_n31277__, new_new_n31278__, new_new_n31279__,
    new_new_n31281__, new_new_n31282__, new_new_n31283__, new_new_n31284__,
    new_new_n31285__, new_new_n31286__, new_new_n31287__, new_new_n31288__,
    new_new_n31289__, new_new_n31290__, new_new_n31291__, new_new_n31292__,
    new_new_n31293__, new_new_n31294__, new_new_n31296__, new_new_n31297__,
    new_new_n31298__, new_new_n31299__, new_new_n31300__, new_new_n31301__,
    new_new_n31302__, new_new_n31303__, new_new_n31304__, new_new_n31305__,
    new_new_n31306__, new_new_n31307__, new_new_n31308__, new_new_n31309__,
    new_new_n31311__, new_new_n31312__, new_new_n31313__, new_new_n31314__,
    new_new_n31315__, new_new_n31316__, new_new_n31317__, new_new_n31318__,
    new_new_n31319__, new_new_n31320__, new_new_n31321__, new_new_n31322__,
    new_new_n31323__, new_new_n31324__, new_new_n31326__, new_new_n31327__,
    new_new_n31328__, new_new_n31329__, new_new_n31330__, new_new_n31331__,
    new_new_n31332__, new_new_n31333__, new_new_n31334__, new_new_n31335__,
    new_new_n31336__, new_new_n31337__, new_new_n31338__, new_new_n31339__,
    new_new_n31341__, new_new_n31342__, new_new_n31343__, new_new_n31344__,
    new_new_n31345__, new_new_n31346__, new_new_n31347__, new_new_n31348__,
    new_new_n31349__, new_new_n31350__, new_new_n31351__, new_new_n31352__,
    new_new_n31353__, new_new_n31354__, new_new_n31356__, new_new_n31357__,
    new_new_n31358__, new_new_n31359__, new_new_n31360__, new_new_n31361__,
    new_new_n31362__, new_new_n31363__, new_new_n31364__, new_new_n31365__,
    new_new_n31366__, new_new_n31367__, new_new_n31368__, new_new_n31369__,
    new_new_n31371__, new_new_n31372__, new_new_n31373__, new_new_n31374__,
    new_new_n31375__, new_new_n31376__, new_new_n31377__, new_new_n31378__,
    new_new_n31379__, new_new_n31380__, new_new_n31381__, new_new_n31382__,
    new_new_n31383__, new_new_n31384__, new_new_n31386__, new_new_n31387__,
    new_new_n31388__, new_new_n31389__, new_new_n31390__, new_new_n31391__,
    new_new_n31392__, new_new_n31393__, new_new_n31394__, new_new_n31395__,
    new_new_n31396__, new_new_n31397__, new_new_n31398__, new_new_n31399__,
    new_new_n31401__, new_new_n31402__, new_new_n31403__, new_new_n31404__,
    new_new_n31405__, new_new_n31406__, new_new_n31407__, new_new_n31408__,
    new_new_n31409__, new_new_n31410__, new_new_n31411__, new_new_n31412__,
    new_new_n31413__, new_new_n31414__, new_new_n31416__, new_new_n31417__,
    new_new_n31418__, new_new_n31419__, new_new_n31420__, new_new_n31421__,
    new_new_n31422__, new_new_n31423__, new_new_n31424__, new_new_n31425__,
    new_new_n31426__, new_new_n31427__, new_new_n31428__, new_new_n31429__,
    new_new_n31431__, new_new_n31432__, new_new_n31433__, new_new_n31434__,
    new_new_n31435__, new_new_n31436__, new_new_n31437__, new_new_n31438__,
    new_new_n31439__, new_new_n31440__, new_new_n31441__, new_new_n31442__,
    new_new_n31443__, new_new_n31444__, new_new_n31446__, new_new_n31447__,
    new_new_n31448__, new_new_n31449__, new_new_n31450__, new_new_n31451__,
    new_new_n31452__, new_new_n31453__, new_new_n31454__, new_new_n31455__,
    new_new_n31456__, new_new_n31457__, new_new_n31458__, new_new_n31459__,
    new_new_n31461__, new_new_n31462__, new_new_n31463__, new_new_n31464__,
    new_new_n31465__, new_new_n31466__, new_new_n31467__, new_new_n31468__,
    new_new_n31469__, new_new_n31470__, new_new_n31471__, new_new_n31472__,
    new_new_n31473__, new_new_n31474__, new_new_n31476__, new_new_n31477__,
    new_new_n31478__, new_new_n31479__, new_new_n31480__, new_new_n31481__,
    new_new_n31482__, new_new_n31483__, new_new_n31484__, new_new_n31485__,
    new_new_n31486__, new_new_n31487__, new_new_n31488__, new_new_n31489__,
    new_new_n31491__, new_new_n31492__, new_new_n31493__, new_new_n31494__,
    new_new_n31495__, new_new_n31496__, new_new_n31497__, new_new_n31498__,
    new_new_n31499__, new_new_n31500__, new_new_n31501__, new_new_n31502__,
    new_new_n31503__, new_new_n31504__, new_new_n31506__, new_new_n31507__,
    new_new_n31508__, new_new_n31509__, new_new_n31510__, new_new_n31511__,
    new_new_n31512__, new_new_n31513__, new_new_n31514__, new_new_n31515__,
    new_new_n31516__, new_new_n31517__, new_new_n31518__, new_new_n31519__,
    new_new_n31521__, new_new_n31522__, new_new_n31523__, new_new_n31524__,
    new_new_n31525__, new_new_n31526__, new_new_n31527__, new_new_n31528__,
    new_new_n31529__, new_new_n31530__, new_new_n31531__, new_new_n31532__,
    new_new_n31533__, new_new_n31534__, new_new_n31536__, new_new_n31537__,
    new_new_n31538__, new_new_n31539__, new_new_n31540__, new_new_n31541__,
    new_new_n31542__, new_new_n31543__, new_new_n31544__, new_new_n31545__,
    new_new_n31546__, new_new_n31547__, new_new_n31548__, new_new_n31549__,
    new_new_n31551__, new_new_n31552__, new_new_n31553__, new_new_n31554__,
    new_new_n31555__, new_new_n31556__, new_new_n31557__, new_new_n31558__,
    new_new_n31559__, new_new_n31560__, new_new_n31561__, new_new_n31562__,
    new_new_n31563__, new_new_n31564__, new_new_n31566__, new_new_n31567__,
    new_new_n31568__, new_new_n31569__, new_new_n31570__, new_new_n31571__,
    new_new_n31572__, new_new_n31573__, new_new_n31574__, new_new_n31575__,
    new_new_n31576__, new_new_n31577__, new_new_n31578__, new_new_n31579__,
    new_new_n31581__, new_new_n31582__, new_new_n31583__, new_new_n31584__,
    new_new_n31585__, new_new_n31586__, new_new_n31587__, new_new_n31588__,
    new_new_n31589__, new_new_n31590__, new_new_n31591__, new_new_n31592__,
    new_new_n31593__, new_new_n31594__, new_new_n32232__, new_new_n32233__,
    new_new_n32234__, new_new_n32235__, new_new_n32236__, new_new_n32237__,
    new_new_n32238__, new_new_n32239__, new_new_n32240__, new_new_n32241__,
    new_new_n32242__, new_new_n32243__, new_new_n32244__, new_new_n32245__,
    new_new_n32246__, new_new_n32247__, new_new_n32248__, new_new_n32249__,
    new_new_n32250__, new_new_n32251__, new_new_n32252__, new_new_n32253__,
    new_new_n32254__, new_new_n32255__, new_new_n32256__, new_new_n32257__,
    new_new_n32258__, new_new_n32259__, new_new_n32260__, new_new_n32261__,
    new_new_n32262__, new_new_n32263__, new_new_n32264__, new_new_n32265__,
    new_new_n32266__, new_new_n32267__, new_new_n32268__, new_new_n32269__,
    new_new_n32270__, new_new_n32271__, new_new_n32272__, new_new_n32273__,
    new_new_n32274__, new_new_n32275__, new_new_n32276__, new_new_n32277__,
    new_new_n32278__, new_new_n32279__, new_new_n32280__, new_new_n32281__,
    new_new_n32282__, new_new_n32283__, new_new_n32284__, new_new_n32285__,
    new_new_n32286__, new_new_n32287__, new_new_n32288__, new_new_n32289__,
    new_new_n32290__, new_new_n32291__, new_new_n32292__, new_new_n32293__,
    new_new_n32294__, new_new_n32295__, new_new_n32296__, new_new_n32297__,
    new_new_n32298__, new_new_n32299__, new_new_n32300__, new_new_n32301__,
    new_new_n32302__, new_new_n32303__, new_new_n32304__, new_new_n32305__,
    new_new_n32306__, new_new_n32307__, new_new_n32308__, new_new_n32309__,
    new_new_n32310__, new_new_n32311__, new_new_n32312__, new_new_n32313__,
    new_new_n32314__, new_new_n32315__, new_new_n32316__, new_new_n32317__,
    new_new_n32318__, new_new_n32319__, new_new_n32320__, new_new_n32321__,
    new_new_n32322__, new_new_n32323__, new_new_n32324__, new_new_n32325__,
    new_new_n32326__, new_new_n32327__, new_new_n32328__, new_new_n32329__,
    new_new_n32330__, new_new_n32331__, new_new_n32332__, new_new_n32333__,
    new_new_n32334__, new_new_n32335__, new_new_n32336__, new_new_n32337__,
    new_new_n32338__, new_new_n32339__, new_new_n32340__, new_new_n32341__,
    new_new_n32342__, new_new_n32343__, new_new_n32344__, new_new_n32345__,
    new_new_n32346__, new_new_n32347__, new_new_n32348__, new_new_n32349__,
    new_new_n32350__, new_new_n32351__, new_new_n32352__, new_new_n32353__,
    new_new_n32354__, new_new_n32355__, new_new_n32356__, new_new_n32357__,
    new_new_n32358__, new_new_n32359__, new_new_n32360__, new_new_n32361__,
    new_new_n32362__, new_new_n32363__, new_new_n32364__, new_new_n32365__,
    new_new_n32366__, new_new_n32367__, new_new_n32368__, new_new_n32369__,
    new_new_n32370__, new_new_n32371__, new_new_n32372__, new_new_n32373__,
    new_new_n32374__, new_new_n32375__, new_new_n32376__, new_new_n32377__,
    new_new_n32378__, new_new_n32379__, new_new_n32380__, new_new_n32381__,
    new_new_n32382__, new_new_n32383__, new_new_n32384__, new_new_n32385__,
    new_new_n32386__, new_new_n32387__, new_new_n32388__, new_new_n32389__,
    new_new_n32390__, new_new_n32391__, new_new_n32392__, new_new_n32393__,
    new_new_n32394__, new_new_n32395__, new_new_n32396__, new_new_n32397__,
    new_new_n32398__, new_new_n32399__, new_new_n32400__, new_new_n32401__,
    new_new_n32402__, new_new_n32403__, new_new_n32404__, new_new_n32405__,
    new_new_n32406__, new_new_n32407__, new_new_n32408__, new_new_n32409__,
    new_new_n32410__, new_new_n32411__, new_new_n32412__, new_new_n32413__,
    new_new_n32414__, new_new_n32415__, new_new_n32416__, new_new_n32417__,
    new_new_n32418__, new_new_n32419__, new_new_n32420__, new_new_n32421__,
    new_new_n32422__, new_new_n32423__, new_new_n32424__, new_new_n32425__,
    new_new_n32426__, new_new_n32427__, new_new_n32428__, new_new_n32429__,
    new_new_n32430__, new_new_n32431__, new_new_n32432__, new_new_n32433__,
    new_new_n32434__, new_new_n32435__, new_new_n32436__, new_new_n32437__,
    new_new_n32438__, new_new_n32439__, new_new_n32440__, new_new_n32441__,
    new_new_n32442__, new_new_n32443__, new_new_n32444__, new_new_n32445__,
    new_new_n32446__, new_new_n32447__, new_new_n32448__, new_new_n32449__,
    new_new_n32450__, new_new_n32451__, new_new_n32452__, new_new_n32453__,
    new_new_n32454__, new_new_n32455__, new_new_n32456__, new_new_n32457__,
    new_new_n32458__, new_new_n32459__, new_new_n32460__, new_new_n32461__,
    new_new_n32462__, new_new_n32463__, new_new_n32464__, new_new_n32465__,
    new_new_n32466__, new_new_n32467__, new_new_n32468__, new_new_n32469__,
    new_new_n32470__, new_new_n32471__, new_new_n32472__, new_new_n32473__,
    new_new_n32474__, new_new_n32475__, new_new_n32476__, new_new_n32477__,
    new_new_n32478__, new_new_n32479__, new_new_n32480__, new_new_n32481__,
    new_new_n32482__, new_new_n32483__, new_new_n32484__, new_new_n32485__,
    new_new_n32486__, new_new_n32487__, new_new_n32488__, new_new_n32489__,
    new_new_n32490__, new_new_n32491__, new_new_n32492__, new_new_n32493__,
    new_new_n32494__, new_new_n32495__, new_new_n32496__, new_new_n32497__,
    new_new_n32498__, new_new_n32499__, new_new_n32500__, new_new_n32501__,
    new_new_n32502__, new_new_n32503__, new_new_n32504__, new_new_n32505__,
    new_new_n32506__, new_new_n32507__, new_new_n32508__, new_new_n32509__,
    new_new_n32510__, new_new_n32511__, new_new_n32512__, new_new_n32513__,
    new_new_n32514__, new_new_n32515__, new_new_n32516__, new_new_n32517__,
    new_new_n32518__, new_new_n32519__, new_new_n32520__, new_new_n32521__,
    new_new_n32522__, new_new_n32523__, new_new_n32524__, new_new_n32525__,
    new_new_n32526__, new_new_n32527__, new_new_n32528__, new_new_n32529__,
    new_new_n32530__, new_new_n32531__, new_new_n32532__, new_new_n32533__,
    new_new_n32534__, new_new_n32535__, new_new_n32536__, new_new_n32537__,
    new_new_n32538__, new_new_n32539__, new_new_n32540__, new_new_n32541__,
    new_new_n32542__, new_new_n32543__, new_new_n32544__, new_new_n32545__,
    new_new_n32546__, new_new_n32547__, new_new_n32548__, new_new_n32549__,
    new_new_n32550__, new_new_n32551__, new_new_n32552__, new_new_n32553__,
    new_new_n32554__, new_new_n32555__, new_new_n32556__, new_new_n32557__,
    new_new_n32558__, new_new_n32559__, new_new_n32560__, new_new_n32561__,
    new_new_n32562__, new_new_n32563__, new_new_n32564__, new_new_n32565__,
    new_new_n32566__, new_new_n32568__, new_new_n32569__, new_new_n32570__,
    new_new_n32571__, new_new_n32572__, new_new_n32573__, new_new_n32574__,
    new_new_n32575__, new_new_n32576__, new_new_n32577__, new_new_n32578__,
    new_new_n32579__, new_new_n32580__, new_new_n32581__, new_new_n32582__,
    new_new_n32583__, new_new_n32584__, new_new_n32585__, new_new_n32586__,
    new_new_n32587__, new_new_n32588__, new_new_n32589__, new_new_n32590__,
    new_new_n32591__, new_new_n32592__, new_new_n32593__, new_new_n32594__,
    new_new_n32595__, new_new_n32596__, new_new_n32597__, new_new_n32598__,
    new_new_n32599__, new_new_n32600__, new_new_n32601__, new_new_n32602__,
    new_new_n32603__, new_new_n32604__, new_new_n32605__, new_new_n32606__,
    new_new_n32607__, new_new_n32608__, new_new_n32609__, new_new_n32610__,
    new_new_n32611__, new_new_n32612__, new_new_n32613__, new_new_n32614__,
    new_new_n32615__, new_new_n32616__, new_new_n32617__, new_new_n32618__,
    new_new_n32619__, new_new_n32620__, new_new_n32621__, new_new_n32622__,
    new_new_n32623__, new_new_n32624__, new_new_n32625__, new_new_n32626__,
    new_new_n32627__, new_new_n32628__, new_new_n32629__, new_new_n32630__,
    new_new_n32631__, new_new_n32632__, new_new_n32633__, new_new_n32634__,
    new_new_n32635__, new_new_n32636__, new_new_n32637__, new_new_n32638__,
    new_new_n32639__, new_new_n32640__, new_new_n32641__, new_new_n32642__,
    new_new_n32643__, new_new_n32644__, new_new_n32645__, new_new_n32646__,
    new_new_n32647__, new_new_n32648__, new_new_n32649__, new_new_n32650__,
    new_new_n32651__, new_new_n32652__, new_new_n32653__, new_new_n32654__,
    new_new_n32655__, new_new_n32656__, new_new_n32657__, new_new_n32658__,
    new_new_n32659__, new_new_n32660__, new_new_n32661__, new_new_n32662__,
    new_new_n32663__, new_new_n32664__, new_new_n32665__, new_new_n32666__,
    new_new_n32667__, new_new_n32668__, new_new_n32669__, new_new_n32670__,
    new_new_n32671__, new_new_n32672__, new_new_n32673__, new_new_n32674__,
    new_new_n32675__, new_new_n32676__, new_new_n32677__, new_new_n32678__,
    new_new_n32679__, new_new_n32680__, new_new_n32681__, new_new_n32682__,
    new_new_n32683__, new_new_n32684__, new_new_n32685__, new_new_n32686__,
    new_new_n32687__, new_new_n32688__, new_new_n32689__, new_new_n32690__,
    new_new_n32691__, new_new_n32692__, new_new_n32693__, new_new_n32694__,
    new_new_n32695__, new_new_n32696__, new_new_n32697__, new_new_n32698__,
    new_new_n32699__, new_new_n32700__, new_new_n32701__, new_new_n32702__,
    new_new_n32703__, new_new_n32704__, new_new_n32705__, new_new_n32706__,
    new_new_n32707__, new_new_n32708__, new_new_n32709__, new_new_n32710__,
    new_new_n32711__, new_new_n32712__, new_new_n32713__, new_new_n32714__,
    new_new_n32715__, new_new_n32716__, new_new_n32717__, new_new_n32718__,
    new_new_n32719__, new_new_n32720__, new_new_n32721__, new_new_n32722__,
    new_new_n32723__, new_new_n32724__, new_new_n32725__, new_new_n32726__,
    new_new_n32727__, new_new_n32728__, new_new_n32729__, new_new_n32730__,
    new_new_n32731__, new_new_n32732__, new_new_n32733__, new_new_n32734__,
    new_new_n32735__, new_new_n32736__, new_new_n32737__, new_new_n32738__,
    new_new_n32739__, new_new_n32740__, new_new_n32741__, new_new_n32742__,
    new_new_n32743__, new_new_n32744__, new_new_n32745__, new_new_n32746__,
    new_new_n32747__, new_new_n32748__, new_new_n32749__, new_new_n32750__,
    new_new_n32751__, new_new_n32752__, new_new_n32753__, new_new_n32754__,
    new_new_n32755__, new_new_n32756__, new_new_n32757__, new_new_n32758__,
    new_new_n32759__, new_new_n32760__, new_new_n32761__, new_new_n32762__,
    new_new_n32763__, new_new_n32764__, new_new_n32765__, new_new_n32766__,
    new_new_n32767__, new_new_n32768__, new_new_n32769__, new_new_n32770__,
    new_new_n32771__, new_new_n32772__, new_new_n32773__, new_new_n32774__,
    new_new_n32775__, new_new_n32776__, new_new_n32777__, new_new_n32778__,
    new_new_n32779__, new_new_n32780__, new_new_n32781__, new_new_n32782__,
    new_new_n32783__, new_new_n32784__, new_new_n32785__, new_new_n32786__,
    new_new_n32787__, new_new_n32788__, new_new_n32789__, new_new_n32790__,
    new_new_n32791__, new_new_n32792__, new_new_n32793__, new_new_n32794__,
    new_new_n32795__, new_new_n32796__, new_new_n32797__, new_new_n32798__,
    new_new_n32799__, new_new_n32800__, new_new_n32801__, new_new_n32802__,
    new_new_n32803__, new_new_n32804__, new_new_n32805__, new_new_n32806__,
    new_new_n32807__, new_new_n32808__, new_new_n32809__, new_new_n32810__,
    new_new_n32811__, new_new_n32812__, new_new_n32813__, new_new_n32814__,
    new_new_n32815__, new_new_n32816__, new_new_n32817__, new_new_n32818__,
    new_new_n32819__, new_new_n32820__, new_new_n32821__, new_new_n32822__,
    new_new_n32823__, new_new_n32824__, new_new_n32825__, new_new_n32826__,
    new_new_n32827__, new_new_n32828__, new_new_n32829__, new_new_n32830__,
    new_new_n32831__, new_new_n32832__, new_new_n32833__, new_new_n32834__,
    new_new_n32835__, new_new_n32836__, new_new_n32837__, new_new_n32838__,
    new_new_n32839__, new_new_n32840__, new_new_n32841__, new_new_n32842__,
    new_new_n32843__, new_new_n32844__, new_new_n32845__, new_new_n32846__,
    new_new_n32847__, new_new_n32848__, new_new_n32849__, new_new_n32850__,
    new_new_n32851__, new_new_n32852__, new_new_n32853__, new_new_n32854__,
    new_new_n32855__, new_new_n32856__, new_new_n32857__, new_new_n32858__,
    new_new_n32859__, new_new_n32860__, new_new_n32861__, new_new_n32862__,
    new_new_n32863__, new_new_n32864__, new_new_n32865__, new_new_n32866__,
    new_new_n32867__, new_new_n32868__, new_new_n32869__, new_new_n32870__,
    new_new_n32871__, new_new_n32872__, new_new_n32873__, new_new_n32874__,
    new_new_n32875__, new_new_n32876__, new_new_n32877__, new_new_n32878__,
    new_new_n32879__, new_new_n32880__, new_new_n32881__, new_new_n32882__,
    new_new_n32883__, new_new_n32884__, new_new_n32885__, new_new_n32886__,
    new_new_n32887__, new_new_n32888__, new_new_n32889__, new_new_n32890__,
    new_new_n32891__, new_new_n32892__, new_new_n32893__, new_new_n32895__,
    new_new_n32896__, new_new_n32897__, new_new_n32898__, new_new_n32899__,
    new_new_n32900__, new_new_n32901__, new_new_n32902__, new_new_n32903__,
    new_new_n32904__, new_new_n32905__, new_new_n32906__, new_new_n32907__,
    new_new_n32908__, new_new_n32909__, new_new_n32910__, new_new_n32911__,
    new_new_n32912__, new_new_n32913__, new_new_n32914__, new_new_n32915__,
    new_new_n32916__, new_new_n32917__, new_new_n32918__, new_new_n32919__,
    new_new_n32920__, new_new_n32921__, new_new_n32922__, new_new_n32923__,
    new_new_n32924__, new_new_n32925__, new_new_n32926__, new_new_n32927__,
    new_new_n32928__, new_new_n32929__, new_new_n32930__, new_new_n32931__,
    new_new_n32932__, new_new_n32933__, new_new_n32934__, new_new_n32935__,
    new_new_n32936__, new_new_n32937__, new_new_n32938__, new_new_n32939__,
    new_new_n32940__, new_new_n32941__, new_new_n32942__, new_new_n32943__,
    new_new_n32944__, new_new_n32945__, new_new_n32946__, new_new_n32947__,
    new_new_n32948__, new_new_n32949__, new_new_n32950__, new_new_n32951__,
    new_new_n32952__, new_new_n32953__, new_new_n32954__, new_new_n32955__,
    new_new_n32956__, new_new_n32957__, new_new_n32958__, new_new_n32959__,
    new_new_n32960__, new_new_n32961__, new_new_n32962__, new_new_n32963__,
    new_new_n32964__, new_new_n32965__, new_new_n32966__, new_new_n32967__,
    new_new_n32968__, new_new_n32969__, new_new_n32970__, new_new_n32971__,
    new_new_n32972__, new_new_n32973__, new_new_n32974__, new_new_n32975__,
    new_new_n32976__, new_new_n32977__, new_new_n32978__, new_new_n32979__,
    new_new_n32980__, new_new_n32981__, new_new_n32982__, new_new_n32983__,
    new_new_n32984__, new_new_n32985__, new_new_n32986__, new_new_n32987__,
    new_new_n32988__, new_new_n32989__, new_new_n32990__, new_new_n32991__,
    new_new_n32992__, new_new_n32993__, new_new_n32994__, new_new_n32995__,
    new_new_n32996__, new_new_n32997__, new_new_n32998__, new_new_n32999__,
    new_new_n33000__, new_new_n33001__, new_new_n33002__, new_new_n33003__,
    new_new_n33004__, new_new_n33005__, new_new_n33006__, new_new_n33007__,
    new_new_n33008__, new_new_n33009__, new_new_n33010__, new_new_n33011__,
    new_new_n33012__, new_new_n33013__, new_new_n33014__, new_new_n33015__,
    new_new_n33016__, new_new_n33017__, new_new_n33018__, new_new_n33019__,
    new_new_n33020__, new_new_n33021__, new_new_n33022__, new_new_n33023__,
    new_new_n33024__, new_new_n33025__, new_new_n33026__, new_new_n33027__,
    new_new_n33028__, new_new_n33029__, new_new_n33030__, new_new_n33031__,
    new_new_n33032__, new_new_n33033__, new_new_n33034__, new_new_n33035__,
    new_new_n33036__, new_new_n33037__, new_new_n33038__, new_new_n33039__,
    new_new_n33040__, new_new_n33041__, new_new_n33042__, new_new_n33043__,
    new_new_n33044__, new_new_n33045__, new_new_n33046__, new_new_n33047__,
    new_new_n33048__, new_new_n33049__, new_new_n33050__, new_new_n33051__,
    new_new_n33052__, new_new_n33053__, new_new_n33054__, new_new_n33055__,
    new_new_n33056__, new_new_n33057__, new_new_n33058__, new_new_n33059__,
    new_new_n33060__, new_new_n33061__, new_new_n33062__, new_new_n33063__,
    new_new_n33064__, new_new_n33065__, new_new_n33066__, new_new_n33067__,
    new_new_n33068__, new_new_n33069__, new_new_n33070__, new_new_n33071__,
    new_new_n33072__, new_new_n33073__, new_new_n33074__, new_new_n33075__,
    new_new_n33076__, new_new_n33077__, new_new_n33078__, new_new_n33079__,
    new_new_n33080__, new_new_n33081__, new_new_n33082__, new_new_n33083__,
    new_new_n33084__, new_new_n33085__, new_new_n33086__, new_new_n33087__,
    new_new_n33088__, new_new_n33089__, new_new_n33090__, new_new_n33091__,
    new_new_n33092__, new_new_n33093__, new_new_n33094__, new_new_n33095__,
    new_new_n33096__, new_new_n33097__, new_new_n33098__, new_new_n33099__,
    new_new_n33100__, new_new_n33101__, new_new_n33102__, new_new_n33103__,
    new_new_n33104__, new_new_n33105__, new_new_n33106__, new_new_n33107__,
    new_new_n33108__, new_new_n33109__, new_new_n33110__, new_new_n33111__,
    new_new_n33112__, new_new_n33113__, new_new_n33114__, new_new_n33115__,
    new_new_n33116__, new_new_n33117__, new_new_n33118__, new_new_n33119__,
    new_new_n33120__, new_new_n33121__, new_new_n33122__, new_new_n33123__,
    new_new_n33124__, new_new_n33125__, new_new_n33126__, new_new_n33127__,
    new_new_n33128__, new_new_n33129__, new_new_n33130__, new_new_n33131__,
    new_new_n33132__, new_new_n33133__, new_new_n33134__, new_new_n33135__,
    new_new_n33136__, new_new_n33137__, new_new_n33138__, new_new_n33139__,
    new_new_n33140__, new_new_n33141__, new_new_n33142__, new_new_n33143__,
    new_new_n33144__, new_new_n33145__, new_new_n33146__, new_new_n33147__,
    new_new_n33148__, new_new_n33149__, new_new_n33150__, new_new_n33151__,
    new_new_n33152__, new_new_n33153__, new_new_n33154__, new_new_n33155__,
    new_new_n33156__, new_new_n33157__, new_new_n33158__, new_new_n33159__,
    new_new_n33160__, new_new_n33161__, new_new_n33162__, new_new_n33163__,
    new_new_n33164__, new_new_n33165__, new_new_n33166__, new_new_n33167__,
    new_new_n33168__, new_new_n33169__, new_new_n33170__, new_new_n33171__,
    new_new_n33172__, new_new_n33173__, new_new_n33174__, new_new_n33175__,
    new_new_n33176__, new_new_n33177__, new_new_n33178__, new_new_n33179__,
    new_new_n33180__, new_new_n33181__, new_new_n33182__, new_new_n33183__,
    new_new_n33184__, new_new_n33185__, new_new_n33186__, new_new_n33187__,
    new_new_n33188__, new_new_n33189__, new_new_n33190__, new_new_n33191__,
    new_new_n33192__, new_new_n33193__, new_new_n33194__, new_new_n33195__,
    new_new_n33196__, new_new_n33197__, new_new_n33198__, new_new_n33199__,
    new_new_n33200__, new_new_n33201__, new_new_n33202__, new_new_n33203__,
    new_new_n33204__, new_new_n33205__, new_new_n33206__, new_new_n33207__,
    new_new_n33208__, new_new_n33209__, new_new_n33210__, new_new_n33211__,
    new_new_n33212__, new_new_n33213__, new_new_n33214__, new_new_n33215__,
    new_new_n33216__, new_new_n33217__, new_new_n33218__, new_new_n33219__,
    new_new_n33220__, new_new_n33222__, new_new_n33223__, new_new_n33224__,
    new_new_n33225__, new_new_n33226__, new_new_n33227__, new_new_n33228__,
    new_new_n33229__, new_new_n33230__, new_new_n33231__, new_new_n33232__,
    new_new_n33233__, new_new_n33234__, new_new_n33235__, new_new_n33236__,
    new_new_n33237__, new_new_n33238__, new_new_n33239__, new_new_n33240__,
    new_new_n33241__, new_new_n33242__, new_new_n33243__, new_new_n33244__,
    new_new_n33245__, new_new_n33246__, new_new_n33247__, new_new_n33248__,
    new_new_n33249__, new_new_n33250__, new_new_n33251__, new_new_n33252__,
    new_new_n33253__, new_new_n33254__, new_new_n33255__, new_new_n33256__,
    new_new_n33257__, new_new_n33258__, new_new_n33259__, new_new_n33260__,
    new_new_n33261__, new_new_n33262__, new_new_n33263__, new_new_n33264__,
    new_new_n33265__, new_new_n33266__, new_new_n33267__, new_new_n33268__,
    new_new_n33269__, new_new_n33270__, new_new_n33271__, new_new_n33272__,
    new_new_n33273__, new_new_n33274__, new_new_n33275__, new_new_n33276__,
    new_new_n33277__, new_new_n33278__, new_new_n33279__, new_new_n33280__,
    new_new_n33281__, new_new_n33282__, new_new_n33283__, new_new_n33284__,
    new_new_n33285__, new_new_n33286__, new_new_n33287__, new_new_n33288__,
    new_new_n33289__, new_new_n33290__, new_new_n33291__, new_new_n33292__,
    new_new_n33293__, new_new_n33294__, new_new_n33295__, new_new_n33296__,
    new_new_n33297__, new_new_n33298__, new_new_n33299__, new_new_n33300__,
    new_new_n33301__, new_new_n33302__, new_new_n33303__, new_new_n33304__,
    new_new_n33305__, new_new_n33306__, new_new_n33307__, new_new_n33308__,
    new_new_n33309__, new_new_n33310__, new_new_n33311__, new_new_n33312__,
    new_new_n33313__, new_new_n33314__, new_new_n33315__, new_new_n33316__,
    new_new_n33317__, new_new_n33318__, new_new_n33319__, new_new_n33320__,
    new_new_n33321__, new_new_n33322__, new_new_n33323__, new_new_n33324__,
    new_new_n33325__, new_new_n33326__, new_new_n33327__, new_new_n33328__,
    new_new_n33329__, new_new_n33330__, new_new_n33331__, new_new_n33332__,
    new_new_n33333__, new_new_n33334__, new_new_n33335__, new_new_n33336__,
    new_new_n33337__, new_new_n33338__, new_new_n33339__, new_new_n33340__,
    new_new_n33341__, new_new_n33342__, new_new_n33343__, new_new_n33344__,
    new_new_n33345__, new_new_n33346__, new_new_n33347__, new_new_n33348__,
    new_new_n33349__, new_new_n33350__, new_new_n33351__, new_new_n33352__,
    new_new_n33353__, new_new_n33354__, new_new_n33355__, new_new_n33356__,
    new_new_n33357__, new_new_n33358__, new_new_n33359__, new_new_n33360__,
    new_new_n33361__, new_new_n33362__, new_new_n33363__, new_new_n33364__,
    new_new_n33365__, new_new_n33366__, new_new_n33367__, new_new_n33368__,
    new_new_n33369__, new_new_n33370__, new_new_n33371__, new_new_n33372__,
    new_new_n33373__, new_new_n33374__, new_new_n33375__, new_new_n33376__,
    new_new_n33377__, new_new_n33378__, new_new_n33379__, new_new_n33380__,
    new_new_n33381__, new_new_n33382__, new_new_n33383__, new_new_n33384__,
    new_new_n33385__, new_new_n33386__, new_new_n33387__, new_new_n33388__,
    new_new_n33389__, new_new_n33390__, new_new_n33391__, new_new_n33392__,
    new_new_n33393__, new_new_n33394__, new_new_n33395__, new_new_n33396__,
    new_new_n33397__, new_new_n33398__, new_new_n33399__, new_new_n33400__,
    new_new_n33401__, new_new_n33402__, new_new_n33403__, new_new_n33404__,
    new_new_n33405__, new_new_n33406__, new_new_n33407__, new_new_n33408__,
    new_new_n33409__, new_new_n33410__, new_new_n33411__, new_new_n33412__,
    new_new_n33413__, new_new_n33414__, new_new_n33415__, new_new_n33416__,
    new_new_n33417__, new_new_n33418__, new_new_n33419__, new_new_n33420__,
    new_new_n33421__, new_new_n33422__, new_new_n33423__, new_new_n33424__,
    new_new_n33425__, new_new_n33426__, new_new_n33427__, new_new_n33428__,
    new_new_n33429__, new_new_n33430__, new_new_n33431__, new_new_n33432__,
    new_new_n33433__, new_new_n33434__, new_new_n33435__, new_new_n33436__,
    new_new_n33437__, new_new_n33438__, new_new_n33439__, new_new_n33440__,
    new_new_n33441__, new_new_n33442__, new_new_n33443__, new_new_n33444__,
    new_new_n33445__, new_new_n33446__, new_new_n33447__, new_new_n33448__,
    new_new_n33449__, new_new_n33450__, new_new_n33451__, new_new_n33452__,
    new_new_n33453__, new_new_n33454__, new_new_n33455__, new_new_n33456__,
    new_new_n33457__, new_new_n33458__, new_new_n33459__, new_new_n33460__,
    new_new_n33461__, new_new_n33462__, new_new_n33463__, new_new_n33464__,
    new_new_n33465__, new_new_n33466__, new_new_n33467__, new_new_n33468__,
    new_new_n33469__, new_new_n33470__, new_new_n33471__, new_new_n33472__,
    new_new_n33473__, new_new_n33474__, new_new_n33475__, new_new_n33476__,
    new_new_n33477__, new_new_n33478__, new_new_n33479__, new_new_n33480__,
    new_new_n33481__, new_new_n33482__, new_new_n33483__, new_new_n33484__,
    new_new_n33485__, new_new_n33486__, new_new_n33487__, new_new_n33488__,
    new_new_n33489__, new_new_n33490__, new_new_n33491__, new_new_n33492__,
    new_new_n33493__, new_new_n33494__, new_new_n33495__, new_new_n33496__,
    new_new_n33497__, new_new_n33498__, new_new_n33499__, new_new_n33500__,
    new_new_n33501__, new_new_n33502__, new_new_n33503__, new_new_n33504__,
    new_new_n33505__, new_new_n33506__, new_new_n33507__, new_new_n33508__,
    new_new_n33509__, new_new_n33510__, new_new_n33511__, new_new_n33512__,
    new_new_n33513__, new_new_n33514__, new_new_n33515__, new_new_n33516__,
    new_new_n33517__, new_new_n33518__, new_new_n33519__, new_new_n33520__,
    new_new_n33521__, new_new_n33522__, new_new_n33523__, new_new_n33524__,
    new_new_n33525__, new_new_n33526__, new_new_n33527__, new_new_n33528__,
    new_new_n33529__, new_new_n33530__, new_new_n33531__, new_new_n33532__,
    new_new_n33533__, new_new_n33534__, new_new_n33535__, new_new_n33536__,
    new_new_n33537__, new_new_n33538__, new_new_n33539__, new_new_n33540__,
    new_new_n33541__, new_new_n33542__, new_new_n33543__, new_new_n33544__,
    new_new_n33545__, new_new_n33546__, new_new_n33547__, new_new_n33548__,
    new_new_n33549__, new_new_n33550__, new_new_n33551__, new_new_n33553__,
    new_new_n33554__, new_new_n33555__, new_new_n33556__, new_new_n33557__,
    new_new_n33558__, new_new_n33559__, new_new_n33560__, new_new_n33561__,
    new_new_n33562__, new_new_n33563__, new_new_n33565__, new_new_n33566__,
    new_new_n33567__, new_new_n33568__, new_new_n33569__, new_new_n33570__,
    new_new_n33571__, new_new_n33572__, new_new_n33573__, new_new_n33574__,
    new_new_n33575__, new_new_n33576__, new_new_n33577__, new_new_n33578__,
    new_new_n33579__, new_new_n33581__, new_new_n33582__, new_new_n33583__,
    new_new_n33584__, new_new_n33585__, new_new_n33587__, new_new_n33588__,
    new_new_n33590__, new_new_n33591__, new_new_n33593__, new_new_n33594__,
    new_new_n33595__, new_new_n33596__, new_new_n33597__, new_new_n33598__,
    new_new_n33600__, new_new_n33601__, new_new_n33603__, new_new_n33604__,
    new_new_n33606__, new_new_n33607__, new_new_n33609__, new_new_n33610__,
    new_new_n33612__, new_new_n33613__, new_new_n33615__, new_new_n33616__,
    new_new_n33618__, new_new_n33619__, new_new_n33621__, new_new_n33622__,
    new_new_n33624__, new_new_n33625__, new_new_n33627__, new_new_n33628__,
    new_new_n33630__, new_new_n33631__, new_new_n33633__, new_new_n33634__,
    new_new_n33636__, new_new_n33637__, new_new_n33639__, new_new_n33640__,
    new_new_n33642__, new_new_n33643__, new_new_n33645__, new_new_n33646__,
    new_new_n33648__, new_new_n33649__, new_new_n33651__, new_new_n33652__,
    new_new_n33654__, new_new_n33655__, new_new_n33657__, new_new_n33658__,
    new_new_n33660__, new_new_n33661__, new_new_n33663__, new_new_n33664__,
    new_new_n33666__, new_new_n33667__, new_new_n33669__, new_new_n33670__,
    new_new_n33672__, new_new_n33673__, new_new_n33675__, new_new_n33676__,
    new_new_n33678__, new_new_n33679__, new_new_n33681__, new_new_n33682__,
    new_new_n33684__, new_new_n33685__, new_new_n33687__, new_new_n33688__,
    new_new_n33690__, new_new_n33691__, new_new_n33693__, new_new_n33694__,
    new_new_n33695__, new_new_n33697__, new_new_n33698__, new_new_n33700__,
    new_new_n33701__, new_new_n33703__, new_new_n33704__, new_new_n33706__,
    new_new_n33707__, new_new_n33709__, new_new_n33710__, new_new_n33712__,
    new_new_n33713__, new_new_n33715__, new_new_n33716__, new_new_n33718__,
    new_new_n33719__, new_new_n33721__, new_new_n33722__, new_new_n33724__,
    new_new_n33725__, new_new_n33727__, new_new_n33728__, new_new_n33730__,
    new_new_n33731__, new_new_n33733__, new_new_n33734__, new_new_n33736__,
    new_new_n33737__, new_new_n33739__, new_new_n33740__, new_new_n33742__,
    new_new_n33743__, new_new_n33745__, new_new_n33746__, new_new_n33748__,
    new_new_n33749__, new_new_n33751__, new_new_n33752__, new_new_n33754__,
    new_new_n33755__, new_new_n33757__, new_new_n33758__, new_new_n33760__,
    new_new_n33761__, new_new_n33763__, new_new_n33764__, new_new_n33766__,
    new_new_n33767__, new_new_n33769__, new_new_n33770__, new_new_n33772__,
    new_new_n33773__, new_new_n33775__, new_new_n33776__, new_new_n33778__,
    new_new_n33779__, new_new_n33781__, new_new_n33782__, new_new_n33784__,
    new_new_n33785__, new_new_n33787__, new_new_n33788__, new_new_n33791__,
    new_new_n33792__, new_new_n33796__, new_new_n33797__, new_new_n33799__,
    new_new_n33800__, new_new_n33802__, new_new_n33803__, new_new_n33805__,
    new_new_n33806__, new_new_n33807__, new_new_n33809__, new_new_n33810__,
    new_new_n33811__, new_new_n33812__, new_new_n33813__, new_new_n33815__,
    new_new_n33816__, new_new_n33817__, new_new_n33819__, new_new_n33820__,
    new_new_n33821__, new_new_n33823__, new_new_n33824__, new_new_n33825__,
    new_new_n33826__, new_new_n33828__, new_new_n33829__, new_new_n33831__,
    new_new_n33832__, new_new_n33834__, new_new_n33835__, new_new_n33837__,
    new_new_n33838__, new_new_n33839__, new_new_n33841__, new_new_n33842__,
    new_new_n33844__, new_new_n33845__, new_new_n33847__, new_new_n33848__,
    new_new_n33850__, new_new_n33851__, new_new_n33852__, new_new_n33854__,
    new_new_n33855__, new_new_n33857__, new_new_n33858__, new_new_n33860__,
    new_new_n33861__, new_new_n33863__, new_new_n33864__, new_new_n33865__,
    new_new_n33867__, new_new_n33869__, new_new_n33871__, new_new_n33873__,
    new_new_n33875__, new_new_n33877__, new_new_n33879__, new_new_n33881__,
    new_new_n33883__, new_new_n33885__, new_new_n33887__, new_new_n33889__,
    new_new_n33891__, new_new_n33893__, new_new_n33895__, new_new_n33897__,
    new_new_n33898__, new_new_n33900__, new_new_n33901__, new_new_n33902__,
    new_new_n33903__, new_new_n33904__, new_new_n33906__, new_new_n33907__,
    new_new_n33908__, new_new_n33909__, new_new_n33910__, new_new_n33911__,
    new_new_n33912__, new_new_n33913__, new_new_n33914__, new_new_n33915__,
    new_new_n33916__, new_new_n33917__, new_new_n33918__, new_new_n33919__,
    new_new_n33921__, new_new_n33922__, new_new_n33923__, new_new_n33924__,
    new_new_n33925__, new_new_n33926__, new_new_n33927__, new_new_n33928__,
    new_new_n33929__, new_new_n33930__, new_new_n33931__, new_new_n33932__,
    new_new_n33933__, new_new_n33934__, new_new_n33935__, new_new_n33936__,
    new_new_n33937__, new_new_n33938__, new_new_n33939__, new_new_n33940__,
    new_new_n33941__, new_new_n33942__, new_new_n33944__, new_new_n33945__,
    new_new_n33946__, new_new_n33947__, new_new_n33948__, new_new_n33950__,
    new_new_n33951__, new_new_n33952__, new_new_n33953__, new_new_n33954__,
    new_new_n33955__, new_new_n33956__, new_new_n33957__, new_new_n33958__,
    new_new_n33959__, new_new_n33960__, new_new_n33961__, new_new_n33962__,
    new_new_n33963__, new_new_n33964__, new_new_n33965__, new_new_n33966__,
    new_new_n33967__, new_new_n33968__, new_new_n33970__, new_new_n33971__,
    new_new_n33972__, new_new_n33973__, new_new_n33974__, new_new_n33975__,
    new_new_n33976__, new_new_n33978__, new_new_n33979__, new_new_n33980__,
    new_new_n33981__, new_new_n33982__, new_new_n33983__, new_new_n33984__,
    new_new_n33985__, new_new_n33986__, new_new_n33987__, new_new_n33988__,
    new_new_n33989__, new_new_n33990__, new_new_n33991__, new_new_n33992__,
    new_new_n33993__, new_new_n33994__, new_new_n33995__, new_new_n33996__,
    new_new_n33997__, new_new_n33999__, new_new_n34000__, new_new_n34001__,
    new_new_n34002__, new_new_n34003__, new_new_n34004__, new_new_n34005__,
    new_new_n34007__, new_new_n34008__, new_new_n34009__, new_new_n34010__,
    new_new_n34011__, new_new_n34012__, new_new_n34013__, new_new_n34014__,
    new_new_n34015__, new_new_n34016__, new_new_n34017__, new_new_n34018__,
    new_new_n34019__, new_new_n34020__, new_new_n34021__, new_new_n34022__,
    new_new_n34023__, new_new_n34024__, new_new_n34025__, new_new_n34026__,
    new_new_n34027__, new_new_n34028__, new_new_n34030__, new_new_n34031__,
    new_new_n34032__, new_new_n34033__, new_new_n34034__, new_new_n34035__,
    new_new_n34037__, new_new_n34038__, new_new_n34039__, new_new_n34040__,
    new_new_n34041__, new_new_n34042__, new_new_n34043__, new_new_n34044__,
    new_new_n34045__, new_new_n34046__, new_new_n34047__, new_new_n34048__,
    new_new_n34049__, new_new_n34050__, new_new_n34051__, new_new_n34052__,
    new_new_n34053__, new_new_n34054__, new_new_n34055__, new_new_n34056__,
    new_new_n34058__, new_new_n34059__, new_new_n34060__, new_new_n34061__,
    new_new_n34062__, new_new_n34063__, new_new_n34065__, new_new_n34066__,
    new_new_n34067__, new_new_n34068__, new_new_n34069__, new_new_n34070__,
    new_new_n34071__, new_new_n34072__, new_new_n34073__, new_new_n34074__,
    new_new_n34075__, new_new_n34076__, new_new_n34077__, new_new_n34078__,
    new_new_n34079__, new_new_n34080__, new_new_n34081__, new_new_n34082__,
    new_new_n34083__, new_new_n34084__, new_new_n34086__, new_new_n34087__,
    new_new_n34088__, new_new_n34089__, new_new_n34090__, new_new_n34091__,
    new_new_n34092__, new_new_n34093__, new_new_n34094__, new_new_n34095__,
    new_new_n34096__, new_new_n34097__, new_new_n34098__, new_new_n34100__,
    new_new_n34101__, new_new_n34102__, new_new_n34103__, new_new_n34104__,
    new_new_n34105__, new_new_n34106__, new_new_n34107__, new_new_n34108__,
    new_new_n34109__, new_new_n34110__, new_new_n34111__, new_new_n34112__,
    new_new_n34113__, new_new_n34114__, new_new_n34115__, new_new_n34116__,
    new_new_n34118__, new_new_n34119__, new_new_n34120__, new_new_n34121__,
    new_new_n34122__, new_new_n34123__, new_new_n34124__, new_new_n34125__,
    new_new_n34126__, new_new_n34127__, new_new_n34128__, new_new_n34129__,
    new_new_n34130__, new_new_n34131__, new_new_n34132__, new_new_n34133__,
    new_new_n34134__, new_new_n34135__, new_new_n34136__, new_new_n34137__,
    new_new_n34138__, new_new_n34139__, new_new_n34141__, new_new_n34142__,
    new_new_n34143__, new_new_n34144__, new_new_n34145__, new_new_n34146__,
    new_new_n34147__, new_new_n34148__, new_new_n34149__, new_new_n34150__,
    new_new_n34151__, new_new_n34152__, new_new_n34153__, new_new_n34154__,
    new_new_n34156__, new_new_n34157__, new_new_n34158__, new_new_n34159__,
    new_new_n34160__, new_new_n34161__, new_new_n34162__, new_new_n34163__,
    new_new_n34164__, new_new_n34165__, new_new_n34166__, new_new_n34167__,
    new_new_n34168__, new_new_n34169__, new_new_n34171__, new_new_n34172__,
    new_new_n34173__, new_new_n34174__, new_new_n34175__, new_new_n34176__,
    new_new_n34177__, new_new_n34178__, new_new_n34179__, new_new_n34180__,
    new_new_n34181__, new_new_n34182__, new_new_n34183__, new_new_n34184__,
    new_new_n34186__, new_new_n34187__, new_new_n34188__, new_new_n34189__,
    new_new_n34190__, new_new_n34191__, new_new_n34192__, new_new_n34193__,
    new_new_n34194__, new_new_n34195__, new_new_n34196__, new_new_n34197__,
    new_new_n34198__, new_new_n34199__, new_new_n34200__, new_new_n34201__,
    new_new_n34202__, new_new_n34204__, new_new_n34205__, new_new_n34206__,
    new_new_n34207__, new_new_n34208__, new_new_n34209__, new_new_n34210__,
    new_new_n34211__, new_new_n34212__, new_new_n34213__, new_new_n34214__,
    new_new_n34215__, new_new_n34216__, new_new_n34217__, new_new_n34219__,
    new_new_n34220__, new_new_n34221__, new_new_n34222__, new_new_n34223__,
    new_new_n34224__, new_new_n34225__, new_new_n34226__, new_new_n34227__,
    new_new_n34228__, new_new_n34229__, new_new_n34230__, new_new_n34231__,
    new_new_n34232__, new_new_n34233__, new_new_n34234__, new_new_n34236__,
    new_new_n34237__, new_new_n34238__, new_new_n34239__, new_new_n34240__,
    new_new_n34241__, new_new_n34242__, new_new_n34243__, new_new_n34244__,
    new_new_n34245__, new_new_n34246__, new_new_n34247__, new_new_n34248__,
    new_new_n34249__, new_new_n34250__, new_new_n34251__, new_new_n34253__,
    new_new_n34254__, new_new_n34255__, new_new_n34256__, new_new_n34257__,
    new_new_n34258__, new_new_n34259__, new_new_n34260__, new_new_n34261__,
    new_new_n34262__, new_new_n34263__, new_new_n34264__, new_new_n34266__,
    new_new_n34267__, new_new_n34268__, new_new_n34269__, new_new_n34270__,
    new_new_n34271__, new_new_n34272__, new_new_n34273__, new_new_n34274__,
    new_new_n34276__, new_new_n34277__, new_new_n34278__, new_new_n34279__,
    new_new_n34280__, new_new_n34281__, new_new_n34282__, new_new_n34283__,
    new_new_n34284__, new_new_n34285__, new_new_n34286__, new_new_n34288__,
    new_new_n34289__, new_new_n34290__, new_new_n34291__, new_new_n34292__,
    new_new_n34293__, new_new_n34294__, new_new_n34295__, new_new_n34296__,
    new_new_n34297__, new_new_n34298__, new_new_n34300__, new_new_n34301__,
    new_new_n34302__, new_new_n34303__, new_new_n34304__, new_new_n34305__,
    new_new_n34306__, new_new_n34307__, new_new_n34308__, new_new_n34310__,
    new_new_n34311__, new_new_n34312__, new_new_n34313__, new_new_n34314__,
    new_new_n34315__, new_new_n34316__, new_new_n34317__, new_new_n34318__,
    new_new_n34320__, new_new_n34321__, new_new_n34322__, new_new_n34323__,
    new_new_n34324__, new_new_n34325__, new_new_n34326__, new_new_n34327__,
    new_new_n34328__, new_new_n34329__, new_new_n34330__, new_new_n34331__,
    new_new_n34332__, new_new_n34334__, new_new_n34335__, new_new_n34336__,
    new_new_n34337__, new_new_n34338__, new_new_n34339__, new_new_n34340__,
    new_new_n34341__, new_new_n34342__, new_new_n34344__, new_new_n34345__,
    new_new_n34346__, new_new_n34347__, new_new_n34348__, new_new_n34349__,
    new_new_n34350__, new_new_n34351__, new_new_n34352__, new_new_n34354__,
    new_new_n34355__, new_new_n34356__, new_new_n34357__, new_new_n34358__,
    new_new_n34359__, new_new_n34360__, new_new_n34361__, new_new_n34362__,
    new_new_n34364__, new_new_n34365__, new_new_n34366__, new_new_n34367__,
    new_new_n34368__, new_new_n34369__, new_new_n34370__, new_new_n34371__,
    new_new_n34372__, new_new_n34374__, new_new_n34375__, new_new_n34376__,
    new_new_n34377__, new_new_n34378__, new_new_n34379__, new_new_n34380__,
    new_new_n34381__, new_new_n34382__, new_new_n34384__, new_new_n34385__,
    new_new_n34386__, new_new_n34387__, new_new_n34388__, new_new_n34389__,
    new_new_n34390__, new_new_n34391__, new_new_n34392__, new_new_n34393__,
    new_new_n34394__, new_new_n34395__, new_new_n34396__, new_new_n34397__,
    new_new_n34399__, new_new_n34400__, new_new_n34401__, new_new_n34402__,
    new_new_n34403__, new_new_n34404__, new_new_n34405__, new_new_n34406__,
    new_new_n34407__, new_new_n34408__, new_new_n34409__, new_new_n34410__,
    new_new_n34411__, new_new_n34412__, new_new_n34413__, new_new_n34414__,
    new_new_n34416__, new_new_n34417__, new_new_n34418__, new_new_n34419__,
    new_new_n34420__, new_new_n34421__, new_new_n34422__, new_new_n34423__,
    new_new_n34424__, new_new_n34425__, new_new_n34426__, new_new_n34427__,
    new_new_n34428__, new_new_n34429__, new_new_n34431__, new_new_n34432__,
    new_new_n34433__, new_new_n34434__, new_new_n34435__, new_new_n34436__,
    new_new_n34437__, new_new_n34438__, new_new_n34439__, new_new_n34440__,
    new_new_n34441__, new_new_n34442__, new_new_n34443__, new_new_n34444__,
    new_new_n34445__, new_new_n34446__, new_new_n34447__, new_new_n34449__,
    new_new_n34450__, new_new_n34451__, new_new_n34452__, new_new_n34453__,
    new_new_n34454__, new_new_n34455__, new_new_n34457__, new_new_n34458__,
    new_new_n34460__, new_new_n34461__, new_new_n34463__, new_new_n34464__,
    new_new_n34466__, new_new_n34467__, new_new_n34469__, new_new_n34470__,
    new_new_n34472__, new_new_n34473__, new_new_n34475__, new_new_n34476__,
    new_new_n34478__, new_new_n34479__, new_new_n34481__, new_new_n34482__,
    new_new_n34484__, new_new_n34485__, new_new_n34487__, new_new_n34488__,
    new_new_n34490__, new_new_n34491__, new_new_n34493__, new_new_n34494__,
    new_new_n34496__, new_new_n34497__, new_new_n34499__, new_new_n34500__,
    new_new_n34502__, new_new_n34503__, new_new_n34505__, new_new_n34506__,
    new_new_n34508__, new_new_n34509__, new_new_n34511__, new_new_n34512__,
    new_new_n34514__, new_new_n34515__, new_new_n34517__, new_new_n34518__,
    new_new_n34520__, new_new_n34521__, new_new_n34523__, new_new_n34524__,
    new_new_n34526__, new_new_n34527__, new_new_n34529__, new_new_n34530__,
    new_new_n34532__, new_new_n34533__, new_new_n34535__, new_new_n34536__,
    new_new_n34538__, new_new_n34539__, new_new_n34541__, new_new_n34542__,
    new_new_n34544__, new_new_n34545__, new_new_n34547__, new_new_n34548__,
    new_new_n34550__, new_new_n34551__, new_new_n34552__, new_new_n34553__,
    new_new_n34554__, new_new_n34555__, new_new_n34556__, new_new_n34557__,
    new_new_n34558__, new_new_n34559__, new_new_n34560__, new_new_n34561__,
    new_new_n34562__, new_new_n34563__, new_new_n34564__, new_new_n34565__,
    new_new_n34566__, new_new_n34567__, new_new_n34568__, new_new_n34569__,
    new_new_n34571__, new_new_n34572__, new_new_n34573__, new_new_n34574__,
    new_new_n34575__, new_new_n34576__, new_new_n34577__, new_new_n34578__,
    new_new_n34579__, new_new_n34580__, new_new_n34581__, new_new_n34582__,
    new_new_n34583__, new_new_n34584__, new_new_n34585__, new_new_n34586__,
    new_new_n34587__, new_new_n34588__, new_new_n34589__, new_new_n34590__,
    new_new_n34591__, new_new_n34592__, new_new_n34593__, new_new_n34595__,
    new_new_n34596__, new_new_n34597__, new_new_n34598__, new_new_n34599__,
    new_new_n34600__, new_new_n34601__, new_new_n34602__, new_new_n34603__,
    new_new_n34604__, new_new_n34605__, new_new_n34606__, new_new_n34607__,
    new_new_n34608__, new_new_n34609__, new_new_n34610__, new_new_n34611__,
    new_new_n34612__, new_new_n34613__, new_new_n34614__, new_new_n34615__,
    new_new_n34616__, new_new_n34617__, new_new_n34618__, new_new_n34619__,
    new_new_n34620__, new_new_n34621__, new_new_n34622__, new_new_n34624__,
    new_new_n34625__, new_new_n34626__, new_new_n34627__, new_new_n34628__,
    new_new_n34629__, new_new_n34630__, new_new_n34631__, new_new_n34632__,
    new_new_n34633__, new_new_n34634__, new_new_n34635__, new_new_n34636__,
    new_new_n34637__, new_new_n34638__, new_new_n34639__, new_new_n34640__,
    new_new_n34641__, new_new_n34642__, new_new_n34643__, new_new_n34644__,
    new_new_n34645__, new_new_n34646__, new_new_n34647__, new_new_n34648__,
    new_new_n34649__, new_new_n34650__, new_new_n34651__, new_new_n34653__,
    new_new_n34654__, new_new_n34655__, new_new_n34656__, new_new_n34657__,
    new_new_n34658__, new_new_n34659__, new_new_n34660__, new_new_n34661__,
    new_new_n34662__, new_new_n34663__, new_new_n34664__, new_new_n34665__,
    new_new_n34666__, new_new_n34667__, new_new_n34668__, new_new_n34669__,
    new_new_n34670__, new_new_n34671__, new_new_n34672__, new_new_n34673__,
    new_new_n34674__, new_new_n34675__, new_new_n34676__, new_new_n34677__,
    new_new_n34678__, new_new_n34679__, new_new_n34680__, new_new_n34682__,
    new_new_n34683__, new_new_n34684__, new_new_n34685__, new_new_n34686__,
    new_new_n34687__, new_new_n34688__, new_new_n34689__, new_new_n34690__,
    new_new_n34691__, new_new_n34692__, new_new_n34693__, new_new_n34694__,
    new_new_n34695__, new_new_n34696__, new_new_n34697__, new_new_n34698__,
    new_new_n34699__, new_new_n34700__, new_new_n34701__, new_new_n34702__,
    new_new_n34703__, new_new_n34704__, new_new_n34705__, new_new_n34706__,
    new_new_n34707__, new_new_n34708__, new_new_n34709__, new_new_n34711__,
    new_new_n34712__, new_new_n34713__, new_new_n34714__, new_new_n34715__,
    new_new_n34716__, new_new_n34717__, new_new_n34718__, new_new_n34719__,
    new_new_n34720__, new_new_n34721__, new_new_n34722__, new_new_n34723__,
    new_new_n34724__, new_new_n34725__, new_new_n34726__, new_new_n34727__,
    new_new_n34728__, new_new_n34729__, new_new_n34730__, new_new_n34731__,
    new_new_n34732__, new_new_n34733__, new_new_n34734__, new_new_n34735__,
    new_new_n34736__, new_new_n34737__, new_new_n34738__, new_new_n34740__,
    new_new_n34741__, new_new_n34742__, new_new_n34743__, new_new_n34744__,
    new_new_n34745__, new_new_n34746__, new_new_n34747__, new_new_n34748__,
    new_new_n34749__, new_new_n34750__, new_new_n34751__, new_new_n34752__,
    new_new_n34753__, new_new_n34754__, new_new_n34755__, new_new_n34756__,
    new_new_n34757__, new_new_n34758__, new_new_n34759__, new_new_n34760__,
    new_new_n34761__, new_new_n34762__, new_new_n34763__, new_new_n34764__,
    new_new_n34765__, new_new_n34766__, new_new_n34767__, new_new_n34769__,
    new_new_n34770__, new_new_n34771__, new_new_n34772__, new_new_n34773__,
    new_new_n34774__, new_new_n34775__, new_new_n34776__, new_new_n34777__,
    new_new_n34778__, new_new_n34779__, new_new_n34780__, new_new_n34781__,
    new_new_n34782__, new_new_n34783__, new_new_n34784__, new_new_n34785__,
    new_new_n34786__, new_new_n34787__, new_new_n34788__, new_new_n34789__,
    new_new_n34790__, new_new_n34791__, new_new_n34792__, new_new_n34793__,
    new_new_n34794__, new_new_n34795__, new_new_n34796__, new_new_n34798__,
    new_new_n34799__, new_new_n34800__, new_new_n34801__, new_new_n34802__,
    new_new_n34803__, new_new_n34804__, new_new_n34805__, new_new_n34806__,
    new_new_n34807__, new_new_n34808__, new_new_n34809__, new_new_n34810__,
    new_new_n34811__, new_new_n34812__, new_new_n34813__, new_new_n34814__,
    new_new_n34815__, new_new_n34816__, new_new_n34817__, new_new_n34818__,
    new_new_n34819__, new_new_n34820__, new_new_n34821__, new_new_n34822__,
    new_new_n34823__, new_new_n34825__, new_new_n34826__, new_new_n34827__,
    new_new_n34828__, new_new_n34829__, new_new_n34830__, new_new_n34831__,
    new_new_n34832__, new_new_n34833__, new_new_n34834__, new_new_n34835__,
    new_new_n34836__, new_new_n34837__, new_new_n34838__, new_new_n34839__,
    new_new_n34840__, new_new_n34841__, new_new_n34842__, new_new_n34843__,
    new_new_n34844__, new_new_n34845__, new_new_n34846__, new_new_n34847__,
    new_new_n34848__, new_new_n34849__, new_new_n34850__, new_new_n34851__,
    new_new_n34852__, new_new_n34854__, new_new_n34855__, new_new_n34856__,
    new_new_n34857__, new_new_n34858__, new_new_n34859__, new_new_n34860__,
    new_new_n34861__, new_new_n34862__, new_new_n34863__, new_new_n34864__,
    new_new_n34865__, new_new_n34866__, new_new_n34867__, new_new_n34868__,
    new_new_n34869__, new_new_n34870__, new_new_n34871__, new_new_n34872__,
    new_new_n34873__, new_new_n34874__, new_new_n34875__, new_new_n34876__,
    new_new_n34877__, new_new_n34878__, new_new_n34879__, new_new_n34880__,
    new_new_n34881__, new_new_n34882__, new_new_n34883__, new_new_n34884__,
    new_new_n34885__, new_new_n34886__, new_new_n34887__, new_new_n34888__,
    new_new_n34890__, new_new_n34891__, new_new_n34892__, new_new_n34893__,
    new_new_n34894__, new_new_n34895__, new_new_n34896__, new_new_n34897__,
    new_new_n34898__, new_new_n34899__, new_new_n34900__, new_new_n34901__,
    new_new_n34902__, new_new_n34903__, new_new_n34904__, new_new_n34905__,
    new_new_n34906__, new_new_n34907__, new_new_n34908__, new_new_n34909__,
    new_new_n34910__, new_new_n34911__, new_new_n34912__, new_new_n34913__,
    new_new_n34914__, new_new_n34915__, new_new_n34916__, new_new_n34917__,
    new_new_n34918__, new_new_n34919__, new_new_n34920__, new_new_n34921__,
    new_new_n34922__, new_new_n34923__, new_new_n34924__, new_new_n34925__,
    new_new_n34926__, new_new_n34928__, new_new_n34929__, new_new_n34930__,
    new_new_n34931__, new_new_n34932__, new_new_n34933__, new_new_n34934__,
    new_new_n34935__, new_new_n34936__, new_new_n34937__, new_new_n34938__,
    new_new_n34939__, new_new_n34940__, new_new_n34941__, new_new_n34942__,
    new_new_n34943__, new_new_n34944__, new_new_n34945__, new_new_n34946__,
    new_new_n34947__, new_new_n34948__, new_new_n34949__, new_new_n34950__,
    new_new_n34951__, new_new_n34952__, new_new_n34953__, new_new_n34954__,
    new_new_n34955__, new_new_n34956__, new_new_n34957__, new_new_n34958__,
    new_new_n34959__, new_new_n34960__, new_new_n34961__, new_new_n34962__,
    new_new_n34963__, new_new_n34964__, new_new_n34965__, new_new_n34966__,
    new_new_n34967__, new_new_n34969__, new_new_n34970__, new_new_n34971__,
    new_new_n34972__, new_new_n34973__, new_new_n34974__, new_new_n34975__,
    new_new_n34976__, new_new_n34977__, new_new_n34978__, new_new_n34979__,
    new_new_n34980__, new_new_n34981__, new_new_n34982__, new_new_n34983__,
    new_new_n34984__, new_new_n34985__, new_new_n34986__, new_new_n34987__,
    new_new_n34988__, new_new_n34989__, new_new_n34990__, new_new_n34991__,
    new_new_n34992__, new_new_n34993__, new_new_n34994__, new_new_n34995__,
    new_new_n34996__, new_new_n34997__, new_new_n34998__, new_new_n34999__,
    new_new_n35000__, new_new_n35001__, new_new_n35002__, new_new_n35003__,
    new_new_n35004__, new_new_n35005__, new_new_n35006__, new_new_n35007__,
    new_new_n35008__, new_new_n35010__, new_new_n35011__, new_new_n35012__,
    new_new_n35013__, new_new_n35014__, new_new_n35015__, new_new_n35016__,
    new_new_n35017__, new_new_n35018__, new_new_n35019__, new_new_n35020__,
    new_new_n35021__, new_new_n35022__, new_new_n35023__, new_new_n35024__,
    new_new_n35025__, new_new_n35026__, new_new_n35027__, new_new_n35028__,
    new_new_n35029__, new_new_n35030__, new_new_n35031__, new_new_n35032__,
    new_new_n35033__, new_new_n35034__, new_new_n35035__, new_new_n35036__,
    new_new_n35037__, new_new_n35038__, new_new_n35039__, new_new_n35040__,
    new_new_n35041__, new_new_n35042__, new_new_n35043__, new_new_n35044__,
    new_new_n35045__, new_new_n35046__, new_new_n35047__, new_new_n35048__,
    new_new_n35049__, new_new_n35050__, new_new_n35051__, new_new_n35052__,
    new_new_n35053__, new_new_n35054__, new_new_n35055__, new_new_n35056__,
    new_new_n35057__, new_new_n35059__, new_new_n35060__, new_new_n35061__,
    new_new_n35062__, new_new_n35063__, new_new_n35064__, new_new_n35065__,
    new_new_n35066__, new_new_n35067__, new_new_n35068__, new_new_n35069__,
    new_new_n35070__, new_new_n35071__, new_new_n35072__, new_new_n35073__,
    new_new_n35074__, new_new_n35075__, new_new_n35076__, new_new_n35077__,
    new_new_n35078__, new_new_n35079__, new_new_n35080__, new_new_n35081__,
    new_new_n35082__, new_new_n35083__, new_new_n35084__, new_new_n35085__,
    new_new_n35086__, new_new_n35087__, new_new_n35088__, new_new_n35089__,
    new_new_n35090__, new_new_n35091__, new_new_n35092__, new_new_n35093__,
    new_new_n35094__, new_new_n35095__, new_new_n35096__, new_new_n35097__,
    new_new_n35098__, new_new_n35099__, new_new_n35100__, new_new_n35101__,
    new_new_n35103__, new_new_n35104__, new_new_n35105__, new_new_n35106__,
    new_new_n35107__, new_new_n35108__, new_new_n35109__, new_new_n35110__,
    new_new_n35111__, new_new_n35112__, new_new_n35113__, new_new_n35114__,
    new_new_n35115__, new_new_n35116__, new_new_n35117__, new_new_n35118__,
    new_new_n35119__, new_new_n35120__, new_new_n35121__, new_new_n35122__,
    new_new_n35123__, new_new_n35124__, new_new_n35125__, new_new_n35126__,
    new_new_n35127__, new_new_n35128__, new_new_n35129__, new_new_n35130__,
    new_new_n35131__, new_new_n35132__, new_new_n35133__, new_new_n35134__,
    new_new_n35135__, new_new_n35136__, new_new_n35137__, new_new_n35138__,
    new_new_n35139__, new_new_n35140__, new_new_n35141__, new_new_n35142__,
    new_new_n35143__, new_new_n35144__, new_new_n35145__, new_new_n35147__,
    new_new_n35148__, new_new_n35149__, new_new_n35150__, new_new_n35151__,
    new_new_n35152__, new_new_n35153__, new_new_n35154__, new_new_n35155__,
    new_new_n35156__, new_new_n35157__, new_new_n35158__, new_new_n35159__,
    new_new_n35160__, new_new_n35161__, new_new_n35162__, new_new_n35163__,
    new_new_n35164__, new_new_n35165__, new_new_n35166__, new_new_n35167__,
    new_new_n35168__, new_new_n35169__, new_new_n35170__, new_new_n35171__,
    new_new_n35172__, new_new_n35173__, new_new_n35174__, new_new_n35175__,
    new_new_n35176__, new_new_n35177__, new_new_n35178__, new_new_n35179__,
    new_new_n35180__, new_new_n35181__, new_new_n35182__, new_new_n35183__,
    new_new_n35184__, new_new_n35185__, new_new_n35186__, new_new_n35188__,
    new_new_n35189__, new_new_n35190__, new_new_n35191__, new_new_n35192__,
    new_new_n35193__, new_new_n35194__, new_new_n35195__, new_new_n35196__,
    new_new_n35197__, new_new_n35198__, new_new_n35199__, new_new_n35200__,
    new_new_n35201__, new_new_n35202__, new_new_n35203__, new_new_n35204__,
    new_new_n35205__, new_new_n35206__, new_new_n35207__, new_new_n35208__,
    new_new_n35209__, new_new_n35210__, new_new_n35211__, new_new_n35212__,
    new_new_n35213__, new_new_n35214__, new_new_n35215__, new_new_n35216__,
    new_new_n35217__, new_new_n35218__, new_new_n35219__, new_new_n35220__,
    new_new_n35221__, new_new_n35222__, new_new_n35223__, new_new_n35224__,
    new_new_n35225__, new_new_n35226__, new_new_n35227__, new_new_n35228__,
    new_new_n35229__, new_new_n35230__, new_new_n35232__, new_new_n35233__,
    new_new_n35234__, new_new_n35235__, new_new_n35236__, new_new_n35237__,
    new_new_n35238__, new_new_n35239__, new_new_n35240__, new_new_n35241__,
    new_new_n35242__, new_new_n35243__, new_new_n35244__, new_new_n35245__,
    new_new_n35246__, new_new_n35247__, new_new_n35248__, new_new_n35249__,
    new_new_n35250__, new_new_n35251__, new_new_n35252__, new_new_n35253__,
    new_new_n35254__, new_new_n35255__, new_new_n35256__, new_new_n35257__,
    new_new_n35258__, new_new_n35259__, new_new_n35260__, new_new_n35261__,
    new_new_n35262__, new_new_n35263__, new_new_n35264__, new_new_n35265__,
    new_new_n35266__, new_new_n35267__, new_new_n35268__, new_new_n35269__,
    new_new_n35270__, new_new_n35271__, new_new_n35272__, new_new_n35273__,
    new_new_n35274__, new_new_n35276__, new_new_n35277__, new_new_n35278__,
    new_new_n35279__, new_new_n35280__, new_new_n35281__, new_new_n35282__,
    new_new_n35283__, new_new_n35284__, new_new_n35285__, new_new_n35286__,
    new_new_n35287__, new_new_n35288__, new_new_n35289__, new_new_n35290__,
    new_new_n35291__, new_new_n35292__, new_new_n35293__, new_new_n35294__,
    new_new_n35295__, new_new_n35296__, new_new_n35297__, new_new_n35298__,
    new_new_n35299__, new_new_n35300__, new_new_n35301__, new_new_n35302__,
    new_new_n35303__, new_new_n35304__, new_new_n35305__, new_new_n35306__,
    new_new_n35307__, new_new_n35308__, new_new_n35309__, new_new_n35310__,
    new_new_n35311__, new_new_n35312__, new_new_n35313__, new_new_n35314__,
    new_new_n35315__, new_new_n35319__, new_new_n35320__, new_new_n35321__,
    new_new_n35322__, new_new_n35323__, new_new_n35324__, new_new_n35325__,
    new_new_n35326__, new_new_n35327__, new_new_n35328__, new_new_n35329__,
    new_new_n35330__, new_new_n35331__, new_new_n35332__, new_new_n35333__,
    new_new_n35334__, new_new_n35335__, new_new_n35336__, new_new_n35337__,
    new_new_n35338__, new_new_n35339__, new_new_n35340__, new_new_n35341__,
    new_new_n35342__, new_new_n35343__, new_new_n35344__, new_new_n35345__,
    new_new_n35346__, new_new_n35347__, new_new_n35348__, new_new_n35349__,
    new_new_n35350__, new_new_n35351__, new_new_n35352__, new_new_n35353__,
    new_new_n35354__, new_new_n35355__, new_new_n35356__, new_new_n35357__,
    new_new_n35358__, new_new_n35359__, new_new_n35360__, new_new_n35361__,
    new_new_n35362__, new_new_n35363__, new_new_n35364__, new_new_n35365__,
    new_new_n35366__, new_new_n35367__, new_new_n35368__, new_new_n35369__,
    new_new_n35370__, new_new_n35371__, new_new_n35372__, new_new_n35373__,
    new_new_n35374__, new_new_n35375__, new_new_n35376__, new_new_n35377__,
    new_new_n35378__, new_new_n35379__, new_new_n35380__, new_new_n35381__,
    new_new_n35382__, new_new_n35383__, new_new_n35384__, new_new_n35385__,
    new_new_n35386__, new_new_n35387__, new_new_n35388__, new_new_n35389__,
    new_new_n35390__, new_new_n35391__, new_new_n35392__, new_new_n35393__,
    new_new_n35394__, new_new_n35395__, new_new_n35396__, new_new_n35397__,
    new_new_n35398__, new_new_n35399__, new_new_n35400__, new_new_n35401__,
    new_new_n35402__, new_new_n35403__, new_new_n35404__, new_new_n35405__,
    new_new_n35406__, new_new_n35407__, new_new_n35408__, new_new_n35409__,
    new_new_n35410__, new_new_n35411__, new_new_n35412__, new_new_n35413__,
    new_new_n35414__, new_new_n35415__, new_new_n35416__, new_new_n35417__,
    new_new_n35418__, new_new_n35419__, new_new_n35420__, new_new_n35421__,
    new_new_n35422__, new_new_n35423__, new_new_n35424__, new_new_n35425__,
    new_new_n35426__, new_new_n35427__, new_new_n35428__, new_new_n35429__,
    new_new_n35430__, new_new_n35431__, new_new_n35432__, new_new_n35434__,
    new_new_n35435__, new_new_n35436__, new_new_n35437__, new_new_n35438__,
    new_new_n35439__, new_new_n35440__, new_new_n35441__, new_new_n35442__,
    new_new_n35443__, new_new_n35444__, new_new_n35445__, new_new_n35446__,
    new_new_n35447__, new_new_n35448__, new_new_n35449__, new_new_n35450__,
    new_new_n35451__, new_new_n35452__, new_new_n35453__, new_new_n35454__,
    new_new_n35455__, new_new_n35456__, new_new_n35457__, new_new_n35458__,
    new_new_n35460__, new_new_n35461__, new_new_n35462__, new_new_n35463__,
    new_new_n35464__, new_new_n35465__, new_new_n35466__, new_new_n35467__,
    new_new_n35468__, new_new_n35469__, new_new_n35470__, new_new_n35471__,
    new_new_n35472__, new_new_n35473__, new_new_n35474__, new_new_n35475__,
    new_new_n35476__, new_new_n35477__, new_new_n35478__, new_new_n35479__,
    new_new_n35480__, new_new_n35481__, new_new_n35482__, new_new_n35483__,
    new_new_n35484__, new_new_n35485__, new_new_n35486__, new_new_n35487__,
    new_new_n35488__, new_new_n35489__, new_new_n35491__, new_new_n35492__,
    new_new_n35493__, new_new_n35494__, new_new_n35495__, new_new_n35496__,
    new_new_n35497__, new_new_n35498__, new_new_n35499__, new_new_n35500__,
    new_new_n35501__, new_new_n35502__, new_new_n35503__, new_new_n35504__,
    new_new_n35505__, new_new_n35506__, new_new_n35507__, new_new_n35508__,
    new_new_n35509__, new_new_n35510__, new_new_n35511__, new_new_n35512__,
    new_new_n35513__, new_new_n35514__, new_new_n35515__, new_new_n35516__,
    new_new_n35517__, new_new_n35518__, new_new_n35519__, new_new_n35520__,
    new_new_n35521__, new_new_n35522__, new_new_n35523__, new_new_n35524__,
    new_new_n35525__, new_new_n35526__, new_new_n35528__, new_new_n35529__,
    new_new_n35530__, new_new_n35531__, new_new_n35532__, new_new_n35533__,
    new_new_n35534__, new_new_n35535__, new_new_n35536__, new_new_n35537__,
    new_new_n35538__, new_new_n35539__, new_new_n35540__, new_new_n35541__,
    new_new_n35542__, new_new_n35543__, new_new_n35544__, new_new_n35545__,
    new_new_n35546__, new_new_n35547__, new_new_n35548__, new_new_n35549__,
    new_new_n35550__, new_new_n35551__, new_new_n35552__, new_new_n35553__,
    new_new_n35554__, new_new_n35555__, new_new_n35556__, new_new_n35557__,
    new_new_n35558__, new_new_n35559__, new_new_n35560__, new_new_n35561__,
    new_new_n35562__, new_new_n35563__, new_new_n35564__, new_new_n35565__,
    new_new_n35566__, new_new_n35567__, new_new_n35569__, new_new_n35570__,
    new_new_n35571__, new_new_n35572__, new_new_n35573__, new_new_n35574__,
    new_new_n35575__, new_new_n35576__, new_new_n35577__, new_new_n35578__,
    new_new_n35579__, new_new_n35580__, new_new_n35581__, new_new_n35582__,
    new_new_n35583__, new_new_n35584__, new_new_n35585__, new_new_n35586__,
    new_new_n35587__, new_new_n35588__, new_new_n35589__, new_new_n35590__,
    new_new_n35591__, new_new_n35592__, new_new_n35593__, new_new_n35594__,
    new_new_n35595__, new_new_n35596__, new_new_n35597__, new_new_n35598__,
    new_new_n35599__, new_new_n35600__, new_new_n35601__, new_new_n35602__,
    new_new_n35603__, new_new_n35604__, new_new_n35605__, new_new_n35606__,
    new_new_n35607__, new_new_n35608__, new_new_n35609__, new_new_n35610__,
    new_new_n35612__, new_new_n35613__, new_new_n35614__, new_new_n35615__,
    new_new_n35616__, new_new_n35617__, new_new_n35618__, new_new_n35619__,
    new_new_n35620__, new_new_n35621__, new_new_n35622__, new_new_n35623__,
    new_new_n35624__, new_new_n35625__, new_new_n35626__, new_new_n35627__,
    new_new_n35628__, new_new_n35629__, new_new_n35630__, new_new_n35631__,
    new_new_n35632__, new_new_n35633__, new_new_n35634__, new_new_n35635__,
    new_new_n35636__, new_new_n35637__, new_new_n35638__, new_new_n35639__,
    new_new_n35640__, new_new_n35641__, new_new_n35642__, new_new_n35643__,
    new_new_n35644__, new_new_n35645__, new_new_n35646__, new_new_n35647__,
    new_new_n35648__, new_new_n35649__, new_new_n35650__, new_new_n35651__,
    new_new_n35652__, new_new_n35653__, new_new_n35655__, new_new_n35656__,
    new_new_n35657__, new_new_n35658__, new_new_n35659__, new_new_n35660__,
    new_new_n35661__, new_new_n35662__, new_new_n35663__, new_new_n35664__,
    new_new_n35665__, new_new_n35666__, new_new_n35667__, new_new_n35668__,
    new_new_n35669__, new_new_n35670__, new_new_n35671__, new_new_n35672__,
    new_new_n35673__, new_new_n35674__, new_new_n35675__, new_new_n35676__,
    new_new_n35677__, new_new_n35678__, new_new_n35679__, new_new_n35680__,
    new_new_n35681__, new_new_n35682__, new_new_n35683__, new_new_n35684__,
    new_new_n35685__, new_new_n35687__, new_new_n35688__, new_new_n35689__,
    new_new_n35690__, new_new_n35691__, new_new_n35692__, new_new_n35693__,
    new_new_n35694__, new_new_n35695__, new_new_n35696__, new_new_n35697__,
    new_new_n35698__, new_new_n35699__, new_new_n35700__, new_new_n35701__,
    new_new_n35702__, new_new_n35703__, new_new_n35704__, new_new_n35705__,
    new_new_n35706__, new_new_n35707__, new_new_n35708__, new_new_n35709__,
    new_new_n35710__, new_new_n35711__, new_new_n35712__, new_new_n35713__,
    new_new_n35714__, new_new_n35715__, new_new_n35716__, new_new_n35717__,
    new_new_n35719__, new_new_n35720__, new_new_n35721__, new_new_n35722__,
    new_new_n35723__, new_new_n35724__, new_new_n35725__, new_new_n35726__,
    new_new_n35727__, new_new_n35728__, new_new_n35729__, new_new_n35730__,
    new_new_n35731__, new_new_n35732__, new_new_n35733__, new_new_n35734__,
    new_new_n35735__, new_new_n35736__, new_new_n35737__, new_new_n35738__,
    new_new_n35739__, new_new_n35740__, new_new_n35741__, new_new_n35742__,
    new_new_n35743__, new_new_n35744__, new_new_n35745__, new_new_n35746__,
    new_new_n35747__, new_new_n35748__, new_new_n35749__, new_new_n35751__,
    new_new_n35752__, new_new_n35753__, new_new_n35754__, new_new_n35755__,
    new_new_n35756__, new_new_n35757__, new_new_n35758__, new_new_n35759__,
    new_new_n35760__, new_new_n35761__, new_new_n35762__, new_new_n35763__,
    new_new_n35764__, new_new_n35765__, new_new_n35766__, new_new_n35767__,
    new_new_n35768__, new_new_n35769__, new_new_n35770__, new_new_n35771__,
    new_new_n35772__, new_new_n35773__, new_new_n35774__, new_new_n35775__,
    new_new_n35776__, new_new_n35777__, new_new_n35778__, new_new_n35779__,
    new_new_n35780__, new_new_n35781__, new_new_n35783__, new_new_n35784__,
    new_new_n35785__, new_new_n35786__, new_new_n35787__, new_new_n35788__,
    new_new_n35789__, new_new_n35790__, new_new_n35791__, new_new_n35792__,
    new_new_n35793__, new_new_n35794__, new_new_n35795__, new_new_n35796__,
    new_new_n35797__, new_new_n35798__, new_new_n35799__, new_new_n35800__,
    new_new_n35801__, new_new_n35802__, new_new_n35803__, new_new_n35804__,
    new_new_n35805__, new_new_n35806__, new_new_n35807__, new_new_n35808__,
    new_new_n35809__, new_new_n35810__, new_new_n35811__, new_new_n35812__,
    new_new_n35813__, new_new_n35815__, new_new_n35816__, new_new_n35817__,
    new_new_n35818__, new_new_n35819__, new_new_n35820__, new_new_n35821__,
    new_new_n35822__, new_new_n35823__, new_new_n35824__, new_new_n35825__,
    new_new_n35826__, new_new_n35827__, new_new_n35828__, new_new_n35829__,
    new_new_n35830__, new_new_n35831__, new_new_n35832__, new_new_n35833__,
    new_new_n35834__, new_new_n35835__, new_new_n35836__, new_new_n35837__,
    new_new_n35838__, new_new_n35839__, new_new_n35840__, new_new_n35841__,
    new_new_n35842__, new_new_n35843__, new_new_n35844__, new_new_n35845__,
    new_new_n35847__, new_new_n35848__, new_new_n35849__, new_new_n35850__,
    new_new_n35851__, new_new_n35852__, new_new_n35853__, new_new_n35854__,
    new_new_n35855__, new_new_n35856__, new_new_n35857__, new_new_n35858__,
    new_new_n35859__, new_new_n35860__, new_new_n35861__, new_new_n35862__,
    new_new_n35863__, new_new_n35864__, new_new_n35865__, new_new_n35866__,
    new_new_n35867__, new_new_n35868__, new_new_n35869__, new_new_n35870__,
    new_new_n35871__, new_new_n35872__, new_new_n35873__, new_new_n35874__,
    new_new_n35875__, new_new_n35876__, new_new_n35877__, new_new_n35879__,
    new_new_n35880__, new_new_n35881__, new_new_n35882__, new_new_n35883__,
    new_new_n35884__, new_new_n35885__, new_new_n35886__, new_new_n35887__,
    new_new_n35888__, new_new_n35889__, new_new_n35890__, new_new_n35891__,
    new_new_n35892__, new_new_n35893__, new_new_n35894__, new_new_n35895__,
    new_new_n35896__, new_new_n35897__, new_new_n35898__, new_new_n35899__,
    new_new_n35900__, new_new_n35901__, new_new_n35903__, new_new_n35904__,
    new_new_n35905__, new_new_n35906__, new_new_n35907__, new_new_n35908__,
    new_new_n35909__, new_new_n35910__, new_new_n35911__, new_new_n35912__,
    new_new_n35913__, new_new_n35914__, new_new_n35915__, new_new_n35916__,
    new_new_n35917__, new_new_n35918__, new_new_n35919__, new_new_n35920__,
    new_new_n35921__, new_new_n35922__, new_new_n35923__, new_new_n35924__,
    new_new_n35925__, new_new_n35927__, new_new_n35928__, new_new_n35929__,
    new_new_n35930__, new_new_n35931__, new_new_n35932__, new_new_n35933__,
    new_new_n35934__, new_new_n35935__, new_new_n35936__, new_new_n35937__,
    new_new_n35938__, new_new_n35939__, new_new_n35940__, new_new_n35941__,
    new_new_n35942__, new_new_n35943__, new_new_n35944__, new_new_n35945__,
    new_new_n35946__, new_new_n35947__, new_new_n35948__, new_new_n35949__,
    new_new_n35951__, new_new_n35952__, new_new_n35953__, new_new_n35954__,
    new_new_n35955__, new_new_n35956__, new_new_n35957__, new_new_n35958__,
    new_new_n35959__, new_new_n35960__, new_new_n35961__, new_new_n35962__,
    new_new_n35963__, new_new_n35964__, new_new_n35965__, new_new_n35966__,
    new_new_n35967__, new_new_n35968__, new_new_n35969__, new_new_n35970__,
    new_new_n35971__, new_new_n35972__, new_new_n35973__, new_new_n35975__,
    new_new_n35976__, new_new_n35977__, new_new_n35978__, new_new_n35979__,
    new_new_n35980__, new_new_n35981__, new_new_n35982__, new_new_n35983__,
    new_new_n35984__, new_new_n35985__, new_new_n35986__, new_new_n35987__,
    new_new_n35988__, new_new_n35989__, new_new_n35990__, new_new_n35991__,
    new_new_n35992__, new_new_n35993__, new_new_n35994__, new_new_n35995__,
    new_new_n35996__, new_new_n35997__, new_new_n35999__, new_new_n36000__,
    new_new_n36001__, new_new_n36002__, new_new_n36003__, new_new_n36004__,
    new_new_n36005__, new_new_n36006__, new_new_n36007__, new_new_n36008__,
    new_new_n36009__, new_new_n36010__, new_new_n36011__, new_new_n36012__,
    new_new_n36013__, new_new_n36014__, new_new_n36015__, new_new_n36016__,
    new_new_n36017__, new_new_n36018__, new_new_n36019__, new_new_n36020__,
    new_new_n36021__, new_new_n36023__, new_new_n36024__, new_new_n36025__,
    new_new_n36026__, new_new_n36027__, new_new_n36028__, new_new_n36029__,
    new_new_n36030__, new_new_n36031__, new_new_n36032__, new_new_n36033__,
    new_new_n36034__, new_new_n36035__, new_new_n36036__, new_new_n36037__,
    new_new_n36038__, new_new_n36039__, new_new_n36040__, new_new_n36041__,
    new_new_n36042__, new_new_n36043__, new_new_n36044__, new_new_n36045__,
    new_new_n36047__, new_new_n36048__, new_new_n36049__, new_new_n36050__,
    new_new_n36051__, new_new_n36052__, new_new_n36053__, new_new_n36054__,
    new_new_n36055__, new_new_n36056__, new_new_n36057__, new_new_n36058__,
    new_new_n36059__, new_new_n36060__, new_new_n36061__, new_new_n36062__,
    new_new_n36063__, new_new_n36064__, new_new_n36065__, new_new_n36066__,
    new_new_n36067__, new_new_n36068__, new_new_n36069__, new_new_n36071__,
    new_new_n36072__, new_new_n36073__, new_new_n36074__, new_new_n36075__,
    new_new_n36076__, new_new_n36077__, new_new_n36078__, new_new_n36079__,
    new_new_n36080__, new_new_n36081__, new_new_n36082__, new_new_n36083__,
    new_new_n36084__, new_new_n36085__, new_new_n36086__, new_new_n36087__,
    new_new_n36088__, new_new_n36089__, new_new_n36090__, new_new_n36091__,
    new_new_n36092__, new_new_n36093__, new_new_n36095__, new_new_n36096__,
    new_new_n36097__, new_new_n36098__, new_new_n36099__, new_new_n36100__,
    new_new_n36101__, new_new_n36102__, new_new_n36103__, new_new_n36104__,
    new_new_n36105__, new_new_n36106__, new_new_n36107__, new_new_n36108__,
    new_new_n36109__, new_new_n36110__, new_new_n36111__, new_new_n36112__,
    new_new_n36113__, new_new_n36114__, new_new_n36115__, new_new_n36116__,
    new_new_n36117__, new_new_n36119__, new_new_n36120__, new_new_n36121__,
    new_new_n36122__, new_new_n36123__, new_new_n36124__, new_new_n36125__,
    new_new_n36126__, new_new_n36127__, new_new_n36128__, new_new_n36129__,
    new_new_n36130__, new_new_n36131__, new_new_n36132__, new_new_n36133__,
    new_new_n36134__, new_new_n36135__, new_new_n36136__, new_new_n36137__,
    new_new_n36138__, new_new_n36139__, new_new_n36140__, new_new_n36141__,
    new_new_n36143__, new_new_n36144__, new_new_n36145__, new_new_n36146__,
    new_new_n36147__, new_new_n36148__, new_new_n36149__, new_new_n36150__,
    new_new_n36151__, new_new_n36152__, new_new_n36153__, new_new_n36154__,
    new_new_n36155__, new_new_n36156__, new_new_n36157__, new_new_n36158__,
    new_new_n36159__, new_new_n36160__, new_new_n36161__, new_new_n36162__,
    new_new_n36163__, new_new_n36164__, new_new_n36165__, new_new_n36167__,
    new_new_n36168__, new_new_n36169__, new_new_n36170__, new_new_n36171__,
    new_new_n36172__, new_new_n36173__, new_new_n36174__, new_new_n36175__,
    new_new_n36176__, new_new_n36177__, new_new_n36178__, new_new_n36179__,
    new_new_n36180__, new_new_n36181__, new_new_n36182__, new_new_n36183__,
    new_new_n36184__, new_new_n36185__, new_new_n36186__, new_new_n36187__,
    new_new_n36188__, new_new_n36189__, new_new_n36191__, new_new_n36192__,
    new_new_n36193__, new_new_n36194__, new_new_n36195__, new_new_n36196__,
    new_new_n36197__, new_new_n36198__, new_new_n36199__, new_new_n36200__,
    new_new_n36201__, new_new_n36202__, new_new_n36203__, new_new_n36204__,
    new_new_n36205__, new_new_n36206__, new_new_n36207__, new_new_n36208__,
    new_new_n36209__, new_new_n36210__, new_new_n36211__, new_new_n36212__,
    new_new_n36213__, new_new_n36215__, new_new_n36216__, new_new_n36217__,
    new_new_n36218__, new_new_n36219__, new_new_n36220__, new_new_n36221__,
    new_new_n36222__, new_new_n36223__, new_new_n36224__, new_new_n36225__,
    new_new_n36226__, new_new_n36227__, new_new_n36228__, new_new_n36229__,
    new_new_n36230__, new_new_n36231__, new_new_n36232__, new_new_n36233__,
    new_new_n36234__, new_new_n36235__, new_new_n36236__, new_new_n36237__,
    new_new_n36239__, new_new_n36240__, new_new_n36241__, new_new_n36242__,
    new_new_n36243__, new_new_n36244__, new_new_n36245__, new_new_n36246__,
    new_new_n36247__, new_new_n36248__, new_new_n36249__, new_new_n36250__,
    new_new_n36251__, new_new_n36252__, new_new_n36253__, new_new_n36254__,
    new_new_n36255__, new_new_n36256__, new_new_n36257__, new_new_n36258__,
    new_new_n36259__, new_new_n36260__, new_new_n36261__, new_new_n36263__,
    new_new_n36264__, new_new_n36265__, new_new_n36266__, new_new_n36267__,
    new_new_n36268__, new_new_n36269__, new_new_n36270__, new_new_n36271__,
    new_new_n36272__, new_new_n36273__, new_new_n36274__, new_new_n36275__,
    new_new_n36276__, new_new_n36277__, new_new_n36278__, new_new_n36279__,
    new_new_n36280__, new_new_n36281__, new_new_n36282__, new_new_n36283__,
    new_new_n36284__, new_new_n36285__, new_new_n36287__, new_new_n36288__,
    new_new_n36289__, new_new_n36290__, new_new_n36291__, new_new_n36292__,
    new_new_n36293__, new_new_n36294__, new_new_n36295__, new_new_n36296__,
    new_new_n36297__, new_new_n36298__, new_new_n36299__, new_new_n36300__,
    new_new_n36301__, new_new_n36302__, new_new_n36303__, new_new_n36304__,
    new_new_n36305__, new_new_n36306__, new_new_n36307__, new_new_n36308__,
    new_new_n36309__, new_new_n36311__, new_new_n36312__, new_new_n36313__,
    new_new_n36314__, new_new_n36315__, new_new_n36316__, new_new_n36317__,
    new_new_n36318__, new_new_n36319__, new_new_n36320__, new_new_n36321__,
    new_new_n36322__, new_new_n36323__, new_new_n36324__, new_new_n36325__,
    new_new_n36326__, new_new_n36327__, new_new_n36328__, new_new_n36329__,
    new_new_n36330__, new_new_n36331__, new_new_n36332__, new_new_n36333__,
    new_new_n36335__, new_new_n36336__, new_new_n36337__, new_new_n36338__,
    new_new_n36339__, new_new_n36340__, new_new_n36341__, new_new_n36342__,
    new_new_n36343__, new_new_n36344__, new_new_n36345__, new_new_n36346__,
    new_new_n36347__, new_new_n36348__, new_new_n36349__, new_new_n36350__,
    new_new_n36351__, new_new_n36352__, new_new_n36353__, new_new_n36354__,
    new_new_n36355__, new_new_n36356__, new_new_n36357__, new_new_n36359__,
    new_new_n36360__, new_new_n36361__, new_new_n36362__, new_new_n36363__,
    new_new_n36364__, new_new_n36365__, new_new_n36366__, new_new_n36367__,
    new_new_n36368__, new_new_n36369__, new_new_n36370__, new_new_n36371__,
    new_new_n36372__, new_new_n36373__, new_new_n36374__, new_new_n36375__,
    new_new_n36376__, new_new_n36377__, new_new_n36378__, new_new_n36379__,
    new_new_n36380__, new_new_n36381__, new_new_n36383__, new_new_n36384__,
    new_new_n36385__, new_new_n36386__, new_new_n36387__, new_new_n36388__,
    new_new_n36389__, new_new_n36390__, new_new_n36391__, new_new_n36392__,
    new_new_n36393__, new_new_n36394__, new_new_n36395__, new_new_n36396__,
    new_new_n36397__, new_new_n36398__, new_new_n36399__, new_new_n36400__,
    new_new_n36401__, new_new_n36402__, new_new_n36403__, new_new_n36404__,
    new_new_n36405__, new_new_n36407__, new_new_n36408__, new_new_n36409__,
    new_new_n36410__, new_new_n36411__, new_new_n36412__, new_new_n36413__,
    new_new_n36414__, new_new_n36415__, new_new_n36416__, new_new_n36417__,
    new_new_n36418__, new_new_n36419__, new_new_n36420__, new_new_n36421__,
    new_new_n36422__, new_new_n36423__, new_new_n36424__, new_new_n36425__,
    new_new_n36426__, new_new_n36427__, new_new_n36428__, new_new_n36429__,
    new_new_n36431__, new_new_n36432__, new_new_n36433__, new_new_n36434__,
    new_new_n36435__, new_new_n36436__, new_new_n36437__, new_new_n36438__,
    new_new_n36439__, new_new_n36440__, new_new_n36441__, new_new_n36442__,
    new_new_n36443__, new_new_n36444__, new_new_n36445__, new_new_n36446__,
    new_new_n36447__, new_new_n36448__, new_new_n36449__, new_new_n36451__,
    new_new_n36452__, new_new_n36453__, new_new_n36454__, new_new_n36455__,
    new_new_n36456__, new_new_n36457__, new_new_n36458__, new_new_n36459__,
    new_new_n36460__, new_new_n36461__, new_new_n36462__, new_new_n36463__,
    new_new_n36465__, new_new_n36466__, new_new_n36467__, new_new_n36468__,
    new_new_n36469__, new_new_n36470__, new_new_n36471__, new_new_n36472__,
    new_new_n36473__, new_new_n36474__, new_new_n36475__, new_new_n36476__,
    new_new_n36477__, new_new_n36479__, new_new_n36480__, new_new_n36481__,
    new_new_n36482__, new_new_n36483__, new_new_n36484__, new_new_n36485__,
    new_new_n36486__, new_new_n36487__, new_new_n36488__, new_new_n36489__,
    new_new_n36490__, new_new_n36491__, new_new_n36493__, new_new_n36494__,
    new_new_n36495__, new_new_n36496__, new_new_n36497__, new_new_n36498__,
    new_new_n36499__, new_new_n36500__, new_new_n36501__, new_new_n36502__,
    new_new_n36503__, new_new_n36504__, new_new_n36505__, new_new_n36507__,
    new_new_n36508__, new_new_n36509__, new_new_n36510__, new_new_n36511__,
    new_new_n36512__, new_new_n36513__, new_new_n36514__, new_new_n36515__,
    new_new_n36516__, new_new_n36517__, new_new_n36518__, new_new_n36520__,
    new_new_n36521__, new_new_n36522__, new_new_n36523__, new_new_n36524__,
    new_new_n36525__, new_new_n36526__, new_new_n36527__, new_new_n36528__,
    new_new_n36529__, new_new_n36530__, new_new_n36531__, new_new_n36533__,
    new_new_n36534__, new_new_n36535__, new_new_n36536__, new_new_n36537__,
    new_new_n36538__, new_new_n36539__, new_new_n36540__, new_new_n36541__,
    new_new_n36542__, new_new_n36544__, new_new_n36545__, new_new_n36546__,
    new_new_n36547__, new_new_n36548__, new_new_n36549__, new_new_n36550__,
    new_new_n36551__, new_new_n36552__, new_new_n36553__, new_new_n36555__,
    new_new_n36556__, new_new_n36557__, new_new_n36558__, new_new_n36559__,
    new_new_n36560__, new_new_n36561__, new_new_n36562__, new_new_n36563__,
    new_new_n36564__, new_new_n36565__, new_new_n36566__, new_new_n36567__,
    new_new_n36568__, new_new_n36569__, new_new_n36570__, new_new_n36571__,
    new_new_n36572__, new_new_n36573__, new_new_n36574__, new_new_n36575__,
    new_new_n36577__, new_new_n36578__, new_new_n36579__, new_new_n36580__,
    new_new_n36581__, new_new_n36582__, new_new_n36583__, new_new_n36584__,
    new_new_n36585__, new_new_n36586__, new_new_n36587__, new_new_n36588__,
    new_new_n36589__, new_new_n36590__, new_new_n36591__, new_new_n36592__,
    new_new_n36593__, new_new_n36594__, new_new_n36595__, new_new_n36596__,
    new_new_n36597__, new_new_n36599__, new_new_n36600__, new_new_n36601__,
    new_new_n36602__, new_new_n36603__, new_new_n36604__, new_new_n36605__,
    new_new_n36606__, new_new_n36607__, new_new_n36608__, new_new_n36609__,
    new_new_n36610__, new_new_n36611__, new_new_n36612__, new_new_n36613__,
    new_new_n36614__, new_new_n36615__, new_new_n36616__, new_new_n36617__,
    new_new_n36618__, new_new_n36619__, new_new_n36621__, new_new_n36622__,
    new_new_n36623__, new_new_n36624__, new_new_n36625__, new_new_n36626__,
    new_new_n36627__, new_new_n36628__, new_new_n36629__, new_new_n36630__,
    new_new_n36631__, new_new_n36632__, new_new_n36633__, new_new_n36634__,
    new_new_n36635__, new_new_n36636__, new_new_n36637__, new_new_n36638__,
    new_new_n36639__, new_new_n36640__, new_new_n36641__, new_new_n36643__,
    new_new_n36644__, new_new_n36645__, new_new_n36646__, new_new_n36647__,
    new_new_n36648__, new_new_n36649__, new_new_n36650__, new_new_n36651__,
    new_new_n36652__, new_new_n36653__, new_new_n36654__, new_new_n36655__,
    new_new_n36656__, new_new_n36657__, new_new_n36658__, new_new_n36659__,
    new_new_n36660__, new_new_n36661__, new_new_n36662__, new_new_n36663__,
    new_new_n36665__, new_new_n36666__, new_new_n36667__, new_new_n36668__,
    new_new_n36669__, new_new_n36670__, new_new_n36671__, new_new_n36672__,
    new_new_n36673__, new_new_n36674__, new_new_n36675__, new_new_n36676__,
    new_new_n36677__, new_new_n36678__, new_new_n36679__, new_new_n36680__,
    new_new_n36681__, new_new_n36682__, new_new_n36683__, new_new_n36684__,
    new_new_n36685__, new_new_n36687__, new_new_n36688__, new_new_n36689__,
    new_new_n36690__, new_new_n36691__, new_new_n36692__, new_new_n36693__,
    new_new_n36694__, new_new_n36695__, new_new_n36696__, new_new_n36697__,
    new_new_n36698__, new_new_n36699__, new_new_n36700__, new_new_n36701__,
    new_new_n36702__, new_new_n36703__, new_new_n36704__, new_new_n36705__,
    new_new_n36706__, new_new_n36707__, new_new_n36709__, new_new_n36710__,
    new_new_n36711__, new_new_n36712__, new_new_n36713__, new_new_n36714__,
    new_new_n36715__, new_new_n36716__, new_new_n36717__, new_new_n36718__,
    new_new_n36719__, new_new_n36720__, new_new_n36721__, new_new_n36722__,
    new_new_n36723__, new_new_n36724__, new_new_n36725__, new_new_n36726__,
    new_new_n36727__, new_new_n36728__, new_new_n36729__, new_new_n36730__,
    new_new_n36731__, new_new_n36732__, new_new_n36733__, new_new_n36734__,
    new_new_n36735__, new_new_n36736__, new_new_n36737__, new_new_n36738__,
    new_new_n36739__, new_new_n36740__, new_new_n36741__, new_new_n36742__,
    new_new_n36743__, new_new_n36744__, new_new_n36745__, new_new_n36746__,
    new_new_n36747__, new_new_n36748__, new_new_n36749__, new_new_n36750__,
    new_new_n36751__, new_new_n36752__, new_new_n36753__, new_new_n36754__,
    new_new_n36755__, new_new_n36756__, new_new_n36757__, new_new_n36758__,
    new_new_n36760__, new_new_n36761__, new_new_n36762__, new_new_n36763__,
    new_new_n36764__, new_new_n36765__, new_new_n36766__, new_new_n36767__,
    new_new_n36768__, new_new_n36769__, new_new_n36770__, new_new_n36771__,
    new_new_n36772__, new_new_n36773__, new_new_n36775__, new_new_n36776__,
    new_new_n36777__, new_new_n36778__, new_new_n36779__, new_new_n36780__,
    new_new_n36781__, new_new_n36782__, new_new_n36783__, new_new_n36784__,
    new_new_n36785__, new_new_n36786__, new_new_n36787__, new_new_n36788__,
    new_new_n36790__, new_new_n36791__, new_new_n36792__, new_new_n36793__,
    new_new_n36794__, new_new_n36795__, new_new_n36796__, new_new_n36797__,
    new_new_n36798__, new_new_n36799__, new_new_n36800__, new_new_n36801__,
    new_new_n36802__, new_new_n36803__, new_new_n36805__, new_new_n36806__,
    new_new_n36807__, new_new_n36808__, new_new_n36809__, new_new_n36810__,
    new_new_n36811__, new_new_n36812__, new_new_n36813__, new_new_n36814__,
    new_new_n36815__, new_new_n36816__, new_new_n36817__, new_new_n36818__,
    new_new_n36820__, new_new_n36821__, new_new_n36822__, new_new_n36823__,
    new_new_n36824__, new_new_n36825__, new_new_n36826__, new_new_n36827__,
    new_new_n36828__, new_new_n36829__, new_new_n36830__, new_new_n36831__,
    new_new_n36832__, new_new_n36833__, new_new_n36835__, new_new_n36836__,
    new_new_n36837__, new_new_n36838__, new_new_n36839__, new_new_n36840__,
    new_new_n36841__, new_new_n36842__, new_new_n36843__, new_new_n36844__,
    new_new_n36845__, new_new_n36846__, new_new_n36847__, new_new_n36848__,
    new_new_n36850__, new_new_n36851__, new_new_n36852__, new_new_n36853__,
    new_new_n36854__, new_new_n36855__, new_new_n36856__, new_new_n36857__,
    new_new_n36858__, new_new_n36859__, new_new_n36860__, new_new_n36861__,
    new_new_n36862__, new_new_n36863__, new_new_n36865__, new_new_n36866__,
    new_new_n36867__, new_new_n36868__, new_new_n36869__, new_new_n36870__,
    new_new_n36871__, new_new_n36872__, new_new_n36873__, new_new_n36874__,
    new_new_n36875__, new_new_n36876__, new_new_n36877__, new_new_n36878__,
    new_new_n36879__, new_new_n36880__, new_new_n36881__, new_new_n36882__,
    new_new_n36884__, new_new_n36885__, new_new_n36886__, new_new_n36887__,
    new_new_n36888__, new_new_n36889__, new_new_n36890__, new_new_n36891__,
    new_new_n36892__, new_new_n36893__, new_new_n36894__, new_new_n36895__,
    new_new_n36896__, new_new_n36897__, new_new_n36899__, new_new_n36900__,
    new_new_n36901__, new_new_n36902__, new_new_n36903__, new_new_n36904__,
    new_new_n36905__, new_new_n36906__, new_new_n36907__, new_new_n36908__,
    new_new_n36909__, new_new_n36910__, new_new_n36911__, new_new_n36912__,
    new_new_n36914__, new_new_n36915__, new_new_n36916__, new_new_n36917__,
    new_new_n36918__, new_new_n36919__, new_new_n36920__, new_new_n36921__,
    new_new_n36922__, new_new_n36923__, new_new_n36924__, new_new_n36925__,
    new_new_n36926__, new_new_n36927__, new_new_n36929__, new_new_n36930__,
    new_new_n36931__, new_new_n36932__, new_new_n36933__, new_new_n36934__,
    new_new_n36935__, new_new_n36936__, new_new_n36937__, new_new_n36938__,
    new_new_n36939__, new_new_n36940__, new_new_n36941__, new_new_n36942__,
    new_new_n36944__, new_new_n36945__, new_new_n36946__, new_new_n36947__,
    new_new_n36948__, new_new_n36949__, new_new_n36950__, new_new_n36951__,
    new_new_n36952__, new_new_n36953__, new_new_n36954__, new_new_n36955__,
    new_new_n36956__, new_new_n36957__, new_new_n36959__, new_new_n36960__,
    new_new_n36961__, new_new_n36962__, new_new_n36963__, new_new_n36964__,
    new_new_n36965__, new_new_n36966__, new_new_n36967__, new_new_n36968__,
    new_new_n36969__, new_new_n36970__, new_new_n36971__, new_new_n36972__,
    new_new_n36974__, new_new_n36975__, new_new_n36976__, new_new_n36977__,
    new_new_n36978__, new_new_n36979__, new_new_n36980__, new_new_n36981__,
    new_new_n36982__, new_new_n36983__, new_new_n36984__, new_new_n36985__,
    new_new_n36986__, new_new_n36987__, new_new_n36989__, new_new_n36990__,
    new_new_n36991__, new_new_n36992__, new_new_n36993__, new_new_n36994__,
    new_new_n36995__, new_new_n36996__, new_new_n36997__, new_new_n36998__,
    new_new_n36999__, new_new_n37000__, new_new_n37001__, new_new_n37002__,
    new_new_n37004__, new_new_n37005__, new_new_n37006__, new_new_n37007__,
    new_new_n37008__, new_new_n37009__, new_new_n37010__, new_new_n37011__,
    new_new_n37012__, new_new_n37013__, new_new_n37014__, new_new_n37015__,
    new_new_n37016__, new_new_n37017__, new_new_n37019__, new_new_n37020__,
    new_new_n37021__, new_new_n37022__, new_new_n37023__, new_new_n37024__,
    new_new_n37025__, new_new_n37026__, new_new_n37027__, new_new_n37028__,
    new_new_n37029__, new_new_n37030__, new_new_n37031__, new_new_n37032__,
    new_new_n37034__, new_new_n37035__, new_new_n37036__, new_new_n37037__,
    new_new_n37038__, new_new_n37039__, new_new_n37040__, new_new_n37041__,
    new_new_n37042__, new_new_n37043__, new_new_n37044__, new_new_n37045__,
    new_new_n37046__, new_new_n37047__, new_new_n37049__, new_new_n37050__,
    new_new_n37051__, new_new_n37052__, new_new_n37053__, new_new_n37054__,
    new_new_n37055__, new_new_n37056__, new_new_n37057__, new_new_n37058__,
    new_new_n37059__, new_new_n37060__, new_new_n37061__, new_new_n37062__,
    new_new_n37064__, new_new_n37065__, new_new_n37066__, new_new_n37067__,
    new_new_n37068__, new_new_n37069__, new_new_n37070__, new_new_n37071__,
    new_new_n37072__, new_new_n37073__, new_new_n37074__, new_new_n37075__,
    new_new_n37076__, new_new_n37077__, new_new_n37079__, new_new_n37080__,
    new_new_n37081__, new_new_n37082__, new_new_n37083__, new_new_n37084__,
    new_new_n37085__, new_new_n37086__, new_new_n37087__, new_new_n37088__,
    new_new_n37089__, new_new_n37090__, new_new_n37091__, new_new_n37092__,
    new_new_n37094__, new_new_n37095__, new_new_n37096__, new_new_n37097__,
    new_new_n37098__, new_new_n37099__, new_new_n37100__, new_new_n37101__,
    new_new_n37102__, new_new_n37103__, new_new_n37104__, new_new_n37105__,
    new_new_n37106__, new_new_n37107__, new_new_n37109__, new_new_n37110__,
    new_new_n37111__, new_new_n37112__, new_new_n37113__, new_new_n37114__,
    new_new_n37115__, new_new_n37116__, new_new_n37117__, new_new_n37119__,
    new_new_n37120__, new_new_n37124__, new_new_n37125__, new_new_n37126__,
    new_new_n37127__, new_new_n37128__, new_new_n37137__, new_new_n37139__,
    new_new_n37140__, new_new_n37142__, new_new_n37143__, new_new_n37144__,
    new_new_n37145__, new_new_n37147__, new_new_n37148__, new_new_n37150__,
    new_new_n37151__, new_new_n37152__, new_new_n37153__, new_new_n37154__,
    new_new_n37155__, new_new_n37156__, new_new_n37157__, new_new_n37158__,
    new_new_n37159__, new_new_n37161__, new_new_n37162__, new_new_n37163__,
    new_new_n37164__, new_new_n37165__, new_new_n37166__, new_new_n37167__,
    new_new_n37169__, new_new_n37170__, new_new_n37171__, new_new_n37172__,
    new_new_n37173__, new_new_n37174__, new_new_n37175__, new_new_n37177__,
    new_new_n37178__, new_new_n37179__, new_new_n37180__, new_new_n37181__,
    new_new_n37182__, new_new_n37183__, new_new_n37185__, new_new_n37186__,
    new_new_n37187__, new_new_n37188__, new_new_n37189__, new_new_n37190__,
    new_new_n37191__, new_new_n37193__, new_new_n37194__, new_new_n37195__,
    new_new_n37196__, new_new_n37197__, new_new_n37198__, new_new_n37199__,
    new_new_n37201__, new_new_n37202__, new_new_n37203__, new_new_n37204__,
    new_new_n37205__, new_new_n37206__, new_new_n37207__, new_new_n37209__,
    new_new_n37210__, new_new_n37211__, new_new_n37212__, new_new_n37213__,
    new_new_n37214__, new_new_n37215__, new_new_n37217__, new_new_n37218__,
    new_new_n37219__, new_new_n37220__, new_new_n37221__, new_new_n37222__,
    new_new_n37223__, new_new_n37225__, new_new_n37226__, new_new_n37227__,
    new_new_n37228__, new_new_n37229__, new_new_n37230__, new_new_n37231__,
    new_new_n37233__, new_new_n37234__, new_new_n37235__, new_new_n37236__,
    new_new_n37237__, new_new_n37238__, new_new_n37239__, new_new_n37241__,
    new_new_n37242__, new_new_n37243__, new_new_n37244__, new_new_n37245__,
    new_new_n37246__, new_new_n37247__, new_new_n37249__, new_new_n37250__,
    new_new_n37251__, new_new_n37252__, new_new_n37253__, new_new_n37254__,
    new_new_n37255__, new_new_n37257__, new_new_n37258__, new_new_n37259__,
    new_new_n37260__, new_new_n37261__, new_new_n37262__, new_new_n37263__,
    new_new_n37265__, new_new_n37266__, new_new_n37267__, new_new_n37268__,
    new_new_n37269__, new_new_n37270__, new_new_n37271__, new_new_n37273__,
    new_new_n37274__, new_new_n37275__, new_new_n37276__, new_new_n37277__,
    new_new_n37278__, new_new_n37279__, new_new_n37281__, new_new_n37282__,
    new_new_n37283__, new_new_n37284__, new_new_n37285__, new_new_n37286__,
    new_new_n37287__, new_new_n37289__, new_new_n37290__, new_new_n37291__,
    new_new_n37292__, new_new_n37293__, new_new_n37294__, new_new_n37295__,
    new_new_n37297__, new_new_n37298__, new_new_n37299__, new_new_n37300__,
    new_new_n37301__, new_new_n37302__, new_new_n37303__, new_new_n37305__,
    new_new_n37306__, new_new_n37307__, new_new_n37308__, new_new_n37309__,
    new_new_n37310__, new_new_n37311__, new_new_n37313__, new_new_n37314__,
    new_new_n37315__, new_new_n37316__, new_new_n37317__, new_new_n37318__,
    new_new_n37319__, new_new_n37321__, new_new_n37322__, new_new_n37323__,
    new_new_n37324__, new_new_n37325__, new_new_n37326__, new_new_n37327__,
    new_new_n37329__, new_new_n37330__, new_new_n37331__, new_new_n37332__,
    new_new_n37333__, new_new_n37334__, new_new_n37335__, new_new_n37337__,
    new_new_n37338__, new_new_n37339__, new_new_n37340__, new_new_n37341__,
    new_new_n37342__, new_new_n37343__, new_new_n37345__, new_new_n37346__,
    new_new_n37347__, new_new_n37348__, new_new_n37349__, new_new_n37350__,
    new_new_n37351__, new_new_n37353__, new_new_n37354__, new_new_n37355__,
    new_new_n37356__, new_new_n37357__, new_new_n37358__, new_new_n37359__,
    new_new_n37361__, new_new_n37362__, new_new_n37363__, new_new_n37364__,
    new_new_n37365__, new_new_n37366__, new_new_n37367__, new_new_n37369__,
    new_new_n37370__, new_new_n37371__, new_new_n37372__, new_new_n37373__,
    new_new_n37374__, new_new_n37375__, new_new_n37377__, new_new_n37378__,
    new_new_n37379__, new_new_n37380__, new_new_n37381__, new_new_n37382__,
    new_new_n37383__, new_new_n37385__, new_new_n37386__, new_new_n37387__,
    new_new_n37388__, new_new_n37389__, new_new_n37390__, new_new_n37391__,
    new_new_n37393__, new_new_n37394__, new_new_n37395__, new_new_n37396__,
    new_new_n37397__, new_new_n37398__, new_new_n37399__, new_new_n37401__,
    new_new_n37402__, new_new_n37403__, new_new_n37404__, new_new_n37405__,
    new_new_n37406__, new_new_n37407__, new_new_n37409__, new_new_n37410__,
    new_new_n37411__, new_new_n37412__, new_new_n37413__, new_new_n37414__,
    new_new_n37415__, new_new_n37416__, new_new_n37418__, new_new_n37419__,
    new_new_n37423__, new_new_n37424__, new_new_n37425__, new_new_n37426__,
    new_new_n37435__, new_new_n37437__, new_new_n37438__, new_new_n37440__,
    new_new_n37441__, new_new_n37442__, new_new_n37443__, new_new_n37445__,
    new_new_n37446__, new_new_n37448__, new_new_n37449__, new_new_n37450__,
    new_new_n37451__, new_new_n37452__, new_new_n37453__, new_new_n37454__,
    new_new_n37455__, new_new_n37456__, new_new_n37457__, new_new_n37459__,
    new_new_n37460__, new_new_n37461__, new_new_n37462__, new_new_n37463__,
    new_new_n37464__, new_new_n37465__, new_new_n37467__, new_new_n37468__,
    new_new_n37469__, new_new_n37470__, new_new_n37471__, new_new_n37472__,
    new_new_n37473__, new_new_n37475__, new_new_n37476__, new_new_n37477__,
    new_new_n37478__, new_new_n37479__, new_new_n37480__, new_new_n37481__,
    new_new_n37483__, new_new_n37484__, new_new_n37485__, new_new_n37486__,
    new_new_n37487__, new_new_n37488__, new_new_n37489__, new_new_n37491__,
    new_new_n37492__, new_new_n37493__, new_new_n37494__, new_new_n37495__,
    new_new_n37496__, new_new_n37497__, new_new_n37499__, new_new_n37500__,
    new_new_n37501__, new_new_n37502__, new_new_n37503__, new_new_n37504__,
    new_new_n37505__, new_new_n37507__, new_new_n37508__, new_new_n37509__,
    new_new_n37510__, new_new_n37511__, new_new_n37512__, new_new_n37513__,
    new_new_n37515__, new_new_n37516__, new_new_n37517__, new_new_n37518__,
    new_new_n37519__, new_new_n37520__, new_new_n37521__, new_new_n37523__,
    new_new_n37524__, new_new_n37525__, new_new_n37526__, new_new_n37527__,
    new_new_n37528__, new_new_n37529__, new_new_n37531__, new_new_n37532__,
    new_new_n37533__, new_new_n37534__, new_new_n37535__, new_new_n37536__,
    new_new_n37537__, new_new_n37539__, new_new_n37540__, new_new_n37541__,
    new_new_n37542__, new_new_n37543__, new_new_n37544__, new_new_n37545__,
    new_new_n37547__, new_new_n37548__, new_new_n37549__, new_new_n37550__,
    new_new_n37551__, new_new_n37552__, new_new_n37553__, new_new_n37555__,
    new_new_n37556__, new_new_n37557__, new_new_n37558__, new_new_n37559__,
    new_new_n37560__, new_new_n37561__, new_new_n37563__, new_new_n37564__,
    new_new_n37565__, new_new_n37566__, new_new_n37567__, new_new_n37568__,
    new_new_n37569__, new_new_n37571__, new_new_n37572__, new_new_n37573__,
    new_new_n37574__, new_new_n37575__, new_new_n37576__, new_new_n37577__,
    new_new_n37579__, new_new_n37580__, new_new_n37581__, new_new_n37582__,
    new_new_n37583__, new_new_n37584__, new_new_n37585__, new_new_n37587__,
    new_new_n37588__, new_new_n37589__, new_new_n37590__, new_new_n37591__,
    new_new_n37592__, new_new_n37593__, new_new_n37595__, new_new_n37596__,
    new_new_n37597__, new_new_n37598__, new_new_n37599__, new_new_n37600__,
    new_new_n37601__, new_new_n37603__, new_new_n37604__, new_new_n37605__,
    new_new_n37606__, new_new_n37607__, new_new_n37608__, new_new_n37609__,
    new_new_n37611__, new_new_n37612__, new_new_n37613__, new_new_n37614__,
    new_new_n37615__, new_new_n37616__, new_new_n37617__, new_new_n37619__,
    new_new_n37620__, new_new_n37621__, new_new_n37622__, new_new_n37623__,
    new_new_n37624__, new_new_n37625__, new_new_n37627__, new_new_n37628__,
    new_new_n37629__, new_new_n37630__, new_new_n37631__, new_new_n37632__,
    new_new_n37633__, new_new_n37635__, new_new_n37636__, new_new_n37637__,
    new_new_n37638__, new_new_n37639__, new_new_n37640__, new_new_n37641__,
    new_new_n37643__, new_new_n37644__, new_new_n37645__, new_new_n37646__,
    new_new_n37647__, new_new_n37648__, new_new_n37649__, new_new_n37651__,
    new_new_n37652__, new_new_n37653__, new_new_n37654__, new_new_n37655__,
    new_new_n37656__, new_new_n37657__, new_new_n37659__, new_new_n37660__,
    new_new_n37661__, new_new_n37662__, new_new_n37663__, new_new_n37664__,
    new_new_n37665__, new_new_n37667__, new_new_n37668__, new_new_n37669__,
    new_new_n37670__, new_new_n37671__, new_new_n37672__, new_new_n37673__,
    new_new_n37675__, new_new_n37676__, new_new_n37677__, new_new_n37678__,
    new_new_n37679__, new_new_n37680__, new_new_n37681__, new_new_n37683__,
    new_new_n37684__, new_new_n37685__, new_new_n37686__, new_new_n37687__,
    new_new_n37688__, new_new_n37689__, new_new_n37691__, new_new_n37692__,
    new_new_n37693__, new_new_n37694__, new_new_n37695__, new_new_n37696__,
    new_new_n37697__, new_new_n37699__, new_new_n37700__, new_new_n37701__,
    new_new_n37702__, new_new_n37703__, new_new_n37704__, new_new_n37705__,
    new_new_n37707__, new_new_n37708__, new_new_n37709__, new_new_n37710__,
    new_new_n37711__, new_new_n37712__, new_new_n37713__, new_new_n37714__,
    new_new_n37716__, new_new_n37717__, new_new_n37721__, new_new_n37722__,
    new_new_n37723__, new_new_n37724__, new_new_n37733__, new_new_n37735__,
    new_new_n37736__, new_new_n37738__, new_new_n37739__, new_new_n37740__,
    new_new_n37741__, new_new_n37743__, new_new_n37744__, new_new_n37746__,
    new_new_n37747__, new_new_n37749__, new_new_n37750__, new_new_n37752__,
    new_new_n37754__, new_new_n37755__, new_new_n37757__, new_new_n37758__,
    new_new_n37760__, new_new_n37761__, new_new_n37763__, new_new_n37764__,
    new_new_n37766__, new_new_n37767__, new_new_n37769__, new_new_n37770__,
    new_new_n37772__, new_new_n37773__, new_new_n37775__, new_new_n37776__,
    new_new_n37778__, new_new_n37779__, new_new_n37781__, new_new_n37782__,
    new_new_n37784__, new_new_n37785__, new_new_n37787__, new_new_n37788__,
    new_new_n37790__, new_new_n37791__, new_new_n37793__, new_new_n37794__,
    new_new_n37796__, new_new_n37797__, new_new_n37799__, new_new_n37800__,
    new_new_n37802__, new_new_n37803__, new_new_n37805__, new_new_n37806__,
    new_new_n37808__, new_new_n37809__, new_new_n37811__, new_new_n37812__,
    new_new_n37814__, new_new_n37815__, new_new_n37817__, new_new_n37818__,
    new_new_n37820__, new_new_n37821__, new_new_n37823__, new_new_n37824__,
    new_new_n37826__, new_new_n37827__, new_new_n37829__, new_new_n37830__,
    new_new_n37832__, new_new_n37833__, new_new_n37835__, new_new_n37836__,
    new_new_n37838__, new_new_n37839__, new_new_n37841__, new_new_n37842__,
    new_new_n37844__, new_new_n37845__, new_new_n37847__, new_new_n37848__,
    new_new_n37849__, new_new_n37850__, new_new_n37851__, new_new_n37852__,
    new_new_n37854__, new_new_n37855__, new_new_n37856__, new_new_n37857__,
    new_new_n37858__, new_new_n37860__, new_new_n37861__, new_new_n37862__,
    new_new_n37863__, new_new_n37864__, new_new_n37866__, new_new_n37867__,
    new_new_n37868__, new_new_n37869__, new_new_n37870__, new_new_n37872__,
    new_new_n37873__, new_new_n37874__, new_new_n37875__, new_new_n37876__,
    new_new_n37878__, new_new_n37879__, new_new_n37880__, new_new_n37881__,
    new_new_n37882__, new_new_n37884__, new_new_n37885__, new_new_n37886__,
    new_new_n37887__, new_new_n37888__, new_new_n37890__, new_new_n37891__,
    new_new_n37892__, new_new_n37893__, new_new_n37894__, new_new_n37896__,
    new_new_n37897__, new_new_n37898__, new_new_n37899__, new_new_n37900__,
    new_new_n37902__, new_new_n37903__, new_new_n37904__, new_new_n37905__,
    new_new_n37906__, new_new_n37908__, new_new_n37909__, new_new_n37910__,
    new_new_n37911__, new_new_n37912__, new_new_n37914__, new_new_n37915__,
    new_new_n37916__, new_new_n37917__, new_new_n37918__, new_new_n37920__,
    new_new_n37921__, new_new_n37922__, new_new_n37923__, new_new_n37924__,
    new_new_n37926__, new_new_n37927__, new_new_n37928__, new_new_n37929__,
    new_new_n37930__, new_new_n37932__, new_new_n37933__, new_new_n37934__,
    new_new_n37935__, new_new_n37936__, new_new_n37938__, new_new_n37939__,
    new_new_n37940__, new_new_n37941__, new_new_n37942__, new_new_n37944__,
    new_new_n37945__, new_new_n37946__, new_new_n37947__, new_new_n37948__,
    new_new_n37950__, new_new_n37951__, new_new_n37952__, new_new_n37953__,
    new_new_n37954__, new_new_n37956__, new_new_n37957__, new_new_n37958__,
    new_new_n37959__, new_new_n37960__, new_new_n37962__, new_new_n37963__,
    new_new_n37964__, new_new_n37965__, new_new_n37966__, new_new_n37968__,
    new_new_n37969__, new_new_n37970__, new_new_n37971__, new_new_n37972__,
    new_new_n37974__, new_new_n37975__, new_new_n37976__, new_new_n37977__,
    new_new_n37978__, new_new_n37980__, new_new_n37981__, new_new_n37982__,
    new_new_n37983__, new_new_n37984__, new_new_n37986__, new_new_n37987__,
    new_new_n37988__, new_new_n37989__, new_new_n37990__, new_new_n37992__,
    new_new_n37993__, new_new_n37994__, new_new_n37995__, new_new_n37996__,
    new_new_n37998__, new_new_n37999__, new_new_n38000__, new_new_n38001__,
    new_new_n38002__, new_new_n38004__, new_new_n38005__, new_new_n38006__,
    new_new_n38007__, new_new_n38008__, new_new_n38010__, new_new_n38011__,
    new_new_n38012__, new_new_n38013__, new_new_n38014__, new_new_n38016__,
    new_new_n38017__, new_new_n38018__, new_new_n38019__, new_new_n38020__,
    new_new_n38022__, new_new_n38023__, new_new_n38024__, new_new_n38025__,
    new_new_n38026__, new_new_n38028__, new_new_n38029__, new_new_n38030__,
    new_new_n38031__, new_new_n38032__, new_new_n38034__, new_new_n38035__,
    new_new_n38036__, new_new_n38037__, new_new_n38038__, new_new_n38040__,
    new_new_n38041__, new_new_n38042__, new_new_n38045__, new_new_n38047__,
    new_new_n38048__, new_new_n38049__, new_new_n38050__, new_new_n38051__,
    new_new_n38052__, new_new_n38053__, new_new_n38054__, new_new_n38055__,
    new_new_n38056__, new_new_n38057__, new_new_n38058__, new_new_n38059__,
    new_new_n38060__, new_new_n38061__, new_new_n38062__, new_new_n38063__,
    new_new_n38064__, new_new_n38065__, new_new_n38066__, new_new_n38067__,
    new_new_n38068__, new_new_n38069__, new_new_n38070__, new_new_n38071__,
    new_new_n38072__, new_new_n38073__, new_new_n38074__, new_new_n38075__,
    new_new_n38076__, new_new_n38077__, new_new_n38078__, new_new_n38079__,
    new_new_n38080__, new_new_n38081__, new_new_n38082__, new_new_n38083__,
    new_new_n38084__, new_new_n38085__, new_new_n38086__, new_new_n38087__,
    new_new_n38088__, new_new_n38089__, new_new_n38090__, new_new_n38091__,
    new_new_n38092__, new_new_n38093__, new_new_n38094__, new_new_n38095__,
    new_new_n38096__, new_new_n38097__, new_new_n38098__, new_new_n38099__,
    new_new_n38100__, new_new_n38101__, new_new_n38102__, new_new_n38103__,
    new_new_n38104__, new_new_n38105__, new_new_n38106__, new_new_n38107__,
    new_new_n38108__, new_new_n38109__, new_new_n38110__, new_new_n38111__,
    new_new_n38112__, new_new_n38113__, new_new_n38114__, new_new_n38115__,
    new_new_n38116__, new_new_n38117__, new_new_n38118__, new_new_n38119__,
    new_new_n38120__, new_new_n38121__, new_new_n38122__, new_new_n38123__,
    new_new_n38124__, new_new_n38125__, new_new_n38126__, new_new_n38127__,
    new_new_n38128__, new_new_n38129__, new_new_n38130__, new_new_n38131__,
    new_new_n38132__, new_new_n38133__, new_new_n38134__, new_new_n38135__,
    new_new_n38136__, new_new_n38137__, new_new_n38138__, new_new_n38139__,
    new_new_n38140__, new_new_n38141__, new_new_n38142__, new_new_n38143__,
    new_new_n38144__, new_new_n38145__, new_new_n38146__, new_new_n38147__,
    new_new_n38148__, new_new_n38149__, new_new_n38150__, new_new_n38151__,
    new_new_n38152__, new_new_n38153__, new_new_n38154__, new_new_n38155__,
    new_new_n38156__, new_new_n38157__, new_new_n38158__, new_new_n38159__,
    new_new_n38160__, new_new_n38161__, new_new_n38162__, new_new_n38163__,
    new_new_n38164__, new_new_n38165__, new_new_n38166__, new_new_n38167__,
    new_new_n38168__, new_new_n38169__, new_new_n38170__, new_new_n38171__,
    new_new_n38172__, new_new_n38173__, new_new_n38174__, new_new_n38175__,
    new_new_n38176__, new_new_n38177__, new_new_n38178__, new_new_n38179__,
    new_new_n38180__, new_new_n38181__, new_new_n38182__, new_new_n38183__,
    new_new_n38184__, new_new_n38185__, new_new_n38186__, new_new_n38187__,
    new_new_n38188__, new_new_n38189__, new_new_n38190__, new_new_n38191__,
    new_new_n38192__, new_new_n38193__, new_new_n38194__, new_new_n38195__,
    new_new_n38196__, new_new_n38197__, new_new_n38198__, new_new_n38199__,
    new_new_n38200__, new_new_n38201__, new_new_n38202__, new_new_n38203__,
    new_new_n38204__, new_new_n38205__, new_new_n38206__, new_new_n38207__,
    new_new_n38208__, new_new_n38209__, new_new_n38210__, new_new_n38211__,
    new_new_n38212__, new_new_n38213__, new_new_n38214__, new_new_n38215__,
    new_new_n38216__, new_new_n38217__, new_new_n38218__, new_new_n38219__,
    new_new_n38220__, new_new_n38221__, new_new_n38222__, new_new_n38223__,
    new_new_n38224__, new_new_n38225__, new_new_n38226__, new_new_n38227__,
    new_new_n38228__, new_new_n38229__, new_new_n38230__, new_new_n38231__,
    new_new_n38232__, new_new_n38233__, new_new_n38234__, new_new_n38235__,
    new_new_n38236__, new_new_n38237__, new_new_n38238__, new_new_n38239__,
    new_new_n38240__, new_new_n38241__, new_new_n38242__, new_new_n38243__,
    new_new_n38244__, new_new_n38245__, new_new_n38246__, new_new_n38247__,
    new_new_n38248__, new_new_n38249__, new_new_n38250__, new_new_n38251__,
    new_new_n38252__, new_new_n38253__, new_new_n38254__, new_new_n38255__,
    new_new_n38256__, new_new_n38257__, new_new_n38258__, new_new_n38259__,
    new_new_n38260__, new_new_n38261__, new_new_n38262__, new_new_n38263__,
    new_new_n38264__, new_new_n38265__, new_new_n38266__, new_new_n38267__,
    new_new_n38268__, new_new_n38269__, new_new_n38270__, new_new_n38271__,
    new_new_n38272__, new_new_n38273__, new_new_n38274__, new_new_n38275__,
    new_new_n38276__, new_new_n38277__, new_new_n38278__, new_new_n38279__,
    new_new_n38280__, new_new_n38281__, new_new_n38282__, new_new_n38283__,
    new_new_n38284__, new_new_n38285__, new_new_n38286__, new_new_n38287__,
    new_new_n38288__, new_new_n38289__, new_new_n38290__, new_new_n38291__,
    new_new_n38292__, new_new_n38293__, new_new_n38294__, new_new_n38295__,
    new_new_n38296__, new_new_n38297__, new_new_n38298__, new_new_n38299__,
    new_new_n38300__, new_new_n38301__, new_new_n38302__, new_new_n38303__,
    new_new_n38304__, new_new_n38305__, new_new_n38306__, new_new_n38307__,
    new_new_n38308__, new_new_n38309__, new_new_n38310__, new_new_n38311__,
    new_new_n38312__, new_new_n38313__, new_new_n38314__, new_new_n38315__,
    new_new_n38316__, new_new_n38317__, new_new_n38318__, new_new_n38319__,
    new_new_n38320__, new_new_n38321__, new_new_n38322__, new_new_n38323__,
    new_new_n38324__, new_new_n38325__, new_new_n38326__, new_new_n38327__,
    new_new_n38328__, new_new_n38329__, new_new_n38330__, new_new_n38331__,
    new_new_n38332__, new_new_n38333__, new_new_n38334__, new_new_n38335__,
    new_new_n38336__, new_new_n38337__, new_new_n38338__, new_new_n38339__,
    new_new_n38340__, new_new_n38341__, new_new_n38342__, new_new_n38343__,
    new_new_n38344__, new_new_n38345__, new_new_n38346__, new_new_n38347__,
    new_new_n38348__, new_new_n38349__, new_new_n38350__, new_new_n38351__,
    new_new_n38352__, new_new_n38353__, new_new_n38354__, new_new_n38355__,
    new_new_n38356__, new_new_n38357__, new_new_n38358__, new_new_n38359__,
    new_new_n38360__, new_new_n38361__, new_new_n38362__, new_new_n38363__,
    new_new_n38364__, new_new_n38365__, new_new_n38366__, new_new_n38367__,
    new_new_n38368__, new_new_n38369__, new_new_n38370__, new_new_n38371__,
    new_new_n38372__, new_new_n38373__, new_new_n38374__, new_new_n38375__,
    new_new_n38376__, new_new_n38377__, new_new_n38378__, new_new_n38379__,
    new_new_n38380__, new_new_n38381__, new_new_n38382__, new_new_n38383__,
    new_new_n38384__, new_new_n38385__, new_new_n38386__, new_new_n38387__,
    new_new_n38388__, new_new_n38389__, new_new_n38390__, new_new_n38391__,
    new_new_n38392__, new_new_n38393__, new_new_n38394__, new_new_n38395__,
    new_new_n38396__, new_new_n38397__, new_new_n38398__, new_new_n38399__,
    new_new_n38400__, new_new_n38401__, new_new_n38402__, new_new_n38403__,
    new_new_n38404__, new_new_n38405__, new_new_n38406__, new_new_n38407__,
    new_new_n38408__, new_new_n38409__, new_new_n38410__, new_new_n38411__,
    new_new_n38412__, new_new_n38413__, new_new_n38414__, new_new_n38415__,
    new_new_n38416__, new_new_n38417__, new_new_n38418__, new_new_n38419__,
    new_new_n38420__, new_new_n38421__, new_new_n38422__, new_new_n38423__,
    new_new_n38424__, new_new_n38425__, new_new_n38426__, new_new_n38427__,
    new_new_n38428__, new_new_n38429__, new_new_n38430__, new_new_n38431__,
    new_new_n38432__, new_new_n38433__, new_new_n38434__, new_new_n38435__,
    new_new_n38436__, new_new_n38437__, new_new_n38438__, new_new_n38439__,
    new_new_n38440__, new_new_n38441__, new_new_n38442__, new_new_n38443__,
    new_new_n38444__, new_new_n38445__, new_new_n38446__, new_new_n38447__,
    new_new_n38448__, new_new_n38449__, new_new_n38450__, new_new_n38451__,
    new_new_n38452__, new_new_n38453__, new_new_n38454__, new_new_n38455__,
    new_new_n38456__, new_new_n38457__, new_new_n38458__, new_new_n38459__,
    new_new_n38460__, new_new_n38461__, new_new_n38462__, new_new_n38463__,
    new_new_n38464__, new_new_n38465__, new_new_n38466__, new_new_n38467__,
    new_new_n38468__, new_new_n38469__, new_new_n38470__, new_new_n38471__,
    new_new_n38472__, new_new_n38473__, new_new_n38474__, new_new_n38475__,
    new_new_n38476__, new_new_n38477__, new_new_n38478__, new_new_n38479__,
    new_new_n38480__, new_new_n38481__, new_new_n38482__, new_new_n38483__,
    new_new_n38484__, new_new_n38485__, new_new_n38486__, new_new_n38487__,
    new_new_n38488__, new_new_n38489__, new_new_n38490__, new_new_n38491__,
    new_new_n38492__, new_new_n38493__, new_new_n38494__, new_new_n38495__,
    new_new_n38496__, new_new_n38497__, new_new_n38498__, new_new_n38499__,
    new_new_n38500__, new_new_n38501__, new_new_n38502__, new_new_n38503__,
    new_new_n38504__, new_new_n38505__, new_new_n38506__, new_new_n38507__,
    new_new_n38508__, new_new_n38509__, new_new_n38510__, new_new_n38511__,
    new_new_n38512__, new_new_n38513__, new_new_n38514__, new_new_n38515__,
    new_new_n38516__, new_new_n38517__, new_new_n38518__, new_new_n38519__,
    new_new_n38520__, new_new_n38521__, new_new_n38522__, new_new_n38523__,
    new_new_n38524__, new_new_n38525__, new_new_n38526__, new_new_n38527__,
    new_new_n38528__, new_new_n38529__, new_new_n38530__, new_new_n38531__,
    new_new_n38532__, new_new_n38533__, new_new_n38534__, new_new_n38535__,
    new_new_n38536__, new_new_n38537__, new_new_n38538__, new_new_n38539__,
    new_new_n38540__, new_new_n38541__, new_new_n38542__, new_new_n38543__,
    new_new_n38544__, new_new_n38545__, new_new_n38546__, new_new_n38547__,
    new_new_n38548__, new_new_n38549__, new_new_n38550__, new_new_n38551__,
    new_new_n38552__, new_new_n38553__, new_new_n38554__, new_new_n38555__,
    new_new_n38556__, new_new_n38557__, new_new_n38558__, new_new_n38559__,
    new_new_n38560__, new_new_n38561__, new_new_n38562__, new_new_n38563__,
    new_new_n38564__, new_new_n38565__, new_new_n38566__, new_new_n38567__,
    new_new_n38568__, new_new_n38569__, new_new_n38570__, new_new_n38571__,
    new_new_n38572__, new_new_n38573__, new_new_n38574__, new_new_n38575__,
    new_new_n38576__, new_new_n38577__, new_new_n38578__, new_new_n38579__,
    new_new_n38580__, new_new_n38581__, new_new_n38582__, new_new_n38583__,
    new_new_n38584__, new_new_n38585__, new_new_n38586__, new_new_n38587__,
    new_new_n38588__, new_new_n38589__, new_new_n38590__, new_new_n38591__,
    new_new_n38592__, new_new_n38593__, new_new_n38594__, new_new_n38595__,
    new_new_n38596__, new_new_n38597__, new_new_n38598__, new_new_n38599__,
    new_new_n38600__, new_new_n38601__, new_new_n38602__, new_new_n38603__,
    new_new_n38604__, new_new_n38605__, new_new_n38606__, new_new_n38607__,
    new_new_n38608__, new_new_n38609__, new_new_n38610__, new_new_n38611__,
    new_new_n38612__, new_new_n38613__, new_new_n38614__, new_new_n38615__,
    new_new_n38616__, new_new_n38617__, new_new_n38618__, new_new_n38619__,
    new_new_n38620__, new_new_n38621__, new_new_n38622__, new_new_n38623__,
    new_new_n38624__, new_new_n38625__, new_new_n38626__, new_new_n38627__,
    new_new_n38628__, new_new_n38629__, new_new_n38630__, new_new_n38631__,
    new_new_n38632__, new_new_n38633__, new_new_n38634__, new_new_n38635__,
    new_new_n38636__, new_new_n38637__, new_new_n38638__, new_new_n38639__,
    new_new_n38640__, new_new_n38641__, new_new_n38642__, new_new_n38643__,
    new_new_n38644__, new_new_n38645__, new_new_n38646__, new_new_n38647__,
    new_new_n38648__, new_new_n38649__, new_new_n38650__, new_new_n38651__,
    new_new_n38652__, new_new_n38653__, new_new_n38654__, new_new_n38655__,
    new_new_n38656__, new_new_n38657__, new_new_n38658__, new_new_n38659__,
    new_new_n38660__, new_new_n38661__, new_new_n38662__, new_new_n38663__,
    new_new_n38664__, new_new_n38665__, new_new_n38666__, new_new_n38667__,
    new_new_n38668__, new_new_n38669__, new_new_n38670__, new_new_n38671__,
    new_new_n38672__, new_new_n38673__, new_new_n38674__, new_new_n38675__,
    new_new_n38676__, new_new_n38677__, new_new_n38678__, new_new_n38679__,
    new_new_n38680__, new_new_n38681__, new_new_n38682__, new_new_n38683__,
    new_new_n38684__, new_new_n38685__, new_new_n38686__, new_new_n38687__,
    new_new_n38688__, new_new_n38689__, new_new_n38690__, new_new_n38691__,
    new_new_n38692__, new_new_n38693__, new_new_n38694__, new_new_n38695__,
    new_new_n38696__, new_new_n38697__, new_new_n38698__, new_new_n38699__,
    new_new_n38700__, new_new_n38701__, new_new_n38702__, new_new_n38703__,
    new_new_n38704__, new_new_n38705__, new_new_n38706__, new_new_n38707__,
    new_new_n38708__, new_new_n38709__, new_new_n38710__, new_new_n38711__,
    new_new_n38712__, new_new_n38713__, new_new_n38714__, new_new_n38715__,
    new_new_n38716__, new_new_n38717__, new_new_n38718__, new_new_n38719__,
    new_new_n38720__, new_new_n38721__, new_new_n38722__, new_new_n38723__,
    new_new_n38724__, new_new_n38725__, new_new_n38726__, new_new_n38727__,
    new_new_n38728__, new_new_n38729__, new_new_n38730__, new_new_n38731__,
    new_new_n38732__, new_new_n38733__, new_new_n38734__, new_new_n38735__,
    new_new_n38736__, new_new_n38737__, new_new_n38738__, new_new_n38739__,
    new_new_n38740__, new_new_n38741__, new_new_n38742__, new_new_n38743__,
    new_new_n38744__, new_new_n38745__, new_new_n38746__, new_new_n38747__,
    new_new_n38748__, new_new_n38749__, new_new_n38750__, new_new_n38751__,
    new_new_n38752__, new_new_n38753__, new_new_n38754__, new_new_n38755__,
    new_new_n38756__, new_new_n38757__, new_new_n38758__, new_new_n38759__,
    new_new_n38760__, new_new_n38761__, new_new_n38762__, new_new_n38763__,
    new_new_n38764__, new_new_n38765__, new_new_n38766__, new_new_n38767__,
    new_new_n38768__, new_new_n38769__, new_new_n38770__, new_new_n38771__,
    new_new_n38772__, new_new_n38773__, new_new_n38774__, new_new_n38775__,
    new_new_n38776__, new_new_n38777__, new_new_n38778__, new_new_n38779__,
    new_new_n38780__, new_new_n38781__, new_new_n38782__, new_new_n38783__,
    new_new_n38784__, new_new_n38785__, new_new_n38786__, new_new_n38787__,
    new_new_n38788__, new_new_n38789__, new_new_n38790__, new_new_n38791__,
    new_new_n38792__, new_new_n38793__, new_new_n38794__, new_new_n38795__,
    new_new_n38796__, new_new_n38797__, new_new_n38798__, new_new_n38799__,
    new_new_n38800__, new_new_n38801__, new_new_n38802__, new_new_n38803__,
    new_new_n38804__, new_new_n38805__, new_new_n38806__, new_new_n38807__,
    new_new_n38808__, new_new_n38809__, new_new_n38810__, new_new_n38811__,
    new_new_n38812__, new_new_n38813__, new_new_n38814__, new_new_n38815__,
    new_new_n38816__, new_new_n38817__, new_new_n38818__, new_new_n38819__,
    new_new_n38820__, new_new_n38821__, new_new_n38822__, new_new_n38823__,
    new_new_n38824__, new_new_n38825__, new_new_n38826__, new_new_n38827__,
    new_new_n38828__, new_new_n38829__, new_new_n38830__, new_new_n38831__,
    new_new_n38832__, new_new_n38833__, new_new_n38834__, new_new_n38835__,
    new_new_n38836__, new_new_n38837__, new_new_n38838__, new_new_n38839__,
    new_new_n38840__, new_new_n38841__, new_new_n38842__, new_new_n38843__,
    new_new_n38844__, new_new_n38845__, new_new_n38846__, new_new_n38847__,
    new_new_n38848__, new_new_n38849__, new_new_n38850__, new_new_n38851__,
    new_new_n38852__, new_new_n38853__, new_new_n38854__, new_new_n38855__,
    new_new_n38856__, new_new_n38857__, new_new_n38858__, new_new_n38859__,
    new_new_n38860__, new_new_n38861__, new_new_n38862__, new_new_n38863__,
    new_new_n38864__, new_new_n38865__, new_new_n38866__, new_new_n38867__,
    new_new_n38868__, new_new_n38869__, new_new_n38870__, new_new_n38871__,
    new_new_n38872__, new_new_n38873__, new_new_n38874__, new_new_n38875__,
    new_new_n38876__, new_new_n38877__, new_new_n38878__, new_new_n38879__,
    new_new_n38880__, new_new_n38881__, new_new_n38882__, new_new_n38883__,
    new_new_n38884__, new_new_n38885__, new_new_n38886__, new_new_n38887__,
    new_new_n38888__, new_new_n38889__, new_new_n38890__, new_new_n38891__,
    new_new_n38892__, new_new_n38893__, new_new_n38894__, new_new_n38895__,
    new_new_n38896__, new_new_n38897__, new_new_n38898__, new_new_n38899__,
    new_new_n38900__, new_new_n38901__, new_new_n38902__, new_new_n38903__,
    new_new_n38904__, new_new_n38905__, new_new_n38906__, new_new_n38907__,
    new_new_n38908__, new_new_n38909__, new_new_n38910__, new_new_n38911__,
    new_new_n38912__, new_new_n38913__, new_new_n38914__, new_new_n38915__,
    new_new_n38916__, new_new_n38917__, new_new_n38918__, new_new_n38919__,
    new_new_n38920__, new_new_n38921__, new_new_n38922__, new_new_n38923__,
    new_new_n38924__, new_new_n38925__, new_new_n38926__, new_new_n38927__,
    new_new_n38928__, new_new_n38929__, new_new_n38930__, new_new_n38931__,
    new_new_n38932__, new_new_n38933__, new_new_n38934__, new_new_n38935__,
    new_new_n38936__, new_new_n38937__, new_new_n38938__, new_new_n38939__,
    new_new_n38940__, new_new_n38941__, new_new_n38942__, new_new_n38943__,
    new_new_n38944__, new_new_n38945__, new_new_n38946__, new_new_n38947__,
    new_new_n38948__, new_new_n38949__, new_new_n38950__, new_new_n38951__,
    new_new_n38952__, new_new_n38953__, new_new_n38954__, new_new_n38955__,
    new_new_n38956__, new_new_n38957__, new_new_n38958__, new_new_n38959__,
    new_new_n38960__, new_new_n38961__, new_new_n38962__, new_new_n38963__,
    new_new_n38964__, new_new_n38965__, new_new_n38966__, new_new_n38967__,
    new_new_n38968__, new_new_n38969__, new_new_n38970__, new_new_n38971__,
    new_new_n38972__, new_new_n38973__, new_new_n38974__, new_new_n38975__,
    new_new_n38976__, new_new_n38977__, new_new_n38978__, new_new_n38979__,
    new_new_n38980__, new_new_n38981__, new_new_n38982__, new_new_n38983__,
    new_new_n38984__, new_new_n38985__, new_new_n38986__, new_new_n38987__,
    new_new_n38988__, new_new_n38989__, new_new_n38990__, new_new_n38991__,
    new_new_n38992__, new_new_n38993__, new_new_n38994__, new_new_n38995__,
    new_new_n38996__, new_new_n38997__, new_new_n38998__, new_new_n38999__,
    new_new_n39000__, new_new_n39001__, new_new_n39002__, new_new_n39003__,
    new_new_n39004__, new_new_n39005__, new_new_n39006__, new_new_n39007__,
    new_new_n39008__, new_new_n39009__, new_new_n39010__, new_new_n39011__,
    new_new_n39012__, new_new_n39013__, new_new_n39014__, new_new_n39015__,
    new_new_n39016__, new_new_n39017__, new_new_n39018__, new_new_n39019__,
    new_new_n39020__, new_new_n39021__, new_new_n39022__, new_new_n39023__,
    new_new_n39024__, new_new_n39025__, new_new_n39026__, new_new_n39027__,
    new_new_n39028__, new_new_n39029__, new_new_n39030__, new_new_n39031__,
    new_new_n39032__, new_new_n39033__, new_new_n39034__, new_new_n39035__,
    new_new_n39036__, new_new_n39037__, new_new_n39038__, new_new_n39039__,
    new_new_n39040__, new_new_n39041__, new_new_n39042__, new_new_n39043__,
    new_new_n39044__, new_new_n39045__, new_new_n39046__, new_new_n39047__,
    new_new_n39048__, new_new_n39049__, new_new_n39050__, new_new_n39051__,
    new_new_n39052__, new_new_n39053__, new_new_n39054__, new_new_n39055__,
    new_new_n39056__, new_new_n39057__, new_new_n39058__, new_new_n39059__,
    new_new_n39060__, new_new_n39061__, new_new_n39062__, new_new_n39063__,
    new_new_n39064__, new_new_n39065__, new_new_n39066__, new_new_n39067__,
    new_new_n39068__, new_new_n39069__, new_new_n39070__, new_new_n39071__,
    new_new_n39072__, new_new_n39073__, new_new_n39074__, new_new_n39075__,
    new_new_n39076__, new_new_n39077__, new_new_n39078__, new_new_n39079__,
    new_new_n39080__, new_new_n39081__, new_new_n39082__, new_new_n39083__,
    new_new_n39084__, new_new_n39085__, new_new_n39086__, new_new_n39087__,
    new_new_n39088__, new_new_n39089__, new_new_n39090__, new_new_n39091__,
    new_new_n39092__, new_new_n39093__, new_new_n39094__, new_new_n39095__,
    new_new_n39096__, new_new_n39097__, new_new_n39098__, new_new_n39099__,
    new_new_n39100__, new_new_n39101__, new_new_n39102__, new_new_n39103__,
    new_new_n39104__, new_new_n39105__, new_new_n39106__, new_new_n39107__,
    new_new_n39108__, new_new_n39109__, new_new_n39110__, new_new_n39111__,
    new_new_n39112__, new_new_n39113__, new_new_n39114__, new_new_n39115__,
    new_new_n39116__, new_new_n39117__, new_new_n39118__, new_new_n39119__,
    new_new_n39120__, new_new_n39121__, new_new_n39122__, new_new_n39123__,
    new_new_n39124__, new_new_n39125__, new_new_n39126__, new_new_n39127__,
    new_new_n39128__, new_new_n39129__, new_new_n39130__, new_new_n39131__,
    new_new_n39132__, new_new_n39133__, new_new_n39134__, new_new_n39135__,
    new_new_n39136__, new_new_n39137__, new_new_n39138__, new_new_n39139__,
    new_new_n39140__, new_new_n39141__, new_new_n39142__, new_new_n39143__,
    new_new_n39144__, new_new_n39145__, new_new_n39146__, new_new_n39147__,
    new_new_n39148__, new_new_n39149__, new_new_n39150__, new_new_n39151__,
    new_new_n39152__, new_new_n39153__, new_new_n39154__, new_new_n39155__,
    new_new_n39156__, new_new_n39157__, new_new_n39158__, new_new_n39159__,
    new_new_n39160__, new_new_n39161__, new_new_n39162__, new_new_n39163__,
    new_new_n39164__, new_new_n39165__, new_new_n39166__, new_new_n39167__,
    new_new_n39168__, new_new_n39169__, new_new_n39170__, new_new_n39171__,
    new_new_n39172__, new_new_n39173__, new_new_n39174__, new_new_n39175__,
    new_new_n39176__, new_new_n39177__, new_new_n39178__, new_new_n39179__,
    new_new_n39180__, new_new_n39181__, new_new_n39182__, new_new_n39183__,
    new_new_n39184__, new_new_n39185__, new_new_n39186__, new_new_n39187__,
    new_new_n39188__, new_new_n39189__, new_new_n39190__, new_new_n39191__,
    new_new_n39192__, new_new_n39193__, new_new_n39194__, new_new_n39195__,
    new_new_n39196__, new_new_n39197__, new_new_n39198__, new_new_n39199__,
    new_new_n39200__, new_new_n39201__, new_new_n39202__, new_new_n39203__,
    new_new_n39204__, new_new_n39205__, new_new_n39206__, new_new_n39207__,
    new_new_n39208__, new_new_n39209__, new_new_n39210__, new_new_n39211__,
    new_new_n39212__, new_new_n39213__, new_new_n39214__, new_new_n39215__,
    new_new_n39216__, new_new_n39217__, new_new_n39218__, new_new_n39219__,
    new_new_n39220__, new_new_n39221__, new_new_n39222__, new_new_n39223__,
    new_new_n39224__, new_new_n39225__, new_new_n39226__, new_new_n39227__,
    new_new_n39228__, new_new_n39229__, new_new_n39230__, new_new_n39231__,
    new_new_n39232__, new_new_n39233__, new_new_n39234__, new_new_n39235__,
    new_new_n39236__, new_new_n39237__, new_new_n39238__, new_new_n39239__,
    new_new_n39240__, new_new_n39241__, new_new_n39242__, new_new_n39243__,
    new_new_n39244__, new_new_n39245__, new_new_n39246__, new_new_n39247__,
    new_new_n39248__, new_new_n39249__, new_new_n39250__, new_new_n39251__,
    new_new_n39252__, new_new_n39253__, new_new_n39254__, new_new_n39255__,
    new_new_n39256__, new_new_n39257__, new_new_n39258__, new_new_n39259__,
    new_new_n39260__, new_new_n39261__, new_new_n39262__, new_new_n39263__,
    new_new_n39264__, new_new_n39265__, new_new_n39266__, new_new_n39267__,
    new_new_n39268__, new_new_n39269__, new_new_n39270__, new_new_n39271__,
    new_new_n39272__, new_new_n39273__, new_new_n39274__, new_new_n39275__,
    new_new_n39276__, new_new_n39277__, new_new_n39278__, new_new_n39279__,
    new_new_n39280__, new_new_n39281__, new_new_n39282__, new_new_n39283__,
    new_new_n39284__, new_new_n39285__, new_new_n39286__, new_new_n39287__,
    new_new_n39288__, new_new_n39289__, new_new_n39290__, new_new_n39291__,
    new_new_n39292__, new_new_n39293__, new_new_n39294__, new_new_n39295__,
    new_new_n39296__, new_new_n39297__, new_new_n39298__, new_new_n39299__,
    new_new_n39300__, new_new_n39301__, new_new_n39302__, new_new_n39303__,
    new_new_n39304__, new_new_n39305__, new_new_n39306__, new_new_n39307__,
    new_new_n39308__, new_new_n39309__, new_new_n39310__, new_new_n39311__,
    new_new_n39312__, new_new_n39313__, new_new_n39314__, new_new_n39315__,
    new_new_n39316__, new_new_n39317__, new_new_n39318__, new_new_n39319__,
    new_new_n39320__, new_new_n39321__, new_new_n39322__, new_new_n39323__,
    new_new_n39324__, new_new_n39325__, new_new_n39326__, new_new_n39327__,
    new_new_n39328__, new_new_n39329__, new_new_n39330__, new_new_n39331__,
    new_new_n39332__, new_new_n39333__, new_new_n39334__, new_new_n39335__,
    new_new_n39336__, new_new_n39337__, new_new_n39338__, new_new_n39339__,
    new_new_n39340__, new_new_n39341__, new_new_n39342__, new_new_n39343__,
    new_new_n39344__, new_new_n39345__, new_new_n39346__, new_new_n39347__,
    new_new_n39348__, new_new_n39349__, new_new_n39350__, new_new_n39351__,
    new_new_n39352__, new_new_n39353__, new_new_n39354__, new_new_n39355__,
    new_new_n39356__, new_new_n39357__, new_new_n39358__, new_new_n39359__,
    new_new_n39360__, new_new_n39361__, new_new_n39362__, new_new_n39363__,
    new_new_n39364__, new_new_n39365__, new_new_n39366__, new_new_n39367__,
    new_new_n39368__, new_new_n39369__, new_new_n39370__, new_new_n39371__,
    new_new_n39372__, new_new_n39373__, new_new_n39374__, new_new_n39375__,
    new_new_n39376__, new_new_n39377__, new_new_n39378__, new_new_n39379__,
    new_new_n39380__, new_new_n39381__, new_new_n39382__, new_new_n39383__,
    new_new_n39384__, new_new_n39385__, new_new_n39386__, new_new_n39387__,
    new_new_n39388__, new_new_n39389__, new_new_n39390__, new_new_n39391__,
    new_new_n39392__, new_new_n39393__, new_new_n39394__, new_new_n39395__,
    new_new_n39396__, new_new_n39397__, new_new_n39398__, new_new_n39399__,
    new_new_n39400__, new_new_n39401__, new_new_n39402__, new_new_n39403__,
    new_new_n39404__, new_new_n39405__, new_new_n39406__, new_new_n39407__,
    new_new_n39408__, new_new_n39409__, new_new_n39410__, new_new_n39411__,
    new_new_n39412__, new_new_n39413__, new_new_n39414__, new_new_n39415__,
    new_new_n39416__, new_new_n39417__, new_new_n39418__, new_new_n39419__,
    new_new_n39420__, new_new_n39421__, new_new_n39422__, new_new_n39423__,
    new_new_n39424__, new_new_n39425__, new_new_n39426__, new_new_n39427__,
    new_new_n39428__, new_new_n39429__, new_new_n39430__, new_new_n39431__,
    new_new_n39432__, new_new_n39433__, new_new_n39434__, new_new_n39435__,
    new_new_n39436__, new_new_n39437__, new_new_n39438__, new_new_n39439__,
    new_new_n39440__, new_new_n39441__, new_new_n39442__, new_new_n39443__,
    new_new_n39444__, new_new_n39445__, new_new_n39446__, new_new_n39447__,
    new_new_n39448__, new_new_n39449__, new_new_n39450__, new_new_n39451__,
    new_new_n39452__, new_new_n39453__, new_new_n39454__, new_new_n39455__,
    new_new_n39456__, new_new_n39457__, new_new_n39458__, new_new_n39459__,
    new_new_n39460__, new_new_n39461__, new_new_n39462__, new_new_n39463__,
    new_new_n39464__, new_new_n39465__, new_new_n39466__, new_new_n39467__,
    new_new_n39468__, new_new_n39469__, new_new_n39470__, new_new_n39471__,
    new_new_n39472__, new_new_n39473__, new_new_n39474__, new_new_n39475__,
    new_new_n39476__, new_new_n39477__, new_new_n39478__, new_new_n39479__,
    new_new_n39480__, new_new_n39481__, new_new_n39482__, new_new_n39483__,
    new_new_n39484__, new_new_n39485__, new_new_n39486__, new_new_n39487__,
    new_new_n39488__, new_new_n39489__, new_new_n39490__, new_new_n39491__,
    new_new_n39492__, new_new_n39493__, new_new_n39494__, new_new_n39495__,
    new_new_n39496__, new_new_n39497__, new_new_n39498__, new_new_n39499__,
    new_new_n39500__, new_new_n39501__, new_new_n39502__, new_new_n39503__,
    new_new_n39504__, new_new_n39505__, new_new_n39506__, new_new_n39507__,
    new_new_n39508__, new_new_n39509__, new_new_n39510__, new_new_n39511__,
    new_new_n39512__, new_new_n39513__, new_new_n39514__, new_new_n39515__,
    new_new_n39516__, new_new_n39517__, new_new_n39518__, new_new_n39519__,
    new_new_n39520__, new_new_n39521__, new_new_n39522__, new_new_n39523__,
    new_new_n39524__, new_new_n39525__, new_new_n39526__, new_new_n39527__,
    new_new_n39528__, new_new_n39529__, new_new_n39530__, new_new_n39531__,
    new_new_n39532__, new_new_n39533__, new_new_n39534__, new_new_n39535__,
    new_new_n39536__, new_new_n39537__, new_new_n39538__, new_new_n39539__,
    new_new_n39540__, new_new_n39541__, new_new_n39542__, new_new_n39543__,
    new_new_n39544__, new_new_n39545__, new_new_n39546__, new_new_n39547__,
    new_new_n39548__, new_new_n39549__, new_new_n39550__, new_new_n39551__,
    new_new_n39552__, new_new_n39553__, new_new_n39554__, new_new_n39555__,
    new_new_n39556__, new_new_n39557__, new_new_n39558__, new_new_n39559__,
    new_new_n39560__, new_new_n39561__, new_new_n39562__, new_new_n39563__,
    new_new_n39564__, new_new_n39565__, new_new_n39566__, new_new_n39567__,
    new_new_n39568__, new_new_n39569__, new_new_n39570__, new_new_n39571__,
    new_new_n39572__, new_new_n39573__, new_new_n39574__, new_new_n39575__,
    new_new_n39576__, new_new_n39577__, new_new_n39578__, new_new_n39579__,
    new_new_n39580__, new_new_n39581__, new_new_n39582__, new_new_n39583__,
    new_new_n39584__, new_new_n39585__, new_new_n39586__, new_new_n39587__,
    new_new_n39588__, new_new_n39589__, new_new_n39590__, new_new_n39591__,
    new_new_n39592__, new_new_n39593__, new_new_n39594__, new_new_n39595__,
    new_new_n39596__, new_new_n39597__, new_new_n39598__, new_new_n39599__,
    new_new_n39600__, new_new_n39601__, new_new_n39602__, new_new_n39603__,
    new_new_n39604__, new_new_n39605__, new_new_n39606__, new_new_n39607__,
    new_new_n39608__, new_new_n39609__, new_new_n39610__, new_new_n39611__,
    new_new_n39612__, new_new_n39613__, new_new_n39614__, new_new_n39615__,
    new_new_n39616__, new_new_n39617__, new_new_n39618__, new_new_n39619__,
    new_new_n39620__, new_new_n39621__, new_new_n39622__, new_new_n39623__,
    new_new_n39624__, new_new_n39625__, new_new_n39626__, new_new_n39627__,
    new_new_n39628__, new_new_n39629__, new_new_n39630__, new_new_n39632__,
    new_new_n39633__, new_new_n39634__, new_new_n39635__, new_new_n39636__,
    new_new_n39637__, new_new_n39638__, new_new_n39639__, new_new_n39640__,
    new_new_n39641__, new_new_n39642__, new_new_n39643__, new_new_n39644__,
    new_new_n39645__, new_new_n39646__, new_new_n39647__, new_new_n39648__,
    new_new_n39649__, new_new_n39650__, new_new_n39651__, new_new_n39652__,
    new_new_n39653__, new_new_n39654__, new_new_n39655__, new_new_n39656__,
    new_new_n39657__, new_new_n39659__, new_new_n39660__, new_new_n39661__,
    new_new_n39662__, new_new_n39663__, new_new_n39664__, new_new_n39665__,
    new_new_n39666__, new_new_n39667__, new_new_n39668__, new_new_n39669__,
    new_new_n39670__, new_new_n39671__, new_new_n39672__, new_new_n39673__,
    new_new_n39674__, new_new_n39675__, new_new_n39676__, new_new_n39677__,
    new_new_n39678__, new_new_n39679__, new_new_n39680__, new_new_n39681__,
    new_new_n39682__, new_new_n39683__, new_new_n39685__, new_new_n39686__,
    new_new_n39687__, new_new_n39688__, new_new_n39689__, new_new_n39690__,
    new_new_n39691__, new_new_n39692__, new_new_n39693__, new_new_n39694__,
    new_new_n39695__, new_new_n39696__, new_new_n39697__, new_new_n39698__,
    new_new_n39699__, new_new_n39700__, new_new_n39701__, new_new_n39702__,
    new_new_n39703__, new_new_n39704__, new_new_n39705__, new_new_n39706__,
    new_new_n39707__, new_new_n39708__, new_new_n39709__, new_new_n39711__,
    new_new_n39712__, new_new_n39713__, new_new_n39714__, new_new_n39715__,
    new_new_n39716__, new_new_n39717__, new_new_n39718__, new_new_n39719__,
    new_new_n39720__, new_new_n39721__, new_new_n39722__, new_new_n39723__,
    new_new_n39724__, new_new_n39725__, new_new_n39726__, new_new_n39727__,
    new_new_n39728__, new_new_n39729__, new_new_n39730__, new_new_n39731__,
    new_new_n39732__, new_new_n39733__, new_new_n39734__, new_new_n39736__,
    new_new_n39737__, new_new_n39738__, new_new_n39739__, new_new_n39740__,
    new_new_n39741__, new_new_n39742__, new_new_n39743__, new_new_n39744__,
    new_new_n39745__, new_new_n39746__, new_new_n39747__, new_new_n39748__,
    new_new_n39749__, new_new_n39750__, new_new_n39751__, new_new_n39752__,
    new_new_n39753__, new_new_n39754__, new_new_n39755__, new_new_n39756__,
    new_new_n39757__, new_new_n39758__, new_new_n39759__, new_new_n39760__,
    new_new_n39761__, new_new_n39762__, new_new_n39764__, new_new_n39765__,
    new_new_n39766__, new_new_n39767__, new_new_n39768__, new_new_n39769__,
    new_new_n39770__, new_new_n39771__, new_new_n39772__, new_new_n39773__,
    new_new_n39774__, new_new_n39775__, new_new_n39776__, new_new_n39777__,
    new_new_n39778__, new_new_n39779__, new_new_n39780__, new_new_n39781__,
    new_new_n39782__, new_new_n39783__, new_new_n39784__, new_new_n39785__,
    new_new_n39786__, new_new_n39787__, new_new_n39788__, new_new_n39789__,
    new_new_n39790__, new_new_n39791__, new_new_n39793__, new_new_n39794__,
    new_new_n39795__, new_new_n39796__, new_new_n39797__, new_new_n39798__,
    new_new_n39799__, new_new_n39800__, new_new_n39801__, new_new_n39802__,
    new_new_n39803__, new_new_n39804__, new_new_n39805__, new_new_n39806__,
    new_new_n39807__, new_new_n39808__, new_new_n39809__, new_new_n39810__,
    new_new_n39811__, new_new_n39812__, new_new_n39813__, new_new_n39814__,
    new_new_n39815__, new_new_n39816__, new_new_n39817__, new_new_n39818__,
    new_new_n39819__, new_new_n39820__, new_new_n39822__, new_new_n39823__,
    new_new_n39824__, new_new_n39825__, new_new_n39826__, new_new_n39827__,
    new_new_n39828__, new_new_n39829__, new_new_n39830__, new_new_n39831__,
    new_new_n39832__, new_new_n39833__, new_new_n39834__, new_new_n39835__,
    new_new_n39836__, new_new_n39837__, new_new_n39838__, new_new_n39839__,
    new_new_n39840__, new_new_n39841__, new_new_n39842__, new_new_n39843__,
    new_new_n39844__, new_new_n39845__, new_new_n39846__, new_new_n39848__,
    new_new_n39849__, new_new_n39850__, new_new_n39851__, new_new_n39852__,
    new_new_n39853__, new_new_n39854__, new_new_n39855__, new_new_n39856__,
    new_new_n39857__, new_new_n39858__, new_new_n39859__, new_new_n39860__,
    new_new_n39861__, new_new_n39862__, new_new_n39863__, new_new_n39864__,
    new_new_n39865__, new_new_n39866__, new_new_n39867__, new_new_n39868__,
    new_new_n39869__, new_new_n39870__, new_new_n39871__, new_new_n39872__,
    new_new_n39873__, new_new_n39874__, new_new_n39876__, new_new_n39877__,
    new_new_n39878__, new_new_n39879__, new_new_n39880__, new_new_n39881__,
    new_new_n39882__, new_new_n39883__, new_new_n39884__, new_new_n39885__,
    new_new_n39886__, new_new_n39887__, new_new_n39888__, new_new_n39889__,
    new_new_n39890__, new_new_n39891__, new_new_n39892__, new_new_n39893__,
    new_new_n39894__, new_new_n39895__, new_new_n39896__, new_new_n39897__,
    new_new_n39898__, new_new_n39899__, new_new_n39900__, new_new_n39901__,
    new_new_n39902__, new_new_n39903__, new_new_n39905__, new_new_n39906__,
    new_new_n39907__, new_new_n39908__, new_new_n39909__, new_new_n39910__,
    new_new_n39911__, new_new_n39912__, new_new_n39913__, new_new_n39914__,
    new_new_n39915__, new_new_n39916__, new_new_n39917__, new_new_n39918__,
    new_new_n39919__, new_new_n39920__, new_new_n39921__, new_new_n39922__,
    new_new_n39923__, new_new_n39924__, new_new_n39925__, new_new_n39926__,
    new_new_n39927__, new_new_n39928__, new_new_n39929__, new_new_n39930__,
    new_new_n39931__, new_new_n39932__, new_new_n39934__, new_new_n39935__,
    new_new_n39936__, new_new_n39937__, new_new_n39938__, new_new_n39939__,
    new_new_n39940__, new_new_n39941__, new_new_n39942__, new_new_n39943__,
    new_new_n39944__, new_new_n39945__, new_new_n39946__, new_new_n39947__,
    new_new_n39948__, new_new_n39949__, new_new_n39950__, new_new_n39951__,
    new_new_n39952__, new_new_n39953__, new_new_n39954__, new_new_n39955__,
    new_new_n39956__, new_new_n39957__, new_new_n39958__, new_new_n39959__,
    new_new_n39960__, new_new_n39961__, new_new_n39963__, new_new_n39964__,
    new_new_n39965__, new_new_n39966__, new_new_n39967__, new_new_n39968__,
    new_new_n39969__, new_new_n39970__, new_new_n39971__, new_new_n39972__,
    new_new_n39973__, new_new_n39974__, new_new_n39975__, new_new_n39976__,
    new_new_n39977__, new_new_n39978__, new_new_n39979__, new_new_n39980__,
    new_new_n39981__, new_new_n39982__, new_new_n39983__, new_new_n39984__,
    new_new_n39985__, new_new_n39986__, new_new_n39987__, new_new_n39988__,
    new_new_n39989__, new_new_n39990__, new_new_n39992__, new_new_n39993__,
    new_new_n39994__, new_new_n39995__, new_new_n39996__, new_new_n39997__,
    new_new_n39998__, new_new_n39999__, new_new_n40000__, new_new_n40001__,
    new_new_n40002__, new_new_n40003__, new_new_n40004__, new_new_n40005__,
    new_new_n40006__, new_new_n40007__, new_new_n40008__, new_new_n40009__,
    new_new_n40010__, new_new_n40011__, new_new_n40012__, new_new_n40013__,
    new_new_n40014__, new_new_n40015__, new_new_n40016__, new_new_n40017__,
    new_new_n40018__, new_new_n40019__, new_new_n40021__, new_new_n40022__,
    new_new_n40023__, new_new_n40024__, new_new_n40025__, new_new_n40026__,
    new_new_n40027__, new_new_n40028__, new_new_n40029__, new_new_n40030__,
    new_new_n40031__, new_new_n40032__, new_new_n40033__, new_new_n40034__,
    new_new_n40035__, new_new_n40036__, new_new_n40037__, new_new_n40038__,
    new_new_n40039__, new_new_n40040__, new_new_n40041__, new_new_n40042__,
    new_new_n40043__, new_new_n40044__, new_new_n40045__, new_new_n40046__,
    new_new_n40047__, new_new_n40048__, new_new_n40050__, new_new_n40051__,
    new_new_n40052__, new_new_n40053__, new_new_n40054__, new_new_n40055__,
    new_new_n40056__, new_new_n40057__, new_new_n40058__, new_new_n40059__,
    new_new_n40060__, new_new_n40061__, new_new_n40062__, new_new_n40063__,
    new_new_n40064__, new_new_n40065__, new_new_n40066__, new_new_n40067__,
    new_new_n40068__, new_new_n40069__, new_new_n40070__, new_new_n40071__,
    new_new_n40072__, new_new_n40073__, new_new_n40074__, new_new_n40076__,
    new_new_n40077__, new_new_n40078__, new_new_n40079__, new_new_n40080__,
    new_new_n40081__, new_new_n40082__, new_new_n40083__, new_new_n40084__,
    new_new_n40085__, new_new_n40086__, new_new_n40087__, new_new_n40088__,
    new_new_n40089__, new_new_n40090__, new_new_n40091__, new_new_n40092__,
    new_new_n40093__, new_new_n40094__, new_new_n40095__, new_new_n40096__,
    new_new_n40097__, new_new_n40098__, new_new_n40099__, new_new_n40100__,
    new_new_n40101__, new_new_n40102__, new_new_n40103__, new_new_n40104__,
    new_new_n40105__, new_new_n40106__, new_new_n40108__, new_new_n40109__,
    new_new_n40110__, new_new_n40111__, new_new_n40112__, new_new_n40113__,
    new_new_n40114__, new_new_n40115__, new_new_n40116__, new_new_n40117__,
    new_new_n40118__, new_new_n40119__, new_new_n40120__, new_new_n40121__,
    new_new_n40122__, new_new_n40123__, new_new_n40124__, new_new_n40125__,
    new_new_n40126__, new_new_n40127__, new_new_n40128__, new_new_n40129__,
    new_new_n40130__, new_new_n40131__, new_new_n40132__, new_new_n40133__,
    new_new_n40134__, new_new_n40135__, new_new_n40136__, new_new_n40137__,
    new_new_n40138__, new_new_n40139__, new_new_n40140__, new_new_n40141__,
    new_new_n40143__, new_new_n40144__, new_new_n40145__, new_new_n40146__,
    new_new_n40147__, new_new_n40148__, new_new_n40149__, new_new_n40150__,
    new_new_n40151__, new_new_n40152__, new_new_n40153__, new_new_n40154__,
    new_new_n40155__, new_new_n40156__, new_new_n40157__, new_new_n40158__,
    new_new_n40159__, new_new_n40160__, new_new_n40161__, new_new_n40162__,
    new_new_n40163__, new_new_n40164__, new_new_n40165__, new_new_n40166__,
    new_new_n40167__, new_new_n40168__, new_new_n40169__, new_new_n40170__,
    new_new_n40171__, new_new_n40172__, new_new_n40173__, new_new_n40174__,
    new_new_n40175__, new_new_n40176__, new_new_n40178__, new_new_n40179__,
    new_new_n40180__, new_new_n40181__, new_new_n40182__, new_new_n40183__,
    new_new_n40184__, new_new_n40185__, new_new_n40186__, new_new_n40187__,
    new_new_n40188__, new_new_n40189__, new_new_n40190__, new_new_n40191__,
    new_new_n40192__, new_new_n40193__, new_new_n40194__, new_new_n40195__,
    new_new_n40196__, new_new_n40197__, new_new_n40198__, new_new_n40199__,
    new_new_n40200__, new_new_n40201__, new_new_n40202__, new_new_n40203__,
    new_new_n40204__, new_new_n40205__, new_new_n40206__, new_new_n40207__,
    new_new_n40208__, new_new_n40209__, new_new_n40210__, new_new_n40211__,
    new_new_n40213__, new_new_n40214__, new_new_n40215__, new_new_n40216__,
    new_new_n40217__, new_new_n40218__, new_new_n40219__, new_new_n40220__,
    new_new_n40221__, new_new_n40222__, new_new_n40223__, new_new_n40224__,
    new_new_n40225__, new_new_n40226__, new_new_n40227__, new_new_n40228__,
    new_new_n40229__, new_new_n40230__, new_new_n40231__, new_new_n40232__,
    new_new_n40233__, new_new_n40234__, new_new_n40235__, new_new_n40236__,
    new_new_n40237__, new_new_n40238__, new_new_n40239__, new_new_n40240__,
    new_new_n40241__, new_new_n40242__, new_new_n40243__, new_new_n40244__,
    new_new_n40245__, new_new_n40246__, new_new_n40247__, new_new_n40248__,
    new_new_n40250__, new_new_n40251__, new_new_n40252__, new_new_n40253__,
    new_new_n40254__, new_new_n40255__, new_new_n40256__, new_new_n40257__,
    new_new_n40258__, new_new_n40259__, new_new_n40260__, new_new_n40261__,
    new_new_n40262__, new_new_n40263__, new_new_n40264__, new_new_n40265__,
    new_new_n40266__, new_new_n40267__, new_new_n40268__, new_new_n40269__,
    new_new_n40270__, new_new_n40271__, new_new_n40272__, new_new_n40273__,
    new_new_n40274__, new_new_n40275__, new_new_n40276__, new_new_n40277__,
    new_new_n40278__, new_new_n40279__, new_new_n40280__, new_new_n40281__,
    new_new_n40282__, new_new_n40283__, new_new_n40284__, new_new_n40285__,
    new_new_n40286__, new_new_n40288__, new_new_n40289__, new_new_n40290__,
    new_new_n40291__, new_new_n40292__, new_new_n40293__, new_new_n40294__,
    new_new_n40295__, new_new_n40296__, new_new_n40297__, new_new_n40298__,
    new_new_n40299__, new_new_n40300__, new_new_n40301__, new_new_n40302__,
    new_new_n40303__, new_new_n40304__, new_new_n40305__, new_new_n40306__,
    new_new_n40307__, new_new_n40308__, new_new_n40309__, new_new_n40310__,
    new_new_n40311__, new_new_n40312__, new_new_n40313__, new_new_n40314__,
    new_new_n40315__, new_new_n40316__, new_new_n40317__, new_new_n40318__,
    new_new_n40319__, new_new_n40320__, new_new_n40321__, new_new_n40322__,
    new_new_n40323__, new_new_n40324__, new_new_n40326__, new_new_n40327__,
    new_new_n40328__, new_new_n40329__, new_new_n40330__, new_new_n40331__,
    new_new_n40332__, new_new_n40333__, new_new_n40334__, new_new_n40335__,
    new_new_n40336__, new_new_n40337__, new_new_n40338__, new_new_n40339__,
    new_new_n40340__, new_new_n40341__, new_new_n40342__, new_new_n40343__,
    new_new_n40344__, new_new_n40345__, new_new_n40346__, new_new_n40347__,
    new_new_n40348__, new_new_n40349__, new_new_n40350__, new_new_n40351__,
    new_new_n40352__, new_new_n40353__, new_new_n40354__, new_new_n40355__,
    new_new_n40356__, new_new_n40357__, new_new_n40358__, new_new_n40359__,
    new_new_n40360__, new_new_n40362__, new_new_n40363__, new_new_n40364__,
    new_new_n40365__, new_new_n40366__, new_new_n40367__, new_new_n40368__,
    new_new_n40369__, new_new_n40370__, new_new_n40371__, new_new_n40372__,
    new_new_n40373__, new_new_n40374__, new_new_n40375__, new_new_n40376__,
    new_new_n40377__, new_new_n40378__, new_new_n40379__, new_new_n40380__,
    new_new_n40381__, new_new_n40382__, new_new_n40383__, new_new_n40384__,
    new_new_n40385__, new_new_n40386__, new_new_n40387__, new_new_n40388__,
    new_new_n40389__, new_new_n40390__, new_new_n40391__, new_new_n40392__,
    new_new_n40393__, new_new_n40394__, new_new_n40395__, new_new_n40396__,
    new_new_n40397__, new_new_n40399__, new_new_n40400__, new_new_n40401__,
    new_new_n40402__, new_new_n40403__, new_new_n40404__, new_new_n40405__,
    new_new_n40406__, new_new_n40407__, new_new_n40408__, new_new_n40409__,
    new_new_n40410__, new_new_n40411__, new_new_n40412__, new_new_n40413__,
    new_new_n40414__, new_new_n40415__, new_new_n40416__, new_new_n40417__,
    new_new_n40418__, new_new_n40419__, new_new_n40420__, new_new_n40421__,
    new_new_n40422__, new_new_n40423__, new_new_n40424__, new_new_n40425__,
    new_new_n40426__, new_new_n40427__, new_new_n40428__, new_new_n40429__,
    new_new_n40430__, new_new_n40431__, new_new_n40432__, new_new_n40433__,
    new_new_n40434__, new_new_n40435__, new_new_n40437__, new_new_n40438__,
    new_new_n40439__, new_new_n40440__, new_new_n40441__, new_new_n40442__,
    new_new_n40443__, new_new_n40444__, new_new_n40445__, new_new_n40446__,
    new_new_n40447__, new_new_n40448__, new_new_n40449__, new_new_n40450__,
    new_new_n40451__, new_new_n40452__, new_new_n40453__, new_new_n40454__,
    new_new_n40455__, new_new_n40456__, new_new_n40457__, new_new_n40458__,
    new_new_n40459__, new_new_n40460__, new_new_n40461__, new_new_n40462__,
    new_new_n40463__, new_new_n40464__, new_new_n40465__, new_new_n40466__,
    new_new_n40467__, new_new_n40468__, new_new_n40469__, new_new_n40470__,
    new_new_n40471__, new_new_n40472__, new_new_n40473__, new_new_n40475__,
    new_new_n40476__, new_new_n40477__, new_new_n40478__, new_new_n40479__,
    new_new_n40480__, new_new_n40481__, new_new_n40482__, new_new_n40483__,
    new_new_n40484__, new_new_n40485__, new_new_n40486__, new_new_n40487__,
    new_new_n40488__, new_new_n40489__, new_new_n40490__, new_new_n40491__,
    new_new_n40492__, new_new_n40493__, new_new_n40494__, new_new_n40495__,
    new_new_n40496__, new_new_n40497__, new_new_n40498__, new_new_n40499__,
    new_new_n40500__, new_new_n40501__, new_new_n40502__, new_new_n40503__,
    new_new_n40504__, new_new_n40505__, new_new_n40506__, new_new_n40507__,
    new_new_n40508__, new_new_n40509__, new_new_n40510__, new_new_n40511__,
    new_new_n40513__, new_new_n40514__, new_new_n40515__, new_new_n40516__,
    new_new_n40517__, new_new_n40518__, new_new_n40519__, new_new_n40520__,
    new_new_n40521__, new_new_n40522__, new_new_n40523__, new_new_n40524__,
    new_new_n40525__, new_new_n40526__, new_new_n40527__, new_new_n40528__,
    new_new_n40529__, new_new_n40530__, new_new_n40531__, new_new_n40532__,
    new_new_n40533__, new_new_n40534__, new_new_n40535__, new_new_n40536__,
    new_new_n40537__, new_new_n40538__, new_new_n40539__, new_new_n40540__,
    new_new_n40541__, new_new_n40542__, new_new_n40543__, new_new_n40544__,
    new_new_n40545__, new_new_n40546__, new_new_n40547__, new_new_n40548__,
    new_new_n40550__, new_new_n40551__, new_new_n40552__, new_new_n40553__,
    new_new_n40554__, new_new_n40555__, new_new_n40556__, new_new_n40557__,
    new_new_n40558__, new_new_n40559__, new_new_n40560__, new_new_n40561__,
    new_new_n40562__, new_new_n40563__, new_new_n40564__, new_new_n40565__,
    new_new_n40566__, new_new_n40567__, new_new_n40568__, new_new_n40569__,
    new_new_n40570__, new_new_n40571__, new_new_n40572__, new_new_n40573__,
    new_new_n40574__, new_new_n40575__, new_new_n40576__, new_new_n40577__,
    new_new_n40578__, new_new_n40579__, new_new_n40580__, new_new_n40581__,
    new_new_n40582__, new_new_n40583__, new_new_n40584__, new_new_n40585__,
    new_new_n40586__, new_new_n40588__, new_new_n40589__, new_new_n40590__,
    new_new_n40591__, new_new_n40592__, new_new_n40593__, new_new_n40594__,
    new_new_n40595__, new_new_n40596__, new_new_n40597__, new_new_n40598__,
    new_new_n40599__, new_new_n40600__, new_new_n40601__, new_new_n40602__,
    new_new_n40603__, new_new_n40604__, new_new_n40605__, new_new_n40606__,
    new_new_n40607__, new_new_n40608__, new_new_n40609__, new_new_n40610__,
    new_new_n40611__, new_new_n40612__, new_new_n40613__, new_new_n40614__,
    new_new_n40615__, new_new_n40616__, new_new_n40617__, new_new_n40618__,
    new_new_n40619__, new_new_n40620__, new_new_n40621__, new_new_n40622__,
    new_new_n40623__, new_new_n40626__, new_new_n40627__, new_new_n40628__,
    new_new_n40629__, new_new_n40630__, new_new_n40631__, new_new_n40632__,
    new_new_n40633__, new_new_n40634__, new_new_n40635__, new_new_n40636__,
    new_new_n40637__, new_new_n40638__, new_new_n40639__, new_new_n40640__,
    new_new_n40641__, new_new_n40642__, new_new_n40643__, new_new_n40644__,
    new_new_n40646__, new_new_n40647__, new_new_n40648__, new_new_n40649__,
    new_new_n40650__, new_new_n40651__, new_new_n40652__, new_new_n40653__,
    new_new_n40654__, new_new_n40656__, new_new_n40657__, new_new_n40658__,
    new_new_n40659__, new_new_n40660__, new_new_n40661__, new_new_n40662__,
    new_new_n40663__, new_new_n40665__, new_new_n40666__, new_new_n40667__,
    new_new_n40668__, new_new_n40669__, new_new_n40671__, new_new_n40672__,
    new_new_n40673__, new_new_n40674__, new_new_n40675__, new_new_n40676__,
    new_new_n40677__, new_new_n40678__, new_new_n40680__, new_new_n40681__,
    new_new_n40682__, new_new_n40683__, new_new_n40684__, new_new_n40685__,
    new_new_n40686__, new_new_n40687__, new_new_n40689__, new_new_n40690__,
    new_new_n40691__, new_new_n40692__, new_new_n40693__, new_new_n40694__,
    new_new_n40695__, new_new_n40696__, new_new_n40697__, new_new_n40698__,
    new_new_n40699__, new_new_n40700__, new_new_n40701__, new_new_n40703__,
    new_new_n40704__, new_new_n40705__, new_new_n40706__, new_new_n40707__,
    new_new_n40709__, new_new_n40710__, new_new_n40711__, new_new_n40712__,
    new_new_n40713__, new_new_n40714__, new_new_n40715__, new_new_n40716__,
    new_new_n40718__, new_new_n40719__, new_new_n40720__, new_new_n40721__,
    new_new_n40722__, new_new_n40723__, new_new_n40724__, new_new_n40725__,
    new_new_n40726__, new_new_n40728__, new_new_n40729__, new_new_n40730__,
    new_new_n40731__, new_new_n40732__, new_new_n40733__, new_new_n40734__,
    new_new_n40735__, new_new_n40736__, new_new_n40737__, new_new_n40738__,
    new_new_n40739__, new_new_n40740__, new_new_n40741__, new_new_n40742__,
    new_new_n40743__, new_new_n40744__, new_new_n40745__, new_new_n40746__,
    new_new_n40747__, new_new_n40748__, new_new_n40749__, new_new_n40750__,
    new_new_n40751__, new_new_n40752__, new_new_n40754__, new_new_n40755__,
    new_new_n40756__, new_new_n40757__, new_new_n40758__, new_new_n40759__,
    new_new_n40760__, new_new_n40761__, new_new_n40763__, new_new_n40764__,
    new_new_n40765__, new_new_n40766__, new_new_n40767__, new_new_n40768__,
    new_new_n40769__, new_new_n40770__, new_new_n40771__, new_new_n40773__,
    new_new_n40774__, new_new_n40775__, new_new_n40776__, new_new_n40777__,
    new_new_n40778__, new_new_n40779__, new_new_n40780__, new_new_n40782__,
    new_new_n40783__, new_new_n40784__, new_new_n40785__, new_new_n40786__,
    new_new_n40787__, new_new_n40788__, new_new_n40789__, new_new_n40790__,
    new_new_n40791__, new_new_n40793__, new_new_n40794__, new_new_n40795__,
    new_new_n40796__, new_new_n40797__, new_new_n40798__, new_new_n40799__,
    new_new_n40800__, new_new_n40802__, new_new_n40803__, new_new_n40804__,
    new_new_n40805__, new_new_n40806__, new_new_n40807__, new_new_n40808__,
    new_new_n40809__, new_new_n40810__, new_new_n40812__, new_new_n40813__,
    new_new_n40814__, new_new_n40815__, new_new_n40816__, new_new_n40817__,
    new_new_n40818__, new_new_n40819__, new_new_n40820__, new_new_n40821__,
    new_new_n40822__, new_new_n40823__, new_new_n40824__, new_new_n40825__,
    new_new_n40826__, new_new_n40827__, new_new_n40828__, new_new_n40829__,
    new_new_n40830__, new_new_n40831__, new_new_n40832__, new_new_n40833__,
    new_new_n40834__, new_new_n40835__, new_new_n40836__, new_new_n40837__,
    new_new_n40838__, new_new_n40839__, new_new_n40840__, new_new_n40841__,
    new_new_n40842__, new_new_n40843__, new_new_n40844__, new_new_n40845__,
    new_new_n40846__, new_new_n40848__, new_new_n40849__, new_new_n40850__,
    new_new_n40851__, new_new_n40852__, new_new_n40853__, new_new_n40854__,
    new_new_n40855__, new_new_n40856__, new_new_n40858__, new_new_n40859__,
    new_new_n40860__, new_new_n40861__, new_new_n40862__, new_new_n40863__,
    new_new_n40864__, new_new_n40865__, new_new_n40866__, new_new_n40867__,
    new_new_n40868__, new_new_n40869__, new_new_n40871__, new_new_n40872__,
    new_new_n40873__, new_new_n40874__, new_new_n40875__, new_new_n40876__,
    new_new_n40877__, new_new_n40878__, new_new_n40879__, new_new_n40881__,
    new_new_n40882__, new_new_n40883__, new_new_n40884__, new_new_n40885__,
    new_new_n40886__, new_new_n40887__, new_new_n40888__, new_new_n40889__,
    new_new_n40890__, new_new_n40891__, new_new_n40892__, new_new_n40893__,
    new_new_n40894__, new_new_n40895__, new_new_n40897__, new_new_n40898__,
    new_new_n40899__, new_new_n40900__, new_new_n40901__, new_new_n40902__,
    new_new_n40903__, new_new_n40904__, new_new_n40905__, new_new_n40907__,
    new_new_n40908__, new_new_n40909__, new_new_n40910__, new_new_n40911__,
    new_new_n40912__, new_new_n40913__, new_new_n40914__, new_new_n40915__,
    new_new_n40916__, new_new_n40917__, new_new_n40918__, new_new_n40919__,
    new_new_n40920__, new_new_n40921__, new_new_n40923__, new_new_n40924__,
    new_new_n40925__, new_new_n40926__, new_new_n40927__, new_new_n40928__,
    new_new_n40929__, new_new_n40930__, new_new_n40931__, new_new_n40933__,
    new_new_n40934__, new_new_n40935__, new_new_n40936__, new_new_n40937__,
    new_new_n40938__, new_new_n40939__, new_new_n40940__, new_new_n40941__,
    new_new_n40942__, new_new_n40943__, new_new_n40944__, new_new_n40945__,
    new_new_n40946__, new_new_n40947__, new_new_n40948__, new_new_n40949__,
    new_new_n40950__, new_new_n40952__, new_new_n40953__, new_new_n40954__,
    new_new_n40955__, new_new_n40956__, new_new_n40957__, new_new_n40958__,
    new_new_n40959__, new_new_n40960__, new_new_n40962__, new_new_n40963__,
    new_new_n40964__, new_new_n40965__, new_new_n40966__, new_new_n40967__,
    new_new_n40968__, new_new_n40969__, new_new_n40970__, new_new_n40971__,
    new_new_n40972__, new_new_n40973__, new_new_n40974__, new_new_n40975__,
    new_new_n40976__, new_new_n40978__, new_new_n40979__, new_new_n40980__,
    new_new_n40981__, new_new_n40982__, new_new_n40983__, new_new_n40984__,
    new_new_n40985__, new_new_n40986__, new_new_n40988__, new_new_n40989__,
    new_new_n40990__, new_new_n40991__, new_new_n40992__, new_new_n40993__,
    new_new_n40994__, new_new_n40995__, new_new_n40996__, new_new_n40997__,
    new_new_n40998__, new_new_n40999__, new_new_n41000__, new_new_n41001__,
    new_new_n41002__, new_new_n41003__, new_new_n41004__, new_new_n41005__,
    new_new_n41006__, new_new_n41008__, new_new_n41009__, new_new_n41010__,
    new_new_n41011__, new_new_n41012__, new_new_n41013__, new_new_n41014__,
    new_new_n41015__, new_new_n41016__, new_new_n41018__, new_new_n41019__,
    new_new_n41020__, new_new_n41021__, new_new_n41022__, new_new_n41023__,
    new_new_n41024__, new_new_n41025__, new_new_n41026__, new_new_n41027__,
    new_new_n41028__, new_new_n41029__, new_new_n41030__, new_new_n41031__,
    new_new_n41032__, new_new_n41034__, new_new_n41035__, new_new_n41036__,
    new_new_n41037__, new_new_n41038__, new_new_n41039__, new_new_n41040__,
    new_new_n41041__, new_new_n41042__, new_new_n41044__, new_new_n41045__,
    new_new_n41046__, new_new_n41047__, new_new_n41048__, new_new_n41049__,
    new_new_n41050__, new_new_n41051__, new_new_n41052__, new_new_n41053__,
    new_new_n41054__, new_new_n41055__, new_new_n41056__, new_new_n41057__,
    new_new_n41058__, new_new_n41059__, new_new_n41060__, new_new_n41061__,
    new_new_n41062__, new_new_n41063__, new_new_n41064__, new_new_n41065__,
    new_new_n41066__, new_new_n41068__, new_new_n41069__, new_new_n41070__,
    new_new_n41071__, new_new_n41072__, new_new_n41073__, new_new_n41074__,
    new_new_n41075__, new_new_n41076__, new_new_n41078__, new_new_n41079__,
    new_new_n41080__, new_new_n41081__, new_new_n41082__, new_new_n41083__,
    new_new_n41084__, new_new_n41085__, new_new_n41086__, new_new_n41087__,
    new_new_n41088__, new_new_n41089__, new_new_n41090__, new_new_n41091__,
    new_new_n41092__, new_new_n41094__, new_new_n41095__, new_new_n41096__,
    new_new_n41097__, new_new_n41098__, new_new_n41099__, new_new_n41100__,
    new_new_n41101__, new_new_n41102__, new_new_n41104__, new_new_n41105__,
    new_new_n41106__, new_new_n41107__, new_new_n41108__, new_new_n41109__,
    new_new_n41110__, new_new_n41111__, new_new_n41112__, new_new_n41113__,
    new_new_n41114__, new_new_n41115__, new_new_n41116__, new_new_n41117__,
    new_new_n41118__, new_new_n41119__, new_new_n41120__, new_new_n41121__,
    new_new_n41122__, new_new_n41124__, new_new_n41125__, new_new_n41126__,
    new_new_n41127__, new_new_n41128__, new_new_n41129__, new_new_n41130__,
    new_new_n41131__, new_new_n41132__, new_new_n41134__, new_new_n41135__,
    new_new_n41136__, new_new_n41137__, new_new_n41138__, new_new_n41139__,
    new_new_n41140__, new_new_n41141__, new_new_n41142__, new_new_n41143__,
    new_new_n41144__, new_new_n41145__, new_new_n41146__, new_new_n41147__,
    new_new_n41148__, new_new_n41150__, new_new_n41151__, new_new_n41152__,
    new_new_n41153__, new_new_n41154__, new_new_n41155__, new_new_n41156__,
    new_new_n41157__, new_new_n41158__, new_new_n41160__, new_new_n41161__,
    new_new_n41162__, new_new_n41163__, new_new_n41164__, new_new_n41165__,
    new_new_n41166__, new_new_n41167__, new_new_n41168__, new_new_n41169__,
    new_new_n41170__, new_new_n41171__, new_new_n41172__, new_new_n41173__,
    new_new_n41174__, new_new_n41175__, new_new_n41176__, new_new_n41177__,
    new_new_n41178__, new_new_n41179__, new_new_n41180__, new_new_n41181__,
    new_new_n41182__, new_new_n41184__, new_new_n41185__, new_new_n41186__,
    new_new_n41187__, new_new_n41188__, new_new_n41189__, new_new_n41190__,
    new_new_n41191__, new_new_n41192__, new_new_n41194__, new_new_n41195__,
    new_new_n41196__, new_new_n41197__, new_new_n41198__, new_new_n41199__,
    new_new_n41200__, new_new_n41201__, new_new_n41202__, new_new_n41203__,
    new_new_n41204__, new_new_n41205__, new_new_n41206__, new_new_n41207__,
    new_new_n41208__, new_new_n41210__, new_new_n41211__, new_new_n41212__,
    new_new_n41213__, new_new_n41214__, new_new_n41215__, new_new_n41216__,
    new_new_n41217__, new_new_n41218__, new_new_n41220__, new_new_n41221__,
    new_new_n41222__, new_new_n41223__, new_new_n41224__, new_new_n41225__,
    new_new_n41226__, new_new_n41227__, new_new_n41228__, new_new_n41229__,
    new_new_n41230__, new_new_n41231__, new_new_n41232__, new_new_n41233__,
    new_new_n41234__, new_new_n41235__, new_new_n41236__, new_new_n41237__,
    new_new_n41238__, new_new_n41240__, new_new_n41241__, new_new_n41242__,
    new_new_n41243__, new_new_n41244__, new_new_n41245__, new_new_n41246__,
    new_new_n41247__, new_new_n41248__, new_new_n41250__, new_new_n41251__,
    new_new_n41252__, new_new_n41253__, new_new_n41254__, new_new_n41255__,
    new_new_n41256__, new_new_n41257__, new_new_n41258__, new_new_n41259__,
    new_new_n41260__, new_new_n41261__, new_new_n41262__, new_new_n41263__,
    new_new_n41264__, new_new_n41266__, new_new_n41267__, new_new_n41269__,
    new_new_n41270__, new_new_n41271__, new_new_n41272__, new_new_n41273__,
    new_new_n41274__, new_new_n41275__, new_new_n41276__, new_new_n41277__,
    new_new_n41278__, new_new_n41279__, new_new_n41280__, new_new_n41281__,
    new_new_n41282__, new_new_n41283__, new_new_n41284__, new_new_n41285__,
    new_new_n41286__, new_new_n41287__, new_new_n41288__, new_new_n41289__,
    new_new_n41290__, new_new_n41291__, new_new_n41292__, new_new_n41293__,
    new_new_n41294__, new_new_n41295__, new_new_n41297__, new_new_n41298__,
    new_new_n41299__, new_new_n41300__, new_new_n41301__, new_new_n41302__,
    new_new_n41303__, new_new_n41304__, new_new_n41305__, new_new_n41307__,
    new_new_n41308__, new_new_n41309__, new_new_n41310__, new_new_n41311__,
    new_new_n41312__, new_new_n41313__, new_new_n41315__, new_new_n41316__,
    new_new_n41318__, new_new_n41319__, new_new_n41321__, new_new_n41322__,
    new_new_n41324__, new_new_n41325__, new_new_n41327__, new_new_n41328__,
    new_new_n41330__, new_new_n41331__, new_new_n41333__, new_new_n41334__,
    new_new_n41336__, new_new_n41337__, new_new_n41339__, new_new_n41340__,
    new_new_n41342__, new_new_n41343__, new_new_n41345__, new_new_n41346__,
    new_new_n41348__, new_new_n41349__, new_new_n41351__, new_new_n41352__,
    new_new_n41354__, new_new_n41355__, new_new_n41357__, new_new_n41358__,
    new_new_n41360__, new_new_n41361__, new_new_n41363__, new_new_n41364__,
    new_new_n41366__, new_new_n41367__, new_new_n41368__, new_new_n41369__,
    new_new_n41370__, new_new_n41371__, new_new_n41372__, new_new_n41373__,
    new_new_n41374__, new_new_n41375__, new_new_n41376__, new_new_n41377__,
    new_new_n41378__, new_new_n41379__, new_new_n41380__, new_new_n41381__,
    new_new_n41382__, new_new_n41383__, new_new_n41384__, new_new_n41385__,
    new_new_n41386__, new_new_n41387__, new_new_n41388__, new_new_n41389__,
    new_new_n41390__, new_new_n41391__, new_new_n41392__, new_new_n41393__,
    new_new_n41394__, new_new_n41395__, new_new_n41396__, new_new_n41397__,
    new_new_n41398__, new_new_n41399__, new_new_n41400__, new_new_n41401__,
    new_new_n41402__, new_new_n41403__, new_new_n41404__, new_new_n41405__,
    new_new_n41406__, new_new_n41408__, new_new_n41409__, new_new_n41410__,
    new_new_n41411__, new_new_n41412__, new_new_n41413__, new_new_n41415__,
    new_new_n41416__, new_new_n41418__, new_new_n41419__, new_new_n41420__,
    new_new_n41422__, new_new_n41423__, new_new_n41424__, new_new_n41426__,
    new_new_n41427__, new_new_n41428__, new_new_n41430__, new_new_n41431__,
    new_new_n41432__, new_new_n41437__, new_new_n41443__, new_new_n41445__,
    new_new_n41452__, new_new_n41453__, new_new_n41454__, new_new_n41455__,
    new_new_n41456__, new_new_n41457__, new_new_n41458__, new_new_n41459__,
    new_new_n41460__, new_new_n41461__, new_new_n41462__, new_new_n41463__,
    new_new_n41464__, new_new_n41465__, new_new_n41466__, new_new_n41467__,
    new_new_n41468__, new_new_n41469__, new_new_n41470__, new_new_n41471__,
    new_new_n41472__, new_new_n41473__, new_new_n41474__, new_new_n41475__,
    new_new_n41476__, new_new_n41477__, new_new_n41478__, new_new_n41479__,
    new_new_n41480__, new_new_n41481__, new_new_n41483__, new_new_n41484__,
    new_new_n41485__, new_new_n41486__, new_new_n41487__, new_new_n41489__,
    new_new_n41490__, new_new_n41491__, new_new_n41492__, new_new_n41493__,
    new_new_n41494__, new_new_n41495__, new_new_n41496__, new_new_n41497__,
    new_new_n41498__, new_new_n41499__, new_new_n41500__, new_new_n41501__,
    new_new_n41502__, new_new_n41503__, new_new_n41504__, new_new_n41505__,
    new_new_n41506__, new_new_n41507__, new_new_n41508__, new_new_n41509__,
    new_new_n41510__, new_new_n41511__, new_new_n41512__, new_new_n41513__,
    new_new_n41514__, new_new_n41515__, new_new_n41516__, new_new_n41517__,
    new_new_n41518__, new_new_n41519__, new_new_n41520__, new_new_n41521__,
    new_new_n41522__, new_new_n41523__, new_new_n41525__, new_new_n41526__,
    new_new_n41527__, new_new_n41528__, new_new_n41529__, new_new_n41530__,
    new_new_n41531__, new_new_n41532__, new_new_n41533__, new_new_n41534__,
    new_new_n41535__, new_new_n41536__, new_new_n41537__, new_new_n41538__,
    new_new_n41539__, new_new_n41540__, new_new_n41541__, new_new_n41542__,
    new_new_n41543__, new_new_n41544__, new_new_n41545__, new_new_n41546__,
    new_new_n41547__, new_new_n41548__, new_new_n41550__, new_new_n41551__,
    new_new_n41552__, new_new_n41553__, new_new_n41554__, new_new_n41555__,
    new_new_n41556__, new_new_n41557__, new_new_n41558__, new_new_n41559__,
    new_new_n41560__, new_new_n41561__, new_new_n41562__, new_new_n41563__,
    new_new_n41564__, new_new_n41565__, new_new_n41566__, new_new_n41567__,
    new_new_n41568__, new_new_n41569__, new_new_n41570__, new_new_n41572__,
    new_new_n41573__, new_new_n41574__, new_new_n41575__, new_new_n41576__,
    new_new_n41577__, new_new_n41578__, new_new_n41579__, new_new_n41580__,
    new_new_n41581__, new_new_n41582__, new_new_n41583__, new_new_n41584__,
    new_new_n41585__, new_new_n41586__, new_new_n41587__, new_new_n41588__,
    new_new_n41589__, new_new_n41590__, new_new_n41591__, new_new_n41592__,
    new_new_n41594__, new_new_n41595__, new_new_n41596__, new_new_n41597__,
    new_new_n41598__, new_new_n41599__, new_new_n41600__, new_new_n41601__,
    new_new_n41602__, new_new_n41603__, new_new_n41604__, new_new_n41605__,
    new_new_n41606__, new_new_n41607__, new_new_n41608__, new_new_n41609__,
    new_new_n41610__, new_new_n41611__, new_new_n41612__, new_new_n41613__,
    new_new_n41614__, new_new_n41615__, new_new_n41617__, new_new_n41618__,
    new_new_n41619__, new_new_n41620__, new_new_n41621__, new_new_n41622__,
    new_new_n41623__, new_new_n41624__, new_new_n41625__, new_new_n41626__,
    new_new_n41627__, new_new_n41628__, new_new_n41629__, new_new_n41630__,
    new_new_n41631__, new_new_n41632__, new_new_n41633__, new_new_n41634__,
    new_new_n41635__, new_new_n41636__, new_new_n41637__, new_new_n41639__,
    new_new_n41640__, new_new_n41641__, new_new_n41642__, new_new_n41643__,
    new_new_n41644__, new_new_n41645__, new_new_n41646__, new_new_n41647__,
    new_new_n41648__, new_new_n41649__, new_new_n41650__, new_new_n41651__,
    new_new_n41652__, new_new_n41653__, new_new_n41654__, new_new_n41655__,
    new_new_n41656__, new_new_n41657__, new_new_n41658__, new_new_n41659__,
    new_new_n41660__, new_new_n41662__, new_new_n41663__, new_new_n41664__,
    new_new_n41665__, new_new_n41666__, new_new_n41667__, new_new_n41668__,
    new_new_n41669__, new_new_n41670__, new_new_n41671__, new_new_n41672__,
    new_new_n41673__, new_new_n41674__, new_new_n41675__, new_new_n41676__,
    new_new_n41677__, new_new_n41678__, new_new_n41679__, new_new_n41680__,
    new_new_n41681__, new_new_n41682__, new_new_n41684__, new_new_n41685__,
    new_new_n41686__, new_new_n41687__, new_new_n41688__, new_new_n41689__,
    new_new_n41690__, new_new_n41691__, new_new_n41692__, new_new_n41693__,
    new_new_n41694__, new_new_n41695__, new_new_n41696__, new_new_n41697__,
    new_new_n41698__, new_new_n41699__, new_new_n41700__, new_new_n41701__,
    new_new_n41702__, new_new_n41703__, new_new_n41704__, new_new_n41705__,
    new_new_n41706__, new_new_n41708__, new_new_n41709__, new_new_n41710__,
    new_new_n41711__, new_new_n41712__, new_new_n41713__, new_new_n41714__,
    new_new_n41715__, new_new_n41716__, new_new_n41717__, new_new_n41718__,
    new_new_n41719__, new_new_n41720__, new_new_n41721__, new_new_n41722__,
    new_new_n41723__, new_new_n41724__, new_new_n41725__, new_new_n41726__,
    new_new_n41727__, new_new_n41728__, new_new_n41730__, new_new_n41731__,
    new_new_n41732__, new_new_n41733__, new_new_n41734__, new_new_n41735__,
    new_new_n41736__, new_new_n41737__, new_new_n41738__, new_new_n41739__,
    new_new_n41740__, new_new_n41741__, new_new_n41742__, new_new_n41743__,
    new_new_n41744__, new_new_n41745__, new_new_n41746__, new_new_n41747__,
    new_new_n41748__, new_new_n41749__, new_new_n41750__, new_new_n41751__,
    new_new_n41753__, new_new_n41754__, new_new_n41755__, new_new_n41756__,
    new_new_n41757__, new_new_n41758__, new_new_n41759__, new_new_n41760__,
    new_new_n41761__, new_new_n41762__, new_new_n41763__, new_new_n41764__,
    new_new_n41765__, new_new_n41766__, new_new_n41767__, new_new_n41768__,
    new_new_n41769__, new_new_n41770__, new_new_n41771__, new_new_n41772__,
    new_new_n41773__, new_new_n41775__, new_new_n41776__, new_new_n41777__,
    new_new_n41778__, new_new_n41779__, new_new_n41780__, new_new_n41781__,
    new_new_n41782__, new_new_n41783__, new_new_n41784__, new_new_n41785__,
    new_new_n41786__, new_new_n41787__, new_new_n41788__, new_new_n41789__,
    new_new_n41790__, new_new_n41791__, new_new_n41792__, new_new_n41793__,
    new_new_n41794__, new_new_n41795__, new_new_n41796__, new_new_n41797__,
    new_new_n41799__, new_new_n41800__, new_new_n41801__, new_new_n41802__,
    new_new_n41803__, new_new_n41804__, new_new_n41805__, new_new_n41806__,
    new_new_n41807__, new_new_n41808__, new_new_n41809__, new_new_n41810__,
    new_new_n41811__, new_new_n41812__, new_new_n41813__, new_new_n41814__,
    new_new_n41815__, new_new_n41816__, new_new_n41817__, new_new_n41818__,
    new_new_n41819__, new_new_n41821__, new_new_n41822__, new_new_n41823__,
    new_new_n41824__, new_new_n41825__, new_new_n41826__, new_new_n41827__,
    new_new_n41828__, new_new_n41829__, new_new_n41830__, new_new_n41831__,
    new_new_n41832__, new_new_n41833__, new_new_n41834__, new_new_n41835__,
    new_new_n41836__, new_new_n41837__, new_new_n41838__, new_new_n41839__,
    new_new_n41840__, new_new_n41841__, new_new_n41842__, new_new_n41844__,
    new_new_n41845__, new_new_n41846__, new_new_n41847__, new_new_n41848__,
    new_new_n41849__, new_new_n41850__, new_new_n41851__, new_new_n41852__,
    new_new_n41853__, new_new_n41854__, new_new_n41855__, new_new_n41856__,
    new_new_n41857__, new_new_n41858__, new_new_n41859__, new_new_n41860__,
    new_new_n41861__, new_new_n41862__, new_new_n41863__, new_new_n41864__,
    new_new_n41866__, new_new_n41867__, new_new_n41868__, new_new_n41869__,
    new_new_n41870__, new_new_n41871__, new_new_n41872__, new_new_n41873__,
    new_new_n41874__, new_new_n41875__, new_new_n41876__, new_new_n41877__,
    new_new_n41878__, new_new_n41879__, new_new_n41880__, new_new_n41881__,
    new_new_n41882__, new_new_n41883__, new_new_n41884__, new_new_n41885__,
    new_new_n41886__, new_new_n41887__, new_new_n41888__, new_new_n41889__,
    new_new_n41891__, new_new_n41892__, new_new_n41893__, new_new_n41894__,
    new_new_n41895__, new_new_n41896__, new_new_n41897__, new_new_n41898__,
    new_new_n41899__, new_new_n41900__, new_new_n41901__, new_new_n41902__,
    new_new_n41903__, new_new_n41904__, new_new_n41905__, new_new_n41906__,
    new_new_n41907__, new_new_n41908__, new_new_n41909__, new_new_n41910__,
    new_new_n41911__, new_new_n41913__, new_new_n41914__, new_new_n41915__,
    new_new_n41916__, new_new_n41917__, new_new_n41918__, new_new_n41919__,
    new_new_n41920__, new_new_n41921__, new_new_n41922__, new_new_n41923__,
    new_new_n41924__, new_new_n41925__, new_new_n41926__, new_new_n41927__,
    new_new_n41928__, new_new_n41929__, new_new_n41930__, new_new_n41931__,
    new_new_n41932__, new_new_n41933__, new_new_n41934__, new_new_n41936__,
    new_new_n41937__, new_new_n41938__, new_new_n41939__, new_new_n41940__,
    new_new_n41941__, new_new_n41942__, new_new_n41943__, new_new_n41944__,
    new_new_n41945__, new_new_n41946__, new_new_n41947__, new_new_n41948__,
    new_new_n41949__, new_new_n41950__, new_new_n41951__, new_new_n41952__,
    new_new_n41953__, new_new_n41954__, new_new_n41955__, new_new_n41956__,
    new_new_n41958__, new_new_n41959__, new_new_n41960__, new_new_n41961__,
    new_new_n41962__, new_new_n41963__, new_new_n41964__, new_new_n41965__,
    new_new_n41966__, new_new_n41967__, new_new_n41968__, new_new_n41969__,
    new_new_n41970__, new_new_n41971__, new_new_n41972__, new_new_n41973__,
    new_new_n41974__, new_new_n41975__, new_new_n41976__, new_new_n41977__,
    new_new_n41978__, new_new_n41979__, new_new_n41980__, new_new_n41982__,
    new_new_n41983__, new_new_n41984__, new_new_n41985__, new_new_n41986__,
    new_new_n41987__, new_new_n41988__, new_new_n41989__, new_new_n41990__,
    new_new_n41991__, new_new_n41992__, new_new_n41993__, new_new_n41994__,
    new_new_n41995__, new_new_n41996__, new_new_n41997__, new_new_n41998__,
    new_new_n41999__, new_new_n42000__, new_new_n42001__, new_new_n42002__,
    new_new_n42004__, new_new_n42005__, new_new_n42006__, new_new_n42007__,
    new_new_n42008__, new_new_n42009__, new_new_n42010__, new_new_n42011__,
    new_new_n42012__, new_new_n42013__, new_new_n42014__, new_new_n42015__,
    new_new_n42016__, new_new_n42017__, new_new_n42018__, new_new_n42019__,
    new_new_n42020__, new_new_n42021__, new_new_n42022__, new_new_n42023__,
    new_new_n42024__, new_new_n42025__, new_new_n42027__, new_new_n42028__,
    new_new_n42029__, new_new_n42030__, new_new_n42031__, new_new_n42032__,
    new_new_n42033__, new_new_n42034__, new_new_n42035__, new_new_n42036__,
    new_new_n42037__, new_new_n42038__, new_new_n42039__, new_new_n42040__,
    new_new_n42041__, new_new_n42042__, new_new_n42043__, new_new_n42044__,
    new_new_n42045__, new_new_n42046__, new_new_n42047__, new_new_n42049__,
    new_new_n42050__, new_new_n42051__, new_new_n42052__, new_new_n42053__,
    new_new_n42054__, new_new_n42055__, new_new_n42056__, new_new_n42057__,
    new_new_n42058__, new_new_n42059__, new_new_n42060__, new_new_n42061__,
    new_new_n42062__, new_new_n42063__, new_new_n42064__, new_new_n42065__,
    new_new_n42066__, new_new_n42067__, new_new_n42068__, new_new_n42069__,
    new_new_n42070__, new_new_n42071__, new_new_n42072__, new_new_n42074__,
    new_new_n42075__, new_new_n42076__, new_new_n42077__, new_new_n42078__,
    new_new_n42079__, new_new_n42080__, new_new_n42081__, new_new_n42082__,
    new_new_n42083__, new_new_n42084__, new_new_n42085__, new_new_n42086__,
    new_new_n42087__, new_new_n42088__, new_new_n42089__, new_new_n42090__,
    new_new_n42091__, new_new_n42092__, new_new_n42093__, new_new_n42094__,
    new_new_n42096__, new_new_n42097__, new_new_n42098__, new_new_n42099__,
    new_new_n42100__, new_new_n42101__, new_new_n42102__, new_new_n42103__,
    new_new_n42104__, new_new_n42105__, new_new_n42106__, new_new_n42107__,
    new_new_n42108__, new_new_n42109__, new_new_n42110__, new_new_n42111__,
    new_new_n42112__, new_new_n42113__, new_new_n42114__, new_new_n42115__,
    new_new_n42116__, new_new_n42117__, new_new_n42119__, new_new_n42120__,
    new_new_n42121__, new_new_n42122__, new_new_n42123__, new_new_n42124__,
    new_new_n42125__, new_new_n42126__, new_new_n42127__, new_new_n42128__,
    new_new_n42129__, new_new_n42130__, new_new_n42131__, new_new_n42132__,
    new_new_n42133__, new_new_n42134__, new_new_n42135__, new_new_n42136__,
    new_new_n42137__, new_new_n42138__, new_new_n42139__, new_new_n42141__,
    new_new_n42142__, new_new_n42143__, new_new_n42144__, new_new_n42145__,
    new_new_n42146__, new_new_n42147__, new_new_n42148__, new_new_n42149__,
    new_new_n42150__, new_new_n42151__, new_new_n42152__, new_new_n42153__,
    new_new_n42154__, new_new_n42155__, new_new_n42156__, new_new_n42157__,
    new_new_n42158__, new_new_n42159__, new_new_n42160__, new_new_n42161__,
    new_new_n42162__, new_new_n42163__, new_new_n42165__, new_new_n42166__,
    new_new_n42167__, new_new_n42168__, new_new_n42169__, new_new_n42170__,
    new_new_n42171__, new_new_n42172__, new_new_n42173__, new_new_n42174__,
    new_new_n42175__, new_new_n42176__, new_new_n42177__, new_new_n42178__,
    new_new_n42179__, new_new_n42180__, new_new_n42181__, new_new_n42182__,
    new_new_n42183__, new_new_n42184__, new_new_n42185__, new_new_n42187__,
    new_new_n42188__, new_new_n42189__, new_new_n42190__, new_new_n42191__,
    new_new_n42192__, new_new_n42193__, new_new_n42194__, new_new_n42195__,
    new_new_n42196__, new_new_n42197__, new_new_n42198__, new_new_n42200__,
    new_new_n42201__, new_new_n42202__, new_new_n42203__, new_new_n42204__,
    new_new_n42205__, new_new_n42206__, new_new_n42207__, new_new_n42208__,
    new_new_n42210__, new_new_n42211__, new_new_n42212__, new_new_n42213__,
    new_new_n42214__, new_new_n42215__, new_new_n42216__, new_new_n42217__,
    new_new_n42218__, new_new_n42219__, new_new_n42220__, new_new_n42222__,
    new_new_n42223__, new_new_n42224__, new_new_n42225__, new_new_n42226__,
    new_new_n42227__, new_new_n42228__, new_new_n42229__, new_new_n42230__,
    new_new_n42232__, new_new_n42233__, new_new_n42234__, new_new_n42235__,
    new_new_n42236__, new_new_n42237__, new_new_n42238__, new_new_n42239__,
    new_new_n42241__, new_new_n42242__, new_new_n42243__, new_new_n42245__,
    new_new_n42246__, new_new_n42247__, new_new_n42249__, new_new_n42250__,
    new_new_n42251__, new_new_n42253__, new_new_n42254__, new_new_n42255__,
    new_new_n42257__, new_new_n42258__, new_new_n42259__, new_new_n42261__,
    new_new_n42262__, new_new_n42263__, new_new_n42265__, new_new_n42266__,
    new_new_n42267__, new_new_n42269__, new_new_n42270__, new_new_n42271__,
    new_new_n42273__, new_new_n42274__, new_new_n42275__, new_new_n42277__,
    new_new_n42278__, new_new_n42279__, new_new_n42281__, new_new_n42282__,
    new_new_n42283__, new_new_n42285__, new_new_n42286__, new_new_n42287__,
    new_new_n42289__, new_new_n42290__, new_new_n42291__, new_new_n42293__,
    new_new_n42294__, new_new_n42295__, new_new_n42297__, new_new_n42298__,
    new_new_n42299__, new_new_n42301__, new_new_n42302__, new_new_n42303__,
    new_new_n42305__, new_new_n42306__, new_new_n42307__, new_new_n42309__,
    new_new_n42310__, new_new_n42311__, new_new_n42313__, new_new_n42314__,
    new_new_n42315__, new_new_n42317__, new_new_n42318__, new_new_n42319__,
    new_new_n42321__, new_new_n42322__, new_new_n42323__, new_new_n42325__,
    new_new_n42326__, new_new_n42327__, new_new_n42329__, new_new_n42330__,
    new_new_n42331__, new_new_n42333__, new_new_n42334__, new_new_n42335__,
    new_new_n42337__, new_new_n42338__, new_new_n42339__, new_new_n42341__,
    new_new_n42342__, new_new_n42343__, new_new_n42345__, new_new_n42346__,
    new_new_n42347__, new_new_n42349__, new_new_n42350__, new_new_n42351__,
    new_new_n42353__, new_new_n42354__, new_new_n42355__, new_new_n42357__,
    new_new_n42358__, new_new_n42359__, new_new_n42361__, new_new_n42362__,
    new_new_n42363__, new_new_n42365__, new_new_n42366__, new_new_n42367__,
    new_new_n42369__, new_new_n42370__, new_new_n42371__, new_new_n42373__,
    new_new_n42374__, new_new_n42375__, new_new_n42377__, new_new_n42378__,
    new_new_n42379__, new_new_n42380__, new_new_n42381__, new_new_n42382__,
    new_new_n42383__, new_new_n42384__, new_new_n42386__, new_new_n42387__,
    new_new_n42388__, new_new_n42390__, new_new_n42391__, new_new_n42392__,
    new_new_n42394__, new_new_n42395__, new_new_n42396__, new_new_n42398__,
    new_new_n42399__, new_new_n42400__, new_new_n42402__, new_new_n42403__,
    new_new_n42404__, new_new_n42406__, new_new_n42407__, new_new_n42408__,
    new_new_n42410__, new_new_n42411__, new_new_n42412__, new_new_n42414__,
    new_new_n42415__, new_new_n42416__, new_new_n42418__, new_new_n42419__,
    new_new_n42420__, new_new_n42422__, new_new_n42423__, new_new_n42424__,
    new_new_n42426__, new_new_n42427__, new_new_n42428__, new_new_n42430__,
    new_new_n42431__, new_new_n42432__, new_new_n42434__, new_new_n42435__,
    new_new_n42436__, new_new_n42438__, new_new_n42439__, new_new_n42440__,
    new_new_n42442__, new_new_n42443__, new_new_n42444__, new_new_n42446__,
    new_new_n42447__, new_new_n42448__, new_new_n42450__, new_new_n42451__,
    new_new_n42452__, new_new_n42454__, new_new_n42455__, new_new_n42456__,
    new_new_n42458__, new_new_n42459__, new_new_n42460__, new_new_n42462__,
    new_new_n42463__, new_new_n42464__, new_new_n42466__, new_new_n42467__,
    new_new_n42468__, new_new_n42470__, new_new_n42471__, new_new_n42472__,
    new_new_n42474__, new_new_n42475__, new_new_n42476__, new_new_n42478__,
    new_new_n42479__, new_new_n42480__, new_new_n42482__, new_new_n42483__,
    new_new_n42484__, new_new_n42486__, new_new_n42487__, new_new_n42488__,
    new_new_n42490__, new_new_n42491__, new_new_n42492__, new_new_n42494__,
    new_new_n42495__, new_new_n42496__, new_new_n42498__, new_new_n42499__,
    new_new_n42500__, new_new_n42502__, new_new_n42503__, new_new_n42504__,
    new_new_n42506__, new_new_n42507__, new_new_n42508__, new_new_n42510__,
    new_new_n42511__, new_new_n42512__, new_new_n42514__, new_new_n42515__,
    new_new_n42516__, new_new_n42518__, new_new_n42519__, new_new_n42520__,
    new_new_n42522__, new_new_n42523__, new_new_n42524__, new_new_n42525__,
    new_new_n42526__, new_new_n42527__, new_new_n42528__, new_new_n42529__,
    new_new_n42531__, new_new_n42532__, new_new_n42533__, new_new_n42535__,
    new_new_n42536__, new_new_n42537__, new_new_n42539__, new_new_n42540__,
    new_new_n42541__, new_new_n42543__, new_new_n42544__, new_new_n42545__,
    new_new_n42547__, new_new_n42548__, new_new_n42549__, new_new_n42551__,
    new_new_n42552__, new_new_n42553__, new_new_n42555__, new_new_n42556__,
    new_new_n42557__, new_new_n42559__, new_new_n42560__, new_new_n42561__,
    new_new_n42563__, new_new_n42564__, new_new_n42565__, new_new_n42567__,
    new_new_n42568__, new_new_n42569__, new_new_n42571__, new_new_n42572__,
    new_new_n42573__, new_new_n42575__, new_new_n42576__, new_new_n42577__,
    new_new_n42579__, new_new_n42580__, new_new_n42581__, new_new_n42583__,
    new_new_n42584__, new_new_n42585__, new_new_n42587__, new_new_n42588__,
    new_new_n42589__, new_new_n42591__, new_new_n42592__, new_new_n42593__,
    new_new_n42595__, new_new_n42596__, new_new_n42597__, new_new_n42599__,
    new_new_n42600__, new_new_n42601__, new_new_n42603__, new_new_n42604__,
    new_new_n42605__, new_new_n42607__, new_new_n42608__, new_new_n42609__,
    new_new_n42611__, new_new_n42612__, new_new_n42613__, new_new_n42615__,
    new_new_n42616__, new_new_n42617__, new_new_n42619__, new_new_n42620__,
    new_new_n42621__, new_new_n42623__, new_new_n42624__, new_new_n42625__,
    new_new_n42627__, new_new_n42628__, new_new_n42629__, new_new_n42631__,
    new_new_n42632__, new_new_n42633__, new_new_n42635__, new_new_n42636__,
    new_new_n42637__, new_new_n42639__, new_new_n42640__, new_new_n42641__,
    new_new_n42643__, new_new_n42644__, new_new_n42645__, new_new_n42647__,
    new_new_n42648__, new_new_n42649__, new_new_n42651__, new_new_n42652__,
    new_new_n42653__, new_new_n42655__, new_new_n42656__, new_new_n42657__,
    new_new_n42659__, new_new_n42660__, new_new_n42661__, new_new_n42663__,
    new_new_n42664__, new_new_n42665__, new_new_n42667__, new_new_n42668__,
    new_new_n42669__, new_new_n42670__, new_new_n42671__, new_new_n42672__,
    new_new_n42673__, new_new_n42674__, new_new_n42675__, new_new_n42676__,
    new_new_n42677__, new_new_n42678__, new_new_n42680__, new_new_n42681__,
    new_new_n42682__, new_new_n42683__, new_new_n42684__, new_new_n42685__,
    new_new_n42686__, new_new_n42687__, new_new_n42688__, new_new_n42689__,
    new_new_n42690__, new_new_n42691__, new_new_n42692__, new_new_n42693__,
    new_new_n42694__, new_new_n42695__, new_new_n42696__, new_new_n42697__,
    new_new_n42698__, new_new_n42699__, new_new_n42700__, new_new_n42702__,
    new_new_n42703__, new_new_n42704__, new_new_n42705__, new_new_n42706__,
    new_new_n42707__, new_new_n42708__, new_new_n42710__, new_new_n42711__,
    new_new_n42712__, new_new_n42713__, new_new_n42714__, new_new_n42715__,
    new_new_n42716__, new_new_n42718__, new_new_n42719__, new_new_n42720__,
    new_new_n42722__, new_new_n42723__, new_new_n42724__, new_new_n42725__,
    new_new_n42726__, new_new_n42727__, new_new_n42728__, new_new_n42730__,
    new_new_n42731__, new_new_n42732__, new_new_n42734__, new_new_n42735__,
    new_new_n42736__, new_new_n42738__, new_new_n42739__, new_new_n42740__,
    new_new_n42742__, new_new_n42743__, new_new_n42744__, new_new_n42746__,
    new_new_n42747__, new_new_n42748__, new_new_n42750__, new_new_n42751__,
    new_new_n42752__, new_new_n42753__, new_new_n42754__, new_new_n42755__,
    new_new_n42756__, new_new_n42757__, new_new_n42759__, new_new_n42760__,
    new_new_n42761__, new_new_n42763__, new_new_n42764__, new_new_n42765__,
    new_new_n42767__, new_new_n42768__, new_new_n42769__, new_new_n42771__,
    new_new_n42772__, new_new_n42773__, new_new_n42775__, new_new_n42776__,
    new_new_n42777__, new_new_n42779__, new_new_n42780__, new_new_n42781__,
    new_new_n42783__, new_new_n42784__, new_new_n42785__, new_new_n42787__,
    new_new_n42788__, new_new_n42789__, new_new_n42791__, new_new_n42792__,
    new_new_n42793__, new_new_n42795__, new_new_n42796__, new_new_n42797__,
    new_new_n42799__, new_new_n42800__, new_new_n42801__, new_new_n42803__,
    new_new_n42804__, new_new_n42805__, new_new_n42807__, new_new_n42808__,
    new_new_n42809__, new_new_n42811__, new_new_n42812__, new_new_n42813__,
    new_new_n42815__, new_new_n42816__, new_new_n42817__, new_new_n42819__,
    new_new_n42820__, new_new_n42821__, new_new_n42823__, new_new_n42824__,
    new_new_n42825__, new_new_n42827__, new_new_n42828__, new_new_n42829__,
    new_new_n42831__, new_new_n42832__, new_new_n42833__, new_new_n42835__,
    new_new_n42836__, new_new_n42837__, new_new_n42839__, new_new_n42840__,
    new_new_n42841__, new_new_n42843__, new_new_n42844__, new_new_n42845__,
    new_new_n42847__, new_new_n42848__, new_new_n42849__, new_new_n42851__,
    new_new_n42852__, new_new_n42853__, new_new_n42855__, new_new_n42856__,
    new_new_n42857__, new_new_n42859__, new_new_n42860__, new_new_n42861__,
    new_new_n42863__, new_new_n42864__, new_new_n42865__, new_new_n42867__,
    new_new_n42868__, new_new_n42869__, new_new_n42871__, new_new_n42872__,
    new_new_n42873__, new_new_n42875__, new_new_n42876__, new_new_n42877__,
    new_new_n42879__, new_new_n42880__, new_new_n42881__, new_new_n42883__,
    new_new_n42884__, new_new_n42885__, new_new_n42887__, new_new_n42888__,
    new_new_n42889__, new_new_n42891__, new_new_n42892__, new_new_n42893__,
    new_new_n42895__, new_new_n42896__, new_new_n42897__, new_new_n42898__,
    new_new_n42899__, new_new_n42900__, new_new_n42901__, new_new_n42902__,
    new_new_n42904__, new_new_n42905__, new_new_n42906__, new_new_n42908__,
    new_new_n42909__, new_new_n42910__, new_new_n42912__, new_new_n42913__,
    new_new_n42914__, new_new_n42916__, new_new_n42917__, new_new_n42918__,
    new_new_n42920__, new_new_n42921__, new_new_n42922__, new_new_n42924__,
    new_new_n42925__, new_new_n42926__, new_new_n42928__, new_new_n42929__,
    new_new_n42930__, new_new_n42932__, new_new_n42933__, new_new_n42934__,
    new_new_n42936__, new_new_n42937__, new_new_n42938__, new_new_n42940__,
    new_new_n42941__, new_new_n42942__, new_new_n42944__, new_new_n42945__,
    new_new_n42946__, new_new_n42948__, new_new_n42949__, new_new_n42950__,
    new_new_n42952__, new_new_n42953__, new_new_n42954__, new_new_n42956__,
    new_new_n42957__, new_new_n42958__, new_new_n42960__, new_new_n42961__,
    new_new_n42962__, new_new_n42964__, new_new_n42965__, new_new_n42966__,
    new_new_n42968__, new_new_n42969__, new_new_n42970__, new_new_n42972__,
    new_new_n42973__, new_new_n42974__, new_new_n42976__, new_new_n42977__,
    new_new_n42978__, new_new_n42980__, new_new_n42981__, new_new_n42982__,
    new_new_n42984__, new_new_n42985__, new_new_n42986__, new_new_n42988__,
    new_new_n42989__, new_new_n42990__, new_new_n42992__, new_new_n42993__,
    new_new_n42994__, new_new_n42996__, new_new_n42997__, new_new_n42998__,
    new_new_n43000__, new_new_n43001__, new_new_n43002__, new_new_n43004__,
    new_new_n43005__, new_new_n43006__, new_new_n43008__, new_new_n43009__,
    new_new_n43010__, new_new_n43012__, new_new_n43013__, new_new_n43014__,
    new_new_n43016__, new_new_n43017__, new_new_n43018__, new_new_n43020__,
    new_new_n43021__, new_new_n43022__, new_new_n43024__, new_new_n43025__,
    new_new_n43026__, new_new_n43028__, new_new_n43029__, new_new_n43030__,
    new_new_n43032__, new_new_n43033__, new_new_n43034__, new_new_n43036__,
    new_new_n43037__, new_new_n43038__, new_new_n43040__, new_new_n43041__,
    new_new_n43042__, new_new_n43043__, new_new_n43044__, new_new_n43045__,
    new_new_n43046__, new_new_n43047__, new_new_n43049__, new_new_n43050__,
    new_new_n43051__, new_new_n43053__, new_new_n43054__, new_new_n43055__,
    new_new_n43057__, new_new_n43058__, new_new_n43059__, new_new_n43061__,
    new_new_n43062__, new_new_n43063__, new_new_n43065__, new_new_n43066__,
    new_new_n43067__, new_new_n43069__, new_new_n43070__, new_new_n43071__,
    new_new_n43073__, new_new_n43074__, new_new_n43075__, new_new_n43077__,
    new_new_n43078__, new_new_n43079__, new_new_n43081__, new_new_n43082__,
    new_new_n43083__, new_new_n43085__, new_new_n43086__, new_new_n43087__,
    new_new_n43089__, new_new_n43090__, new_new_n43091__, new_new_n43093__,
    new_new_n43094__, new_new_n43095__, new_new_n43097__, new_new_n43098__,
    new_new_n43099__, new_new_n43101__, new_new_n43102__, new_new_n43103__,
    new_new_n43105__, new_new_n43106__, new_new_n43107__, new_new_n43109__,
    new_new_n43110__, new_new_n43111__, new_new_n43113__, new_new_n43114__,
    new_new_n43115__, new_new_n43117__, new_new_n43118__, new_new_n43119__,
    new_new_n43121__, new_new_n43122__, new_new_n43123__, new_new_n43125__,
    new_new_n43126__, new_new_n43127__, new_new_n43129__, new_new_n43130__,
    new_new_n43131__, new_new_n43133__, new_new_n43134__, new_new_n43135__,
    new_new_n43137__, new_new_n43138__, new_new_n43139__, new_new_n43141__,
    new_new_n43142__, new_new_n43143__, new_new_n43145__, new_new_n43146__,
    new_new_n43147__, new_new_n43149__, new_new_n43150__, new_new_n43151__,
    new_new_n43153__, new_new_n43154__, new_new_n43155__, new_new_n43157__,
    new_new_n43158__, new_new_n43159__, new_new_n43161__, new_new_n43162__,
    new_new_n43163__, new_new_n43165__, new_new_n43166__, new_new_n43167__,
    new_new_n43169__, new_new_n43170__, new_new_n43171__, new_new_n43173__,
    new_new_n43174__, new_new_n43175__, new_new_n43177__, new_new_n43178__,
    new_new_n43179__, new_new_n43181__, new_new_n43182__, new_new_n43183__,
    new_new_n43185__, new_new_n43186__, new_new_n43187__, new_new_n43188__,
    new_new_n43189__, new_new_n43190__, new_new_n43191__, new_new_n43192__,
    new_new_n43193__, new_new_n43194__, new_new_n43195__, new_new_n43196__,
    new_new_n43198__, new_new_n43199__, new_new_n43200__, new_new_n43202__,
    new_new_n43203__, new_new_n43204__, new_new_n43205__, new_new_n43206__,
    new_new_n43207__, new_new_n43208__, new_new_n43210__, new_new_n43212__,
    new_new_n43214__, new_new_n43215__, new_new_n43216__, new_new_n43217__,
    new_new_n43219__, new_new_n43220__, new_new_n43221__, new_new_n43222__,
    new_new_n43223__, new_new_n43224__, new_new_n43225__, new_new_n43226__,
    new_new_n43228__, new_new_n43229__, new_new_n43230__, new_new_n43232__,
    new_new_n43233__, new_new_n43234__, new_new_n43236__, new_new_n43237__,
    new_new_n43238__, new_new_n43240__, new_new_n43241__, new_new_n43242__,
    new_new_n43244__, new_new_n43245__, new_new_n43246__, new_new_n43248__,
    new_new_n43249__, new_new_n43250__, new_new_n43252__, new_new_n43253__,
    new_new_n43254__, new_new_n43256__, new_new_n43257__, new_new_n43258__,
    new_new_n43260__, new_new_n43261__, new_new_n43262__, new_new_n43264__,
    new_new_n43265__, new_new_n43266__, new_new_n43268__, new_new_n43269__,
    new_new_n43270__, new_new_n43272__, new_new_n43273__, new_new_n43274__,
    new_new_n43276__, new_new_n43277__, new_new_n43278__, new_new_n43280__,
    new_new_n43281__, new_new_n43282__, new_new_n43284__, new_new_n43285__,
    new_new_n43286__, new_new_n43288__, new_new_n43289__, new_new_n43290__,
    new_new_n43292__, new_new_n43293__, new_new_n43294__, new_new_n43296__,
    new_new_n43297__, new_new_n43298__, new_new_n43300__, new_new_n43301__,
    new_new_n43302__, new_new_n43304__, new_new_n43305__, new_new_n43306__,
    new_new_n43308__, new_new_n43309__, new_new_n43310__, new_new_n43312__,
    new_new_n43313__, new_new_n43314__, new_new_n43316__, new_new_n43317__,
    new_new_n43318__, new_new_n43320__, new_new_n43321__, new_new_n43322__,
    new_new_n43324__, new_new_n43325__, new_new_n43326__, new_new_n43328__,
    new_new_n43329__, new_new_n43330__, new_new_n43332__, new_new_n43333__,
    new_new_n43334__, new_new_n43336__, new_new_n43337__, new_new_n43338__,
    new_new_n43340__, new_new_n43341__, new_new_n43342__, new_new_n43344__,
    new_new_n43345__, new_new_n43346__, new_new_n43348__, new_new_n43349__,
    new_new_n43350__, new_new_n43352__, new_new_n43353__, new_new_n43354__,
    new_new_n43356__, new_new_n43357__, new_new_n43358__, new_new_n43360__,
    new_new_n43361__, new_new_n43362__, new_new_n43364__, new_new_n43365__,
    new_new_n43366__, new_new_n43367__, new_new_n43368__, new_new_n43369__,
    new_new_n43370__, new_new_n43371__, new_new_n43373__, new_new_n43374__,
    new_new_n43375__, new_new_n43377__, new_new_n43378__, new_new_n43379__,
    new_new_n43381__, new_new_n43382__, new_new_n43383__, new_new_n43385__,
    new_new_n43386__, new_new_n43387__, new_new_n43389__, new_new_n43390__,
    new_new_n43391__, new_new_n43393__, new_new_n43394__, new_new_n43395__,
    new_new_n43397__, new_new_n43398__, new_new_n43399__, new_new_n43401__,
    new_new_n43402__, new_new_n43403__, new_new_n43405__, new_new_n43406__,
    new_new_n43407__, new_new_n43409__, new_new_n43410__, new_new_n43411__,
    new_new_n43413__, new_new_n43414__, new_new_n43415__, new_new_n43417__,
    new_new_n43418__, new_new_n43419__, new_new_n43421__, new_new_n43422__,
    new_new_n43423__, new_new_n43425__, new_new_n43426__, new_new_n43427__,
    new_new_n43429__, new_new_n43430__, new_new_n43431__, new_new_n43433__,
    new_new_n43434__, new_new_n43435__, new_new_n43437__, new_new_n43438__,
    new_new_n43439__, new_new_n43441__, new_new_n43442__, new_new_n43443__,
    new_new_n43445__, new_new_n43446__, new_new_n43447__, new_new_n43449__,
    new_new_n43450__, new_new_n43451__, new_new_n43453__, new_new_n43454__,
    new_new_n43455__, new_new_n43457__, new_new_n43458__, new_new_n43459__,
    new_new_n43461__, new_new_n43462__, new_new_n43463__, new_new_n43465__,
    new_new_n43466__, new_new_n43467__, new_new_n43469__, new_new_n43470__,
    new_new_n43471__, new_new_n43473__, new_new_n43474__, new_new_n43475__,
    new_new_n43477__, new_new_n43478__, new_new_n43479__, new_new_n43481__,
    new_new_n43482__, new_new_n43483__, new_new_n43485__, new_new_n43486__,
    new_new_n43487__, new_new_n43489__, new_new_n43490__, new_new_n43491__,
    new_new_n43493__, new_new_n43494__, new_new_n43495__, new_new_n43497__,
    new_new_n43498__, new_new_n43499__, new_new_n43501__, new_new_n43502__,
    new_new_n43503__, new_new_n43505__, new_new_n43506__, new_new_n43507__,
    new_new_n43509__, new_new_n43510__, new_new_n43511__, new_new_n43512__,
    new_new_n43513__, new_new_n43514__, new_new_n43515__, new_new_n43516__,
    new_new_n43518__, new_new_n43519__, new_new_n43520__, new_new_n43522__,
    new_new_n43523__, new_new_n43524__, new_new_n43526__, new_new_n43527__,
    new_new_n43528__, new_new_n43530__, new_new_n43531__, new_new_n43532__,
    new_new_n43534__, new_new_n43535__, new_new_n43536__, new_new_n43538__,
    new_new_n43539__, new_new_n43540__, new_new_n43542__, new_new_n43543__,
    new_new_n43544__, new_new_n43546__, new_new_n43547__, new_new_n43548__,
    new_new_n43550__, new_new_n43551__, new_new_n43552__, new_new_n43554__,
    new_new_n43555__, new_new_n43556__, new_new_n43558__, new_new_n43559__,
    new_new_n43560__, new_new_n43562__, new_new_n43563__, new_new_n43564__,
    new_new_n43566__, new_new_n43567__, new_new_n43568__, new_new_n43570__,
    new_new_n43571__, new_new_n43572__, new_new_n43574__, new_new_n43575__,
    new_new_n43576__, new_new_n43578__, new_new_n43579__, new_new_n43580__,
    new_new_n43582__, new_new_n43583__, new_new_n43584__, new_new_n43586__,
    new_new_n43587__, new_new_n43588__, new_new_n43590__, new_new_n43591__,
    new_new_n43592__, new_new_n43594__, new_new_n43595__, new_new_n43596__,
    new_new_n43598__, new_new_n43599__, new_new_n43600__, new_new_n43602__,
    new_new_n43603__, new_new_n43604__, new_new_n43606__, new_new_n43607__,
    new_new_n43608__, new_new_n43610__, new_new_n43611__, new_new_n43612__,
    new_new_n43614__, new_new_n43615__, new_new_n43616__, new_new_n43618__,
    new_new_n43619__, new_new_n43620__, new_new_n43622__, new_new_n43623__,
    new_new_n43624__, new_new_n43626__, new_new_n43627__, new_new_n43628__,
    new_new_n43630__, new_new_n43631__, new_new_n43632__, new_new_n43634__,
    new_new_n43635__, new_new_n43636__, new_new_n43638__, new_new_n43639__,
    new_new_n43640__, new_new_n43642__, new_new_n43643__, new_new_n43644__,
    new_new_n43646__, new_new_n43647__, new_new_n43648__, new_new_n43650__,
    new_new_n43651__, new_new_n43652__, new_new_n43654__, new_new_n43655__,
    new_new_n43656__, new_new_n43657__, new_new_n43658__, new_new_n43659__,
    new_new_n43660__, new_new_n43661__, new_new_n43663__, new_new_n43664__,
    new_new_n43665__, new_new_n43667__, new_new_n43668__, new_new_n43669__,
    new_new_n43671__, new_new_n43672__, new_new_n43673__, new_new_n43675__,
    new_new_n43676__, new_new_n43677__, new_new_n43679__, new_new_n43680__,
    new_new_n43681__, new_new_n43683__, new_new_n43684__, new_new_n43685__,
    new_new_n43687__, new_new_n43688__, new_new_n43689__, new_new_n43691__,
    new_new_n43692__, new_new_n43693__, new_new_n43695__, new_new_n43696__,
    new_new_n43697__, new_new_n43699__, new_new_n43700__, new_new_n43701__,
    new_new_n43703__, new_new_n43704__, new_new_n43705__, new_new_n43707__,
    new_new_n43708__, new_new_n43709__, new_new_n43711__, new_new_n43712__,
    new_new_n43713__, new_new_n43715__, new_new_n43716__, new_new_n43717__,
    new_new_n43719__, new_new_n43720__, new_new_n43721__, new_new_n43723__,
    new_new_n43724__, new_new_n43725__, new_new_n43727__, new_new_n43728__,
    new_new_n43729__, new_new_n43731__, new_new_n43732__, new_new_n43733__,
    new_new_n43735__, new_new_n43736__, new_new_n43737__, new_new_n43739__,
    new_new_n43740__, new_new_n43741__, new_new_n43743__, new_new_n43744__,
    new_new_n43745__, new_new_n43747__, new_new_n43748__, new_new_n43749__,
    new_new_n43751__, new_new_n43752__, new_new_n43753__, new_new_n43755__,
    new_new_n43756__, new_new_n43757__, new_new_n43759__, new_new_n43760__,
    new_new_n43761__, new_new_n43763__, new_new_n43764__, new_new_n43765__,
    new_new_n43767__, new_new_n43768__, new_new_n43769__, new_new_n43771__,
    new_new_n43772__, new_new_n43773__, new_new_n43775__, new_new_n43776__,
    new_new_n43777__, new_new_n43779__, new_new_n43780__, new_new_n43781__,
    new_new_n43783__, new_new_n43784__, new_new_n43785__, new_new_n43787__,
    new_new_n43788__, new_new_n43789__, new_new_n43791__, new_new_n43792__,
    new_new_n43793__, new_new_n43795__, new_new_n43796__, new_new_n43797__,
    new_new_n43799__, new_new_n43800__, new_new_n43801__, new_new_n43802__,
    new_new_n43803__, new_new_n43804__, new_new_n43805__, new_new_n43806__,
    new_new_n43808__, new_new_n43809__, new_new_n43810__, new_new_n43812__,
    new_new_n43813__, new_new_n43814__, new_new_n43816__, new_new_n43817__,
    new_new_n43818__, new_new_n43820__, new_new_n43821__, new_new_n43822__,
    new_new_n43824__, new_new_n43825__, new_new_n43826__, new_new_n43828__,
    new_new_n43829__, new_new_n43830__, new_new_n43832__, new_new_n43833__,
    new_new_n43834__, new_new_n43836__, new_new_n43837__, new_new_n43838__,
    new_new_n43840__, new_new_n43841__, new_new_n43842__, new_new_n43844__,
    new_new_n43845__, new_new_n43846__, new_new_n43848__, new_new_n43849__,
    new_new_n43850__, new_new_n43852__, new_new_n43853__, new_new_n43854__,
    new_new_n43856__, new_new_n43857__, new_new_n43858__, new_new_n43860__,
    new_new_n43861__, new_new_n43862__, new_new_n43864__, new_new_n43865__,
    new_new_n43866__, new_new_n43868__, new_new_n43869__, new_new_n43870__,
    new_new_n43872__, new_new_n43873__, new_new_n43874__, new_new_n43876__,
    new_new_n43877__, new_new_n43878__, new_new_n43880__, new_new_n43881__,
    new_new_n43882__, new_new_n43884__, new_new_n43885__, new_new_n43886__,
    new_new_n43888__, new_new_n43889__, new_new_n43890__, new_new_n43892__,
    new_new_n43893__, new_new_n43894__, new_new_n43896__, new_new_n43897__,
    new_new_n43898__, new_new_n43900__, new_new_n43901__, new_new_n43902__,
    new_new_n43904__, new_new_n43905__, new_new_n43906__, new_new_n43908__,
    new_new_n43909__, new_new_n43910__, new_new_n43912__, new_new_n43913__,
    new_new_n43914__, new_new_n43916__, new_new_n43917__, new_new_n43918__,
    new_new_n43920__, new_new_n43921__, new_new_n43922__, new_new_n43924__,
    new_new_n43925__, new_new_n43926__, new_new_n43928__, new_new_n43929__,
    new_new_n43930__, new_new_n43932__, new_new_n43933__, new_new_n43934__,
    new_new_n43936__, new_new_n43937__, new_new_n43938__, new_new_n43940__,
    new_new_n43941__, new_new_n43942__, new_new_n43944__, new_new_n43945__,
    new_new_n43946__, new_new_n43947__, new_new_n43948__, new_new_n43949__,
    new_new_n43950__, new_new_n43951__, new_new_n43953__, new_new_n43954__,
    new_new_n43955__, new_new_n43957__, new_new_n43958__, new_new_n43959__,
    new_new_n43961__, new_new_n43962__, new_new_n43963__, new_new_n43965__,
    new_new_n43966__, new_new_n43967__, new_new_n43969__, new_new_n43970__,
    new_new_n43971__, new_new_n43973__, new_new_n43974__, new_new_n43975__,
    new_new_n43977__, new_new_n43978__, new_new_n43979__, new_new_n43981__,
    new_new_n43982__, new_new_n43983__, new_new_n43985__, new_new_n43986__,
    new_new_n43987__, new_new_n43989__, new_new_n43990__, new_new_n43991__,
    new_new_n43993__, new_new_n43994__, new_new_n43995__, new_new_n43997__,
    new_new_n43998__, new_new_n43999__, new_new_n44001__, new_new_n44002__,
    new_new_n44003__, new_new_n44005__, new_new_n44006__, new_new_n44007__,
    new_new_n44009__, new_new_n44010__, new_new_n44011__, new_new_n44013__,
    new_new_n44014__, new_new_n44015__, new_new_n44017__, new_new_n44018__,
    new_new_n44019__, new_new_n44021__, new_new_n44022__, new_new_n44023__,
    new_new_n44025__, new_new_n44026__, new_new_n44027__, new_new_n44029__,
    new_new_n44030__, new_new_n44031__, new_new_n44033__, new_new_n44034__,
    new_new_n44035__, new_new_n44037__, new_new_n44038__, new_new_n44039__,
    new_new_n44041__, new_new_n44042__, new_new_n44043__, new_new_n44045__,
    new_new_n44046__, new_new_n44047__, new_new_n44049__, new_new_n44050__,
    new_new_n44051__, new_new_n44053__, new_new_n44054__, new_new_n44055__,
    new_new_n44057__, new_new_n44058__, new_new_n44059__, new_new_n44061__,
    new_new_n44062__, new_new_n44063__, new_new_n44065__, new_new_n44066__,
    new_new_n44067__, new_new_n44069__, new_new_n44070__, new_new_n44071__,
    new_new_n44073__, new_new_n44074__, new_new_n44075__, new_new_n44077__,
    new_new_n44078__, new_new_n44079__, new_new_n44081__, new_new_n44082__,
    new_new_n44083__, new_new_n44085__, new_new_n44086__, new_new_n44087__,
    new_new_n44089__, new_new_n44090__, new_new_n44091__, new_new_n44092__,
    new_new_n44093__, new_new_n44094__, new_new_n44095__, new_new_n44096__,
    new_new_n44097__, new_new_n44098__, new_new_n44099__, new_new_n44100__,
    new_new_n44101__, new_new_n44102__, new_new_n44103__, new_new_n44104__,
    new_new_n44105__, new_new_n44106__, new_new_n44107__, new_new_n44108__,
    new_new_n44109__, new_new_n44110__, new_new_n44111__, new_new_n44112__,
    new_new_n44113__, new_new_n44114__, new_new_n44115__, new_new_n44116__,
    new_new_n44117__, new_new_n44118__, new_new_n44119__, new_new_n44120__,
    new_new_n44121__, new_new_n44122__, new_new_n44123__, new_new_n44124__,
    new_new_n44125__, new_new_n44126__, new_new_n44127__, new_new_n44128__,
    new_new_n44129__, new_new_n44130__, new_new_n44131__, new_new_n44132__,
    new_new_n44133__, new_new_n44134__, new_new_n44135__, new_new_n44136__,
    new_new_n44137__, new_new_n44138__, new_new_n44139__, new_new_n44140__,
    new_new_n44141__, new_new_n44142__, new_new_n44143__, new_new_n44144__,
    new_new_n44145__, new_new_n44146__, new_new_n44147__, new_new_n44148__,
    new_new_n44149__, new_new_n44150__, new_new_n44151__, new_new_n44152__,
    new_new_n44153__, new_new_n44154__, new_new_n44155__, new_new_n44156__,
    new_new_n44157__, new_new_n44158__, new_new_n44159__, new_new_n44160__,
    new_new_n44161__, new_new_n44162__, new_new_n44163__, new_new_n44164__,
    new_new_n44165__, new_new_n44166__, new_new_n44167__, new_new_n44168__,
    new_new_n44169__, new_new_n44170__, new_new_n44171__, new_new_n44172__,
    new_new_n44173__, new_new_n44174__, new_new_n44175__, new_new_n44176__,
    new_new_n44177__, new_new_n44179__, new_new_n44180__, new_new_n44181__,
    new_new_n44182__, new_new_n44183__, new_new_n44184__, new_new_n44185__,
    new_new_n44186__, new_new_n44187__, new_new_n44188__, new_new_n44189__,
    new_new_n44190__, new_new_n44191__, new_new_n44192__, new_new_n44193__,
    new_new_n44194__, new_new_n44195__, new_new_n44196__, new_new_n44197__,
    new_new_n44198__, new_new_n44199__, new_new_n44200__, new_new_n44201__,
    new_new_n44202__, new_new_n44203__, new_new_n44204__, new_new_n44205__,
    new_new_n44206__, new_new_n44207__, new_new_n44208__, new_new_n44209__,
    new_new_n44210__, new_new_n44211__, new_new_n44212__, new_new_n44213__,
    new_new_n44215__, new_new_n44216__, new_new_n44217__, new_new_n44218__,
    new_new_n44219__, new_new_n44220__, new_new_n44221__, new_new_n44222__,
    new_new_n44223__, new_new_n44224__, new_new_n44226__, new_new_n44227__,
    new_new_n44228__, new_new_n44229__, new_new_n44230__, new_new_n44231__,
    new_new_n44232__, new_new_n44233__, new_new_n44234__, new_new_n44236__,
    new_new_n44237__, new_new_n44238__, new_new_n44239__, new_new_n44240__,
    new_new_n44241__, new_new_n44242__, new_new_n44243__, new_new_n44244__,
    new_new_n44245__, new_new_n44246__, new_new_n44248__, new_new_n44249__,
    new_new_n44250__, new_new_n44251__, new_new_n44252__, new_new_n44253__,
    new_new_n44254__, new_new_n44255__, new_new_n44256__, new_new_n44257__,
    new_new_n44259__, new_new_n44260__, new_new_n44261__, new_new_n44262__,
    new_new_n44263__, new_new_n44264__, new_new_n44265__, new_new_n44266__,
    new_new_n44267__, new_new_n44268__, new_new_n44270__, new_new_n44271__,
    new_new_n44272__, new_new_n44273__, new_new_n44274__, new_new_n44275__,
    new_new_n44276__, new_new_n44277__, new_new_n44278__, new_new_n44279__,
    new_new_n44281__, new_new_n44282__, new_new_n44283__, new_new_n44284__,
    new_new_n44285__, new_new_n44286__, new_new_n44287__, new_new_n44288__,
    new_new_n44289__, new_new_n44290__, new_new_n44291__, new_new_n44292__,
    new_new_n44294__, new_new_n44295__, new_new_n44296__, new_new_n44297__,
    new_new_n44298__, new_new_n44299__, new_new_n44300__, new_new_n44301__,
    new_new_n44302__, new_new_n44303__, new_new_n44305__, new_new_n44306__,
    new_new_n44307__, new_new_n44308__, new_new_n44309__, new_new_n44310__,
    new_new_n44311__, new_new_n44312__, new_new_n44313__, new_new_n44314__,
    new_new_n44315__, new_new_n44316__, new_new_n44318__, new_new_n44319__,
    new_new_n44330__, new_new_n44331__, new_new_n44333__, new_new_n44334__,
    new_new_n44336__, new_new_n44337__, new_new_n44338__, new_new_n44339__,
    new_new_n44341__, new_new_n44342__, new_new_n44343__, new_new_n44344__,
    new_new_n44347__, new_new_n44348__, new_new_n44350__, new_new_n44352__,
    new_new_n44354__, new_new_n44356__, new_new_n44357__, new_new_n44358__,
    new_new_n44359__, new_new_n44360__, new_new_n44361__, new_new_n44362__,
    new_new_n44363__, new_new_n44364__, new_new_n44365__, new_new_n44366__,
    new_new_n44367__, new_new_n44368__, new_new_n44369__, new_new_n44370__,
    new_new_n44371__, new_new_n44372__, new_new_n44373__, new_new_n44374__,
    new_new_n44375__, new_new_n44376__, new_new_n44377__, new_new_n44378__,
    new_new_n44379__, new_new_n44380__, new_new_n44381__, new_new_n44385__,
    new_new_n44386__, new_new_n44387__, new_new_n44389__, new_new_n44390__,
    new_new_n44391__, new_new_n44393__, new_new_n44394__, new_new_n44395__,
    new_new_n44397__, new_new_n44398__, new_new_n44399__, new_new_n44401__,
    new_new_n44402__, new_new_n44403__, new_new_n44405__, new_new_n44406__,
    new_new_n44407__, new_new_n44409__, new_new_n44410__, new_new_n44411__,
    new_new_n44413__, new_new_n44414__, new_new_n44415__, new_new_n44417__,
    new_new_n44418__, new_new_n44419__, new_new_n44421__, new_new_n44422__,
    new_new_n44423__, new_new_n44425__, new_new_n44426__, new_new_n44427__,
    new_new_n44429__, new_new_n44430__, new_new_n44431__, new_new_n44433__,
    new_new_n44434__, new_new_n44435__, new_new_n44437__, new_new_n44438__,
    new_new_n44439__, new_new_n44441__, new_new_n44442__, new_new_n44443__,
    new_new_n44445__, new_new_n44446__, new_new_n44447__, new_new_n44449__,
    new_new_n44450__, new_new_n44451__, new_new_n44453__, new_new_n44454__,
    new_new_n44455__, new_new_n44457__, new_new_n44458__, new_new_n44459__,
    new_new_n44461__, new_new_n44462__, new_new_n44463__, new_new_n44465__,
    new_new_n44466__, new_new_n44467__, new_new_n44469__, new_new_n44470__,
    new_new_n44471__, new_new_n44473__, new_new_n44474__, new_new_n44475__,
    new_new_n44477__, new_new_n44478__, new_new_n44479__, new_new_n44481__,
    new_new_n44482__, new_new_n44483__, new_new_n44485__, new_new_n44486__,
    new_new_n44487__, new_new_n44489__, new_new_n44490__, new_new_n44491__,
    new_new_n44493__, new_new_n44494__, new_new_n44495__, new_new_n44497__,
    new_new_n44498__, new_new_n44499__, new_new_n44501__, new_new_n44502__,
    new_new_n44503__, new_new_n44505__, new_new_n44506__, new_new_n44507__,
    new_new_n44509__, new_new_n44510__, new_new_n44511__, new_new_n44513__,
    new_new_n44514__, new_new_n44515__, new_new_n44516__, new_new_n44517__,
    new_new_n44518__, new_new_n44519__, new_new_n44520__, new_new_n44521__,
    new_new_n44522__, new_new_n44523__, new_new_n44524__, new_new_n44525__,
    new_new_n44526__, new_new_n44527__, new_new_n44529__, new_new_n44530__,
    new_new_n44531__, new_new_n44532__, new_new_n44533__, new_new_n44534__,
    new_new_n44535__, new_new_n44537__, new_new_n44538__, new_new_n44539__,
    new_new_n44540__, new_new_n44541__, new_new_n44542__, new_new_n44543__,
    new_new_n44545__, new_new_n44546__, new_new_n44547__, new_new_n44548__,
    new_new_n44549__, new_new_n44550__, new_new_n44551__, new_new_n44553__,
    new_new_n44554__, new_new_n44555__, new_new_n44556__, new_new_n44557__,
    new_new_n44558__, new_new_n44559__, new_new_n44561__, new_new_n44562__,
    new_new_n44563__, new_new_n44564__, new_new_n44565__, new_new_n44566__,
    new_new_n44567__, new_new_n44569__, new_new_n44570__, new_new_n44571__,
    new_new_n44572__, new_new_n44573__, new_new_n44574__, new_new_n44575__,
    new_new_n44577__, new_new_n44578__, new_new_n44579__, new_new_n44580__,
    new_new_n44581__, new_new_n44582__, new_new_n44583__, new_new_n44585__,
    new_new_n44586__, new_new_n44587__, new_new_n44588__, new_new_n44589__,
    new_new_n44590__, new_new_n44591__, new_new_n44593__, new_new_n44594__,
    new_new_n44595__, new_new_n44596__, new_new_n44597__, new_new_n44598__,
    new_new_n44599__, new_new_n44601__, new_new_n44602__, new_new_n44603__,
    new_new_n44604__, new_new_n44605__, new_new_n44606__, new_new_n44607__,
    new_new_n44609__, new_new_n44610__, new_new_n44611__, new_new_n44612__,
    new_new_n44613__, new_new_n44614__, new_new_n44615__, new_new_n44617__,
    new_new_n44618__, new_new_n44619__, new_new_n44620__, new_new_n44621__,
    new_new_n44622__, new_new_n44623__, new_new_n44625__, new_new_n44626__,
    new_new_n44627__, new_new_n44628__, new_new_n44629__, new_new_n44630__,
    new_new_n44631__, new_new_n44633__, new_new_n44634__, new_new_n44635__,
    new_new_n44636__, new_new_n44637__, new_new_n44638__, new_new_n44639__,
    new_new_n44641__, new_new_n44642__, new_new_n44643__, new_new_n44644__,
    new_new_n44645__, new_new_n44646__, new_new_n44647__, new_new_n44649__,
    new_new_n44650__, new_new_n44651__, new_new_n44652__, new_new_n44653__,
    new_new_n44654__, new_new_n44655__, new_new_n44657__, new_new_n44658__,
    new_new_n44659__, new_new_n44660__, new_new_n44661__, new_new_n44662__,
    new_new_n44663__, new_new_n44665__, new_new_n44666__, new_new_n44667__,
    new_new_n44668__, new_new_n44669__, new_new_n44670__, new_new_n44671__,
    new_new_n44673__, new_new_n44674__, new_new_n44675__, new_new_n44676__,
    new_new_n44677__, new_new_n44678__, new_new_n44679__, new_new_n44681__,
    new_new_n44682__, new_new_n44683__, new_new_n44684__, new_new_n44685__,
    new_new_n44686__, new_new_n44687__, new_new_n44689__, new_new_n44690__,
    new_new_n44691__, new_new_n44692__, new_new_n44693__, new_new_n44694__,
    new_new_n44695__, new_new_n44697__, new_new_n44698__, new_new_n44699__,
    new_new_n44700__, new_new_n44701__, new_new_n44702__, new_new_n44703__,
    new_new_n44705__, new_new_n44706__, new_new_n44707__, new_new_n44708__,
    new_new_n44709__, new_new_n44710__, new_new_n44711__, new_new_n44713__,
    new_new_n44714__, new_new_n44715__, new_new_n44716__, new_new_n44717__,
    new_new_n44718__, new_new_n44719__, new_new_n44721__, new_new_n44722__,
    new_new_n44723__, new_new_n44724__, new_new_n44725__, new_new_n44726__,
    new_new_n44727__, new_new_n44729__, new_new_n44730__, new_new_n44731__,
    new_new_n44732__, new_new_n44733__, new_new_n44734__, new_new_n44735__,
    new_new_n44737__, new_new_n44738__, new_new_n44739__, new_new_n44740__,
    new_new_n44741__, new_new_n44742__, new_new_n44743__, new_new_n44745__,
    new_new_n44746__, new_new_n44747__, new_new_n44748__, new_new_n44749__,
    new_new_n44750__, new_new_n44751__, new_new_n44753__, new_new_n44754__,
    new_new_n44755__, new_new_n44756__, new_new_n44757__, new_new_n44758__,
    new_new_n44759__, new_new_n44761__, new_new_n44762__, new_new_n44763__,
    new_new_n44764__, new_new_n44765__, new_new_n44766__, new_new_n44767__,
    new_new_n44769__, new_new_n44770__, new_new_n44771__, new_new_n44772__,
    new_new_n44773__, new_new_n44774__, new_new_n44775__, new_new_n44777__,
    new_new_n44778__, new_new_n44779__, new_new_n44780__, new_new_n44781__,
    new_new_n44782__, new_new_n44783__, new_new_n44784__, new_new_n44785__,
    new_new_n44786__, new_new_n44787__, new_new_n44788__, new_new_n44789__,
    new_new_n44790__, new_new_n44791__, new_new_n44792__, new_new_n44793__,
    new_new_n44794__, new_new_n44795__, new_new_n44796__, new_new_n44797__,
    new_new_n44798__, new_new_n44799__, new_new_n44800__, new_new_n44801__,
    new_new_n44802__, new_new_n44803__, new_new_n44804__, new_new_n44805__,
    new_new_n44806__, new_new_n44807__, new_new_n44808__, new_new_n44809__,
    new_new_n44810__, new_new_n44811__, new_new_n44812__, new_new_n44813__,
    new_new_n44814__, new_new_n44815__, new_new_n44816__, new_new_n44817__,
    new_new_n44818__, new_new_n44819__, new_new_n44820__, new_new_n44821__,
    new_new_n44822__, new_new_n44823__, new_new_n44824__, new_new_n44825__,
    new_new_n44826__, new_new_n44827__, new_new_n44828__, new_new_n44829__,
    new_new_n44830__, new_new_n44831__, new_new_n44832__, new_new_n44833__,
    new_new_n44834__, new_new_n44835__, new_new_n44836__, new_new_n44837__,
    new_new_n44838__, new_new_n44839__, new_new_n44840__, new_new_n44841__,
    new_new_n44842__, new_new_n44843__, new_new_n44844__, new_new_n44845__,
    new_new_n44847__, new_new_n44848__, new_new_n44849__, new_new_n44850__,
    new_new_n44851__, new_new_n44852__, new_new_n44853__, new_new_n44854__,
    new_new_n44855__, new_new_n44856__, new_new_n44857__, new_new_n44858__,
    new_new_n44859__, new_new_n44860__, new_new_n44861__, new_new_n44862__,
    new_new_n44863__, new_new_n44864__, new_new_n44865__, new_new_n44866__,
    new_new_n44867__, new_new_n44868__, new_new_n44869__, new_new_n44870__,
    new_new_n44871__, new_new_n44872__, new_new_n44873__, new_new_n44874__,
    new_new_n44875__, new_new_n44876__, new_new_n44877__, new_new_n44878__,
    new_new_n44879__, new_new_n44880__, new_new_n44881__, new_new_n44882__,
    new_new_n44884__, new_new_n44885__, new_new_n44886__, new_new_n44887__,
    new_new_n44888__, new_new_n44889__, new_new_n44890__, new_new_n44891__,
    new_new_n44892__, new_new_n44893__, new_new_n44894__, new_new_n44895__,
    new_new_n44896__, new_new_n44897__, new_new_n44898__, new_new_n44899__,
    new_new_n44900__, new_new_n44901__, new_new_n44902__, new_new_n44903__,
    new_new_n44904__, new_new_n44905__, new_new_n44906__, new_new_n44907__,
    new_new_n44908__, new_new_n44909__, new_new_n44910__, new_new_n44911__,
    new_new_n44912__, new_new_n44913__, new_new_n44914__, new_new_n44915__,
    new_new_n44916__, new_new_n44917__, new_new_n44918__, new_new_n44919__,
    new_new_n44920__, new_new_n44921__, new_new_n44923__, new_new_n44924__,
    new_new_n44925__, new_new_n44926__, new_new_n44927__, new_new_n44928__,
    new_new_n44929__, new_new_n44930__, new_new_n44931__, new_new_n44932__,
    new_new_n44933__, new_new_n44934__, new_new_n44935__, new_new_n44936__,
    new_new_n44937__, new_new_n44938__, new_new_n44939__, new_new_n44940__,
    new_new_n44941__, new_new_n44942__, new_new_n44943__, new_new_n44944__,
    new_new_n44945__, new_new_n44946__, new_new_n44947__, new_new_n44948__,
    new_new_n44949__, new_new_n44950__, new_new_n44951__, new_new_n44952__,
    new_new_n44953__, new_new_n44954__, new_new_n44955__, new_new_n44956__,
    new_new_n44957__, new_new_n44958__, new_new_n44959__, new_new_n44960__,
    new_new_n44962__, new_new_n44963__, new_new_n44964__, new_new_n44965__,
    new_new_n44966__, new_new_n44967__, new_new_n44968__, new_new_n44969__,
    new_new_n44970__, new_new_n44971__, new_new_n44972__, new_new_n44973__,
    new_new_n44974__, new_new_n44975__, new_new_n44976__, new_new_n44977__,
    new_new_n44978__, new_new_n44979__, new_new_n44980__, new_new_n44981__,
    new_new_n44982__, new_new_n44983__, new_new_n44984__, new_new_n44985__,
    new_new_n44986__, new_new_n44987__, new_new_n44988__, new_new_n44989__,
    new_new_n44990__, new_new_n44991__, new_new_n44992__, new_new_n44993__,
    new_new_n44994__, new_new_n44995__, new_new_n44996__, new_new_n44997__,
    new_new_n44999__, new_new_n45000__, new_new_n45001__, new_new_n45002__,
    new_new_n45003__, new_new_n45004__, new_new_n45005__, new_new_n45006__,
    new_new_n45007__, new_new_n45008__, new_new_n45009__, new_new_n45010__,
    new_new_n45011__, new_new_n45012__, new_new_n45013__, new_new_n45014__,
    new_new_n45015__, new_new_n45016__, new_new_n45017__, new_new_n45018__,
    new_new_n45019__, new_new_n45020__, new_new_n45021__, new_new_n45022__,
    new_new_n45023__, new_new_n45024__, new_new_n45025__, new_new_n45026__,
    new_new_n45027__, new_new_n45028__, new_new_n45030__, new_new_n45031__,
    new_new_n45032__, new_new_n45033__, new_new_n45034__, new_new_n45035__,
    new_new_n45036__, new_new_n45037__, new_new_n45038__, new_new_n45039__,
    new_new_n45040__, new_new_n45041__, new_new_n45042__, new_new_n45043__,
    new_new_n45044__, new_new_n45045__, new_new_n45046__, new_new_n45047__,
    new_new_n45048__, new_new_n45049__, new_new_n45050__, new_new_n45051__,
    new_new_n45052__, new_new_n45053__, new_new_n45054__, new_new_n45055__,
    new_new_n45056__, new_new_n45057__, new_new_n45058__, new_new_n45059__,
    new_new_n45061__, new_new_n45062__, new_new_n45063__, new_new_n45064__,
    new_new_n45065__, new_new_n45066__, new_new_n45067__, new_new_n45068__,
    new_new_n45069__, new_new_n45070__, new_new_n45071__, new_new_n45072__,
    new_new_n45073__, new_new_n45074__, new_new_n45075__, new_new_n45076__,
    new_new_n45077__, new_new_n45078__, new_new_n45079__, new_new_n45080__,
    new_new_n45081__, new_new_n45082__, new_new_n45083__, new_new_n45084__,
    new_new_n45085__, new_new_n45086__, new_new_n45087__, new_new_n45088__,
    new_new_n45089__, new_new_n45090__, new_new_n45092__, new_new_n45093__,
    new_new_n45094__, new_new_n45095__, new_new_n45096__, new_new_n45097__,
    new_new_n45098__, new_new_n45099__, new_new_n45100__, new_new_n45101__,
    new_new_n45102__, new_new_n45103__, new_new_n45104__, new_new_n45105__,
    new_new_n45106__, new_new_n45107__, new_new_n45108__, new_new_n45109__,
    new_new_n45110__, new_new_n45111__, new_new_n45112__, new_new_n45113__,
    new_new_n45114__, new_new_n45115__, new_new_n45116__, new_new_n45117__,
    new_new_n45118__, new_new_n45119__, new_new_n45120__, new_new_n45121__,
    new_new_n45123__, new_new_n45124__, new_new_n45125__, new_new_n45126__,
    new_new_n45127__, new_new_n45128__, new_new_n45129__, new_new_n45130__,
    new_new_n45131__, new_new_n45132__, new_new_n45133__, new_new_n45134__,
    new_new_n45135__, new_new_n45136__, new_new_n45137__, new_new_n45138__,
    new_new_n45139__, new_new_n45140__, new_new_n45141__, new_new_n45142__,
    new_new_n45143__, new_new_n45144__, new_new_n45145__, new_new_n45146__,
    new_new_n45147__, new_new_n45148__, new_new_n45149__, new_new_n45150__,
    new_new_n45151__, new_new_n45152__, new_new_n45154__, new_new_n45155__,
    new_new_n45156__, new_new_n45157__, new_new_n45158__, new_new_n45159__,
    new_new_n45160__, new_new_n45161__, new_new_n45162__, new_new_n45163__,
    new_new_n45164__, new_new_n45165__, new_new_n45166__, new_new_n45167__,
    new_new_n45168__, new_new_n45169__, new_new_n45170__, new_new_n45171__,
    new_new_n45172__, new_new_n45173__, new_new_n45174__, new_new_n45175__,
    new_new_n45176__, new_new_n45177__, new_new_n45178__, new_new_n45179__,
    new_new_n45180__, new_new_n45181__, new_new_n45182__, new_new_n45183__,
    new_new_n45185__, new_new_n45186__, new_new_n45187__, new_new_n45188__,
    new_new_n45189__, new_new_n45190__, new_new_n45191__, new_new_n45192__,
    new_new_n45193__, new_new_n45194__, new_new_n45195__, new_new_n45196__,
    new_new_n45197__, new_new_n45198__, new_new_n45199__, new_new_n45200__,
    new_new_n45201__, new_new_n45202__, new_new_n45203__, new_new_n45204__,
    new_new_n45205__, new_new_n45206__, new_new_n45207__, new_new_n45208__,
    new_new_n45209__, new_new_n45210__, new_new_n45211__, new_new_n45212__,
    new_new_n45213__, new_new_n45214__, new_new_n45216__, new_new_n45217__,
    new_new_n45218__, new_new_n45219__, new_new_n45220__, new_new_n45221__,
    new_new_n45222__, new_new_n45223__, new_new_n45224__, new_new_n45225__,
    new_new_n45226__, new_new_n45227__, new_new_n45228__, new_new_n45229__,
    new_new_n45230__, new_new_n45231__, new_new_n45232__, new_new_n45233__,
    new_new_n45234__, new_new_n45235__, new_new_n45236__, new_new_n45237__,
    new_new_n45238__, new_new_n45239__, new_new_n45240__, new_new_n45241__,
    new_new_n45242__, new_new_n45243__, new_new_n45244__, new_new_n45245__,
    new_new_n45247__, new_new_n45248__, new_new_n45249__, new_new_n45250__,
    new_new_n45251__, new_new_n45252__, new_new_n45253__, new_new_n45254__,
    new_new_n45255__, new_new_n45256__, new_new_n45257__, new_new_n45258__,
    new_new_n45259__, new_new_n45260__, new_new_n45261__, new_new_n45262__,
    new_new_n45263__, new_new_n45264__, new_new_n45265__, new_new_n45266__,
    new_new_n45267__, new_new_n45268__, new_new_n45269__, new_new_n45270__,
    new_new_n45271__, new_new_n45272__, new_new_n45273__, new_new_n45274__,
    new_new_n45275__, new_new_n45276__, new_new_n45278__, new_new_n45279__,
    new_new_n45280__, new_new_n45281__, new_new_n45282__, new_new_n45283__,
    new_new_n45284__, new_new_n45285__, new_new_n45286__, new_new_n45287__,
    new_new_n45288__, new_new_n45289__, new_new_n45290__, new_new_n45291__,
    new_new_n45292__, new_new_n45293__, new_new_n45294__, new_new_n45295__,
    new_new_n45296__, new_new_n45297__, new_new_n45298__, new_new_n45299__,
    new_new_n45300__, new_new_n45301__, new_new_n45302__, new_new_n45303__,
    new_new_n45304__, new_new_n45305__, new_new_n45306__, new_new_n45307__,
    new_new_n45309__, new_new_n45310__, new_new_n45311__, new_new_n45312__,
    new_new_n45313__, new_new_n45314__, new_new_n45315__, new_new_n45316__,
    new_new_n45317__, new_new_n45318__, new_new_n45319__, new_new_n45320__,
    new_new_n45321__, new_new_n45322__, new_new_n45323__, new_new_n45324__,
    new_new_n45325__, new_new_n45326__, new_new_n45327__, new_new_n45328__,
    new_new_n45329__, new_new_n45330__, new_new_n45331__, new_new_n45332__,
    new_new_n45333__, new_new_n45334__, new_new_n45335__, new_new_n45336__,
    new_new_n45337__, new_new_n45338__, new_new_n45340__, new_new_n45341__,
    new_new_n45342__, new_new_n45343__, new_new_n45344__, new_new_n45345__,
    new_new_n45346__, new_new_n45347__, new_new_n45348__, new_new_n45349__,
    new_new_n45350__, new_new_n45351__, new_new_n45352__, new_new_n45353__,
    new_new_n45354__, new_new_n45355__, new_new_n45356__, new_new_n45357__,
    new_new_n45358__, new_new_n45359__, new_new_n45360__, new_new_n45361__,
    new_new_n45362__, new_new_n45363__, new_new_n45364__, new_new_n45365__,
    new_new_n45366__, new_new_n45367__, new_new_n45368__, new_new_n45369__,
    new_new_n45371__, new_new_n45372__, new_new_n45373__, new_new_n45374__,
    new_new_n45375__, new_new_n45376__, new_new_n45377__, new_new_n45378__,
    new_new_n45379__, new_new_n45380__, new_new_n45381__, new_new_n45382__,
    new_new_n45383__, new_new_n45384__, new_new_n45385__, new_new_n45386__,
    new_new_n45387__, new_new_n45388__, new_new_n45389__, new_new_n45390__,
    new_new_n45391__, new_new_n45392__, new_new_n45393__, new_new_n45394__,
    new_new_n45395__, new_new_n45396__, new_new_n45397__, new_new_n45398__,
    new_new_n45399__, new_new_n45400__, new_new_n45402__, new_new_n45403__,
    new_new_n45404__, new_new_n45405__, new_new_n45406__, new_new_n45407__,
    new_new_n45408__, new_new_n45409__, new_new_n45410__, new_new_n45411__,
    new_new_n45412__, new_new_n45413__, new_new_n45414__, new_new_n45415__,
    new_new_n45416__, new_new_n45417__, new_new_n45418__, new_new_n45419__,
    new_new_n45420__, new_new_n45421__, new_new_n45422__, new_new_n45423__,
    new_new_n45424__, new_new_n45425__, new_new_n45426__, new_new_n45427__,
    new_new_n45428__, new_new_n45429__, new_new_n45430__, new_new_n45431__,
    new_new_n45433__, new_new_n45434__, new_new_n45435__, new_new_n45436__,
    new_new_n45437__, new_new_n45438__, new_new_n45439__, new_new_n45440__,
    new_new_n45441__, new_new_n45442__, new_new_n45443__, new_new_n45444__,
    new_new_n45445__, new_new_n45446__, new_new_n45447__, new_new_n45448__,
    new_new_n45449__, new_new_n45450__, new_new_n45451__, new_new_n45452__,
    new_new_n45453__, new_new_n45454__, new_new_n45455__, new_new_n45456__,
    new_new_n45457__, new_new_n45458__, new_new_n45459__, new_new_n45460__,
    new_new_n45461__, new_new_n45462__, new_new_n45464__, new_new_n45465__,
    new_new_n45466__, new_new_n45467__, new_new_n45468__, new_new_n45469__,
    new_new_n45470__, new_new_n45471__, new_new_n45472__, new_new_n45473__,
    new_new_n45474__, new_new_n45475__, new_new_n45476__, new_new_n45477__,
    new_new_n45478__, new_new_n45479__, new_new_n45480__, new_new_n45481__,
    new_new_n45482__, new_new_n45483__, new_new_n45484__, new_new_n45485__,
    new_new_n45486__, new_new_n45487__, new_new_n45488__, new_new_n45489__,
    new_new_n45490__, new_new_n45491__, new_new_n45492__, new_new_n45493__,
    new_new_n45495__, new_new_n45496__, new_new_n45497__, new_new_n45498__,
    new_new_n45499__, new_new_n45500__, new_new_n45501__, new_new_n45502__,
    new_new_n45503__, new_new_n45504__, new_new_n45505__, new_new_n45506__,
    new_new_n45507__, new_new_n45508__, new_new_n45509__, new_new_n45510__,
    new_new_n45511__, new_new_n45512__, new_new_n45513__, new_new_n45514__,
    new_new_n45515__, new_new_n45516__, new_new_n45517__, new_new_n45518__,
    new_new_n45519__, new_new_n45520__, new_new_n45521__, new_new_n45522__,
    new_new_n45523__, new_new_n45524__, new_new_n45526__, new_new_n45527__,
    new_new_n45528__, new_new_n45529__, new_new_n45530__, new_new_n45531__,
    new_new_n45532__, new_new_n45533__, new_new_n45534__, new_new_n45535__,
    new_new_n45536__, new_new_n45537__, new_new_n45538__, new_new_n45539__,
    new_new_n45540__, new_new_n45541__, new_new_n45542__, new_new_n45543__,
    new_new_n45544__, new_new_n45545__, new_new_n45546__, new_new_n45547__,
    new_new_n45548__, new_new_n45549__, new_new_n45550__, new_new_n45551__,
    new_new_n45552__, new_new_n45553__, new_new_n45554__, new_new_n45555__,
    new_new_n45557__, new_new_n45558__, new_new_n45559__, new_new_n45560__,
    new_new_n45561__, new_new_n45562__, new_new_n45563__, new_new_n45564__,
    new_new_n45565__, new_new_n45566__, new_new_n45567__, new_new_n45568__,
    new_new_n45569__, new_new_n45570__, new_new_n45571__, new_new_n45572__,
    new_new_n45573__, new_new_n45574__, new_new_n45575__, new_new_n45576__,
    new_new_n45577__, new_new_n45578__, new_new_n45579__, new_new_n45580__,
    new_new_n45581__, new_new_n45582__, new_new_n45583__, new_new_n45584__,
    new_new_n45585__, new_new_n45586__, new_new_n45588__, new_new_n45589__,
    new_new_n45590__, new_new_n45591__, new_new_n45592__, new_new_n45593__,
    new_new_n45594__, new_new_n45595__, new_new_n45596__, new_new_n45597__,
    new_new_n45598__, new_new_n45599__, new_new_n45600__, new_new_n45601__,
    new_new_n45602__, new_new_n45603__, new_new_n45604__, new_new_n45605__,
    new_new_n45606__, new_new_n45607__, new_new_n45608__, new_new_n45609__,
    new_new_n45610__, new_new_n45611__, new_new_n45612__, new_new_n45613__,
    new_new_n45614__, new_new_n45615__, new_new_n45616__, new_new_n45617__,
    new_new_n45619__, new_new_n45620__, new_new_n45621__, new_new_n45622__,
    new_new_n45623__, new_new_n45624__, new_new_n45625__, new_new_n45626__,
    new_new_n45627__, new_new_n45628__, new_new_n45629__, new_new_n45630__,
    new_new_n45631__, new_new_n45632__, new_new_n45633__, new_new_n45634__,
    new_new_n45635__, new_new_n45636__, new_new_n45637__, new_new_n45638__,
    new_new_n45639__, new_new_n45640__, new_new_n45641__, new_new_n45642__,
    new_new_n45643__, new_new_n45644__, new_new_n45645__, new_new_n45646__,
    new_new_n45647__, new_new_n45648__, new_new_n45650__, new_new_n45651__,
    new_new_n45652__, new_new_n45653__, new_new_n45654__, new_new_n45655__,
    new_new_n45656__, new_new_n45657__, new_new_n45658__, new_new_n45659__,
    new_new_n45660__, new_new_n45661__, new_new_n45662__, new_new_n45663__,
    new_new_n45664__, new_new_n45665__, new_new_n45666__, new_new_n45667__,
    new_new_n45668__, new_new_n45669__, new_new_n45670__, new_new_n45671__,
    new_new_n45672__, new_new_n45673__, new_new_n45674__, new_new_n45675__,
    new_new_n45676__, new_new_n45677__, new_new_n45678__, new_new_n45679__,
    new_new_n45681__, new_new_n45682__, new_new_n45683__, new_new_n45684__,
    new_new_n45685__, new_new_n45686__, new_new_n45687__, new_new_n45688__,
    new_new_n45689__, new_new_n45690__, new_new_n45691__, new_new_n45692__,
    new_new_n45693__, new_new_n45694__, new_new_n45695__, new_new_n45696__,
    new_new_n45697__, new_new_n45698__, new_new_n45699__, new_new_n45700__,
    new_new_n45701__, new_new_n45702__, new_new_n45703__, new_new_n45704__,
    new_new_n45705__, new_new_n45706__, new_new_n45707__, new_new_n45708__,
    new_new_n45709__, new_new_n45710__, new_new_n45712__, new_new_n45713__,
    new_new_n45714__, new_new_n45715__, new_new_n45716__, new_new_n45717__,
    new_new_n45718__, new_new_n45719__, new_new_n45720__, new_new_n45721__,
    new_new_n45722__, new_new_n45723__, new_new_n45724__, new_new_n45725__,
    new_new_n45726__, new_new_n45727__, new_new_n45728__, new_new_n45729__,
    new_new_n45730__, new_new_n45731__, new_new_n45732__, new_new_n45733__,
    new_new_n45734__, new_new_n45735__, new_new_n45736__, new_new_n45737__,
    new_new_n45738__, new_new_n45739__, new_new_n45740__, new_new_n45741__,
    new_new_n45743__, new_new_n45744__, new_new_n45745__, new_new_n45746__,
    new_new_n45747__, new_new_n45748__, new_new_n45749__, new_new_n45750__,
    new_new_n45751__, new_new_n45752__, new_new_n45753__, new_new_n45754__,
    new_new_n45755__, new_new_n45756__, new_new_n45757__, new_new_n45758__,
    new_new_n45759__, new_new_n45760__, new_new_n45761__, new_new_n45762__,
    new_new_n45763__, new_new_n45764__, new_new_n45765__, new_new_n45766__,
    new_new_n45767__, new_new_n45768__, new_new_n45769__, new_new_n45770__,
    new_new_n45771__, new_new_n45772__, new_new_n45774__, new_new_n45775__,
    new_new_n45776__, new_new_n45777__, new_new_n45778__, new_new_n45779__,
    new_new_n45780__, new_new_n45781__, new_new_n45782__, new_new_n45783__,
    new_new_n45784__, new_new_n45785__, new_new_n45786__, new_new_n45787__,
    new_new_n45788__, new_new_n45789__, new_new_n45790__, new_new_n45791__,
    new_new_n45792__, new_new_n45793__, new_new_n45794__, new_new_n45795__,
    new_new_n45796__, new_new_n45797__, new_new_n45798__, new_new_n45799__,
    new_new_n45800__, new_new_n45801__, new_new_n45802__, new_new_n45803__,
    new_new_n45805__, new_new_n45806__, new_new_n45807__, new_new_n45808__,
    new_new_n45809__, new_new_n45810__, new_new_n45811__, new_new_n45812__,
    new_new_n45813__, new_new_n45814__, new_new_n45815__, new_new_n45816__,
    new_new_n45817__, new_new_n45818__, new_new_n45819__, new_new_n45820__,
    new_new_n45821__, new_new_n45822__, new_new_n45823__, new_new_n45824__,
    new_new_n45825__, new_new_n45826__, new_new_n45827__, new_new_n45828__,
    new_new_n45829__, new_new_n45830__, new_new_n45831__, new_new_n45832__,
    new_new_n45833__, new_new_n45834__, new_new_n45836__, new_new_n45837__,
    new_new_n45839__, new_new_n45840__, new_new_n45841__, new_new_n45842__,
    new_new_n45843__, new_new_n45845__, new_new_n45846__, new_new_n45847__,
    new_new_n45848__, new_new_n45849__, new_new_n45850__, new_new_n45851__,
    new_new_n45852__, new_new_n45854__, new_new_n45855__, new_new_n45856__,
    new_new_n45858__, new_new_n45859__, new_new_n45860__, new_new_n45862__,
    new_new_n45863__, new_new_n45864__, new_new_n45866__, new_new_n45867__,
    new_new_n45868__, new_new_n45870__, new_new_n45871__, new_new_n45872__,
    new_new_n45874__, new_new_n45875__, new_new_n45876__, new_new_n45878__,
    new_new_n45879__, new_new_n45880__, new_new_n45882__, new_new_n45883__,
    new_new_n45884__, new_new_n45886__, new_new_n45887__, new_new_n45888__,
    new_new_n45890__, new_new_n45891__, new_new_n45892__, new_new_n45894__,
    new_new_n45895__, new_new_n45896__, new_new_n45898__, new_new_n45899__,
    new_new_n45900__, new_new_n45902__, new_new_n45903__, new_new_n45904__,
    new_new_n45906__, new_new_n45907__, new_new_n45908__, new_new_n45910__,
    new_new_n45911__, new_new_n45912__, new_new_n45914__, new_new_n45915__,
    new_new_n45916__, new_new_n45918__, new_new_n45919__, new_new_n45920__,
    new_new_n45922__, new_new_n45923__, new_new_n45924__, new_new_n45926__,
    new_new_n45927__, new_new_n45928__, new_new_n45930__, new_new_n45931__,
    new_new_n45932__, new_new_n45934__, new_new_n45935__, new_new_n45936__,
    new_new_n45938__, new_new_n45939__, new_new_n45940__, new_new_n45942__,
    new_new_n45943__, new_new_n45944__, new_new_n45946__, new_new_n45947__,
    new_new_n45948__, new_new_n45950__, new_new_n45951__, new_new_n45952__,
    new_new_n45954__, new_new_n45955__, new_new_n45956__, new_new_n45958__,
    new_new_n45959__, new_new_n45960__, new_new_n45962__, new_new_n45963__,
    new_new_n45964__, new_new_n45966__, new_new_n45967__, new_new_n45968__,
    new_new_n45970__, new_new_n45971__, new_new_n45972__, new_new_n45974__,
    new_new_n45975__, new_new_n45976__, new_new_n45978__, new_new_n45979__,
    new_new_n45980__, new_new_n45982__, new_new_n45983__, new_new_n45984__,
    new_new_n45986__, new_new_n45987__, new_new_n45988__, new_new_n45989__,
    new_new_n45990__, new_new_n45991__, new_new_n45992__, new_new_n45993__,
    new_new_n45995__, new_new_n45996__, new_new_n45997__, new_new_n45999__,
    new_new_n46000__, new_new_n46001__, new_new_n46003__, new_new_n46004__,
    new_new_n46005__, new_new_n46007__, new_new_n46008__, new_new_n46009__,
    new_new_n46011__, new_new_n46012__, new_new_n46013__, new_new_n46015__,
    new_new_n46016__, new_new_n46017__, new_new_n46019__, new_new_n46020__,
    new_new_n46021__, new_new_n46023__, new_new_n46024__, new_new_n46025__,
    new_new_n46027__, new_new_n46028__, new_new_n46029__, new_new_n46031__,
    new_new_n46032__, new_new_n46033__, new_new_n46035__, new_new_n46036__,
    new_new_n46037__, new_new_n46039__, new_new_n46040__, new_new_n46041__,
    new_new_n46043__, new_new_n46044__, new_new_n46045__, new_new_n46047__,
    new_new_n46048__, new_new_n46049__, new_new_n46051__, new_new_n46052__,
    new_new_n46053__, new_new_n46055__, new_new_n46056__, new_new_n46057__,
    new_new_n46059__, new_new_n46060__, new_new_n46061__, new_new_n46063__,
    new_new_n46064__, new_new_n46065__, new_new_n46067__, new_new_n46068__,
    new_new_n46069__, new_new_n46071__, new_new_n46072__, new_new_n46073__,
    new_new_n46075__, new_new_n46076__, new_new_n46077__, new_new_n46079__,
    new_new_n46080__, new_new_n46081__, new_new_n46083__, new_new_n46084__,
    new_new_n46085__, new_new_n46087__, new_new_n46088__, new_new_n46089__,
    new_new_n46091__, new_new_n46092__, new_new_n46093__, new_new_n46095__,
    new_new_n46096__, new_new_n46097__, new_new_n46099__, new_new_n46100__,
    new_new_n46101__, new_new_n46103__, new_new_n46104__, new_new_n46105__,
    new_new_n46107__, new_new_n46108__, new_new_n46109__, new_new_n46111__,
    new_new_n46112__, new_new_n46113__, new_new_n46115__, new_new_n46116__,
    new_new_n46117__, new_new_n46119__, new_new_n46120__, new_new_n46121__,
    new_new_n46123__, new_new_n46124__, new_new_n46125__, new_new_n46127__,
    new_new_n46128__, new_new_n46129__, new_new_n46130__, new_new_n46131__,
    new_new_n46132__, new_new_n46133__, new_new_n46134__, new_new_n46136__,
    new_new_n46137__, new_new_n46138__, new_new_n46140__, new_new_n46141__,
    new_new_n46142__, new_new_n46144__, new_new_n46145__, new_new_n46146__,
    new_new_n46148__, new_new_n46149__, new_new_n46150__, new_new_n46152__,
    new_new_n46153__, new_new_n46154__, new_new_n46156__, new_new_n46157__,
    new_new_n46158__, new_new_n46160__, new_new_n46161__, new_new_n46162__,
    new_new_n46164__, new_new_n46165__, new_new_n46166__, new_new_n46168__,
    new_new_n46169__, new_new_n46170__, new_new_n46172__, new_new_n46173__,
    new_new_n46174__, new_new_n46176__, new_new_n46177__, new_new_n46178__,
    new_new_n46180__, new_new_n46181__, new_new_n46182__, new_new_n46184__,
    new_new_n46185__, new_new_n46186__, new_new_n46188__, new_new_n46189__,
    new_new_n46190__, new_new_n46192__, new_new_n46193__, new_new_n46194__,
    new_new_n46196__, new_new_n46197__, new_new_n46198__, new_new_n46200__,
    new_new_n46201__, new_new_n46202__, new_new_n46204__, new_new_n46205__,
    new_new_n46206__, new_new_n46208__, new_new_n46209__, new_new_n46210__,
    new_new_n46212__, new_new_n46213__, new_new_n46214__, new_new_n46216__,
    new_new_n46217__, new_new_n46218__, new_new_n46220__, new_new_n46221__,
    new_new_n46222__, new_new_n46224__, new_new_n46225__, new_new_n46226__,
    new_new_n46228__, new_new_n46229__, new_new_n46230__, new_new_n46232__,
    new_new_n46233__, new_new_n46234__, new_new_n46236__, new_new_n46237__,
    new_new_n46238__, new_new_n46240__, new_new_n46241__, new_new_n46242__,
    new_new_n46244__, new_new_n46245__, new_new_n46246__, new_new_n46248__,
    new_new_n46249__, new_new_n46250__, new_new_n46252__, new_new_n46253__,
    new_new_n46254__, new_new_n46256__, new_new_n46257__, new_new_n46258__,
    new_new_n46260__, new_new_n46261__, new_new_n46262__, new_new_n46264__,
    new_new_n46265__, new_new_n46266__, new_new_n46268__, new_new_n46269__,
    new_new_n46270__, new_new_n46271__, new_new_n46272__, new_new_n46273__,
    new_new_n46274__, new_new_n46275__, new_new_n46277__, new_new_n46278__,
    new_new_n46279__, new_new_n46281__, new_new_n46282__, new_new_n46283__,
    new_new_n46285__, new_new_n46286__, new_new_n46287__, new_new_n46289__,
    new_new_n46290__, new_new_n46291__, new_new_n46293__, new_new_n46294__,
    new_new_n46295__, new_new_n46297__, new_new_n46298__, new_new_n46299__,
    new_new_n46301__, new_new_n46302__, new_new_n46303__, new_new_n46305__,
    new_new_n46306__, new_new_n46307__, new_new_n46309__, new_new_n46310__,
    new_new_n46311__, new_new_n46313__, new_new_n46314__, new_new_n46315__,
    new_new_n46317__, new_new_n46318__, new_new_n46319__, new_new_n46321__,
    new_new_n46322__, new_new_n46323__, new_new_n46325__, new_new_n46326__,
    new_new_n46327__, new_new_n46329__, new_new_n46330__, new_new_n46331__,
    new_new_n46333__, new_new_n46334__, new_new_n46335__, new_new_n46337__,
    new_new_n46338__, new_new_n46339__, new_new_n46341__, new_new_n46342__,
    new_new_n46343__, new_new_n46345__, new_new_n46346__, new_new_n46347__,
    new_new_n46349__, new_new_n46350__, new_new_n46351__, new_new_n46353__,
    new_new_n46354__, new_new_n46355__, new_new_n46357__, new_new_n46358__,
    new_new_n46359__, new_new_n46361__, new_new_n46362__, new_new_n46363__,
    new_new_n46365__, new_new_n46366__, new_new_n46367__, new_new_n46369__,
    new_new_n46370__, new_new_n46371__, new_new_n46373__, new_new_n46374__,
    new_new_n46375__, new_new_n46377__, new_new_n46378__, new_new_n46379__,
    new_new_n46381__, new_new_n46382__, new_new_n46383__, new_new_n46385__,
    new_new_n46386__, new_new_n46387__, new_new_n46389__, new_new_n46390__,
    new_new_n46391__, new_new_n46393__, new_new_n46394__, new_new_n46395__,
    new_new_n46397__, new_new_n46398__, new_new_n46399__, new_new_n46401__,
    new_new_n46402__, new_new_n46403__, new_new_n46405__, new_new_n46406__,
    new_new_n46407__, new_new_n46409__, new_new_n46410__, new_new_n46411__,
    new_new_n46412__, new_new_n46413__, new_new_n46414__, new_new_n46415__,
    new_new_n46416__, new_new_n46418__, new_new_n46419__, new_new_n46420__,
    new_new_n46422__, new_new_n46423__, new_new_n46424__, new_new_n46426__,
    new_new_n46427__, new_new_n46428__, new_new_n46430__, new_new_n46431__,
    new_new_n46432__, new_new_n46434__, new_new_n46435__, new_new_n46436__,
    new_new_n46438__, new_new_n46439__, new_new_n46440__, new_new_n46442__,
    new_new_n46443__, new_new_n46444__, new_new_n46446__, new_new_n46447__,
    new_new_n46448__, new_new_n46450__, new_new_n46451__, new_new_n46452__,
    new_new_n46454__, new_new_n46455__, new_new_n46456__, new_new_n46458__,
    new_new_n46459__, new_new_n46460__, new_new_n46462__, new_new_n46463__,
    new_new_n46464__, new_new_n46466__, new_new_n46467__, new_new_n46468__,
    new_new_n46470__, new_new_n46471__, new_new_n46472__, new_new_n46474__,
    new_new_n46475__, new_new_n46476__, new_new_n46478__, new_new_n46479__,
    new_new_n46480__, new_new_n46482__, new_new_n46483__, new_new_n46484__,
    new_new_n46486__, new_new_n46487__, new_new_n46488__, new_new_n46490__,
    new_new_n46491__, new_new_n46492__, new_new_n46494__, new_new_n46495__,
    new_new_n46496__, new_new_n46498__, new_new_n46499__, new_new_n46500__,
    new_new_n46502__, new_new_n46503__, new_new_n46504__, new_new_n46506__,
    new_new_n46507__, new_new_n46508__, new_new_n46510__, new_new_n46511__,
    new_new_n46512__, new_new_n46514__, new_new_n46515__, new_new_n46516__,
    new_new_n46518__, new_new_n46519__, new_new_n46520__, new_new_n46522__,
    new_new_n46523__, new_new_n46524__, new_new_n46526__, new_new_n46527__,
    new_new_n46528__, new_new_n46530__, new_new_n46531__, new_new_n46532__,
    new_new_n46534__, new_new_n46535__, new_new_n46536__, new_new_n46538__,
    new_new_n46539__, new_new_n46540__, new_new_n46542__, new_new_n46543__,
    new_new_n46544__, new_new_n46546__, new_new_n46547__, new_new_n46548__,
    new_new_n46550__, new_new_n46551__, new_new_n46552__, new_new_n46553__,
    new_new_n46554__, new_new_n46555__, new_new_n46556__, new_new_n46557__,
    new_new_n46559__, new_new_n46560__, new_new_n46561__, new_new_n46563__,
    new_new_n46564__, new_new_n46565__, new_new_n46567__, new_new_n46568__,
    new_new_n46569__, new_new_n46571__, new_new_n46572__, new_new_n46573__,
    new_new_n46575__, new_new_n46576__, new_new_n46577__, new_new_n46579__,
    new_new_n46580__, new_new_n46581__, new_new_n46583__, new_new_n46584__,
    new_new_n46585__, new_new_n46587__, new_new_n46588__, new_new_n46589__,
    new_new_n46591__, new_new_n46592__, new_new_n46593__, new_new_n46595__,
    new_new_n46596__, new_new_n46597__, new_new_n46599__, new_new_n46600__,
    new_new_n46601__, new_new_n46603__, new_new_n46604__, new_new_n46605__,
    new_new_n46607__, new_new_n46608__, new_new_n46609__, new_new_n46611__,
    new_new_n46612__, new_new_n46613__, new_new_n46615__, new_new_n46616__,
    new_new_n46617__, new_new_n46619__, new_new_n46620__, new_new_n46621__,
    new_new_n46623__, new_new_n46624__, new_new_n46625__, new_new_n46627__,
    new_new_n46628__, new_new_n46629__, new_new_n46631__, new_new_n46632__,
    new_new_n46633__, new_new_n46635__, new_new_n46636__, new_new_n46637__,
    new_new_n46639__, new_new_n46640__, new_new_n46641__, new_new_n46643__,
    new_new_n46644__, new_new_n46645__, new_new_n46647__, new_new_n46648__,
    new_new_n46649__, new_new_n46651__, new_new_n46652__, new_new_n46653__,
    new_new_n46655__, new_new_n46656__, new_new_n46657__, new_new_n46659__,
    new_new_n46660__, new_new_n46661__, new_new_n46663__, new_new_n46664__,
    new_new_n46665__, new_new_n46667__, new_new_n46668__, new_new_n46669__,
    new_new_n46671__, new_new_n46672__, new_new_n46673__, new_new_n46675__,
    new_new_n46676__, new_new_n46677__, new_new_n46679__, new_new_n46680__,
    new_new_n46681__, new_new_n46683__, new_new_n46684__, new_new_n46685__,
    new_new_n46687__, new_new_n46688__, new_new_n46689__, new_new_n46691__,
    new_new_n46692__, new_new_n46693__, new_new_n46694__, new_new_n46695__,
    new_new_n46696__, new_new_n46697__, new_new_n46698__, new_new_n46700__,
    new_new_n46701__, new_new_n46702__, new_new_n46704__, new_new_n46705__,
    new_new_n46706__, new_new_n46708__, new_new_n46709__, new_new_n46710__,
    new_new_n46712__, new_new_n46713__, new_new_n46714__, new_new_n46716__,
    new_new_n46717__, new_new_n46718__, new_new_n46720__, new_new_n46721__,
    new_new_n46722__, new_new_n46724__, new_new_n46725__, new_new_n46726__,
    new_new_n46728__, new_new_n46729__, new_new_n46730__, new_new_n46732__,
    new_new_n46733__, new_new_n46734__, new_new_n46736__, new_new_n46737__,
    new_new_n46738__, new_new_n46740__, new_new_n46741__, new_new_n46742__,
    new_new_n46744__, new_new_n46745__, new_new_n46746__, new_new_n46748__,
    new_new_n46749__, new_new_n46750__, new_new_n46752__, new_new_n46753__,
    new_new_n46754__, new_new_n46756__, new_new_n46757__, new_new_n46758__,
    new_new_n46760__, new_new_n46761__, new_new_n46762__, new_new_n46764__,
    new_new_n46765__, new_new_n46766__, new_new_n46768__, new_new_n46769__,
    new_new_n46770__, new_new_n46772__, new_new_n46773__, new_new_n46774__,
    new_new_n46776__, new_new_n46777__, new_new_n46778__, new_new_n46780__,
    new_new_n46781__, new_new_n46782__, new_new_n46784__, new_new_n46785__,
    new_new_n46786__, new_new_n46788__, new_new_n46789__, new_new_n46790__,
    new_new_n46792__, new_new_n46793__, new_new_n46794__, new_new_n46796__,
    new_new_n46797__, new_new_n46798__, new_new_n46800__, new_new_n46801__,
    new_new_n46802__, new_new_n46804__, new_new_n46805__, new_new_n46806__,
    new_new_n46808__, new_new_n46809__, new_new_n46810__, new_new_n46812__,
    new_new_n46813__, new_new_n46814__, new_new_n46816__, new_new_n46817__,
    new_new_n46818__, new_new_n46820__, new_new_n46821__, new_new_n46822__,
    new_new_n46824__, new_new_n46825__, new_new_n46826__, new_new_n46828__,
    new_new_n46829__, new_new_n46830__, new_new_n46832__, new_new_n46833__,
    new_new_n46834__, new_new_n46835__, new_new_n46836__, new_new_n46837__,
    new_new_n46838__, new_new_n46839__, new_new_n46841__, new_new_n46842__,
    new_new_n46843__, new_new_n46845__, new_new_n46846__, new_new_n46847__,
    new_new_n46849__, new_new_n46850__, new_new_n46851__, new_new_n46853__,
    new_new_n46854__, new_new_n46855__, new_new_n46857__, new_new_n46858__,
    new_new_n46859__, new_new_n46861__, new_new_n46862__, new_new_n46863__,
    new_new_n46865__, new_new_n46866__, new_new_n46867__, new_new_n46869__,
    new_new_n46870__, new_new_n46871__, new_new_n46873__, new_new_n46874__,
    new_new_n46875__, new_new_n46877__, new_new_n46878__, new_new_n46879__,
    new_new_n46881__, new_new_n46882__, new_new_n46883__, new_new_n46885__,
    new_new_n46886__, new_new_n46887__, new_new_n46889__, new_new_n46890__,
    new_new_n46891__, new_new_n46893__, new_new_n46894__, new_new_n46895__,
    new_new_n46897__, new_new_n46898__, new_new_n46899__, new_new_n46901__,
    new_new_n46902__, new_new_n46903__, new_new_n46905__, new_new_n46906__,
    new_new_n46907__, new_new_n46909__, new_new_n46910__, new_new_n46911__,
    new_new_n46913__, new_new_n46914__, new_new_n46915__, new_new_n46917__,
    new_new_n46918__, new_new_n46919__, new_new_n46921__, new_new_n46922__,
    new_new_n46923__, new_new_n46925__, new_new_n46926__, new_new_n46927__,
    new_new_n46929__, new_new_n46930__, new_new_n46931__, new_new_n46933__,
    new_new_n46934__, new_new_n46935__, new_new_n46937__, new_new_n46938__,
    new_new_n46939__, new_new_n46941__, new_new_n46942__, new_new_n46943__,
    new_new_n46945__, new_new_n46946__, new_new_n46947__, new_new_n46949__,
    new_new_n46950__, new_new_n46951__, new_new_n46953__, new_new_n46954__,
    new_new_n46955__, new_new_n46957__, new_new_n46958__, new_new_n46959__,
    new_new_n46961__, new_new_n46962__, new_new_n46963__, new_new_n46965__,
    new_new_n46966__, new_new_n46967__, new_new_n46968__, new_new_n46969__,
    new_new_n46970__, new_new_n46971__, new_new_n46972__, new_new_n46974__,
    new_new_n46975__, new_new_n46976__, new_new_n46978__, new_new_n46979__,
    new_new_n46980__, new_new_n46982__, new_new_n46983__, new_new_n46984__,
    new_new_n46986__, new_new_n46987__, new_new_n46988__, new_new_n46990__,
    new_new_n46991__, new_new_n46992__, new_new_n46994__, new_new_n46995__,
    new_new_n46996__, new_new_n46998__, new_new_n46999__, new_new_n47000__,
    new_new_n47002__, new_new_n47003__, new_new_n47004__, new_new_n47006__,
    new_new_n47007__, new_new_n47008__, new_new_n47010__, new_new_n47011__,
    new_new_n47012__, new_new_n47014__, new_new_n47015__, new_new_n47016__,
    new_new_n47018__, new_new_n47019__, new_new_n47020__, new_new_n47022__,
    new_new_n47023__, new_new_n47024__, new_new_n47026__, new_new_n47027__,
    new_new_n47028__, new_new_n47030__, new_new_n47031__, new_new_n47032__,
    new_new_n47034__, new_new_n47035__, new_new_n47036__, new_new_n47038__,
    new_new_n47039__, new_new_n47040__, new_new_n47042__, new_new_n47043__,
    new_new_n47044__, new_new_n47046__, new_new_n47047__, new_new_n47048__,
    new_new_n47050__, new_new_n47051__, new_new_n47052__, new_new_n47054__,
    new_new_n47055__, new_new_n47056__, new_new_n47058__, new_new_n47059__,
    new_new_n47060__, new_new_n47062__, new_new_n47063__, new_new_n47064__,
    new_new_n47066__, new_new_n47067__, new_new_n47068__, new_new_n47070__,
    new_new_n47071__, new_new_n47072__, new_new_n47074__, new_new_n47075__,
    new_new_n47076__, new_new_n47078__, new_new_n47079__, new_new_n47080__,
    new_new_n47082__, new_new_n47083__, new_new_n47084__, new_new_n47086__,
    new_new_n47087__, new_new_n47088__, new_new_n47090__, new_new_n47091__,
    new_new_n47092__, new_new_n47094__, new_new_n47095__, new_new_n47096__,
    new_new_n47098__, new_new_n47099__, new_new_n47100__, new_new_n47101__,
    new_new_n47102__, new_new_n47103__, new_new_n47104__, new_new_n47105__,
    new_new_n47107__, new_new_n47108__, new_new_n47109__, new_new_n47111__,
    new_new_n47112__, new_new_n47113__, new_new_n47115__, new_new_n47116__,
    new_new_n47117__, new_new_n47119__, new_new_n47120__, new_new_n47121__,
    new_new_n47123__, new_new_n47124__, new_new_n47125__, new_new_n47127__,
    new_new_n47128__, new_new_n47129__, new_new_n47131__, new_new_n47132__,
    new_new_n47133__, new_new_n47135__, new_new_n47136__, new_new_n47137__,
    new_new_n47139__, new_new_n47140__, new_new_n47141__, new_new_n47143__,
    new_new_n47144__, new_new_n47145__, new_new_n47147__, new_new_n47148__,
    new_new_n47149__, new_new_n47151__, new_new_n47152__, new_new_n47153__,
    new_new_n47155__, new_new_n47156__, new_new_n47157__, new_new_n47159__,
    new_new_n47160__, new_new_n47161__, new_new_n47163__, new_new_n47164__,
    new_new_n47165__, new_new_n47167__, new_new_n47168__, new_new_n47169__,
    new_new_n47171__, new_new_n47172__, new_new_n47173__, new_new_n47175__,
    new_new_n47176__, new_new_n47177__, new_new_n47179__, new_new_n47180__,
    new_new_n47181__, new_new_n47183__, new_new_n47184__, new_new_n47185__,
    new_new_n47187__, new_new_n47188__, new_new_n47189__, new_new_n47191__,
    new_new_n47192__, new_new_n47193__, new_new_n47195__, new_new_n47196__,
    new_new_n47197__, new_new_n47199__, new_new_n47200__, new_new_n47201__,
    new_new_n47203__, new_new_n47204__, new_new_n47205__, new_new_n47207__,
    new_new_n47208__, new_new_n47209__, new_new_n47211__, new_new_n47212__,
    new_new_n47213__, new_new_n47215__, new_new_n47216__, new_new_n47217__,
    new_new_n47219__, new_new_n47220__, new_new_n47221__, new_new_n47223__,
    new_new_n47224__, new_new_n47225__, new_new_n47227__, new_new_n47228__,
    new_new_n47229__, new_new_n47231__, new_new_n47232__, new_new_n47233__,
    new_new_n47235__, new_new_n47236__, new_new_n47237__, new_new_n47239__,
    new_new_n47240__, new_new_n47241__, new_new_n47243__, new_new_n47244__,
    new_new_n47245__, new_new_n47247__, new_new_n47248__, new_new_n47249__,
    new_new_n47251__, new_new_n47252__, new_new_n47253__, new_new_n47255__,
    new_new_n47256__, new_new_n47257__, new_new_n47259__, new_new_n47260__,
    new_new_n47261__, new_new_n47263__, new_new_n47264__, new_new_n47265__,
    new_new_n47267__, new_new_n47268__, new_new_n47269__, new_new_n47271__,
    new_new_n47272__, new_new_n47273__, new_new_n47275__, new_new_n47276__,
    new_new_n47277__, new_new_n47279__, new_new_n47280__, new_new_n47281__,
    new_new_n47283__, new_new_n47284__, new_new_n47285__, new_new_n47287__,
    new_new_n47288__, new_new_n47289__, new_new_n47291__, new_new_n47292__,
    new_new_n47293__, new_new_n47295__, new_new_n47296__, new_new_n47297__,
    new_new_n47299__, new_new_n47300__, new_new_n47301__, new_new_n47303__,
    new_new_n47304__, new_new_n47305__, new_new_n47307__, new_new_n47308__,
    new_new_n47309__, new_new_n47311__, new_new_n47312__, new_new_n47313__,
    new_new_n47315__, new_new_n47316__, new_new_n47317__, new_new_n47319__,
    new_new_n47320__, new_new_n47321__, new_new_n47323__, new_new_n47324__,
    new_new_n47325__, new_new_n47327__, new_new_n47328__, new_new_n47329__,
    new_new_n47331__, new_new_n47332__, new_new_n47333__, new_new_n47335__,
    new_new_n47336__, new_new_n47337__, new_new_n47339__, new_new_n47340__,
    new_new_n47341__, new_new_n47343__, new_new_n47344__, new_new_n47345__,
    new_new_n47347__, new_new_n47348__, new_new_n47349__, new_new_n47351__,
    new_new_n47352__, new_new_n47353__, new_new_n47355__, new_new_n47356__,
    new_new_n47357__, new_new_n47359__, new_new_n47360__, new_new_n47361__,
    new_new_n47363__, new_new_n47364__, new_new_n47365__, new_new_n47367__,
    new_new_n47368__, new_new_n47369__, new_new_n47371__, new_new_n47372__,
    new_new_n47373__, new_new_n47375__, new_new_n47376__, new_new_n47377__,
    new_new_n47379__, new_new_n47380__, new_new_n47381__, new_new_n47383__,
    new_new_n47384__, new_new_n47385__, new_new_n47387__, new_new_n47388__,
    new_new_n47389__, new_new_n47391__, new_new_n47392__, new_new_n47393__,
    new_new_n47395__, new_new_n47396__, new_new_n47397__, new_new_n47399__,
    new_new_n47400__, new_new_n47401__, new_new_n47403__, new_new_n47404__,
    new_new_n47405__, new_new_n47407__, new_new_n47408__, new_new_n47409__,
    new_new_n47411__, new_new_n47412__, new_new_n47413__, new_new_n47415__,
    new_new_n47416__, new_new_n47417__, new_new_n47419__, new_new_n47420__,
    new_new_n47421__, new_new_n47423__, new_new_n47424__, new_new_n47425__,
    new_new_n47427__, new_new_n47428__, new_new_n47429__, new_new_n47431__,
    new_new_n47432__, new_new_n47433__, new_new_n47435__, new_new_n47436__,
    new_new_n47437__, new_new_n47439__, new_new_n47440__, new_new_n47441__,
    new_new_n47443__, new_new_n47444__, new_new_n47445__, new_new_n47447__,
    new_new_n47448__, new_new_n47449__, new_new_n47451__, new_new_n47452__,
    new_new_n47453__, new_new_n47455__, new_new_n47456__, new_new_n47457__,
    new_new_n47459__, new_new_n47460__, new_new_n47461__, new_new_n47463__,
    new_new_n47464__, new_new_n47465__, new_new_n47467__, new_new_n47468__,
    new_new_n47469__, new_new_n47471__, new_new_n47472__, new_new_n47473__,
    new_new_n47475__, new_new_n47476__, new_new_n47477__, new_new_n47479__,
    new_new_n47480__, new_new_n47481__, new_new_n47483__, new_new_n47484__,
    new_new_n47485__, new_new_n47487__, new_new_n47488__, new_new_n47489__,
    new_new_n47491__, new_new_n47492__, new_new_n47493__, new_new_n47495__,
    new_new_n47496__, new_new_n47497__, new_new_n47499__, new_new_n47500__,
    new_new_n47501__, new_new_n47503__, new_new_n47504__, new_new_n47505__,
    new_new_n47507__, new_new_n47508__, new_new_n47509__, new_new_n47511__,
    new_new_n47512__, new_new_n47513__, new_new_n47515__, new_new_n47516__,
    new_new_n47517__, new_new_n47519__, new_new_n47520__, new_new_n47521__,
    new_new_n47523__, new_new_n47524__, new_new_n47525__, new_new_n47527__,
    new_new_n47528__, new_new_n47529__, new_new_n47531__, new_new_n47532__,
    new_new_n47533__, new_new_n47535__, new_new_n47536__, new_new_n47537__,
    new_new_n47539__, new_new_n47540__, new_new_n47541__, new_new_n47543__,
    new_new_n47544__, new_new_n47545__, new_new_n47547__, new_new_n47548__,
    new_new_n47549__, new_new_n47551__, new_new_n47552__, new_new_n47553__,
    new_new_n47555__, new_new_n47556__, new_new_n47557__, new_new_n47559__,
    new_new_n47560__, new_new_n47561__, new_new_n47563__, new_new_n47564__,
    new_new_n47565__, new_new_n47567__, new_new_n47568__, new_new_n47569__,
    new_new_n47571__, new_new_n47572__, new_new_n47573__, new_new_n47575__,
    new_new_n47576__, new_new_n47577__, new_new_n47579__, new_new_n47580__,
    new_new_n47581__, new_new_n47583__, new_new_n47584__, new_new_n47585__,
    new_new_n47587__, new_new_n47588__, new_new_n47589__, new_new_n47591__,
    new_new_n47592__, new_new_n47593__, new_new_n47595__, new_new_n47596__,
    new_new_n47597__, new_new_n47599__, new_new_n47600__, new_new_n47601__,
    new_new_n47603__, new_new_n47604__, new_new_n47605__, new_new_n47607__,
    new_new_n47608__, new_new_n47609__, new_new_n47611__, new_new_n47612__,
    new_new_n47613__, new_new_n47615__, new_new_n47616__, new_new_n47617__,
    new_new_n47619__, new_new_n47620__, new_new_n47621__, new_new_n47623__,
    new_new_n47624__, new_new_n47625__, new_new_n47627__, new_new_n47628__,
    new_new_n47629__, new_new_n47631__, new_new_n47632__, new_new_n47633__,
    new_new_n47635__, new_new_n47636__, new_new_n47637__, new_new_n47639__,
    new_new_n47640__, new_new_n47641__, new_new_n47643__, new_new_n47644__,
    new_new_n47645__, new_new_n47647__, new_new_n47648__, new_new_n47649__,
    new_new_n47651__, new_new_n47652__, new_new_n47653__, new_new_n47655__,
    new_new_n47656__, new_new_n47657__, new_new_n47659__, new_new_n47660__,
    new_new_n47661__, new_new_n47663__, new_new_n47664__, new_new_n47665__,
    new_new_n47667__, new_new_n47668__, new_new_n47669__, new_new_n47671__,
    new_new_n47672__, new_new_n47673__, new_new_n47675__, new_new_n47676__,
    new_new_n47677__, new_new_n47679__, new_new_n47680__, new_new_n47681__,
    new_new_n47683__, new_new_n47684__, new_new_n47685__, new_new_n47687__,
    new_new_n47688__, new_new_n47689__, new_new_n47691__, new_new_n47692__,
    new_new_n47693__, new_new_n47695__, new_new_n47696__, new_new_n47697__,
    new_new_n47699__, new_new_n47700__, new_new_n47701__, new_new_n47703__,
    new_new_n47704__, new_new_n47705__, new_new_n47707__, new_new_n47708__,
    new_new_n47709__, new_new_n47711__, new_new_n47712__, new_new_n47713__,
    new_new_n47715__, new_new_n47716__, new_new_n47717__, new_new_n47719__,
    new_new_n47720__, new_new_n47721__, new_new_n47723__, new_new_n47724__,
    new_new_n47725__, new_new_n47727__, new_new_n47728__, new_new_n47729__,
    new_new_n47731__, new_new_n47732__, new_new_n47733__, new_new_n47735__,
    new_new_n47736__, new_new_n47737__, new_new_n47739__, new_new_n47740__,
    new_new_n47741__, new_new_n47743__, new_new_n47744__, new_new_n47745__,
    new_new_n47747__, new_new_n47748__, new_new_n47749__, new_new_n47751__,
    new_new_n47752__, new_new_n47753__, new_new_n47755__, new_new_n47756__,
    new_new_n47757__, new_new_n47759__, new_new_n47760__, new_new_n47761__,
    new_new_n47763__, new_new_n47764__, new_new_n47765__, new_new_n47767__,
    new_new_n47768__, new_new_n47769__, new_new_n47771__, new_new_n47772__,
    new_new_n47773__, new_new_n47775__, new_new_n47776__, new_new_n47777__,
    new_new_n47779__, new_new_n47780__, new_new_n47781__, new_new_n47783__,
    new_new_n47784__, new_new_n47785__, new_new_n47787__, new_new_n47788__,
    new_new_n47789__, new_new_n47791__, new_new_n47792__, new_new_n47793__,
    new_new_n47795__, new_new_n47796__, new_new_n47797__, new_new_n47799__,
    new_new_n47800__, new_new_n47801__, new_new_n47803__, new_new_n47804__,
    new_new_n47805__, new_new_n47807__, new_new_n47808__, new_new_n47809__,
    new_new_n47811__, new_new_n47812__, new_new_n47813__, new_new_n47815__,
    new_new_n47816__, new_new_n47817__, new_new_n47819__, new_new_n47820__,
    new_new_n47821__, new_new_n47823__, new_new_n47824__, new_new_n47825__,
    new_new_n47827__, new_new_n47828__, new_new_n47829__, new_new_n47831__,
    new_new_n47832__, new_new_n47833__, new_new_n47835__, new_new_n47836__,
    new_new_n47837__, new_new_n47839__, new_new_n47840__, new_new_n47841__,
    new_new_n47843__, new_new_n47844__, new_new_n47845__, new_new_n47847__,
    new_new_n47848__, new_new_n47849__, new_new_n47851__, new_new_n47852__,
    new_new_n47853__, new_new_n47855__, new_new_n47856__, new_new_n47857__,
    new_new_n47859__, new_new_n47860__, new_new_n47861__, new_new_n47863__,
    new_new_n47864__, new_new_n47865__, new_new_n47867__, new_new_n47868__,
    new_new_n47869__, new_new_n47871__, new_new_n47872__, new_new_n47873__,
    new_new_n47875__, new_new_n47876__, new_new_n47877__, new_new_n47879__,
    new_new_n47880__, new_new_n47881__, new_new_n47883__, new_new_n47884__,
    new_new_n47885__, new_new_n47887__, new_new_n47888__, new_new_n47889__,
    new_new_n47891__, new_new_n47892__, new_new_n47893__, new_new_n47895__,
    new_new_n47896__, new_new_n47897__, new_new_n47899__, new_new_n47900__,
    new_new_n47901__, new_new_n47903__, new_new_n47904__, new_new_n47905__,
    new_new_n47907__, new_new_n47908__, new_new_n47909__, new_new_n47911__,
    new_new_n47912__, new_new_n47913__, new_new_n47915__, new_new_n47916__,
    new_new_n47917__, new_new_n47919__, new_new_n47920__, new_new_n47921__,
    new_new_n47923__, new_new_n47924__, new_new_n47925__, new_new_n47927__,
    new_new_n47928__, new_new_n47929__, new_new_n47931__, new_new_n47932__,
    new_new_n47933__, new_new_n47935__, new_new_n47936__, new_new_n47937__,
    new_new_n47939__, new_new_n47940__, new_new_n47941__, new_new_n47943__,
    new_new_n47944__, new_new_n47945__, new_new_n47947__, new_new_n47948__,
    new_new_n47949__, new_new_n47951__, new_new_n47952__, new_new_n47953__,
    new_new_n47955__, new_new_n47956__, new_new_n47957__, new_new_n47959__,
    new_new_n47960__, new_new_n47961__, new_new_n47963__, new_new_n47964__,
    new_new_n47965__, new_new_n47967__, new_new_n47968__, new_new_n47969__,
    new_new_n47971__, new_new_n47972__, new_new_n47973__, new_new_n47975__,
    new_new_n47976__, new_new_n47977__, new_new_n47979__, new_new_n47980__,
    new_new_n47981__, new_new_n47983__, new_new_n47984__, new_new_n47985__,
    new_new_n47987__, new_new_n47988__, new_new_n47989__, new_new_n47991__,
    new_new_n47992__, new_new_n47993__, new_new_n47995__, new_new_n47996__,
    new_new_n47997__, new_new_n47999__, new_new_n48000__, new_new_n48001__,
    new_new_n48003__, new_new_n48004__, new_new_n48005__, new_new_n48007__,
    new_new_n48008__, new_new_n48009__, new_new_n48011__, new_new_n48012__,
    new_new_n48013__, new_new_n48015__, new_new_n48016__, new_new_n48017__,
    new_new_n48019__, new_new_n48020__, new_new_n48021__, new_new_n48023__,
    new_new_n48024__, new_new_n48025__, new_new_n48027__, new_new_n48028__,
    new_new_n48029__, new_new_n48031__, new_new_n48032__, new_new_n48033__,
    new_new_n48035__, new_new_n48036__, new_new_n48037__, new_new_n48039__,
    new_new_n48040__, new_new_n48041__, new_new_n48043__, new_new_n48044__,
    new_new_n48045__, new_new_n48047__, new_new_n48048__, new_new_n48049__,
    new_new_n48051__, new_new_n48052__, new_new_n48053__, new_new_n48055__,
    new_new_n48056__, new_new_n48057__, new_new_n48059__, new_new_n48060__,
    new_new_n48061__, new_new_n48063__, new_new_n48064__, new_new_n48065__,
    new_new_n48067__, new_new_n48068__, new_new_n48069__, new_new_n48071__,
    new_new_n48072__, new_new_n48073__, new_new_n48075__, new_new_n48076__,
    new_new_n48077__, new_new_n48079__, new_new_n48080__, new_new_n48081__,
    new_new_n48083__, new_new_n48084__, new_new_n48085__, new_new_n48087__,
    new_new_n48088__, new_new_n48089__, new_new_n48091__, new_new_n48092__,
    new_new_n48093__, new_new_n48095__, new_new_n48096__, new_new_n48097__,
    new_new_n48099__, new_new_n48100__, new_new_n48101__, new_new_n48103__,
    new_new_n48104__, new_new_n48105__, new_new_n48107__, new_new_n48108__,
    new_new_n48109__, new_new_n48111__, new_new_n48112__, new_new_n48113__,
    new_new_n48115__, new_new_n48116__, new_new_n48117__, new_new_n48119__,
    new_new_n48120__, new_new_n48121__, new_new_n48123__, new_new_n48124__,
    new_new_n48125__, new_new_n48127__, new_new_n48128__, new_new_n48129__,
    new_new_n48131__, new_new_n48132__, new_new_n48133__, new_new_n48135__,
    new_new_n48136__, new_new_n48137__, new_new_n48139__, new_new_n48140__,
    new_new_n48141__, new_new_n48143__, new_new_n48144__, new_new_n48145__,
    new_new_n48147__, new_new_n48148__, new_new_n48149__, new_new_n48151__,
    new_new_n48152__, new_new_n48153__, new_new_n48155__, new_new_n48156__,
    new_new_n48157__, new_new_n48159__, new_new_n48160__, new_new_n48161__,
    new_new_n48163__, new_new_n48164__, new_new_n48165__, new_new_n48167__,
    new_new_n48168__, new_new_n48169__, new_new_n48171__, new_new_n48172__,
    new_new_n48173__, new_new_n48175__, new_new_n48176__, new_new_n48177__,
    new_new_n48179__, new_new_n48180__, new_new_n48181__, new_new_n48183__,
    new_new_n48184__, new_new_n48185__, new_new_n48187__, new_new_n48188__,
    new_new_n48189__, new_new_n48191__, new_new_n48192__, new_new_n48193__,
    new_new_n48195__, new_new_n48196__, new_new_n48197__, new_new_n48199__,
    new_new_n48200__, new_new_n48201__, new_new_n48203__, new_new_n48204__,
    new_new_n48205__, new_new_n48207__, new_new_n48208__, new_new_n48209__,
    new_new_n48211__, new_new_n48212__, new_new_n48213__, new_new_n48215__,
    new_new_n48216__, new_new_n48217__, new_new_n48219__, new_new_n48220__,
    new_new_n48221__, new_new_n48223__, new_new_n48224__, new_new_n48225__,
    new_new_n48227__, new_new_n48228__, new_new_n48229__, new_new_n48231__,
    new_new_n48232__, new_new_n48233__, new_new_n48235__, new_new_n48236__,
    new_new_n48237__, new_new_n48239__, new_new_n48240__, new_new_n48241__,
    new_new_n48243__, new_new_n48244__, new_new_n48245__, new_new_n48247__,
    new_new_n48248__, new_new_n48249__, new_new_n48251__, new_new_n48252__,
    new_new_n48253__, new_new_n48255__, new_new_n48256__, new_new_n48257__,
    new_new_n48259__, new_new_n48260__, new_new_n48261__, new_new_n48263__,
    new_new_n48264__, new_new_n48265__, new_new_n48267__, new_new_n48268__,
    new_new_n48269__, new_new_n48271__, new_new_n48272__, new_new_n48273__,
    new_new_n48275__, new_new_n48276__, new_new_n48277__, new_new_n48279__,
    new_new_n48280__, new_new_n48281__, new_new_n48283__, new_new_n48284__,
    new_new_n48285__, new_new_n48287__, new_new_n48288__, new_new_n48289__,
    new_new_n48291__, new_new_n48292__, new_new_n48293__, new_new_n48295__,
    new_new_n48296__, new_new_n48297__, new_new_n48299__, new_new_n48300__,
    new_new_n48301__, new_new_n48303__, new_new_n48304__, new_new_n48305__,
    new_new_n48307__, new_new_n48308__, new_new_n48309__, new_new_n48311__,
    new_new_n48312__, new_new_n48313__, new_new_n48315__, new_new_n48316__,
    new_new_n48317__, new_new_n48319__, new_new_n48320__, new_new_n48321__,
    new_new_n48323__, new_new_n48324__, new_new_n48325__, new_new_n48327__,
    new_new_n48328__, new_new_n48329__, new_new_n48331__, new_new_n48332__,
    new_new_n48333__, new_new_n48335__, new_new_n48336__, new_new_n48337__,
    new_new_n48339__, new_new_n48340__, new_new_n48341__, new_new_n48343__,
    new_new_n48344__, new_new_n48345__, new_new_n48347__, new_new_n48348__,
    new_new_n48349__, new_new_n48351__, new_new_n48352__, new_new_n48353__,
    new_new_n48355__, new_new_n48356__, new_new_n48357__, new_new_n48359__,
    new_new_n48360__, new_new_n48361__, new_new_n48363__, new_new_n48364__,
    new_new_n48365__, new_new_n48367__, new_new_n48368__, new_new_n48369__,
    new_new_n48371__, new_new_n48372__, new_new_n48373__, new_new_n48375__,
    new_new_n48376__, new_new_n48377__, new_new_n48379__, new_new_n48380__,
    new_new_n48381__, new_new_n48383__, new_new_n48384__, new_new_n48385__,
    new_new_n48387__, new_new_n48388__, new_new_n48389__, new_new_n48391__,
    new_new_n48392__, new_new_n48393__, new_new_n48395__, new_new_n48396__,
    new_new_n48397__, new_new_n48399__, new_new_n48400__, new_new_n48401__,
    new_new_n48403__, new_new_n48404__, new_new_n48405__, new_new_n48407__,
    new_new_n48408__, new_new_n48409__, new_new_n48411__, new_new_n48412__,
    new_new_n48413__, new_new_n48415__, new_new_n48416__, new_new_n48417__,
    new_new_n48419__, new_new_n48420__, new_new_n48421__, new_new_n48423__,
    new_new_n48424__, new_new_n48425__, new_new_n48427__, new_new_n48428__,
    new_new_n48429__, new_new_n48431__, new_new_n48432__, new_new_n48433__,
    new_new_n48435__, new_new_n48436__, new_new_n48437__, new_new_n48439__,
    new_new_n48440__, new_new_n48441__, new_new_n48443__, new_new_n48444__,
    new_new_n48445__, new_new_n48447__, new_new_n48448__, new_new_n48449__,
    new_new_n48451__, new_new_n48452__, new_new_n48453__, new_new_n48455__,
    new_new_n48456__, new_new_n48457__, new_new_n48459__, new_new_n48460__,
    new_new_n48461__, new_new_n48463__, new_new_n48464__, new_new_n48465__,
    new_new_n48467__, new_new_n48468__, new_new_n48469__, new_new_n48471__,
    new_new_n48472__, new_new_n48473__, new_new_n48475__, new_new_n48476__,
    new_new_n48477__, new_new_n48479__, new_new_n48480__, new_new_n48481__,
    new_new_n48483__, new_new_n48484__, new_new_n48485__, new_new_n48487__,
    new_new_n48488__, new_new_n48489__, new_new_n48491__, new_new_n48492__,
    new_new_n48493__, new_new_n48495__, new_new_n48496__, new_new_n48497__,
    new_new_n48499__, new_new_n48500__, new_new_n48501__, new_new_n48503__,
    new_new_n48504__, new_new_n48505__, new_new_n48507__, new_new_n48508__,
    new_new_n48509__, new_new_n48511__, new_new_n48512__, new_new_n48513__,
    new_new_n48515__, new_new_n48516__, new_new_n48517__, new_new_n48519__,
    new_new_n48520__, new_new_n48521__, new_new_n48523__, new_new_n48524__,
    new_new_n48525__, new_new_n48527__, new_new_n48528__, new_new_n48529__,
    new_new_n48531__, new_new_n48532__, new_new_n48533__, new_new_n48535__,
    new_new_n48536__, new_new_n48537__, new_new_n48539__, new_new_n48540__,
    new_new_n48541__, new_new_n48543__, new_new_n48544__, new_new_n48545__,
    new_new_n48547__, new_new_n48548__, new_new_n48549__, new_new_n48551__,
    new_new_n48552__, new_new_n48553__, new_new_n48555__, new_new_n48556__,
    new_new_n48557__, new_new_n48559__, new_new_n48560__, new_new_n48561__,
    new_new_n48563__, new_new_n48564__, new_new_n48565__, new_new_n48567__,
    new_new_n48568__, new_new_n48569__, new_new_n48571__, new_new_n48572__,
    new_new_n48573__, new_new_n48575__, new_new_n48576__, new_new_n48577__,
    new_new_n48579__, new_new_n48580__, new_new_n48581__, new_new_n48583__,
    new_new_n48584__, new_new_n48585__, new_new_n48587__, new_new_n48588__,
    new_new_n48589__, new_new_n48591__, new_new_n48592__, new_new_n48593__,
    new_new_n48595__, new_new_n48596__, new_new_n48597__, new_new_n48599__,
    new_new_n48600__, new_new_n48601__, new_new_n48603__, new_new_n48604__,
    new_new_n48605__, new_new_n48607__, new_new_n48608__, new_new_n48609__,
    new_new_n48611__, new_new_n48612__, new_new_n48613__, new_new_n48615__,
    new_new_n48616__, new_new_n48617__, new_new_n48619__, new_new_n48620__,
    new_new_n48621__, new_new_n48623__, new_new_n48624__, new_new_n48625__,
    new_new_n48627__, new_new_n48628__, new_new_n48629__, new_new_n48631__,
    new_new_n48632__, new_new_n48633__, new_new_n48635__, new_new_n48636__,
    new_new_n48637__, new_new_n48639__, new_new_n48640__, new_new_n48641__,
    new_new_n48643__, new_new_n48644__, new_new_n48645__, new_new_n48647__,
    new_new_n48648__, new_new_n48649__, new_new_n48651__, new_new_n48652__,
    new_new_n48653__, new_new_n48655__, new_new_n48656__, new_new_n48657__,
    new_new_n48659__, new_new_n48660__, new_new_n48661__, new_new_n48663__,
    new_new_n48664__, new_new_n48665__, new_new_n48667__, new_new_n48668__,
    new_new_n48669__, new_new_n48671__, new_new_n48672__, new_new_n48673__,
    new_new_n48675__, new_new_n48676__, new_new_n48677__, new_new_n48679__,
    new_new_n48680__, new_new_n48681__, new_new_n48683__, new_new_n48684__,
    new_new_n48685__, new_new_n48687__, new_new_n48688__, new_new_n48689__,
    new_new_n48691__, new_new_n48692__, new_new_n48693__, new_new_n48695__,
    new_new_n48696__, new_new_n48697__, new_new_n48699__, new_new_n48700__,
    new_new_n48701__, new_new_n48703__, new_new_n48704__, new_new_n48705__,
    new_new_n48707__, new_new_n48708__, new_new_n48709__, new_new_n48711__,
    new_new_n48712__, new_new_n48713__, new_new_n48715__, new_new_n48716__,
    new_new_n48717__, new_new_n48719__, new_new_n48720__, new_new_n48721__,
    new_new_n48723__, new_new_n48724__, new_new_n48725__, new_new_n48727__,
    new_new_n48728__, new_new_n48729__, new_new_n48731__, new_new_n48732__,
    new_new_n48733__, new_new_n48735__, new_new_n48736__, new_new_n48737__,
    new_new_n48739__, new_new_n48740__, new_new_n48741__, new_new_n48743__,
    new_new_n48744__, new_new_n48745__, new_new_n48747__, new_new_n48748__,
    new_new_n48749__, new_new_n48751__, new_new_n48752__, new_new_n48753__,
    new_new_n48755__, new_new_n48756__, new_new_n48757__, new_new_n48759__,
    new_new_n48760__, new_new_n48761__, new_new_n48763__, new_new_n48764__,
    new_new_n48765__, new_new_n48767__, new_new_n48768__, new_new_n48769__,
    new_new_n48771__, new_new_n48772__, new_new_n48773__, new_new_n48775__,
    new_new_n48776__, new_new_n48777__, new_new_n48779__, new_new_n48780__,
    new_new_n48781__, new_new_n48783__, new_new_n48784__, new_new_n48785__,
    new_new_n48787__, new_new_n48788__, new_new_n48789__, new_new_n48791__,
    new_new_n48792__, new_new_n48793__, new_new_n48795__, new_new_n48796__,
    new_new_n48797__, new_new_n48799__, new_new_n48800__, new_new_n48801__,
    new_new_n48803__, new_new_n48804__, new_new_n48805__, new_new_n48807__,
    new_new_n48808__, new_new_n48809__, new_new_n48811__, new_new_n48812__,
    new_new_n48813__, new_new_n48815__, new_new_n48816__, new_new_n48817__,
    new_new_n48819__, new_new_n48820__, new_new_n48821__, new_new_n48823__,
    new_new_n48824__, new_new_n48825__, new_new_n48827__, new_new_n48828__,
    new_new_n48829__, new_new_n48831__, new_new_n48832__, new_new_n48833__,
    new_new_n48835__, new_new_n48836__, new_new_n48837__, new_new_n48839__,
    new_new_n48840__, new_new_n48841__, new_new_n48843__, new_new_n48844__,
    new_new_n48845__, new_new_n48847__, new_new_n48848__, new_new_n48849__,
    new_new_n48851__, new_new_n48852__, new_new_n48853__, new_new_n48855__,
    new_new_n48856__, new_new_n48857__, new_new_n48859__, new_new_n48860__,
    new_new_n48861__, new_new_n48863__, new_new_n48864__, new_new_n48865__,
    new_new_n48867__, new_new_n48868__, new_new_n48869__, new_new_n48871__,
    new_new_n48872__, new_new_n48873__, new_new_n48875__, new_new_n48876__,
    new_new_n48877__, new_new_n48879__, new_new_n48880__, new_new_n48881__,
    new_new_n48883__, new_new_n48884__, new_new_n48885__, new_new_n48887__,
    new_new_n48888__, new_new_n48889__, new_new_n48891__, new_new_n48892__,
    new_new_n48893__, new_new_n48895__, new_new_n48896__, new_new_n48897__,
    new_new_n48899__, new_new_n48900__, new_new_n48901__, new_new_n48903__,
    new_new_n48904__, new_new_n48905__, new_new_n48907__, new_new_n48908__,
    new_new_n48909__, new_new_n48911__, new_new_n48912__, new_new_n48913__,
    new_new_n48915__, new_new_n48916__, new_new_n48917__, new_new_n48919__,
    new_new_n48920__, new_new_n48921__, new_new_n48923__, new_new_n48924__,
    new_new_n48925__, new_new_n48927__, new_new_n48928__, new_new_n48929__,
    new_new_n48931__, new_new_n48932__, new_new_n48933__, new_new_n48935__,
    new_new_n48936__, new_new_n48937__, new_new_n48939__, new_new_n48940__,
    new_new_n48941__, new_new_n48943__, new_new_n48944__, new_new_n48945__,
    new_new_n48947__, new_new_n48948__, new_new_n48949__, new_new_n48951__,
    new_new_n48952__, new_new_n48953__, new_new_n48955__, new_new_n48956__,
    new_new_n48957__, new_new_n48959__, new_new_n48960__, new_new_n48961__,
    new_new_n48963__, new_new_n48964__, new_new_n48965__, new_new_n48967__,
    new_new_n48968__, new_new_n48969__, new_new_n48971__, new_new_n48972__,
    new_new_n48973__, new_new_n48975__, new_new_n48976__, new_new_n48977__,
    new_new_n48979__, new_new_n48980__, new_new_n48981__, new_new_n48983__,
    new_new_n48984__, new_new_n48985__, new_new_n48987__, new_new_n48988__,
    new_new_n48989__, new_new_n48991__, new_new_n48992__, new_new_n48993__,
    new_new_n48995__, new_new_n48996__, new_new_n48997__, new_new_n48999__,
    new_new_n49000__, new_new_n49001__, new_new_n49003__, new_new_n49004__,
    new_new_n49005__, new_new_n49007__, new_new_n49008__, new_new_n49009__,
    new_new_n49011__, new_new_n49012__, new_new_n49013__, new_new_n49015__,
    new_new_n49016__, new_new_n49017__, new_new_n49019__, new_new_n49020__,
    new_new_n49021__, new_new_n49023__, new_new_n49024__, new_new_n49025__,
    new_new_n49027__, new_new_n49028__, new_new_n49029__, new_new_n49031__,
    new_new_n49032__, new_new_n49033__, new_new_n49035__, new_new_n49036__,
    new_new_n49037__, new_new_n49039__, new_new_n49040__, new_new_n49041__,
    new_new_n49043__, new_new_n49044__, new_new_n49045__, new_new_n49047__,
    new_new_n49048__, new_new_n49049__, new_new_n49051__, new_new_n49052__,
    new_new_n49053__, new_new_n49055__, new_new_n49056__, new_new_n49057__,
    new_new_n49059__, new_new_n49060__, new_new_n49061__, new_new_n49063__,
    new_new_n49064__, new_new_n49065__, new_new_n49067__, new_new_n49068__,
    new_new_n49069__, new_new_n49071__, new_new_n49072__, new_new_n49073__,
    new_new_n49075__, new_new_n49076__, new_new_n49077__, new_new_n49079__,
    new_new_n49080__, new_new_n49081__, new_new_n49083__, new_new_n49084__,
    new_new_n49085__, new_new_n49087__, new_new_n49088__, new_new_n49089__,
    new_new_n49091__, new_new_n49092__, new_new_n49093__, new_new_n49095__,
    new_new_n49096__, new_new_n49097__, new_new_n49099__, new_new_n49100__,
    new_new_n49101__, new_new_n49103__, new_new_n49104__, new_new_n49105__,
    new_new_n49107__, new_new_n49108__, new_new_n49109__, new_new_n49111__,
    new_new_n49112__, new_new_n49113__, new_new_n49115__, new_new_n49116__,
    new_new_n49117__, new_new_n49119__, new_new_n49120__, new_new_n49121__,
    new_new_n49123__, new_new_n49124__, new_new_n49125__, new_new_n49127__,
    new_new_n49128__, new_new_n49129__, new_new_n49131__, new_new_n49132__,
    new_new_n49133__, new_new_n49135__, new_new_n49136__, new_new_n49137__,
    new_new_n49139__, new_new_n49140__, new_new_n49141__, new_new_n49143__,
    new_new_n49144__, new_new_n49145__, new_new_n49147__, new_new_n49148__,
    new_new_n49149__, new_new_n49151__, new_new_n49152__, new_new_n49153__,
    new_new_n49155__, new_new_n49156__, new_new_n49157__, new_new_n49159__,
    new_new_n49160__, new_new_n49161__, new_new_n49163__, new_new_n49164__,
    new_new_n49165__, new_new_n49167__, new_new_n49168__, new_new_n49169__,
    new_new_n49171__, new_new_n49172__, new_new_n49173__, new_new_n49175__,
    new_new_n49176__, new_new_n49177__, new_new_n49179__, new_new_n49180__,
    new_new_n49181__, new_new_n49183__, new_new_n49184__, new_new_n49185__,
    new_new_n49187__, new_new_n49188__, new_new_n49189__, new_new_n49191__,
    new_new_n49192__, new_new_n49193__, new_new_n49195__, new_new_n49196__,
    new_new_n49197__, new_new_n49199__, new_new_n49200__, new_new_n49201__,
    new_new_n49203__, new_new_n49204__, new_new_n49205__, new_new_n49207__,
    new_new_n49208__, new_new_n49209__, new_new_n49211__, new_new_n49212__,
    new_new_n49213__, new_new_n49215__, new_new_n49216__, new_new_n49217__,
    new_new_n49219__, new_new_n49220__, new_new_n49221__, new_new_n49223__,
    new_new_n49224__, new_new_n49225__, new_new_n49227__, new_new_n49228__,
    new_new_n49229__, new_new_n49231__, new_new_n49232__, new_new_n49233__,
    new_new_n49235__, new_new_n49236__, new_new_n49237__, new_new_n49239__,
    new_new_n49240__, new_new_n49241__, new_new_n49243__, new_new_n49244__,
    new_new_n49245__, new_new_n49248__, new_new_n49249__, new_new_n49250__,
    new_new_n49251__, new_new_n49252__, new_new_n49253__, new_new_n49254__,
    new_new_n49255__, new_new_n49256__, new_new_n49257__, new_new_n49258__,
    new_new_n49259__, new_new_n49260__, new_new_n49261__, new_new_n49262__,
    new_new_n49263__, new_new_n49264__, new_new_n49266__, new_new_n49267__,
    new_new_n49268__, new_new_n49269__, new_new_n49270__, new_new_n49271__,
    new_new_n49272__, new_new_n49273__, new_new_n49274__, new_new_n49275__,
    new_new_n49276__, new_new_n49277__, new_new_n49279__, new_new_n49280__,
    new_new_n49281__, new_new_n49282__, new_new_n49283__, new_new_n49284__,
    new_new_n49285__, new_new_n49286__, new_new_n49287__, new_new_n49288__,
    new_new_n49289__, new_new_n49290__, new_new_n49292__, new_new_n49293__,
    new_new_n49294__, new_new_n49295__, new_new_n49296__, new_new_n49297__,
    new_new_n49298__, new_new_n49299__, new_new_n49300__, new_new_n49301__,
    new_new_n49302__, new_new_n49303__, new_new_n49305__, new_new_n49306__,
    new_new_n49307__, new_new_n49308__, new_new_n49309__, new_new_n49310__,
    new_new_n49311__, new_new_n49312__, new_new_n49313__, new_new_n49314__,
    new_new_n49315__, new_new_n49316__, new_new_n49318__, new_new_n49319__,
    new_new_n49320__, new_new_n49321__, new_new_n49322__, new_new_n49323__,
    new_new_n49324__, new_new_n49325__, new_new_n49326__, new_new_n49327__,
    new_new_n49328__, new_new_n49329__, new_new_n49331__, new_new_n49332__,
    new_new_n49333__, new_new_n49334__, new_new_n49335__, new_new_n49336__,
    new_new_n49337__, new_new_n49338__, new_new_n49339__, new_new_n49340__,
    new_new_n49341__, new_new_n49342__, new_new_n49344__, new_new_n49345__,
    new_new_n49346__, new_new_n49347__, new_new_n49348__, new_new_n49349__,
    new_new_n49350__, new_new_n49351__, new_new_n49352__, new_new_n49353__,
    new_new_n49354__, new_new_n49355__, new_new_n49357__, new_new_n49358__,
    new_new_n49359__, new_new_n49360__, new_new_n49361__, new_new_n49362__,
    new_new_n49363__, new_new_n49364__, new_new_n49365__, new_new_n49366__,
    new_new_n49367__, new_new_n49368__, new_new_n49370__, new_new_n49371__,
    new_new_n49372__, new_new_n49373__, new_new_n49374__, new_new_n49375__,
    new_new_n49376__, new_new_n49377__, new_new_n49378__, new_new_n49379__,
    new_new_n49380__, new_new_n49381__, new_new_n49383__, new_new_n49384__,
    new_new_n49385__, new_new_n49386__, new_new_n49387__, new_new_n49388__,
    new_new_n49389__, new_new_n49390__, new_new_n49391__, new_new_n49392__,
    new_new_n49393__, new_new_n49394__, new_new_n49396__, new_new_n49397__,
    new_new_n49398__, new_new_n49399__, new_new_n49400__, new_new_n49401__,
    new_new_n49402__, new_new_n49403__, new_new_n49404__, new_new_n49405__,
    new_new_n49406__, new_new_n49407__, new_new_n49409__, new_new_n49410__,
    new_new_n49411__, new_new_n49412__, new_new_n49413__, new_new_n49414__,
    new_new_n49415__, new_new_n49416__, new_new_n49417__, new_new_n49418__,
    new_new_n49419__, new_new_n49420__, new_new_n49422__, new_new_n49423__,
    new_new_n49424__, new_new_n49425__, new_new_n49426__, new_new_n49427__,
    new_new_n49428__, new_new_n49429__, new_new_n49430__, new_new_n49431__,
    new_new_n49432__, new_new_n49433__, new_new_n49435__, new_new_n49436__,
    new_new_n49437__, new_new_n49438__, new_new_n49439__, new_new_n49440__,
    new_new_n49441__, new_new_n49442__, new_new_n49443__, new_new_n49444__,
    new_new_n49445__, new_new_n49446__, new_new_n49448__, new_new_n49449__,
    new_new_n49450__, new_new_n49451__, new_new_n49452__, new_new_n49453__,
    new_new_n49454__, new_new_n49455__, new_new_n49456__, new_new_n49457__,
    new_new_n49458__, new_new_n49459__, new_new_n49461__, new_new_n49462__,
    new_new_n49463__, new_new_n49464__, new_new_n49465__, new_new_n49466__,
    new_new_n49467__, new_new_n49468__, new_new_n49469__, new_new_n49470__,
    new_new_n49471__, new_new_n49472__, new_new_n49474__, new_new_n49475__,
    new_new_n49476__, new_new_n49477__, new_new_n49478__, new_new_n49479__,
    new_new_n49480__, new_new_n49481__, new_new_n49482__, new_new_n49483__,
    new_new_n49484__, new_new_n49485__, new_new_n49487__, new_new_n49488__,
    new_new_n49489__, new_new_n49490__, new_new_n49491__, new_new_n49492__,
    new_new_n49493__, new_new_n49494__, new_new_n49495__, new_new_n49496__,
    new_new_n49497__, new_new_n49498__, new_new_n49500__, new_new_n49501__,
    new_new_n49502__, new_new_n49503__, new_new_n49504__, new_new_n49505__,
    new_new_n49506__, new_new_n49507__, new_new_n49508__, new_new_n49509__,
    new_new_n49510__, new_new_n49511__, new_new_n49513__, new_new_n49514__,
    new_new_n49515__, new_new_n49516__, new_new_n49517__, new_new_n49518__,
    new_new_n49519__, new_new_n49520__, new_new_n49521__, new_new_n49522__,
    new_new_n49523__, new_new_n49524__, new_new_n49526__, new_new_n49527__,
    new_new_n49528__, new_new_n49529__, new_new_n49531__, new_new_n49532__,
    new_new_n49533__, new_new_n49534__, new_new_n49535__, new_new_n49536__,
    new_new_n49537__, new_new_n49538__, new_new_n49539__, new_new_n49540__,
    new_new_n49541__, new_new_n49542__, new_new_n49543__, new_new_n49545__,
    new_new_n49546__, new_new_n49547__, new_new_n49548__, new_new_n49549__,
    new_new_n49550__, new_new_n49551__, new_new_n49552__, new_new_n49553__,
    new_new_n49555__, new_new_n49556__, new_new_n49557__, new_new_n49558__,
    new_new_n49559__, new_new_n49560__, new_new_n49561__, new_new_n49562__,
    new_new_n49563__, new_new_n49565__, new_new_n49566__, new_new_n49567__,
    new_new_n49568__, new_new_n49569__, new_new_n49570__, new_new_n49571__,
    new_new_n49572__, new_new_n49573__, new_new_n49575__, new_new_n49576__,
    new_new_n49577__, new_new_n49578__, new_new_n49579__, new_new_n49580__,
    new_new_n49581__, new_new_n49582__, new_new_n49583__, new_new_n49585__,
    new_new_n49586__, new_new_n49587__, new_new_n49588__, new_new_n49589__,
    new_new_n49590__, new_new_n49591__, new_new_n49592__, new_new_n49593__,
    new_new_n49595__, new_new_n49596__, new_new_n49597__, new_new_n49598__,
    new_new_n49599__, new_new_n49600__, new_new_n49601__, new_new_n49602__,
    new_new_n49603__, new_new_n49605__, new_new_n49606__, new_new_n49607__,
    new_new_n49608__, new_new_n49609__, new_new_n49610__, new_new_n49611__,
    new_new_n49612__, new_new_n49613__, new_new_n49615__, new_new_n49616__,
    new_new_n49617__, new_new_n49618__, new_new_n49619__, new_new_n49620__,
    new_new_n49621__, new_new_n49622__, new_new_n49623__, new_new_n49625__,
    new_new_n49626__, new_new_n49627__, new_new_n49628__, new_new_n49629__,
    new_new_n49630__, new_new_n49631__, new_new_n49632__, new_new_n49633__,
    new_new_n49635__, new_new_n49636__, new_new_n49637__, new_new_n49638__,
    new_new_n49639__, new_new_n49640__, new_new_n49641__, new_new_n49642__,
    new_new_n49643__, new_new_n49645__, new_new_n49646__, new_new_n49647__,
    new_new_n49648__, new_new_n49649__, new_new_n49650__, new_new_n49651__,
    new_new_n49652__, new_new_n49653__, new_new_n49655__, new_new_n49656__,
    new_new_n49657__, new_new_n49658__, new_new_n49659__, new_new_n49660__,
    new_new_n49661__, new_new_n49662__, new_new_n49663__, new_new_n49665__,
    new_new_n49666__, new_new_n49667__, new_new_n49668__, new_new_n49669__,
    new_new_n49670__, new_new_n49671__, new_new_n49672__, new_new_n49673__,
    new_new_n49675__, new_new_n49676__, new_new_n49677__, new_new_n49678__,
    new_new_n49679__, new_new_n49680__, new_new_n49681__, new_new_n49682__,
    new_new_n49683__, new_new_n49685__, new_new_n49686__, new_new_n49687__,
    new_new_n49688__, new_new_n49689__, new_new_n49690__, new_new_n49691__,
    new_new_n49692__, new_new_n49693__, new_new_n49695__, new_new_n49696__,
    new_new_n49697__, new_new_n49698__, new_new_n49699__, new_new_n49700__,
    new_new_n49701__, new_new_n49702__, new_new_n49703__, new_new_n49705__,
    new_new_n49706__, new_new_n49707__, new_new_n49708__, new_new_n49709__,
    new_new_n49710__, new_new_n49711__, new_new_n49712__, new_new_n49713__,
    new_new_n49715__, new_new_n49716__, new_new_n49717__, new_new_n49718__,
    new_new_n49719__, new_new_n49720__, new_new_n49721__, new_new_n49722__,
    new_new_n49723__, new_new_n49725__, new_new_n49726__, new_new_n49727__,
    new_new_n49728__, new_new_n49729__, new_new_n49730__, new_new_n49731__,
    new_new_n49732__, new_new_n49733__, new_new_n49735__, new_new_n49736__,
    new_new_n49737__, new_new_n49738__, new_new_n49739__, new_new_n49740__,
    new_new_n49741__, new_new_n49742__, new_new_n49743__, new_new_n49745__,
    new_new_n49746__, new_new_n49747__, new_new_n49748__, new_new_n49750__,
    new_new_n49751__, new_new_n49752__, new_new_n49753__, new_new_n49754__,
    new_new_n49755__, new_new_n49756__, new_new_n49757__, new_new_n49758__,
    new_new_n49759__, new_new_n49760__, new_new_n49761__, new_new_n49762__,
    new_new_n49764__, new_new_n49765__, new_new_n49766__, new_new_n49767__,
    new_new_n49768__, new_new_n49769__, new_new_n49770__, new_new_n49771__,
    new_new_n49772__, new_new_n49774__, new_new_n49775__, new_new_n49776__,
    new_new_n49777__, new_new_n49778__, new_new_n49779__, new_new_n49780__,
    new_new_n49781__, new_new_n49782__, new_new_n49784__, new_new_n49785__,
    new_new_n49786__, new_new_n49787__, new_new_n49788__, new_new_n49789__,
    new_new_n49790__, new_new_n49791__, new_new_n49792__, new_new_n49794__,
    new_new_n49795__, new_new_n49796__, new_new_n49797__, new_new_n49798__,
    new_new_n49799__, new_new_n49800__, new_new_n49801__, new_new_n49802__,
    new_new_n49804__, new_new_n49805__, new_new_n49806__, new_new_n49807__,
    new_new_n49808__, new_new_n49809__, new_new_n49810__, new_new_n49811__,
    new_new_n49812__, new_new_n49814__, new_new_n49815__, new_new_n49816__,
    new_new_n49817__, new_new_n49818__, new_new_n49819__, new_new_n49820__,
    new_new_n49821__, new_new_n49822__, new_new_n49824__, new_new_n49825__,
    new_new_n49826__, new_new_n49827__, new_new_n49828__, new_new_n49829__,
    new_new_n49830__, new_new_n49831__, new_new_n49832__, new_new_n49834__,
    new_new_n49835__, new_new_n49836__, new_new_n49837__, new_new_n49838__,
    new_new_n49839__, new_new_n49840__, new_new_n49841__, new_new_n49842__,
    new_new_n49844__, new_new_n49845__, new_new_n49846__, new_new_n49847__,
    new_new_n49848__, new_new_n49849__, new_new_n49850__, new_new_n49851__,
    new_new_n49852__, new_new_n49854__, new_new_n49855__, new_new_n49856__,
    new_new_n49857__, new_new_n49858__, new_new_n49859__, new_new_n49860__,
    new_new_n49861__, new_new_n49862__, new_new_n49864__, new_new_n49865__,
    new_new_n49866__, new_new_n49867__, new_new_n49868__, new_new_n49869__,
    new_new_n49870__, new_new_n49871__, new_new_n49872__, new_new_n49874__,
    new_new_n49875__, new_new_n49876__, new_new_n49877__, new_new_n49878__,
    new_new_n49879__, new_new_n49880__, new_new_n49881__, new_new_n49882__,
    new_new_n49884__, new_new_n49885__, new_new_n49886__, new_new_n49887__,
    new_new_n49888__, new_new_n49889__, new_new_n49890__, new_new_n49891__,
    new_new_n49892__, new_new_n49894__, new_new_n49895__, new_new_n49896__,
    new_new_n49897__, new_new_n49898__, new_new_n49899__, new_new_n49900__,
    new_new_n49901__, new_new_n49902__, new_new_n49904__, new_new_n49905__,
    new_new_n49906__, new_new_n49907__, new_new_n49908__, new_new_n49909__,
    new_new_n49910__, new_new_n49911__, new_new_n49912__, new_new_n49914__,
    new_new_n49915__, new_new_n49916__, new_new_n49917__, new_new_n49918__,
    new_new_n49919__, new_new_n49920__, new_new_n49921__, new_new_n49922__,
    new_new_n49924__, new_new_n49925__, new_new_n49926__, new_new_n49927__,
    new_new_n49928__, new_new_n49929__, new_new_n49930__, new_new_n49931__,
    new_new_n49932__, new_new_n49934__, new_new_n49935__, new_new_n49936__,
    new_new_n49937__, new_new_n49938__, new_new_n49939__, new_new_n49940__,
    new_new_n49941__, new_new_n49942__, new_new_n49944__, new_new_n49945__,
    new_new_n49946__, new_new_n49947__, new_new_n49948__, new_new_n49949__,
    new_new_n49950__, new_new_n49951__, new_new_n49952__, new_new_n49954__,
    new_new_n49955__, new_new_n49956__, new_new_n49957__, new_new_n49958__,
    new_new_n49959__, new_new_n49960__, new_new_n49961__, new_new_n49962__,
    new_new_n49964__, new_new_n49965__, new_new_n49966__, new_new_n49968__,
    new_new_n49969__, new_new_n49970__, new_new_n49971__, new_new_n49972__,
    new_new_n49973__, new_new_n49975__, new_new_n49976__, new_new_n49977__,
    new_new_n49978__, new_new_n49979__, new_new_n49980__, new_new_n49982__,
    new_new_n49983__, new_new_n49984__, new_new_n49985__, new_new_n49986__,
    new_new_n49987__, new_new_n49989__, new_new_n49990__, new_new_n49991__,
    new_new_n49992__, new_new_n49993__, new_new_n49994__, new_new_n49996__,
    new_new_n49997__, new_new_n49998__, new_new_n49999__, new_new_n50000__,
    new_new_n50001__, new_new_n50003__, new_new_n50004__, new_new_n50005__,
    new_new_n50006__, new_new_n50007__, new_new_n50008__, new_new_n50010__,
    new_new_n50011__, new_new_n50012__, new_new_n50013__, new_new_n50014__,
    new_new_n50015__, new_new_n50017__, new_new_n50018__, new_new_n50019__,
    new_new_n50020__, new_new_n50021__, new_new_n50022__, new_new_n50024__,
    new_new_n50025__, new_new_n50026__, new_new_n50027__, new_new_n50028__,
    new_new_n50029__, new_new_n50031__, new_new_n50032__, new_new_n50033__,
    new_new_n50034__, new_new_n50035__, new_new_n50036__, new_new_n50038__,
    new_new_n50039__, new_new_n50040__, new_new_n50041__, new_new_n50042__,
    new_new_n50043__, new_new_n50045__, new_new_n50046__, new_new_n50047__,
    new_new_n50048__, new_new_n50049__, new_new_n50050__, new_new_n50052__,
    new_new_n50053__, new_new_n50054__, new_new_n50055__, new_new_n50056__,
    new_new_n50057__, new_new_n50059__, new_new_n50060__, new_new_n50061__,
    new_new_n50062__, new_new_n50063__, new_new_n50064__, new_new_n50066__,
    new_new_n50067__, new_new_n50068__, new_new_n50069__, new_new_n50070__,
    new_new_n50071__, new_new_n50073__, new_new_n50074__, new_new_n50075__,
    new_new_n50076__, new_new_n50077__, new_new_n50078__, new_new_n50080__,
    new_new_n50081__, new_new_n50082__, new_new_n50083__, new_new_n50084__,
    new_new_n50085__, new_new_n50087__, new_new_n50088__, new_new_n50089__,
    new_new_n50090__, new_new_n50091__, new_new_n50092__, new_new_n50094__,
    new_new_n50095__, new_new_n50096__, new_new_n50097__, new_new_n50098__,
    new_new_n50099__, new_new_n50101__, new_new_n50102__, new_new_n50103__,
    new_new_n50104__, new_new_n50105__, new_new_n50106__, new_new_n50108__,
    new_new_n50109__, new_new_n50110__, new_new_n50111__, new_new_n50112__,
    new_new_n50113__, new_new_n50115__, new_new_n50116__, new_new_n50117__,
    new_new_n50118__, new_new_n50119__, new_new_n50120__, new_new_n50122__,
    new_new_n50123__, new_new_n50124__, new_new_n50125__, new_new_n50126__,
    new_new_n50127__, new_new_n50129__, new_new_n50130__, new_new_n50131__,
    new_new_n50132__, new_new_n50133__, new_new_n50134__, new_new_n50136__,
    new_new_n50137__, new_new_n50138__, new_new_n50139__, new_new_n50140__,
    new_new_n50141__, new_new_n50143__, new_new_n50144__, new_new_n50145__,
    new_new_n50146__, new_new_n50147__, new_new_n50148__, new_new_n50150__,
    new_new_n50151__, new_new_n50152__, new_new_n50153__, new_new_n50154__,
    new_new_n50155__, new_new_n50157__, new_new_n50158__, new_new_n50159__,
    new_new_n50160__, new_new_n50161__, new_new_n50162__, new_new_n50164__,
    new_new_n50165__, new_new_n50166__, new_new_n50167__, new_new_n50168__,
    new_new_n50169__, new_new_n50171__, new_new_n50172__, new_new_n50173__,
    new_new_n50174__, new_new_n50175__, new_new_n50176__, new_new_n50178__,
    new_new_n50179__, new_new_n50180__, new_new_n50181__, new_new_n50182__,
    new_new_n50183__, new_new_n50185__, new_new_n50186__, new_new_n50187__,
    new_new_n50188__, new_new_n50190__, new_new_n50193__, new_new_n50194__,
    new_new_n50195__, new_new_n50196__, new_new_n50197__, new_new_n50198__,
    new_new_n50199__, new_new_n50200__, new_new_n50201__, new_new_n50202__,
    new_new_n50203__, new_new_n50205__, new_new_n50206__, new_new_n50207__,
    new_new_n50208__, new_new_n50209__, new_new_n50213__, new_new_n50215__,
    new_new_n50216__, new_new_n50217__, new_new_n50218__, new_new_n50220__,
    new_new_n50221__, new_new_n50223__, new_new_n50224__, new_new_n50225__,
    new_new_n50227__, new_new_n50228__, new_new_n50229__, new_new_n50231__,
    new_new_n50232__, new_new_n50233__, new_new_n50234__, new_new_n50236__,
    new_new_n50237__, new_new_n50238__, new_new_n50240__, new_new_n50241__,
    new_new_n50242__, new_new_n50243__, new_new_n50245__, new_new_n50246__,
    new_new_n50247__, new_new_n50249__, new_new_n50250__, new_new_n50251__,
    new_new_n50252__, new_new_n50253__, new_new_n50255__, new_new_n50256__,
    new_new_n50257__, new_new_n50259__, new_new_n50260__, new_new_n50261__,
    new_new_n50262__, new_new_n50264__, new_new_n50265__, new_new_n50266__,
    new_new_n50268__, new_new_n50269__, new_new_n50270__, new_new_n50271__,
    new_new_n50272__, new_new_n50274__, new_new_n50275__, new_new_n50276__,
    new_new_n50278__, new_new_n50279__, new_new_n50280__, new_new_n50281__,
    new_new_n50283__, new_new_n50284__, new_new_n50285__, new_new_n50287__,
    new_new_n50288__, new_new_n50289__, new_new_n50290__, new_new_n50291__,
    new_new_n50292__, new_new_n50294__, new_new_n50295__, new_new_n50296__,
    new_new_n50298__, new_new_n50299__, new_new_n50300__, new_new_n50301__,
    new_new_n50303__, new_new_n50304__, new_new_n50305__, new_new_n50307__,
    new_new_n50308__, new_new_n50309__, new_new_n50310__, new_new_n50311__,
    new_new_n50313__, new_new_n50314__, new_new_n50315__, new_new_n50317__,
    new_new_n50318__, new_new_n50319__, new_new_n50320__, new_new_n50322__,
    new_new_n50323__, new_new_n50324__, new_new_n50326__, new_new_n50327__,
    new_new_n50328__, new_new_n50329__, new_new_n50330__, new_new_n50331__,
    new_new_n50333__, new_new_n50334__, new_new_n50335__, new_new_n50337__,
    new_new_n50338__, new_new_n50339__, new_new_n50340__, new_new_n50342__,
    new_new_n50343__, new_new_n50344__, new_new_n50346__, new_new_n50347__,
    new_new_n50348__, new_new_n50349__, new_new_n50350__, new_new_n50352__,
    new_new_n50353__, new_new_n50354__, new_new_n50356__, new_new_n50357__,
    new_new_n50358__, new_new_n50359__, new_new_n50361__, new_new_n50362__,
    new_new_n50363__, new_new_n50365__, new_new_n50366__, new_new_n50367__,
    new_new_n50368__, new_new_n50369__, new_new_n50370__, new_new_n50371__,
    new_new_n50373__, new_new_n50374__, new_new_n50376__, new_new_n50377__,
    new_new_n50379__, new_new_n50380__, new_new_n50381__, new_new_n50383__,
    new_new_n50384__, new_new_n50386__, new_new_n50387__, new_new_n50388__,
    new_new_n50390__, new_new_n50391__, new_new_n50392__, new_new_n50394__,
    new_new_n50395__, new_new_n50397__, new_new_n50398__, new_new_n50400__,
    new_new_n50401__, new_new_n50402__, new_new_n50404__, new_new_n50405__,
    new_new_n50407__, new_new_n50408__, new_new_n50409__, new_new_n50411__,
    new_new_n50412__, new_new_n50413__, new_new_n50415__, new_new_n50416__,
    new_new_n50420__, new_new_n50421__, new_new_n50423__, new_new_n50424__,
    new_new_n50425__, new_new_n50427__, new_new_n50428__, new_new_n50429__,
    new_new_n50430__, new_new_n50432__, new_new_n50433__, new_new_n50438__,
    new_new_n50439__, new_new_n50440__, new_new_n50441__, new_new_n50442__,
    new_new_n50443__, new_new_n50445__, new_new_n50446__, new_new_n50448__,
    new_new_n50449__, new_new_n50450__, new_new_n50452__, new_new_n50453__,
    new_new_n50454__, new_new_n50455__, new_new_n50456__, new_new_n50457__,
    new_new_n50458__, new_new_n50459__, new_new_n50460__, new_new_n50461__,
    new_new_n50462__, new_new_n50463__, new_new_n50464__, new_new_n50465__,
    new_new_n50466__, new_new_n50467__, new_new_n50468__, new_new_n50469__,
    new_new_n50470__, new_new_n50473__, new_new_n50474__, new_new_n50475__,
    new_new_n50476__, new_new_n50477__, new_new_n50481__, new_new_n50482__,
    new_new_n50483__, new_new_n50484__, new_new_n50485__, new_new_n50486__,
    new_new_n50487__, new_new_n50488__, new_new_n50489__, new_new_n50490__,
    new_new_n50491__, new_new_n50492__, new_new_n50494__, new_new_n50495__,
    new_new_n50496__, new_new_n50497__, new_new_n50498__, new_new_n50499__,
    new_new_n50500__, new_new_n50501__, new_new_n50502__, new_new_n50503__,
    new_new_n50504__, new_new_n50505__, new_new_n50506__, new_new_n50507__,
    new_new_n50508__, new_new_n50509__, new_new_n50510__, new_new_n50511__,
    new_new_n50512__, new_new_n50513__, new_new_n50514__, new_new_n50515__,
    new_new_n50516__, new_new_n50517__, new_new_n50518__, new_new_n50519__,
    new_new_n50520__, new_new_n50521__, new_new_n50522__, new_new_n50523__,
    new_new_n50524__, new_new_n50525__, new_new_n50526__, new_new_n50527__,
    new_new_n50528__, new_new_n50529__, new_new_n50530__, new_new_n50531__,
    new_new_n50532__, new_new_n50533__, new_new_n50534__, new_new_n50535__,
    new_new_n50536__, new_new_n50537__, new_new_n50538__, new_new_n50539__,
    new_new_n50540__, new_new_n50541__, new_new_n50542__, new_new_n50543__,
    new_new_n50544__, new_new_n50545__, new_new_n50546__, new_new_n50547__,
    new_new_n50548__, new_new_n50549__, new_new_n50550__, new_new_n50551__,
    new_new_n50552__, new_new_n50553__, new_new_n50554__, new_new_n50555__,
    new_new_n50556__, new_new_n50557__, new_new_n50558__, new_new_n50559__,
    new_new_n50560__, new_new_n50561__, new_new_n50562__, new_new_n50563__,
    new_new_n50564__, new_new_n50565__, new_new_n50566__, new_new_n50567__,
    new_new_n50568__, new_new_n50569__, new_new_n50570__, new_new_n50571__,
    new_new_n50572__, new_new_n50573__, new_new_n50574__, new_new_n50575__,
    new_new_n50576__, new_new_n50577__, new_new_n50578__, new_new_n50579__,
    new_new_n50580__, new_new_n50581__, new_new_n50582__, new_new_n50583__,
    new_new_n50584__, new_new_n50585__, new_new_n50586__, new_new_n50587__,
    new_new_n50588__, new_new_n50589__, new_new_n50590__, new_new_n50591__,
    new_new_n50592__, new_new_n50593__, new_new_n50594__, new_new_n50595__,
    new_new_n50596__, new_new_n50597__, new_new_n50598__, new_new_n50599__,
    new_new_n50600__, new_new_n50601__, new_new_n50602__, new_new_n50603__,
    new_new_n50604__, new_new_n50605__, new_new_n50606__, new_new_n50607__,
    new_new_n50608__, new_new_n50609__, new_new_n50610__, new_new_n50611__,
    new_new_n50612__, new_new_n50613__, new_new_n50614__, new_new_n50615__,
    new_new_n50616__, new_new_n50617__, new_new_n50618__, new_new_n50619__,
    new_new_n50620__, new_new_n50621__, new_new_n50622__, new_new_n50623__,
    new_new_n50624__, new_new_n50625__, new_new_n50626__, new_new_n50627__,
    new_new_n50628__, new_new_n50629__, new_new_n50630__, new_new_n50631__,
    new_new_n50632__, new_new_n50633__, new_new_n50634__, new_new_n50635__,
    new_new_n50636__, new_new_n50637__, new_new_n50638__, new_new_n50639__,
    new_new_n50640__, new_new_n50641__, new_new_n50642__, new_new_n50643__,
    new_new_n50644__, new_new_n50645__, new_new_n50646__, new_new_n50647__,
    new_new_n50648__, new_new_n50649__, new_new_n50650__, new_new_n50651__,
    new_new_n50652__, new_new_n50653__, new_new_n50654__, new_new_n50655__,
    new_new_n50656__, new_new_n50657__, new_new_n50658__, new_new_n50659__,
    new_new_n50660__, new_new_n50661__, new_new_n50662__, new_new_n50663__,
    new_new_n50664__, new_new_n50665__, new_new_n50666__, new_new_n50667__,
    new_new_n50668__, new_new_n50669__, new_new_n50670__, new_new_n50671__,
    new_new_n50672__, new_new_n50673__, new_new_n50674__, new_new_n50675__,
    new_new_n50676__, new_new_n50677__, new_new_n50678__, new_new_n50679__,
    new_new_n50680__, new_new_n50681__, new_new_n50682__, new_new_n50683__,
    new_new_n50684__, new_new_n50685__, new_new_n50686__, new_new_n50687__,
    new_new_n50688__, new_new_n50689__, new_new_n50690__, new_new_n50691__,
    new_new_n50692__, new_new_n50693__, new_new_n50694__, new_new_n50695__,
    new_new_n50696__, new_new_n50697__, new_new_n50698__, new_new_n50699__,
    new_new_n50700__, new_new_n50701__, new_new_n50702__, new_new_n50703__,
    new_new_n50704__, new_new_n50705__, new_new_n50706__, new_new_n50707__,
    new_new_n50708__, new_new_n50709__, new_new_n50710__, new_new_n50711__,
    new_new_n50712__, new_new_n50713__, new_new_n50714__, new_new_n50715__,
    new_new_n50716__, new_new_n50717__, new_new_n50718__, new_new_n50719__,
    new_new_n50720__, new_new_n50721__, new_new_n50722__, new_new_n50723__,
    new_new_n50724__, new_new_n50725__, new_new_n50726__, new_new_n50727__,
    new_new_n50728__, new_new_n50729__, new_new_n50730__, new_new_n50731__,
    new_new_n50732__, new_new_n50733__, new_new_n50734__, new_new_n50735__,
    new_new_n50736__, new_new_n50737__, new_new_n50738__, new_new_n50739__,
    new_new_n50740__, new_new_n50741__, new_new_n50742__, new_new_n50743__,
    new_new_n50744__, new_new_n50745__, new_new_n50746__, new_new_n50747__,
    new_new_n50748__, new_new_n50749__, new_new_n50750__, new_new_n50751__,
    new_new_n50752__, new_new_n50753__, new_new_n50754__, new_new_n50755__,
    new_new_n50756__, new_new_n50757__, new_new_n50758__, new_new_n50759__,
    new_new_n50760__, new_new_n50761__, new_new_n50762__, new_new_n50763__,
    new_new_n50764__, new_new_n50765__, new_new_n50766__, new_new_n50767__,
    new_new_n50768__, new_new_n50769__, new_new_n50770__, new_new_n50771__,
    new_new_n50772__, new_new_n50773__, new_new_n50774__, new_new_n50775__,
    new_new_n50776__, new_new_n50777__, new_new_n50778__, new_new_n50779__,
    new_new_n50780__, new_new_n50781__, new_new_n50782__, new_new_n50783__,
    new_new_n50784__, new_new_n50785__, new_new_n50786__, new_new_n50787__,
    new_new_n50788__, new_new_n50789__, new_new_n50790__, new_new_n50791__,
    new_new_n50792__, new_new_n50793__, new_new_n50794__, new_new_n50795__,
    new_new_n50796__, new_new_n50797__, new_new_n50798__, new_new_n50799__,
    new_new_n50800__, new_new_n50801__, new_new_n50802__, new_new_n50803__,
    new_new_n50804__, new_new_n50805__, new_new_n50806__, new_new_n50807__,
    new_new_n50808__, new_new_n50809__, new_new_n50810__, new_new_n50811__,
    new_new_n50812__, new_new_n50813__, new_new_n50814__, new_new_n50815__,
    new_new_n50816__, new_new_n50817__, new_new_n50818__, new_new_n50819__,
    new_new_n50820__, new_new_n50821__, new_new_n50822__, new_new_n50823__,
    new_new_n50824__, new_new_n50825__, new_new_n50826__, new_new_n50827__,
    new_new_n50828__, new_new_n50829__, new_new_n50830__, new_new_n50831__,
    new_new_n50832__, new_new_n50833__, new_new_n50834__, new_new_n50835__,
    new_new_n50836__, new_new_n50837__, new_new_n50838__, new_new_n50839__,
    new_new_n50840__, new_new_n50841__, new_new_n50842__, new_new_n50843__,
    new_new_n50844__, new_new_n50845__, new_new_n50846__, new_new_n50847__,
    new_new_n50848__, new_new_n50849__, new_new_n50850__, new_new_n50851__,
    new_new_n50852__, new_new_n50853__, new_new_n50854__, new_new_n50855__,
    new_new_n50856__, new_new_n50857__, new_new_n50858__, new_new_n50859__,
    new_new_n50860__, new_new_n50861__, new_new_n50862__, new_new_n50863__,
    new_new_n50864__, new_new_n50865__, new_new_n50866__, new_new_n50867__,
    new_new_n50868__, new_new_n50869__, new_new_n50870__, new_new_n50871__,
    new_new_n50872__, new_new_n50873__, new_new_n50874__, new_new_n50875__,
    new_new_n50876__, new_new_n50877__, new_new_n50878__, new_new_n50879__,
    new_new_n50880__, new_new_n50881__, new_new_n50882__, new_new_n50883__,
    new_new_n50884__, new_new_n50885__, new_new_n50886__, new_new_n50887__,
    new_new_n50888__, new_new_n50889__, new_new_n50890__, new_new_n50891__,
    new_new_n50892__, new_new_n50893__, new_new_n50894__, new_new_n50895__,
    new_new_n50896__, new_new_n50897__, new_new_n50898__, new_new_n50899__,
    new_new_n50900__, new_new_n50901__, new_new_n50902__, new_new_n50903__,
    new_new_n50904__, new_new_n50905__, new_new_n50906__, new_new_n50907__,
    new_new_n50908__, new_new_n50909__, new_new_n50910__, new_new_n50911__,
    new_new_n50912__, new_new_n50913__, new_new_n50914__, new_new_n50915__,
    new_new_n50916__, new_new_n50917__, new_new_n50918__, new_new_n50919__,
    new_new_n50920__, new_new_n50921__, new_new_n50922__, new_new_n50923__,
    new_new_n50924__, new_new_n50925__, new_new_n50926__, new_new_n50927__,
    new_new_n50928__, new_new_n50929__, new_new_n50930__, new_new_n50931__,
    new_new_n50932__, new_new_n50933__, new_new_n50934__, new_new_n50935__,
    new_new_n50936__, new_new_n50937__, new_new_n50938__, new_new_n50939__,
    new_new_n50940__, new_new_n50941__, new_new_n50942__, new_new_n50943__,
    new_new_n50944__, new_new_n50945__, new_new_n50946__, new_new_n50947__,
    new_new_n50948__, new_new_n50949__, new_new_n50950__, new_new_n50951__,
    new_new_n50952__, new_new_n50953__, new_new_n50954__, new_new_n50955__,
    new_new_n50956__, new_new_n50957__, new_new_n50958__, new_new_n50959__,
    new_new_n50960__, new_new_n50961__, new_new_n50962__, new_new_n50963__,
    new_new_n50964__, new_new_n50965__, new_new_n50966__, new_new_n50967__,
    new_new_n50968__, new_new_n50969__, new_new_n50970__, new_new_n50971__,
    new_new_n50972__, new_new_n50973__, new_new_n50974__, new_new_n50975__,
    new_new_n50976__, new_new_n50977__, new_new_n50978__, new_new_n50979__,
    new_new_n50980__, new_new_n50981__, new_new_n50982__, new_new_n50983__,
    new_new_n50984__, new_new_n50985__, new_new_n50986__, new_new_n50987__,
    new_new_n50988__, new_new_n50989__, new_new_n50990__, new_new_n50991__,
    new_new_n50992__, new_new_n50993__, new_new_n50994__, new_new_n50995__,
    new_new_n50996__, new_new_n50997__, new_new_n50998__, new_new_n50999__,
    new_new_n51000__, new_new_n51001__, new_new_n51002__, new_new_n51003__,
    new_new_n51004__, new_new_n51005__, new_new_n51006__, new_new_n51007__,
    new_new_n51008__, new_new_n51009__, new_new_n51010__, new_new_n51011__,
    new_new_n51012__, new_new_n51013__, new_new_n51014__, new_new_n51015__,
    new_new_n51016__, new_new_n51017__, new_new_n51018__, new_new_n51019__,
    new_new_n51020__, new_new_n51021__, new_new_n51022__, new_new_n51023__,
    new_new_n51024__, new_new_n51025__, new_new_n51026__, new_new_n51027__,
    new_new_n51028__, new_new_n51029__, new_new_n51030__, new_new_n51031__,
    new_new_n51032__, new_new_n51033__, new_new_n51034__, new_new_n51035__,
    new_new_n51036__, new_new_n51037__, new_new_n51038__, new_new_n51039__,
    new_new_n51040__, new_new_n51041__, new_new_n51042__, new_new_n51043__,
    new_new_n51044__, new_new_n51045__, new_new_n51046__, new_new_n51047__,
    new_new_n51048__, new_new_n51049__, new_new_n51050__, new_new_n51051__,
    new_new_n51052__, new_new_n51053__, new_new_n51054__, new_new_n51055__,
    new_new_n51056__, new_new_n51057__, new_new_n51058__, new_new_n51059__,
    new_new_n51060__, new_new_n51061__, new_new_n51062__, new_new_n51063__,
    new_new_n51064__, new_new_n51065__, new_new_n51066__, new_new_n51067__,
    new_new_n51068__, new_new_n51069__, new_new_n51070__, new_new_n51071__,
    new_new_n51072__, new_new_n51073__, new_new_n51074__, new_new_n51075__,
    new_new_n51076__, new_new_n51077__, new_new_n51078__, new_new_n51079__,
    new_new_n51080__, new_new_n51081__, new_new_n51082__, new_new_n51083__,
    new_new_n51084__, new_new_n51085__, new_new_n51086__, new_new_n51087__,
    new_new_n51088__, new_new_n51089__, new_new_n51090__, new_new_n51091__,
    new_new_n51092__, new_new_n51093__, new_new_n51094__, new_new_n51095__,
    new_new_n51096__, new_new_n51097__, new_new_n51098__, new_new_n51099__,
    new_new_n51100__, new_new_n51101__, new_new_n51102__, new_new_n51103__,
    new_new_n51104__, new_new_n51105__, new_new_n51106__, new_new_n51107__,
    new_new_n51108__, new_new_n51109__, new_new_n51110__, new_new_n51111__,
    new_new_n51112__, new_new_n51113__, new_new_n51114__, new_new_n51115__,
    new_new_n51116__, new_new_n51117__, new_new_n51118__, new_new_n51119__,
    new_new_n51120__, new_new_n51121__, new_new_n51123__, new_new_n51124__,
    new_new_n51125__, new_new_n51126__, new_new_n51127__, new_new_n51128__,
    new_new_n51129__, new_new_n51130__, new_new_n51131__, new_new_n51134__,
    new_new_n51135__, new_new_n51136__, new_new_n51137__, new_new_n51138__,
    new_new_n51139__, new_new_n51140__, new_new_n51141__, new_new_n51142__,
    new_new_n51143__, new_new_n51144__, new_new_n51145__, new_new_n51146__,
    new_new_n51151__, new_new_n51156__, new_new_n51158__, new_new_n51160__,
    new_new_n51161__, new_new_n51162__, new_new_n51164__, new_new_n51165__,
    new_new_n51166__, new_new_n51169__, new_new_n51174__, new_new_n51175__,
    new_new_n51176__, new_new_n51177__, new_new_n51178__, new_new_n51179__,
    new_new_n51181__, new_new_n51183__, new_new_n51184__, new_new_n51185__,
    new_new_n51186__, new_new_n51187__, new_new_n51189__, new_new_n51190__,
    new_new_n51191__, new_new_n51192__, new_new_n51193__, new_new_n51194__,
    new_new_n51195__, new_new_n51196__, new_new_n51197__, new_new_n51198__,
    new_new_n51199__, new_new_n51201__, new_new_n51202__, new_new_n51203__,
    new_new_n51204__, new_new_n51205__, new_new_n51206__, new_new_n51207__,
    new_new_n51208__, new_new_n51209__, new_new_n51210__, new_new_n51211__,
    new_new_n51212__, new_new_n51213__, new_new_n51214__, new_new_n51215__,
    new_new_n51216__, new_new_n51217__, new_new_n51218__, new_new_n51219__,
    new_new_n51220__, new_new_n51221__, new_new_n51222__, new_new_n51223__,
    new_new_n51224__, new_new_n51228__, new_new_n51229__, new_new_n51230__,
    new_new_n51234__, new_new_n51236__, new_new_n51237__, new_new_n51239__,
    new_new_n51240__, new_new_n51241__, new_new_n51243__, new_new_n51245__,
    new_new_n51246__, new_new_n51247__, new_new_n51249__, new_new_n51250__,
    new_new_n51252__, new_new_n51254__, new_new_n51255__, new_new_n51256__,
    new_new_n51257__, new_new_n51258__, new_new_n51259__, new_new_n51260__,
    new_new_n51261__, new_new_n51262__, new_new_n51264__, new_new_n51265__,
    new_new_n51266__, new_new_n51267__, new_new_n51268__, new_new_n51269__,
    new_new_n51270__, new_new_n51271__, new_new_n51272__, new_new_n51274__,
    new_new_n51275__, new_new_n51276__, new_new_n51277__, new_new_n51280__,
    new_new_n51281__, new_new_n51282__, new_new_n51283__, new_new_n51284__,
    new_new_n51285__, new_new_n51286__, new_new_n51287__, new_new_n51288__,
    new_new_n51289__, new_new_n51290__, new_new_n51291__, new_new_n51292__,
    new_new_n51293__, new_new_n51294__, new_new_n51295__, new_new_n51296__,
    new_new_n51297__, new_new_n51298__, new_new_n51300__, new_new_n51301__,
    new_new_n51302__, new_new_n51304__, new_new_n51306__, new_new_n51307__,
    new_new_n51308__, new_new_n51309__, new_new_n51310__, new_new_n51311__,
    new_new_n51312__, new_new_n51314__, new_new_n51315__, new_new_n51316__,
    new_new_n51317__, new_new_n51318__, new_new_n51320__, new_new_n51321__,
    new_new_n51322__, new_new_n51323__, new_new_n51324__, new_new_n51326__,
    new_new_n51327__, new_new_n51328__, new_new_n51329__, new_new_n51330__,
    new_new_n51331__, new_new_n51332__, new_new_n51333__, new_new_n51334__,
    new_new_n51335__, new_new_n51336__, new_new_n51337__, new_new_n51338__,
    new_new_n51340__, new_new_n51341__, new_new_n51342__, new_new_n51343__,
    new_new_n51344__, new_new_n51345__, new_new_n51346__, new_new_n51347__,
    new_new_n51348__, new_new_n51349__, new_new_n51351__, new_new_n51352__,
    new_new_n51353__, new_new_n51355__, new_new_n51356__, new_new_n51357__,
    new_new_n51358__, new_new_n51359__, new_new_n51360__, new_new_n51361__,
    new_new_n51362__, new_new_n51363__, new_new_n51364__, new_new_n51365__,
    new_new_n51366__, new_new_n51367__, new_new_n51368__, new_new_n51369__,
    new_new_n51370__, new_new_n51371__, new_new_n51372__, new_new_n51373__,
    new_new_n51374__, new_new_n51375__, new_new_n51376__, new_new_n51377__,
    new_new_n51378__, new_new_n51379__, new_new_n51380__, new_new_n51381__,
    new_new_n51382__, new_new_n51383__, new_new_n51384__, new_new_n51385__,
    new_new_n51386__, new_new_n51387__, new_new_n51388__, new_new_n51389__,
    new_new_n51390__, new_new_n51391__, new_new_n51392__, new_new_n51393__,
    new_new_n51394__, new_new_n51395__, new_new_n51396__, new_new_n51397__,
    new_new_n51398__, new_new_n51399__, new_new_n51400__, new_new_n51401__,
    new_new_n51402__, new_new_n51403__, new_new_n51404__, new_new_n51405__,
    new_new_n51406__, new_new_n51407__, new_new_n51408__, new_new_n51409__,
    new_new_n51410__, new_new_n51411__, new_new_n51412__, new_new_n51413__,
    new_new_n51414__, new_new_n51415__, new_new_n51416__, new_new_n51417__,
    new_new_n51418__, new_new_n51419__, new_new_n51420__, new_new_n51421__,
    new_new_n51422__, new_new_n51423__, new_new_n51424__, new_new_n51425__,
    new_new_n51426__, new_new_n51427__, new_new_n51428__, new_new_n51429__,
    new_new_n51430__, new_new_n51431__, new_new_n51432__, new_new_n51433__,
    new_new_n51434__, new_new_n51435__, new_new_n51436__, new_new_n51437__,
    new_new_n51438__, new_new_n51439__, new_new_n51440__, new_new_n51441__,
    new_new_n51442__, new_new_n51443__, new_new_n51444__, new_new_n51445__,
    new_new_n51446__, new_new_n51447__, new_new_n51448__, new_new_n51449__,
    new_new_n51450__, new_new_n51453__, new_new_n51454__, new_new_n51455__,
    new_new_n51457__, new_new_n51458__, new_new_n51459__, new_new_n51460__,
    new_new_n51461__, new_new_n51462__, new_new_n51464__, new_new_n51465__,
    new_new_n51466__, new_new_n51468__, new_new_n51469__, new_new_n51470__,
    new_new_n51472__, new_new_n51473__, new_new_n51474__, new_new_n51476__,
    new_new_n51477__, new_new_n51478__, new_new_n51480__, new_new_n51481__,
    new_new_n51482__, new_new_n51484__, new_new_n51485__, new_new_n51486__,
    new_new_n51488__, new_new_n51489__, new_new_n51490__, new_new_n51492__,
    new_new_n51493__, new_new_n51494__, new_new_n51496__, new_new_n51497__,
    new_new_n51498__, new_new_n51500__, new_new_n51501__, new_new_n51502__,
    new_new_n51510__, new_new_n51511__, new_new_n51512__, new_new_n51513__,
    new_new_n51514__, new_new_n51515__, new_new_n51516__, new_new_n51517__,
    new_new_n51518__, new_new_n51520__, new_new_n51521__, new_new_n51522__,
    new_new_n51523__, new_new_n51524__, new_new_n51526__, new_new_n51527__,
    new_new_n51528__, new_new_n51529__, new_new_n51530__, new_new_n51532__,
    new_new_n51533__, new_new_n51534__, new_new_n51535__, new_new_n51536__,
    new_new_n51538__, new_new_n51539__, new_new_n51540__, new_new_n51541__,
    new_new_n51543__, new_new_n51544__, new_new_n51545__, new_new_n51546__,
    new_new_n51547__, new_new_n51549__, new_new_n51550__, new_new_n51551__,
    new_new_n51552__, new_new_n51553__, new_new_n51554__, new_new_n51555__,
    new_new_n51557__, new_new_n51558__, new_new_n51559__, new_new_n51560__,
    new_new_n51561__, new_new_n51562__, new_new_n51563__, new_new_n51564__,
    new_new_n51565__, new_new_n51566__, new_new_n51567__, new_new_n51568__,
    new_new_n51569__, new_new_n51570__, new_new_n51571__, new_new_n51572__,
    new_new_n51574__, new_new_n51575__, new_new_n51576__, new_new_n51577__,
    new_new_n51578__, new_new_n51579__, new_new_n51581__, new_new_n51582__,
    new_new_n51583__, new_new_n51584__, new_new_n51586__, new_new_n51587__,
    new_new_n51588__, new_new_n51589__, new_new_n51590__, new_new_n51591__,
    new_new_n51592__, new_new_n51593__, new_new_n51594__, new_new_n51595__,
    new_new_n51596__, new_new_n51597__, new_new_n51598__, new_new_n51599__,
    new_new_n51600__, new_new_n51601__, new_new_n51602__, new_new_n51603__,
    new_new_n51604__, new_new_n51605__, new_new_n51606__, new_new_n51607__,
    new_new_n51608__, new_new_n51609__, new_new_n51610__, new_new_n51611__,
    new_new_n51612__, new_new_n51613__, new_new_n51614__, new_new_n51615__,
    new_new_n51616__, new_new_n51617__, new_new_n51618__, new_new_n51620__,
    new_new_n51621__, new_new_n51622__, new_new_n51623__, new_new_n51624__,
    new_new_n51625__, new_new_n51626__, new_new_n51627__, new_new_n51628__,
    new_new_n51629__, new_new_n51631__, new_new_n51632__, new_new_n51633__,
    new_new_n51634__, new_new_n51635__, new_new_n51636__, new_new_n51637__,
    new_new_n51638__, new_new_n51639__, new_new_n51640__, new_new_n51641__,
    new_new_n51642__, new_new_n51643__, new_new_n51644__, new_new_n51648__,
    new_new_n51649__, new_new_n51651__, new_new_n51653__, new_new_n51656__,
    new_new_n51658__, new_new_n51660__, new_new_n51662__, new_new_n51663__,
    new_new_n51664__, new_new_n51666__, new_new_n51667__, new_new_n51670__,
    new_new_n51671__, new_new_n51673__, new_new_n51674__, new_new_n51675__,
    new_new_n51676__, new_new_n51677__, new_new_n51678__, new_new_n51679__,
    new_new_n51682__, new_new_n51684__, new_new_n51686__, new_new_n51688__,
    new_new_n51689__, new_new_n51690__, new_new_n51691__, new_new_n51692__,
    new_new_n51693__, new_new_n51694__, new_new_n51695__, new_new_n51696__,
    new_new_n51698__, new_new_n51699__, new_new_n51700__, new_new_n51701__,
    new_new_n51702__, new_new_n51703__, new_new_n51706__, new_new_n51707__,
    new_new_n51711__, new_new_n51712__, new_new_n51713__, new_new_n51714__,
    new_new_n51715__, new_new_n51716__, new_new_n51717__, new_new_n51718__,
    new_new_n51719__, new_new_n51722__, new_new_n51725__, new_new_n51726__,
    new_new_n51727__, new_new_n51729__, new_new_n51730__, new_new_n51731__,
    new_new_n51733__, new_new_n51735__, new_new_n51736__, new_new_n51737__,
    new_new_n51738__, new_new_n51739__, new_new_n51740__, new_new_n51741__,
    new_new_n51742__, new_new_n51743__, new_new_n51744__, new_new_n51745__,
    new_new_n51747__, new_new_n51748__, new_new_n51751__, new_new_n51752__,
    new_new_n51753__, new_new_n51754__, new_new_n51755__, new_new_n51756__,
    new_new_n51757__, new_new_n51758__, new_new_n51759__, new_new_n51760__,
    new_new_n51761__, new_new_n51762__, new_new_n51763__, new_new_n51764__,
    new_new_n51765__, new_new_n51767__, new_new_n51768__, new_new_n51769__,
    new_new_n51770__, new_new_n51771__, new_new_n51773__, new_new_n51774__,
    new_new_n51775__, new_new_n51776__, new_new_n51777__, new_new_n51778__,
    new_new_n51779__, new_new_n51780__, new_new_n51781__, new_new_n51782__,
    new_new_n51783__, new_new_n51785__, new_new_n51786__, new_new_n51787__,
    new_new_n51788__, new_new_n51789__, new_new_n51791__, new_new_n51792__,
    new_new_n51793__, new_new_n51794__, new_new_n51795__, new_new_n51796__,
    new_new_n51797__, new_new_n51798__, new_new_n51800__, new_new_n51801__,
    new_new_n51802__, new_new_n51803__, new_new_n51804__, new_new_n51806__,
    new_new_n51807__, new_new_n51808__, new_new_n51809__, new_new_n51810__,
    new_new_n51811__, new_new_n51812__, new_new_n51813__, new_new_n51814__,
    new_new_n51815__, new_new_n51816__, new_new_n51817__, new_new_n51818__,
    new_new_n51819__, new_new_n51820__, new_new_n51821__, new_new_n51822__,
    new_new_n51823__, new_new_n51824__, new_new_n51825__, new_new_n51826__,
    new_new_n51827__, new_new_n51828__, new_new_n51829__, new_new_n51830__,
    new_new_n51831__, new_new_n51832__, new_new_n51833__, new_new_n51835__,
    new_new_n51836__, new_new_n51837__, new_new_n51838__, new_new_n51839__,
    new_new_n51840__, new_new_n51841__, new_new_n51843__, new_new_n51844__,
    new_new_n51845__, new_new_n51846__, new_new_n51847__, new_new_n51848__,
    new_new_n51849__, new_new_n51850__, new_new_n51851__, new_new_n51852__,
    new_new_n51853__, new_new_n51854__, new_new_n51856__, new_new_n51857__,
    new_new_n51858__, new_new_n51859__, new_new_n51860__, new_new_n51861__,
    new_new_n51862__, new_new_n51863__, new_new_n51864__, new_new_n51865__,
    new_new_n51866__, new_new_n51867__, new_new_n51868__, new_new_n51870__,
    new_new_n51871__, new_new_n51872__, new_new_n51873__, new_new_n51874__,
    new_new_n51875__, new_new_n51876__, new_new_n51877__, new_new_n51879__,
    new_new_n51880__, new_new_n51882__, new_new_n51883__, new_new_n51884__,
    new_new_n51885__, new_new_n51886__, new_new_n51888__, new_new_n51889__,
    new_new_n51890__, new_new_n51891__, new_new_n51892__, new_new_n51893__,
    new_new_n51894__, new_new_n51895__, new_new_n51896__, new_new_n51898__,
    new_new_n51899__, new_new_n51900__, new_new_n51901__, new_new_n51902__,
    new_new_n51904__, new_new_n51905__, new_new_n51906__, new_new_n51907__,
    new_new_n51908__, new_new_n51909__, new_new_n51910__, new_new_n51911__,
    new_new_n51913__, new_new_n51914__, new_new_n51915__, new_new_n51916__,
    new_new_n51917__, new_new_n51919__, new_new_n51920__, new_new_n51921__,
    new_new_n51922__, new_new_n51923__, new_new_n51924__, new_new_n51925__,
    new_new_n51926__, new_new_n51927__, new_new_n51928__, new_new_n51929__,
    new_new_n51930__, new_new_n51931__, new_new_n51933__, new_new_n51934__,
    new_new_n51935__, new_new_n51936__, new_new_n51937__, new_new_n51938__,
    new_new_n51939__, new_new_n51940__, new_new_n51941__, new_new_n51942__,
    new_new_n51943__, new_new_n51944__, new_new_n51946__, new_new_n51947__,
    new_new_n51948__, new_new_n51949__, new_new_n51950__, new_new_n51951__,
    new_new_n51952__, new_new_n51953__, new_new_n51954__, new_new_n51955__,
    new_new_n51956__, new_new_n51957__, new_new_n51958__, new_new_n51960__,
    new_new_n51961__, new_new_n51962__, new_new_n51963__, new_new_n51964__,
    new_new_n51965__, new_new_n51966__, new_new_n51967__, new_new_n51969__,
    new_new_n51970__, new_new_n51972__, new_new_n51973__, new_new_n51974__,
    new_new_n51975__, new_new_n51976__, new_new_n51978__, new_new_n51979__,
    new_new_n51980__, new_new_n51981__, new_new_n51982__, new_new_n51983__,
    new_new_n51984__, new_new_n51985__, new_new_n51986__, new_new_n51988__,
    new_new_n51989__, new_new_n51990__, new_new_n51991__, new_new_n51992__,
    new_new_n51994__, new_new_n51995__, new_new_n51996__, new_new_n51997__,
    new_new_n51998__, new_new_n51999__, new_new_n52000__, new_new_n52001__,
    new_new_n52003__, new_new_n52004__, new_new_n52005__, new_new_n52006__,
    new_new_n52007__, new_new_n52009__, new_new_n52010__, new_new_n52011__,
    new_new_n52012__, new_new_n52013__, new_new_n52014__, new_new_n52015__,
    new_new_n52016__, new_new_n52017__, new_new_n52018__, new_new_n52019__,
    new_new_n52020__, new_new_n52021__, new_new_n52023__, new_new_n52024__,
    new_new_n52025__, new_new_n52026__, new_new_n52027__, new_new_n52028__,
    new_new_n52029__, new_new_n52030__, new_new_n52031__, new_new_n52032__,
    new_new_n52033__, new_new_n52034__, new_new_n52036__, new_new_n52037__,
    new_new_n52038__, new_new_n52039__, new_new_n52040__, new_new_n52041__,
    new_new_n52042__, new_new_n52043__, new_new_n52044__, new_new_n52045__,
    new_new_n52046__, new_new_n52047__, new_new_n52048__, new_new_n52050__,
    new_new_n52051__, new_new_n52052__, new_new_n52053__, new_new_n52054__,
    new_new_n52055__, new_new_n52056__, new_new_n52057__, new_new_n52059__,
    new_new_n52060__, new_new_n52062__, new_new_n52063__, new_new_n52064__,
    new_new_n52065__, new_new_n52066__, new_new_n52068__, new_new_n52069__,
    new_new_n52070__, new_new_n52071__, new_new_n52072__, new_new_n52073__,
    new_new_n52074__, new_new_n52075__, new_new_n52076__, new_new_n52078__,
    new_new_n52079__, new_new_n52080__, new_new_n52081__, new_new_n52082__,
    new_new_n52084__, new_new_n52085__, new_new_n52086__, new_new_n52087__,
    new_new_n52088__, new_new_n52089__, new_new_n52090__, new_new_n52091__,
    new_new_n52093__, new_new_n52094__, new_new_n52095__, new_new_n52096__,
    new_new_n52097__, new_new_n52099__, new_new_n52100__, new_new_n52101__,
    new_new_n52102__, new_new_n52103__, new_new_n52104__, new_new_n52105__,
    new_new_n52106__, new_new_n52107__, new_new_n52108__, new_new_n52109__,
    new_new_n52110__, new_new_n52111__, new_new_n52113__, new_new_n52114__,
    new_new_n52115__, new_new_n52116__, new_new_n52117__, new_new_n52118__,
    new_new_n52119__, new_new_n52120__, new_new_n52121__, new_new_n52122__,
    new_new_n52123__, new_new_n52124__, new_new_n52126__, new_new_n52127__,
    new_new_n52128__, new_new_n52129__, new_new_n52130__, new_new_n52131__,
    new_new_n52132__, new_new_n52133__, new_new_n52134__, new_new_n52135__,
    new_new_n52136__, new_new_n52137__, new_new_n52138__, new_new_n52140__,
    new_new_n52141__, new_new_n52142__, new_new_n52143__, new_new_n52144__,
    new_new_n52145__, new_new_n52146__, new_new_n52147__, new_new_n52149__,
    new_new_n52150__, new_new_n52152__, new_new_n52153__, new_new_n52154__,
    new_new_n52155__, new_new_n52156__, new_new_n52158__, new_new_n52159__,
    new_new_n52160__, new_new_n52161__, new_new_n52162__, new_new_n52163__,
    new_new_n52164__, new_new_n52165__, new_new_n52166__, new_new_n52168__,
    new_new_n52169__, new_new_n52170__, new_new_n52171__, new_new_n52172__,
    new_new_n52174__, new_new_n52175__, new_new_n52176__, new_new_n52177__,
    new_new_n52178__, new_new_n52179__, new_new_n52180__, new_new_n52181__,
    new_new_n52183__, new_new_n52184__, new_new_n52185__, new_new_n52186__,
    new_new_n52187__, new_new_n52189__, new_new_n52190__, new_new_n52191__,
    new_new_n52192__, new_new_n52193__, new_new_n52194__, new_new_n52195__,
    new_new_n52196__, new_new_n52197__, new_new_n52198__, new_new_n52199__,
    new_new_n52200__, new_new_n52201__, new_new_n52203__, new_new_n52204__,
    new_new_n52205__, new_new_n52206__, new_new_n52207__, new_new_n52208__,
    new_new_n52209__, new_new_n52210__, new_new_n52211__, new_new_n52212__,
    new_new_n52213__, new_new_n52214__, new_new_n52216__, new_new_n52217__,
    new_new_n52218__, new_new_n52219__, new_new_n52220__, new_new_n52221__,
    new_new_n52222__, new_new_n52223__, new_new_n52224__, new_new_n52225__,
    new_new_n52226__, new_new_n52227__, new_new_n52228__, new_new_n52230__,
    new_new_n52231__, new_new_n52232__, new_new_n52233__, new_new_n52234__,
    new_new_n52235__, new_new_n52236__, new_new_n52237__, new_new_n52240__,
    new_new_n52241__, new_new_n52242__, new_new_n52243__, new_new_n52244__,
    new_new_n52245__, new_new_n52246__, new_new_n52248__, new_new_n52249__,
    new_new_n52250__, new_new_n52251__, new_new_n52252__, new_new_n52253__,
    new_new_n52254__, new_new_n52255__, new_new_n52256__, new_new_n52257__,
    new_new_n52258__, new_new_n52259__, new_new_n52260__, new_new_n52261__,
    new_new_n52262__, new_new_n52263__, new_new_n52264__, new_new_n52265__,
    new_new_n52267__, new_new_n52268__, new_new_n52269__, new_new_n52270__,
    new_new_n52271__, new_new_n52272__, new_new_n52273__, new_new_n52274__,
    new_new_n52275__, new_new_n52276__, new_new_n52277__, new_new_n52278__,
    new_new_n52280__, new_new_n52281__, new_new_n52282__, new_new_n52283__,
    new_new_n52284__, new_new_n52285__, new_new_n52286__, new_new_n52287__,
    new_new_n52288__, new_new_n52289__, new_new_n52290__, new_new_n52291__,
    new_new_n52292__, new_new_n52294__, new_new_n52295__, new_new_n52296__,
    new_new_n52297__, new_new_n52298__, new_new_n52300__, new_new_n52301__,
    new_new_n52302__, new_new_n52303__, new_new_n52304__, new_new_n52305__,
    new_new_n52306__, new_new_n52307__, new_new_n52308__, new_new_n52309__,
    new_new_n52310__, new_new_n52311__, new_new_n52312__, new_new_n52313__,
    new_new_n52314__, new_new_n52315__, new_new_n52316__, new_new_n52317__,
    new_new_n52318__, new_new_n52319__, new_new_n52320__, new_new_n52321__,
    new_new_n52322__, new_new_n52323__, new_new_n52324__, new_new_n52325__,
    new_new_n52326__, new_new_n52327__, new_new_n52330__, new_new_n52331__,
    new_new_n52332__, new_new_n52333__, new_new_n52334__, new_new_n52335__,
    new_new_n52336__, new_new_n52337__, new_new_n52338__, new_new_n52339__,
    new_new_n52340__, new_new_n52341__, new_new_n52342__, new_new_n52343__,
    new_new_n52344__, new_new_n52345__, new_new_n52346__, new_new_n52347__,
    new_new_n52348__, new_new_n52349__, new_new_n52350__, new_new_n52351__,
    new_new_n52352__, new_new_n52353__, new_new_n52354__, new_new_n52355__,
    new_new_n52356__, new_new_n52357__, new_new_n52358__, new_new_n52359__,
    new_new_n52360__, new_new_n52361__, new_new_n52362__, new_new_n52363__,
    new_new_n52364__, new_new_n52365__, new_new_n52366__, new_new_n52367__,
    new_new_n52368__, new_new_n52369__, new_new_n52370__, new_new_n52371__,
    new_new_n52372__, new_new_n52373__, new_new_n52374__, new_new_n52375__,
    new_new_n52376__, new_new_n52377__, new_new_n52378__, new_new_n52379__,
    new_new_n52380__, new_new_n52381__, new_new_n52382__, new_new_n52383__,
    new_new_n52384__, new_new_n52385__, new_new_n52386__, new_new_n52387__,
    new_new_n52388__, new_new_n52389__, new_new_n52390__, new_new_n52391__,
    new_new_n52392__, new_new_n52393__, new_new_n52394__, new_new_n52395__,
    new_new_n52396__, new_new_n52397__, new_new_n52398__, new_new_n52399__,
    new_new_n52400__, new_new_n52401__, new_new_n52402__, new_new_n52403__,
    new_new_n52404__, new_new_n52405__, new_new_n52406__, new_new_n52407__,
    new_new_n52408__, new_new_n52409__, new_new_n52410__, new_new_n52411__,
    new_new_n52412__, new_new_n52413__, new_new_n52414__, new_new_n52415__,
    new_new_n52416__, new_new_n52417__, new_new_n52418__, new_new_n52419__,
    new_new_n52420__, new_new_n52421__, new_new_n52422__, new_new_n52423__,
    new_new_n52424__, new_new_n52425__, new_new_n52426__, new_new_n52427__,
    new_new_n52428__, new_new_n52429__, new_new_n52430__, new_new_n52431__,
    new_new_n52432__, new_new_n52433__, new_new_n52434__, new_new_n52435__,
    new_new_n52436__, new_new_n52437__, new_new_n52438__, new_new_n52439__,
    new_new_n52440__, new_new_n52441__, new_new_n52442__, new_new_n52443__,
    new_new_n52444__, new_new_n52445__, new_new_n52446__, new_new_n52447__,
    new_new_n52448__, new_new_n52449__, new_new_n52450__, new_new_n52451__,
    new_new_n52452__, new_new_n52453__, new_new_n52454__, new_new_n52455__,
    new_new_n52456__, new_new_n52457__, new_new_n52458__, new_new_n52459__,
    new_new_n52460__, new_new_n52461__, new_new_n52462__, new_new_n52463__,
    new_new_n52464__, new_new_n52465__, new_new_n52466__, new_new_n52467__,
    new_new_n52468__, new_new_n52469__, new_new_n52470__, new_new_n52471__,
    new_new_n52472__, new_new_n52473__, new_new_n52474__, new_new_n52475__,
    new_new_n52476__, new_new_n52477__, new_new_n52478__, new_new_n52479__,
    new_new_n52480__, new_new_n52481__, new_new_n52482__, new_new_n52483__,
    new_new_n52484__, new_new_n52485__, new_new_n52486__, new_new_n52487__,
    new_new_n52488__, new_new_n52489__, new_new_n52490__, new_new_n52491__,
    new_new_n52492__, new_new_n52493__, new_new_n52494__, new_new_n52495__,
    new_new_n52496__, new_new_n52497__, new_new_n52498__, new_new_n52499__,
    new_new_n52500__, new_new_n52501__, new_new_n52502__, new_new_n52503__,
    new_new_n52504__, new_new_n52505__, new_new_n52506__, new_new_n52507__,
    new_new_n52508__, new_new_n52509__, new_new_n52510__, new_new_n52511__,
    new_new_n52512__, new_new_n52513__, new_new_n52514__, new_new_n52515__,
    new_new_n52516__, new_new_n52517__, new_new_n52518__, new_new_n52519__,
    new_new_n52520__, new_new_n52521__, new_new_n52522__, new_new_n52523__,
    new_new_n52524__, new_new_n52525__, new_new_n52526__, new_new_n52527__,
    new_new_n52528__, new_new_n52529__, new_new_n52530__, new_new_n52531__,
    new_new_n52532__, new_new_n52533__, new_new_n52534__, new_new_n52535__,
    new_new_n52536__, new_new_n52537__, new_new_n52538__, new_new_n52539__,
    new_new_n52540__, new_new_n52542__, new_new_n52543__, new_new_n52544__,
    new_new_n52545__, new_new_n52546__, new_new_n52547__, new_new_n52548__,
    new_new_n52549__, new_new_n52550__, new_new_n52551__, new_new_n52552__,
    new_new_n52553__, new_new_n52554__, new_new_n52555__, new_new_n52556__,
    new_new_n52557__, new_new_n52558__, new_new_n52559__, new_new_n52560__,
    new_new_n52561__, new_new_n52562__, new_new_n52563__, new_new_n52564__,
    new_new_n52565__, new_new_n52566__, new_new_n52567__, new_new_n52568__,
    new_new_n52569__, new_new_n52570__, new_new_n52571__, new_new_n52572__,
    new_new_n52573__, new_new_n52574__, new_new_n52575__, new_new_n52576__,
    new_new_n52577__, new_new_n52578__, new_new_n52579__, new_new_n52580__,
    new_new_n52581__, new_new_n52582__, new_new_n52583__, new_new_n52584__,
    new_new_n52585__, new_new_n52586__, new_new_n52587__, new_new_n52588__,
    new_new_n52589__, new_new_n52590__, new_new_n52591__, new_new_n52592__,
    new_new_n52593__, new_new_n52594__, new_new_n52596__, new_new_n52597__,
    new_new_n52598__, new_new_n52599__, new_new_n52600__, new_new_n52601__,
    new_new_n52602__, new_new_n52603__, new_new_n52604__, new_new_n52606__,
    new_new_n52607__, new_new_n52608__, new_new_n52609__, new_new_n52610__,
    new_new_n52611__, new_new_n52612__, new_new_n52613__, new_new_n52614__,
    new_new_n52615__, new_new_n52616__, new_new_n52617__, new_new_n52618__,
    new_new_n52619__, new_new_n52620__, new_new_n52621__, new_new_n52622__,
    new_new_n52623__, new_new_n52624__, new_new_n52625__, new_new_n52626__,
    new_new_n52627__, new_new_n52628__, new_new_n52629__, new_new_n52630__,
    new_new_n52631__, new_new_n52632__, new_new_n52633__, new_new_n52634__,
    new_new_n52635__, new_new_n52636__, new_new_n52637__, new_new_n52638__,
    new_new_n52639__, new_new_n52640__, new_new_n52641__, new_new_n52642__,
    new_new_n52643__, new_new_n52644__, new_new_n52645__, new_new_n52646__,
    new_new_n52647__, new_new_n52648__, new_new_n52649__, new_new_n52650__,
    new_new_n52651__, new_new_n52652__, new_new_n52653__, new_new_n52654__,
    new_new_n52655__, new_new_n52656__, new_new_n52658__, new_new_n52659__,
    new_new_n52660__, new_new_n52661__, new_new_n52662__, new_new_n52663__,
    new_new_n52664__, new_new_n52665__, new_new_n52666__, new_new_n52668__,
    new_new_n52669__, new_new_n52670__, new_new_n52671__, new_new_n52672__,
    new_new_n52673__, new_new_n52674__, new_new_n52675__, new_new_n52676__,
    new_new_n52677__, new_new_n52678__, new_new_n52679__, new_new_n52680__,
    new_new_n52681__, new_new_n52682__, new_new_n52683__, new_new_n52684__,
    new_new_n52685__, new_new_n52686__, new_new_n52687__, new_new_n52688__,
    new_new_n52689__, new_new_n52690__, new_new_n52691__, new_new_n52692__,
    new_new_n52693__, new_new_n52694__, new_new_n52695__, new_new_n52696__,
    new_new_n52697__, new_new_n52698__, new_new_n52699__, new_new_n52700__,
    new_new_n52701__, new_new_n52702__, new_new_n52703__, new_new_n52704__,
    new_new_n52705__, new_new_n52706__, new_new_n52707__, new_new_n52708__,
    new_new_n52709__, new_new_n52710__, new_new_n52711__, new_new_n52712__,
    new_new_n52713__, new_new_n52714__, new_new_n52715__, new_new_n52716__,
    new_new_n52717__, new_new_n52718__, new_new_n52719__, new_new_n52720__,
    new_new_n52721__, new_new_n52723__, new_new_n52724__, new_new_n52725__,
    new_new_n52726__, new_new_n52727__, new_new_n52728__, new_new_n52729__,
    new_new_n52730__, new_new_n52731__, new_new_n52733__, new_new_n52734__,
    new_new_n52735__, new_new_n52736__, new_new_n52737__, new_new_n52738__,
    new_new_n52739__, new_new_n52740__, new_new_n52741__, new_new_n52742__,
    new_new_n52743__, new_new_n52744__, new_new_n52745__, new_new_n52746__,
    new_new_n52747__, new_new_n52748__, new_new_n52749__, new_new_n52750__,
    new_new_n52751__, new_new_n52752__, new_new_n52753__, new_new_n52754__,
    new_new_n52755__, new_new_n52756__, new_new_n52757__, new_new_n52758__,
    new_new_n52759__, new_new_n52760__, new_new_n52761__, new_new_n52762__,
    new_new_n52763__, new_new_n52764__, new_new_n52765__, new_new_n52766__,
    new_new_n52767__, new_new_n52768__, new_new_n52769__, new_new_n52770__,
    new_new_n52771__, new_new_n52772__, new_new_n52773__, new_new_n52774__,
    new_new_n52775__, new_new_n52776__, new_new_n52777__, new_new_n52778__,
    new_new_n52779__, new_new_n52780__, new_new_n52781__, new_new_n52782__,
    new_new_n52783__, new_new_n52784__, new_new_n52785__, new_new_n52786__,
    new_new_n52787__, new_new_n52788__, new_new_n52789__, new_new_n52790__,
    new_new_n52791__, new_new_n52792__, new_new_n52793__, new_new_n52794__,
    new_new_n52795__, new_new_n52796__, new_new_n52797__, new_new_n52798__,
    new_new_n52799__, new_new_n52800__, new_new_n52802__, new_new_n52803__,
    new_new_n52804__, new_new_n52805__, new_new_n52806__, new_new_n52807__,
    new_new_n52808__, new_new_n52809__, new_new_n52810__, new_new_n52812__,
    new_new_n52813__, new_new_n52814__, new_new_n52815__, new_new_n52816__,
    new_new_n52817__, new_new_n52818__, new_new_n52819__, new_new_n52820__,
    new_new_n52821__, new_new_n52822__, new_new_n52823__, new_new_n52824__,
    new_new_n52825__, new_new_n52826__, new_new_n52827__, new_new_n52828__,
    new_new_n52829__, new_new_n52830__, new_new_n52831__, new_new_n52832__,
    new_new_n52833__, new_new_n52834__, new_new_n52835__, new_new_n52836__,
    new_new_n52837__, new_new_n52838__, new_new_n52839__, new_new_n52840__,
    new_new_n52841__, new_new_n52842__, new_new_n52843__, new_new_n52844__,
    new_new_n52845__, new_new_n52846__, new_new_n52847__, new_new_n52848__,
    new_new_n52849__, new_new_n52850__, new_new_n52851__, new_new_n52852__,
    new_new_n52853__, new_new_n52854__, new_new_n52855__, new_new_n52856__,
    new_new_n52857__, new_new_n52858__, new_new_n52859__, new_new_n52860__,
    new_new_n52861__, new_new_n52862__, new_new_n52863__, new_new_n52864__,
    new_new_n52865__, new_new_n52866__, new_new_n52867__, new_new_n52868__,
    new_new_n52869__, new_new_n52870__, new_new_n52871__, new_new_n52872__,
    new_new_n52873__, new_new_n52874__, new_new_n52875__, new_new_n52876__,
    new_new_n52877__, new_new_n52879__, new_new_n52880__, new_new_n52881__,
    new_new_n52882__, new_new_n52883__, new_new_n52884__, new_new_n52885__,
    new_new_n52886__, new_new_n52887__, new_new_n52889__, new_new_n52890__,
    new_new_n52891__, new_new_n52892__, new_new_n52893__, new_new_n52894__,
    new_new_n52895__, new_new_n52896__, new_new_n52897__, new_new_n52898__,
    new_new_n52899__, new_new_n52900__, new_new_n52901__, new_new_n52902__,
    new_new_n52903__, new_new_n52904__, new_new_n52905__, new_new_n52906__,
    new_new_n52907__, new_new_n52908__, new_new_n52909__, new_new_n52910__,
    new_new_n52911__, new_new_n52912__, new_new_n52913__, new_new_n52914__,
    new_new_n52915__, new_new_n52916__, new_new_n52917__, new_new_n52918__,
    new_new_n52919__, new_new_n52920__, new_new_n52921__, new_new_n52922__,
    new_new_n52923__, new_new_n52924__, new_new_n52925__, new_new_n52926__,
    new_new_n52927__, new_new_n52928__, new_new_n52929__, new_new_n52930__,
    new_new_n52931__, new_new_n52932__, new_new_n52933__, new_new_n52934__,
    new_new_n52935__, new_new_n52936__, new_new_n52937__, new_new_n52938__,
    new_new_n52939__, new_new_n52940__, new_new_n52941__, new_new_n52942__,
    new_new_n52943__, new_new_n52944__, new_new_n52945__, new_new_n52946__,
    new_new_n52947__, new_new_n52948__, new_new_n52949__, new_new_n52950__,
    new_new_n52951__, new_new_n52952__, new_new_n52953__, new_new_n52954__,
    new_new_n52955__, new_new_n52956__, new_new_n52957__, new_new_n52959__,
    new_new_n52960__, new_new_n52961__, new_new_n52962__, new_new_n52963__,
    new_new_n52964__, new_new_n52965__, new_new_n52966__, new_new_n52967__,
    new_new_n52969__, new_new_n52970__, new_new_n52971__, new_new_n52972__,
    new_new_n52973__, new_new_n52974__, new_new_n52975__, new_new_n52976__,
    new_new_n52977__, new_new_n52978__, new_new_n52979__, new_new_n52980__,
    new_new_n52981__, new_new_n52982__, new_new_n52983__, new_new_n52984__,
    new_new_n52985__, new_new_n52986__, new_new_n52987__, new_new_n52988__,
    new_new_n52989__, new_new_n52990__, new_new_n52991__, new_new_n52992__,
    new_new_n52993__, new_new_n52994__, new_new_n52995__, new_new_n52996__,
    new_new_n52997__, new_new_n52998__, new_new_n52999__, new_new_n53000__,
    new_new_n53001__, new_new_n53002__, new_new_n53003__, new_new_n53004__,
    new_new_n53005__, new_new_n53006__, new_new_n53007__, new_new_n53008__,
    new_new_n53009__, new_new_n53010__, new_new_n53011__, new_new_n53012__,
    new_new_n53013__, new_new_n53014__, new_new_n53015__, new_new_n53016__,
    new_new_n53017__, new_new_n53018__, new_new_n53019__, new_new_n53020__,
    new_new_n53021__, new_new_n53022__, new_new_n53023__, new_new_n53024__,
    new_new_n53025__, new_new_n53026__, new_new_n53027__, new_new_n53028__,
    new_new_n53029__, new_new_n53030__, new_new_n53031__, new_new_n53032__,
    new_new_n53033__, new_new_n53034__, new_new_n53035__, new_new_n53036__,
    new_new_n53037__, new_new_n53038__, new_new_n53039__, new_new_n53040__,
    new_new_n53041__, new_new_n53042__, new_new_n53043__, new_new_n53044__,
    new_new_n53045__, new_new_n53046__, new_new_n53047__, new_new_n53048__,
    new_new_n53049__, new_new_n53050__, new_new_n53051__, new_new_n53052__,
    new_new_n53053__, new_new_n53054__, new_new_n53055__, new_new_n53057__,
    new_new_n53058__, new_new_n53059__, new_new_n53060__, new_new_n53061__,
    new_new_n53062__, new_new_n53063__, new_new_n53064__, new_new_n53065__,
    new_new_n53067__, new_new_n53068__, new_new_n53069__, new_new_n53070__,
    new_new_n53071__, new_new_n53072__, new_new_n53073__, new_new_n53074__,
    new_new_n53075__, new_new_n53076__, new_new_n53077__, new_new_n53078__,
    new_new_n53079__, new_new_n53080__, new_new_n53081__, new_new_n53082__,
    new_new_n53083__, new_new_n53084__, new_new_n53085__, new_new_n53086__,
    new_new_n53087__, new_new_n53088__, new_new_n53089__, new_new_n53090__,
    new_new_n53091__, new_new_n53092__, new_new_n53093__, new_new_n53094__,
    new_new_n53095__, new_new_n53096__, new_new_n53097__, new_new_n53098__,
    new_new_n53099__, new_new_n53100__, new_new_n53101__, new_new_n53102__,
    new_new_n53103__, new_new_n53104__, new_new_n53105__, new_new_n53106__,
    new_new_n53107__, new_new_n53108__, new_new_n53109__, new_new_n53110__,
    new_new_n53111__, new_new_n53112__, new_new_n53113__, new_new_n53114__,
    new_new_n53115__, new_new_n53116__, new_new_n53117__, new_new_n53118__,
    new_new_n53119__, new_new_n53120__, new_new_n53121__, new_new_n53122__,
    new_new_n53123__, new_new_n53124__, new_new_n53125__, new_new_n53126__,
    new_new_n53127__, new_new_n53128__, new_new_n53129__, new_new_n53130__,
    new_new_n53131__, new_new_n53132__, new_new_n53133__, new_new_n53134__,
    new_new_n53135__, new_new_n53136__, new_new_n53137__, new_new_n53138__,
    new_new_n53139__, new_new_n53140__, new_new_n53141__, new_new_n53142__,
    new_new_n53143__, new_new_n53144__, new_new_n53145__, new_new_n53146__,
    new_new_n53147__, new_new_n53148__, new_new_n53149__, new_new_n53150__,
    new_new_n53151__, new_new_n53153__, new_new_n53154__, new_new_n53155__,
    new_new_n53156__, new_new_n53157__, new_new_n53158__, new_new_n53159__,
    new_new_n53160__, new_new_n53161__, new_new_n53163__, new_new_n53164__,
    new_new_n53165__, new_new_n53166__, new_new_n53167__, new_new_n53168__,
    new_new_n53169__, new_new_n53170__, new_new_n53171__, new_new_n53172__,
    new_new_n53173__, new_new_n53174__, new_new_n53175__, new_new_n53176__,
    new_new_n53177__, new_new_n53178__, new_new_n53179__, new_new_n53180__,
    new_new_n53181__, new_new_n53182__, new_new_n53183__, new_new_n53184__,
    new_new_n53185__, new_new_n53186__, new_new_n53187__, new_new_n53188__,
    new_new_n53189__, new_new_n53190__, new_new_n53191__, new_new_n53192__,
    new_new_n53193__, new_new_n53194__, new_new_n53195__, new_new_n53196__,
    new_new_n53197__, new_new_n53198__, new_new_n53199__, new_new_n53200__,
    new_new_n53201__, new_new_n53202__, new_new_n53203__, new_new_n53204__,
    new_new_n53205__, new_new_n53206__, new_new_n53207__, new_new_n53208__,
    new_new_n53209__, new_new_n53210__, new_new_n53211__, new_new_n53212__,
    new_new_n53213__, new_new_n53214__, new_new_n53215__, new_new_n53216__,
    new_new_n53217__, new_new_n53218__, new_new_n53219__, new_new_n53220__,
    new_new_n53221__, new_new_n53222__, new_new_n53223__, new_new_n53224__,
    new_new_n53225__, new_new_n53226__, new_new_n53227__, new_new_n53228__,
    new_new_n53229__, new_new_n53230__, new_new_n53231__, new_new_n53232__,
    new_new_n53233__, new_new_n53234__, new_new_n53235__, new_new_n53236__,
    new_new_n53237__, new_new_n53238__, new_new_n53239__, new_new_n53240__,
    new_new_n53241__, new_new_n53242__, new_new_n53243__, new_new_n53244__,
    new_new_n53245__, new_new_n53246__, new_new_n53247__, new_new_n53248__,
    new_new_n53249__, new_new_n53250__, new_new_n53251__, new_new_n53252__,
    new_new_n53253__, new_new_n53254__, new_new_n53255__, new_new_n53256__,
    new_new_n53257__, new_new_n53258__, new_new_n53259__, new_new_n53260__,
    new_new_n53262__, new_new_n53263__, new_new_n53264__, new_new_n53265__,
    new_new_n53266__, new_new_n53267__, new_new_n53268__, new_new_n53269__,
    new_new_n53270__, new_new_n53272__, new_new_n53273__, new_new_n53274__,
    new_new_n53275__, new_new_n53276__, new_new_n53277__, new_new_n53278__,
    new_new_n53279__, new_new_n53280__, new_new_n53281__, new_new_n53282__,
    new_new_n53283__, new_new_n53284__, new_new_n53285__, new_new_n53286__,
    new_new_n53287__, new_new_n53288__, new_new_n53289__, new_new_n53290__,
    new_new_n53291__, new_new_n53292__, new_new_n53293__, new_new_n53294__,
    new_new_n53295__, new_new_n53296__, new_new_n53297__, new_new_n53298__,
    new_new_n53299__, new_new_n53300__, new_new_n53301__, new_new_n53302__,
    new_new_n53303__, new_new_n53304__, new_new_n53305__, new_new_n53306__,
    new_new_n53307__, new_new_n53308__, new_new_n53309__, new_new_n53310__,
    new_new_n53311__, new_new_n53312__, new_new_n53313__, new_new_n53314__,
    new_new_n53315__, new_new_n53316__, new_new_n53317__, new_new_n53318__,
    new_new_n53319__, new_new_n53320__, new_new_n53321__, new_new_n53322__,
    new_new_n53323__, new_new_n53324__, new_new_n53325__, new_new_n53326__,
    new_new_n53327__, new_new_n53328__, new_new_n53329__, new_new_n53330__,
    new_new_n53331__, new_new_n53332__, new_new_n53333__, new_new_n53334__,
    new_new_n53335__, new_new_n53336__, new_new_n53337__, new_new_n53338__,
    new_new_n53339__, new_new_n53340__, new_new_n53341__, new_new_n53342__,
    new_new_n53343__, new_new_n53344__, new_new_n53345__, new_new_n53346__,
    new_new_n53347__, new_new_n53348__, new_new_n53349__, new_new_n53350__,
    new_new_n53351__, new_new_n53352__, new_new_n53353__, new_new_n53354__,
    new_new_n53355__, new_new_n53356__, new_new_n53357__, new_new_n53358__,
    new_new_n53359__, new_new_n53360__, new_new_n53361__, new_new_n53362__,
    new_new_n53363__, new_new_n53364__, new_new_n53365__, new_new_n53366__,
    new_new_n53367__, new_new_n53368__, new_new_n53369__, new_new_n53370__,
    new_new_n53371__, new_new_n53372__, new_new_n53373__, new_new_n53374__,
    new_new_n53375__, new_new_n53376__, new_new_n53377__, new_new_n53378__,
    new_new_n53379__, new_new_n53380__, new_new_n53381__, new_new_n53382__,
    new_new_n53383__, new_new_n53384__, new_new_n53386__, new_new_n53387__,
    new_new_n53388__, new_new_n53389__, new_new_n53390__, new_new_n53391__,
    new_new_n53392__, new_new_n53393__, new_new_n53394__, new_new_n53396__,
    new_new_n53397__, new_new_n53398__, new_new_n53399__, new_new_n53400__,
    new_new_n53401__, new_new_n53402__, new_new_n53403__, new_new_n53404__,
    new_new_n53405__, new_new_n53406__, new_new_n53407__, new_new_n53408__,
    new_new_n53409__, new_new_n53410__, new_new_n53411__, new_new_n53412__,
    new_new_n53413__, new_new_n53414__, new_new_n53415__, new_new_n53416__,
    new_new_n53417__, new_new_n53418__, new_new_n53419__, new_new_n53420__,
    new_new_n53421__, new_new_n53422__, new_new_n53423__, new_new_n53424__,
    new_new_n53425__, new_new_n53426__, new_new_n53427__, new_new_n53428__,
    new_new_n53429__, new_new_n53430__, new_new_n53431__, new_new_n53432__,
    new_new_n53433__, new_new_n53434__, new_new_n53435__, new_new_n53436__,
    new_new_n53437__, new_new_n53438__, new_new_n53439__, new_new_n53440__,
    new_new_n53441__, new_new_n53442__, new_new_n53443__, new_new_n53444__,
    new_new_n53445__, new_new_n53446__, new_new_n53447__, new_new_n53448__,
    new_new_n53449__, new_new_n53450__, new_new_n53451__, new_new_n53452__,
    new_new_n53453__, new_new_n53454__, new_new_n53455__, new_new_n53456__,
    new_new_n53457__, new_new_n53458__, new_new_n53459__, new_new_n53460__,
    new_new_n53461__, new_new_n53462__, new_new_n53463__, new_new_n53464__,
    new_new_n53465__, new_new_n53466__, new_new_n53467__, new_new_n53468__,
    new_new_n53469__, new_new_n53470__, new_new_n53471__, new_new_n53472__,
    new_new_n53473__, new_new_n53474__, new_new_n53475__, new_new_n53476__,
    new_new_n53477__, new_new_n53478__, new_new_n53479__, new_new_n53480__,
    new_new_n53481__, new_new_n53482__, new_new_n53483__, new_new_n53484__,
    new_new_n53485__, new_new_n53486__, new_new_n53487__, new_new_n53488__,
    new_new_n53489__, new_new_n53490__, new_new_n53491__, new_new_n53492__,
    new_new_n53493__, new_new_n53494__, new_new_n53495__, new_new_n53496__,
    new_new_n53497__, new_new_n53498__, new_new_n53499__, new_new_n53500__,
    new_new_n53501__, new_new_n53502__, new_new_n53503__, new_new_n53504__,
    new_new_n53505__, new_new_n53506__, new_new_n53508__, new_new_n53509__,
    new_new_n53510__, new_new_n53511__, new_new_n53512__, new_new_n53513__,
    new_new_n53514__, new_new_n53515__, new_new_n53516__, new_new_n53518__,
    new_new_n53519__, new_new_n53520__, new_new_n53521__, new_new_n53522__,
    new_new_n53523__, new_new_n53524__, new_new_n53525__, new_new_n53526__,
    new_new_n53527__, new_new_n53528__, new_new_n53529__, new_new_n53530__,
    new_new_n53531__, new_new_n53532__, new_new_n53533__, new_new_n53534__,
    new_new_n53535__, new_new_n53536__, new_new_n53537__, new_new_n53538__,
    new_new_n53539__, new_new_n53540__, new_new_n53541__, new_new_n53542__,
    new_new_n53543__, new_new_n53544__, new_new_n53545__, new_new_n53546__,
    new_new_n53547__, new_new_n53548__, new_new_n53549__, new_new_n53550__,
    new_new_n53551__, new_new_n53552__, new_new_n53553__, new_new_n53554__,
    new_new_n53555__, new_new_n53556__, new_new_n53557__, new_new_n53558__,
    new_new_n53559__, new_new_n53560__, new_new_n53561__, new_new_n53562__,
    new_new_n53563__, new_new_n53564__, new_new_n53565__, new_new_n53566__,
    new_new_n53567__, new_new_n53568__, new_new_n53569__, new_new_n53570__,
    new_new_n53571__, new_new_n53572__, new_new_n53573__, new_new_n53574__,
    new_new_n53575__, new_new_n53576__, new_new_n53577__, new_new_n53578__,
    new_new_n53579__, new_new_n53580__, new_new_n53581__, new_new_n53582__,
    new_new_n53583__, new_new_n53584__, new_new_n53585__, new_new_n53586__,
    new_new_n53587__, new_new_n53588__, new_new_n53589__, new_new_n53590__,
    new_new_n53591__, new_new_n53592__, new_new_n53593__, new_new_n53594__,
    new_new_n53595__, new_new_n53596__, new_new_n53597__, new_new_n53598__,
    new_new_n53599__, new_new_n53600__, new_new_n53601__, new_new_n53602__,
    new_new_n53603__, new_new_n53604__, new_new_n53605__, new_new_n53606__,
    new_new_n53607__, new_new_n53608__, new_new_n53609__, new_new_n53610__,
    new_new_n53611__, new_new_n53612__, new_new_n53613__, new_new_n53614__,
    new_new_n53615__, new_new_n53616__, new_new_n53617__, new_new_n53618__,
    new_new_n53619__, new_new_n53620__, new_new_n53621__, new_new_n53622__,
    new_new_n53623__, new_new_n53624__, new_new_n53625__, new_new_n53626__,
    new_new_n53627__, new_new_n53628__, new_new_n53629__, new_new_n53630__,
    new_new_n53631__, new_new_n53633__, new_new_n53634__, new_new_n53635__,
    new_new_n53636__, new_new_n53637__, new_new_n53638__, new_new_n53639__,
    new_new_n53640__, new_new_n53641__, new_new_n53643__, new_new_n53644__,
    new_new_n53645__, new_new_n53646__, new_new_n53647__, new_new_n53648__,
    new_new_n53649__, new_new_n53650__, new_new_n53651__, new_new_n53652__,
    new_new_n53653__, new_new_n53654__, new_new_n53655__, new_new_n53656__,
    new_new_n53657__, new_new_n53658__, new_new_n53659__, new_new_n53660__,
    new_new_n53661__, new_new_n53662__, new_new_n53663__, new_new_n53664__,
    new_new_n53665__, new_new_n53666__, new_new_n53667__, new_new_n53668__,
    new_new_n53669__, new_new_n53670__, new_new_n53671__, new_new_n53672__,
    new_new_n53673__, new_new_n53674__, new_new_n53675__, new_new_n53676__,
    new_new_n53677__, new_new_n53678__, new_new_n53679__, new_new_n53680__,
    new_new_n53681__, new_new_n53682__, new_new_n53683__, new_new_n53684__,
    new_new_n53685__, new_new_n53686__, new_new_n53687__, new_new_n53688__,
    new_new_n53689__, new_new_n53690__, new_new_n53691__, new_new_n53692__,
    new_new_n53693__, new_new_n53694__, new_new_n53695__, new_new_n53696__,
    new_new_n53697__, new_new_n53698__, new_new_n53699__, new_new_n53700__,
    new_new_n53701__, new_new_n53702__, new_new_n53703__, new_new_n53704__,
    new_new_n53705__, new_new_n53706__, new_new_n53707__, new_new_n53708__,
    new_new_n53709__, new_new_n53710__, new_new_n53711__, new_new_n53712__,
    new_new_n53713__, new_new_n53714__, new_new_n53715__, new_new_n53716__,
    new_new_n53717__, new_new_n53718__, new_new_n53719__, new_new_n53720__,
    new_new_n53721__, new_new_n53722__, new_new_n53723__, new_new_n53724__,
    new_new_n53725__, new_new_n53726__, new_new_n53727__, new_new_n53728__,
    new_new_n53729__, new_new_n53730__, new_new_n53731__, new_new_n53732__,
    new_new_n53733__, new_new_n53734__, new_new_n53735__, new_new_n53736__,
    new_new_n53737__, new_new_n53738__, new_new_n53739__, new_new_n53740__,
    new_new_n53741__, new_new_n53742__, new_new_n53743__, new_new_n53744__,
    new_new_n53745__, new_new_n53746__, new_new_n53747__, new_new_n53748__,
    new_new_n53749__, new_new_n53750__, new_new_n53751__, new_new_n53752__,
    new_new_n53753__, new_new_n53754__, new_new_n53755__, new_new_n53756__,
    new_new_n53757__, new_new_n53758__, new_new_n53759__, new_new_n53760__,
    new_new_n53761__, new_new_n53762__, new_new_n53763__, new_new_n53764__,
    new_new_n53765__, new_new_n53766__, new_new_n53767__, new_new_n53768__,
    new_new_n53769__, new_new_n53770__, new_new_n53772__, new_new_n53773__,
    new_new_n53774__, new_new_n53775__, new_new_n53776__, new_new_n53777__,
    new_new_n53778__, new_new_n53779__, new_new_n53780__, new_new_n53782__,
    new_new_n53783__, new_new_n53784__, new_new_n53785__, new_new_n53786__,
    new_new_n53787__, new_new_n53788__, new_new_n53789__, new_new_n53790__,
    new_new_n53791__, new_new_n53792__, new_new_n53793__, new_new_n53794__,
    new_new_n53795__, new_new_n53796__, new_new_n53797__, new_new_n53798__,
    new_new_n53799__, new_new_n53800__, new_new_n53801__, new_new_n53802__,
    new_new_n53803__, new_new_n53804__, new_new_n53805__, new_new_n53806__,
    new_new_n53807__, new_new_n53808__, new_new_n53809__, new_new_n53810__,
    new_new_n53811__, new_new_n53812__, new_new_n53813__, new_new_n53814__,
    new_new_n53815__, new_new_n53816__, new_new_n53817__, new_new_n53818__,
    new_new_n53819__, new_new_n53820__, new_new_n53821__, new_new_n53822__,
    new_new_n53823__, new_new_n53824__, new_new_n53825__, new_new_n53826__,
    new_new_n53827__, new_new_n53828__, new_new_n53829__, new_new_n53830__,
    new_new_n53831__, new_new_n53832__, new_new_n53833__, new_new_n53834__,
    new_new_n53835__, new_new_n53836__, new_new_n53837__, new_new_n53838__,
    new_new_n53839__, new_new_n53840__, new_new_n53841__, new_new_n53842__,
    new_new_n53843__, new_new_n53844__, new_new_n53845__, new_new_n53846__,
    new_new_n53847__, new_new_n53848__, new_new_n53849__, new_new_n53850__,
    new_new_n53851__, new_new_n53852__, new_new_n53853__, new_new_n53854__,
    new_new_n53855__, new_new_n53856__, new_new_n53857__, new_new_n53858__,
    new_new_n53859__, new_new_n53860__, new_new_n53861__, new_new_n53862__,
    new_new_n53863__, new_new_n53864__, new_new_n53865__, new_new_n53866__,
    new_new_n53867__, new_new_n53868__, new_new_n53869__, new_new_n53870__,
    new_new_n53871__, new_new_n53872__, new_new_n53873__, new_new_n53874__,
    new_new_n53875__, new_new_n53876__, new_new_n53877__, new_new_n53878__,
    new_new_n53879__, new_new_n53880__, new_new_n53881__, new_new_n53882__,
    new_new_n53883__, new_new_n53884__, new_new_n53885__, new_new_n53886__,
    new_new_n53887__, new_new_n53888__, new_new_n53889__, new_new_n53890__,
    new_new_n53891__, new_new_n53892__, new_new_n53893__, new_new_n53894__,
    new_new_n53895__, new_new_n53896__, new_new_n53897__, new_new_n53898__,
    new_new_n53899__, new_new_n53900__, new_new_n53901__, new_new_n53902__,
    new_new_n53903__, new_new_n53904__, new_new_n53905__, new_new_n53906__,
    new_new_n53907__, new_new_n53909__, new_new_n53910__, new_new_n53911__,
    new_new_n53912__, new_new_n53913__, new_new_n53914__, new_new_n53915__,
    new_new_n53916__, new_new_n53917__, new_new_n53919__, new_new_n53920__,
    new_new_n53921__, new_new_n53922__, new_new_n53923__, new_new_n53924__,
    new_new_n53925__, new_new_n53926__, new_new_n53927__, new_new_n53928__,
    new_new_n53929__, new_new_n53930__, new_new_n53931__, new_new_n53932__,
    new_new_n53933__, new_new_n53934__, new_new_n53935__, new_new_n53936__,
    new_new_n53937__, new_new_n53938__, new_new_n53939__, new_new_n53940__,
    new_new_n53941__, new_new_n53942__, new_new_n53943__, new_new_n53944__,
    new_new_n53945__, new_new_n53946__, new_new_n53947__, new_new_n53948__,
    new_new_n53949__, new_new_n53950__, new_new_n53951__, new_new_n53952__,
    new_new_n53953__, new_new_n53954__, new_new_n53955__, new_new_n53956__,
    new_new_n53957__, new_new_n53958__, new_new_n53959__, new_new_n53960__,
    new_new_n53961__, new_new_n53962__, new_new_n53963__, new_new_n53964__,
    new_new_n53965__, new_new_n53966__, new_new_n53967__, new_new_n53968__,
    new_new_n53969__, new_new_n53970__, new_new_n53971__, new_new_n53972__,
    new_new_n53973__, new_new_n53974__, new_new_n53975__, new_new_n53976__,
    new_new_n53977__, new_new_n53978__, new_new_n53979__, new_new_n53980__,
    new_new_n53981__, new_new_n53982__, new_new_n53983__, new_new_n53984__,
    new_new_n53985__, new_new_n53986__, new_new_n53987__, new_new_n53988__,
    new_new_n53989__, new_new_n53990__, new_new_n53991__, new_new_n53992__,
    new_new_n53993__, new_new_n53994__, new_new_n53995__, new_new_n53996__,
    new_new_n53997__, new_new_n53998__, new_new_n53999__, new_new_n54000__,
    new_new_n54001__, new_new_n54002__, new_new_n54003__, new_new_n54004__,
    new_new_n54005__, new_new_n54006__, new_new_n54007__, new_new_n54008__,
    new_new_n54009__, new_new_n54010__, new_new_n54011__, new_new_n54012__,
    new_new_n54013__, new_new_n54014__, new_new_n54015__, new_new_n54016__,
    new_new_n54017__, new_new_n54018__, new_new_n54019__, new_new_n54020__,
    new_new_n54021__, new_new_n54022__, new_new_n54023__, new_new_n54024__,
    new_new_n54025__, new_new_n54026__, new_new_n54027__, new_new_n54028__,
    new_new_n54029__, new_new_n54030__, new_new_n54031__, new_new_n54032__,
    new_new_n54033__, new_new_n54034__, new_new_n54035__, new_new_n54036__,
    new_new_n54037__, new_new_n54038__, new_new_n54039__, new_new_n54040__,
    new_new_n54041__, new_new_n54042__, new_new_n54043__, new_new_n54044__,
    new_new_n54045__, new_new_n54046__, new_new_n54047__, new_new_n54049__,
    new_new_n54050__, new_new_n54051__, new_new_n54052__, new_new_n54053__,
    new_new_n54054__, new_new_n54055__, new_new_n54056__, new_new_n54057__,
    new_new_n54059__, new_new_n54060__, new_new_n54061__, new_new_n54062__,
    new_new_n54063__, new_new_n54064__, new_new_n54065__, new_new_n54066__,
    new_new_n54067__, new_new_n54068__, new_new_n54069__, new_new_n54070__,
    new_new_n54071__, new_new_n54072__, new_new_n54073__, new_new_n54074__,
    new_new_n54075__, new_new_n54076__, new_new_n54077__, new_new_n54078__,
    new_new_n54079__, new_new_n54080__, new_new_n54081__, new_new_n54082__,
    new_new_n54083__, new_new_n54084__, new_new_n54085__, new_new_n54086__,
    new_new_n54087__, new_new_n54088__, new_new_n54089__, new_new_n54090__,
    new_new_n54091__, new_new_n54092__, new_new_n54093__, new_new_n54094__,
    new_new_n54095__, new_new_n54096__, new_new_n54097__, new_new_n54098__,
    new_new_n54099__, new_new_n54100__, new_new_n54101__, new_new_n54102__,
    new_new_n54103__, new_new_n54104__, new_new_n54105__, new_new_n54106__,
    new_new_n54107__, new_new_n54108__, new_new_n54109__, new_new_n54110__,
    new_new_n54111__, new_new_n54112__, new_new_n54113__, new_new_n54114__,
    new_new_n54115__, new_new_n54116__, new_new_n54117__, new_new_n54118__,
    new_new_n54119__, new_new_n54120__, new_new_n54121__, new_new_n54122__,
    new_new_n54123__, new_new_n54124__, new_new_n54125__, new_new_n54126__,
    new_new_n54127__, new_new_n54128__, new_new_n54129__, new_new_n54130__,
    new_new_n54131__, new_new_n54132__, new_new_n54133__, new_new_n54134__,
    new_new_n54135__, new_new_n54136__, new_new_n54137__, new_new_n54138__,
    new_new_n54139__, new_new_n54140__, new_new_n54141__, new_new_n54142__,
    new_new_n54143__, new_new_n54144__, new_new_n54145__, new_new_n54146__,
    new_new_n54147__, new_new_n54148__, new_new_n54149__, new_new_n54150__,
    new_new_n54151__, new_new_n54152__, new_new_n54153__, new_new_n54154__,
    new_new_n54155__, new_new_n54156__, new_new_n54157__, new_new_n54158__,
    new_new_n54159__, new_new_n54160__, new_new_n54161__, new_new_n54162__,
    new_new_n54163__, new_new_n54164__, new_new_n54165__, new_new_n54166__,
    new_new_n54167__, new_new_n54168__, new_new_n54169__, new_new_n54170__,
    new_new_n54171__, new_new_n54172__, new_new_n54173__, new_new_n54174__,
    new_new_n54175__, new_new_n54176__, new_new_n54177__, new_new_n54178__,
    new_new_n54179__, new_new_n54180__, new_new_n54181__, new_new_n54182__,
    new_new_n54183__, new_new_n54184__, new_new_n54185__, new_new_n54186__,
    new_new_n54187__, new_new_n54188__, new_new_n54189__, new_new_n54191__,
    new_new_n54192__, new_new_n54193__, new_new_n54194__, new_new_n54195__,
    new_new_n54196__, new_new_n54197__, new_new_n54198__, new_new_n54199__,
    new_new_n54201__, new_new_n54202__, new_new_n54203__, new_new_n54204__,
    new_new_n54205__, new_new_n54206__, new_new_n54207__, new_new_n54208__,
    new_new_n54209__, new_new_n54210__, new_new_n54211__, new_new_n54212__,
    new_new_n54213__, new_new_n54214__, new_new_n54215__, new_new_n54216__,
    new_new_n54217__, new_new_n54218__, new_new_n54219__, new_new_n54220__,
    new_new_n54221__, new_new_n54222__, new_new_n54223__, new_new_n54224__,
    new_new_n54225__, new_new_n54226__, new_new_n54227__, new_new_n54228__,
    new_new_n54229__, new_new_n54230__, new_new_n54231__, new_new_n54232__,
    new_new_n54233__, new_new_n54234__, new_new_n54235__, new_new_n54236__,
    new_new_n54237__, new_new_n54238__, new_new_n54239__, new_new_n54240__,
    new_new_n54241__, new_new_n54242__, new_new_n54243__, new_new_n54244__,
    new_new_n54245__, new_new_n54246__, new_new_n54247__, new_new_n54248__,
    new_new_n54249__, new_new_n54250__, new_new_n54251__, new_new_n54252__,
    new_new_n54253__, new_new_n54254__, new_new_n54255__, new_new_n54256__,
    new_new_n54257__, new_new_n54258__, new_new_n54259__, new_new_n54260__,
    new_new_n54261__, new_new_n54262__, new_new_n54263__, new_new_n54264__,
    new_new_n54265__, new_new_n54266__, new_new_n54267__, new_new_n54268__,
    new_new_n54269__, new_new_n54270__, new_new_n54271__, new_new_n54272__,
    new_new_n54273__, new_new_n54274__, new_new_n54275__, new_new_n54276__,
    new_new_n54277__, new_new_n54278__, new_new_n54279__, new_new_n54280__,
    new_new_n54281__, new_new_n54282__, new_new_n54283__, new_new_n54284__,
    new_new_n54285__, new_new_n54286__, new_new_n54287__, new_new_n54288__,
    new_new_n54289__, new_new_n54290__, new_new_n54291__, new_new_n54292__,
    new_new_n54293__, new_new_n54294__, new_new_n54295__, new_new_n54296__,
    new_new_n54297__, new_new_n54298__, new_new_n54299__, new_new_n54300__,
    new_new_n54301__, new_new_n54302__, new_new_n54303__, new_new_n54304__,
    new_new_n54305__, new_new_n54306__, new_new_n54307__, new_new_n54308__,
    new_new_n54309__, new_new_n54310__, new_new_n54311__, new_new_n54312__,
    new_new_n54313__, new_new_n54314__, new_new_n54315__, new_new_n54316__,
    new_new_n54317__, new_new_n54318__, new_new_n54319__, new_new_n54320__,
    new_new_n54321__, new_new_n54322__, new_new_n54323__, new_new_n54324__,
    new_new_n54325__, new_new_n54326__, new_new_n54327__, new_new_n54328__,
    new_new_n54329__, new_new_n54330__, new_new_n54331__, new_new_n54333__,
    new_new_n54334__, new_new_n54335__, new_new_n54336__, new_new_n54337__,
    new_new_n54338__, new_new_n54339__, new_new_n54340__, new_new_n54341__,
    new_new_n54343__, new_new_n54344__, new_new_n54345__, new_new_n54346__,
    new_new_n54347__, new_new_n54348__, new_new_n54349__, new_new_n54350__,
    new_new_n54351__, new_new_n54352__, new_new_n54353__, new_new_n54354__,
    new_new_n54355__, new_new_n54356__, new_new_n54357__, new_new_n54358__,
    new_new_n54359__, new_new_n54360__, new_new_n54361__, new_new_n54362__,
    new_new_n54363__, new_new_n54364__, new_new_n54365__, new_new_n54366__,
    new_new_n54367__, new_new_n54368__, new_new_n54369__, new_new_n54370__,
    new_new_n54371__, new_new_n54372__, new_new_n54373__, new_new_n54374__,
    new_new_n54375__, new_new_n54376__, new_new_n54377__, new_new_n54378__,
    new_new_n54379__, new_new_n54380__, new_new_n54381__, new_new_n54382__,
    new_new_n54383__, new_new_n54384__, new_new_n54385__, new_new_n54386__,
    new_new_n54387__, new_new_n54388__, new_new_n54389__, new_new_n54390__,
    new_new_n54391__, new_new_n54392__, new_new_n54393__, new_new_n54394__,
    new_new_n54395__, new_new_n54396__, new_new_n54397__, new_new_n54398__,
    new_new_n54399__, new_new_n54400__, new_new_n54401__, new_new_n54402__,
    new_new_n54403__, new_new_n54404__, new_new_n54405__, new_new_n54406__,
    new_new_n54407__, new_new_n54408__, new_new_n54409__, new_new_n54410__,
    new_new_n54411__, new_new_n54412__, new_new_n54413__, new_new_n54414__,
    new_new_n54415__, new_new_n54416__, new_new_n54417__, new_new_n54418__,
    new_new_n54419__, new_new_n54420__, new_new_n54421__, new_new_n54422__,
    new_new_n54423__, new_new_n54424__, new_new_n54425__, new_new_n54426__,
    new_new_n54427__, new_new_n54428__, new_new_n54429__, new_new_n54430__,
    new_new_n54431__, new_new_n54432__, new_new_n54433__, new_new_n54434__,
    new_new_n54435__, new_new_n54436__, new_new_n54437__, new_new_n54438__,
    new_new_n54439__, new_new_n54440__, new_new_n54441__, new_new_n54442__,
    new_new_n54443__, new_new_n54444__, new_new_n54445__, new_new_n54446__,
    new_new_n54447__, new_new_n54448__, new_new_n54449__, new_new_n54450__,
    new_new_n54451__, new_new_n54452__, new_new_n54453__, new_new_n54454__,
    new_new_n54455__, new_new_n54456__, new_new_n54457__, new_new_n54458__,
    new_new_n54459__, new_new_n54460__, new_new_n54461__, new_new_n54462__,
    new_new_n54463__, new_new_n54464__, new_new_n54465__, new_new_n54466__,
    new_new_n54467__, new_new_n54468__, new_new_n54469__, new_new_n54470__,
    new_new_n54471__, new_new_n54472__, new_new_n54473__, new_new_n54475__,
    new_new_n54476__, new_new_n54477__, new_new_n54478__, new_new_n54479__,
    new_new_n54480__, new_new_n54481__, new_new_n54482__, new_new_n54483__,
    new_new_n54485__, new_new_n54486__, new_new_n54487__, new_new_n54488__,
    new_new_n54489__, new_new_n54490__, new_new_n54491__, new_new_n54492__,
    new_new_n54493__, new_new_n54494__, new_new_n54495__, new_new_n54496__,
    new_new_n54497__, new_new_n54498__, new_new_n54499__, new_new_n54500__,
    new_new_n54501__, new_new_n54502__, new_new_n54503__, new_new_n54504__,
    new_new_n54505__, new_new_n54506__, new_new_n54507__, new_new_n54508__,
    new_new_n54509__, new_new_n54510__, new_new_n54511__, new_new_n54512__,
    new_new_n54513__, new_new_n54514__, new_new_n54515__, new_new_n54516__,
    new_new_n54517__, new_new_n54518__, new_new_n54519__, new_new_n54520__,
    new_new_n54521__, new_new_n54522__, new_new_n54523__, new_new_n54524__,
    new_new_n54525__, new_new_n54526__, new_new_n54527__, new_new_n54528__,
    new_new_n54529__, new_new_n54530__, new_new_n54531__, new_new_n54532__,
    new_new_n54533__, new_new_n54534__, new_new_n54535__, new_new_n54536__,
    new_new_n54537__, new_new_n54538__, new_new_n54539__, new_new_n54540__,
    new_new_n54541__, new_new_n54542__, new_new_n54543__, new_new_n54544__,
    new_new_n54545__, new_new_n54546__, new_new_n54547__, new_new_n54548__,
    new_new_n54549__, new_new_n54550__, new_new_n54551__, new_new_n54552__,
    new_new_n54553__, new_new_n54554__, new_new_n54555__, new_new_n54556__,
    new_new_n54557__, new_new_n54558__, new_new_n54559__, new_new_n54560__,
    new_new_n54561__, new_new_n54562__, new_new_n54563__, new_new_n54564__,
    new_new_n54565__, new_new_n54566__, new_new_n54567__, new_new_n54568__,
    new_new_n54569__, new_new_n54570__, new_new_n54571__, new_new_n54572__,
    new_new_n54573__, new_new_n54574__, new_new_n54575__, new_new_n54576__,
    new_new_n54577__, new_new_n54578__, new_new_n54579__, new_new_n54580__,
    new_new_n54581__, new_new_n54582__, new_new_n54583__, new_new_n54584__,
    new_new_n54585__, new_new_n54586__, new_new_n54587__, new_new_n54588__,
    new_new_n54589__, new_new_n54590__, new_new_n54591__, new_new_n54592__,
    new_new_n54593__, new_new_n54594__, new_new_n54595__, new_new_n54596__,
    new_new_n54597__, new_new_n54598__, new_new_n54599__, new_new_n54600__,
    new_new_n54601__, new_new_n54602__, new_new_n54603__, new_new_n54604__,
    new_new_n54605__, new_new_n54606__, new_new_n54607__, new_new_n54608__,
    new_new_n54609__, new_new_n54610__, new_new_n54611__, new_new_n54612__,
    new_new_n54613__, new_new_n54614__, new_new_n54615__, new_new_n54617__,
    new_new_n54618__, new_new_n54619__, new_new_n54620__, new_new_n54621__,
    new_new_n54622__, new_new_n54623__, new_new_n54624__, new_new_n54625__,
    new_new_n54627__, new_new_n54628__, new_new_n54629__, new_new_n54630__,
    new_new_n54631__, new_new_n54632__, new_new_n54633__, new_new_n54634__,
    new_new_n54635__, new_new_n54636__, new_new_n54637__, new_new_n54638__,
    new_new_n54639__, new_new_n54640__, new_new_n54641__, new_new_n54642__,
    new_new_n54643__, new_new_n54644__, new_new_n54645__, new_new_n54646__,
    new_new_n54647__, new_new_n54648__, new_new_n54649__, new_new_n54650__,
    new_new_n54651__, new_new_n54652__, new_new_n54653__, new_new_n54654__,
    new_new_n54655__, new_new_n54656__, new_new_n54657__, new_new_n54658__,
    new_new_n54659__, new_new_n54660__, new_new_n54661__, new_new_n54662__,
    new_new_n54663__, new_new_n54664__, new_new_n54665__, new_new_n54666__,
    new_new_n54667__, new_new_n54668__, new_new_n54669__, new_new_n54670__,
    new_new_n54671__, new_new_n54672__, new_new_n54673__, new_new_n54674__,
    new_new_n54675__, new_new_n54676__, new_new_n54677__, new_new_n54678__,
    new_new_n54679__, new_new_n54680__, new_new_n54681__, new_new_n54682__,
    new_new_n54683__, new_new_n54684__, new_new_n54685__, new_new_n54686__,
    new_new_n54687__, new_new_n54688__, new_new_n54689__, new_new_n54690__,
    new_new_n54691__, new_new_n54692__, new_new_n54693__, new_new_n54694__,
    new_new_n54695__, new_new_n54696__, new_new_n54697__, new_new_n54698__,
    new_new_n54699__, new_new_n54700__, new_new_n54701__, new_new_n54702__,
    new_new_n54703__, new_new_n54704__, new_new_n54705__, new_new_n54706__,
    new_new_n54707__, new_new_n54708__, new_new_n54709__, new_new_n54710__,
    new_new_n54711__, new_new_n54712__, new_new_n54713__, new_new_n54714__,
    new_new_n54715__, new_new_n54716__, new_new_n54717__, new_new_n54718__,
    new_new_n54719__, new_new_n54720__, new_new_n54721__, new_new_n54722__,
    new_new_n54723__, new_new_n54724__, new_new_n54725__, new_new_n54726__,
    new_new_n54727__, new_new_n54728__, new_new_n54729__, new_new_n54730__,
    new_new_n54731__, new_new_n54732__, new_new_n54733__, new_new_n54734__,
    new_new_n54735__, new_new_n54736__, new_new_n54737__, new_new_n54738__,
    new_new_n54739__, new_new_n54740__, new_new_n54741__, new_new_n54742__,
    new_new_n54743__, new_new_n54744__, new_new_n54745__, new_new_n54746__,
    new_new_n54747__, new_new_n54748__, new_new_n54749__, new_new_n54750__,
    new_new_n54751__, new_new_n54752__, new_new_n54753__, new_new_n54754__,
    new_new_n54755__, new_new_n54756__, new_new_n54757__, new_new_n54759__,
    new_new_n54760__, new_new_n54761__, new_new_n54762__, new_new_n54763__,
    new_new_n54764__, new_new_n54765__, new_new_n54766__, new_new_n54767__,
    new_new_n54769__, new_new_n54770__, new_new_n54771__, new_new_n54772__,
    new_new_n54773__, new_new_n54774__, new_new_n54775__, new_new_n54776__,
    new_new_n54777__, new_new_n54778__, new_new_n54779__, new_new_n54780__,
    new_new_n54781__, new_new_n54782__, new_new_n54783__, new_new_n54784__,
    new_new_n54785__, new_new_n54786__, new_new_n54787__, new_new_n54788__,
    new_new_n54789__, new_new_n54790__, new_new_n54791__, new_new_n54792__,
    new_new_n54793__, new_new_n54794__, new_new_n54795__, new_new_n54796__,
    new_new_n54797__, new_new_n54798__, new_new_n54799__, new_new_n54800__,
    new_new_n54801__, new_new_n54802__, new_new_n54803__, new_new_n54804__,
    new_new_n54805__, new_new_n54806__, new_new_n54807__, new_new_n54808__,
    new_new_n54809__, new_new_n54810__, new_new_n54811__, new_new_n54812__,
    new_new_n54813__, new_new_n54814__, new_new_n54815__, new_new_n54816__,
    new_new_n54817__, new_new_n54818__, new_new_n54819__, new_new_n54820__,
    new_new_n54821__, new_new_n54822__, new_new_n54823__, new_new_n54824__,
    new_new_n54825__, new_new_n54826__, new_new_n54827__, new_new_n54828__,
    new_new_n54829__, new_new_n54830__, new_new_n54831__, new_new_n54832__,
    new_new_n54833__, new_new_n54834__, new_new_n54835__, new_new_n54836__,
    new_new_n54837__, new_new_n54838__, new_new_n54839__, new_new_n54840__,
    new_new_n54841__, new_new_n54842__, new_new_n54843__, new_new_n54844__,
    new_new_n54845__, new_new_n54846__, new_new_n54847__, new_new_n54848__,
    new_new_n54849__, new_new_n54850__, new_new_n54851__, new_new_n54852__,
    new_new_n54853__, new_new_n54854__, new_new_n54855__, new_new_n54856__,
    new_new_n54857__, new_new_n54858__, new_new_n54859__, new_new_n54860__,
    new_new_n54861__, new_new_n54862__, new_new_n54863__, new_new_n54864__,
    new_new_n54865__, new_new_n54866__, new_new_n54867__, new_new_n54868__,
    new_new_n54869__, new_new_n54870__, new_new_n54871__, new_new_n54872__,
    new_new_n54873__, new_new_n54874__, new_new_n54875__, new_new_n54876__,
    new_new_n54877__, new_new_n54878__, new_new_n54879__, new_new_n54880__,
    new_new_n54881__, new_new_n54882__, new_new_n54883__, new_new_n54884__,
    new_new_n54885__, new_new_n54886__, new_new_n54887__, new_new_n54888__,
    new_new_n54889__, new_new_n54890__, new_new_n54891__, new_new_n54892__,
    new_new_n54893__, new_new_n54894__, new_new_n54895__, new_new_n54896__,
    new_new_n54897__, new_new_n54898__, new_new_n54899__, new_new_n54901__,
    new_new_n54902__, new_new_n54903__, new_new_n54904__, new_new_n54905__,
    new_new_n54906__, new_new_n54907__, new_new_n54908__, new_new_n54909__,
    new_new_n54911__, new_new_n54912__, new_new_n54913__, new_new_n54914__,
    new_new_n54915__, new_new_n54916__, new_new_n54917__, new_new_n54918__,
    new_new_n54919__, new_new_n54920__, new_new_n54921__, new_new_n54922__,
    new_new_n54923__, new_new_n54924__, new_new_n54925__, new_new_n54926__,
    new_new_n54927__, new_new_n54928__, new_new_n54929__, new_new_n54930__,
    new_new_n54931__, new_new_n54932__, new_new_n54933__, new_new_n54934__,
    new_new_n54935__, new_new_n54936__, new_new_n54937__, new_new_n54938__,
    new_new_n54939__, new_new_n54940__, new_new_n54941__, new_new_n54942__,
    new_new_n54943__, new_new_n54944__, new_new_n54945__, new_new_n54946__,
    new_new_n54947__, new_new_n54948__, new_new_n54949__, new_new_n54950__,
    new_new_n54951__, new_new_n54952__, new_new_n54953__, new_new_n54954__,
    new_new_n54955__, new_new_n54956__, new_new_n54957__, new_new_n54958__,
    new_new_n54959__, new_new_n54960__, new_new_n54961__, new_new_n54962__,
    new_new_n54963__, new_new_n54964__, new_new_n54965__, new_new_n54966__,
    new_new_n54967__, new_new_n54968__, new_new_n54969__, new_new_n54970__,
    new_new_n54971__, new_new_n54972__, new_new_n54973__, new_new_n54974__,
    new_new_n54975__, new_new_n54976__, new_new_n54977__, new_new_n54978__,
    new_new_n54979__, new_new_n54980__, new_new_n54981__, new_new_n54982__,
    new_new_n54983__, new_new_n54984__, new_new_n54985__, new_new_n54986__,
    new_new_n54987__, new_new_n54988__, new_new_n54989__, new_new_n54990__,
    new_new_n54991__, new_new_n54992__, new_new_n54993__, new_new_n54994__,
    new_new_n54995__, new_new_n54996__, new_new_n54997__, new_new_n54998__,
    new_new_n54999__, new_new_n55000__, new_new_n55001__, new_new_n55002__,
    new_new_n55003__, new_new_n55004__, new_new_n55005__, new_new_n55006__,
    new_new_n55007__, new_new_n55008__, new_new_n55009__, new_new_n55010__,
    new_new_n55011__, new_new_n55012__, new_new_n55013__, new_new_n55014__,
    new_new_n55015__, new_new_n55016__, new_new_n55017__, new_new_n55018__,
    new_new_n55019__, new_new_n55020__, new_new_n55021__, new_new_n55022__,
    new_new_n55023__, new_new_n55024__, new_new_n55025__, new_new_n55026__,
    new_new_n55027__, new_new_n55028__, new_new_n55029__, new_new_n55030__,
    new_new_n55031__, new_new_n55032__, new_new_n55033__, new_new_n55034__,
    new_new_n55035__, new_new_n55036__, new_new_n55037__, new_new_n55038__,
    new_new_n55039__, new_new_n55040__, new_new_n55041__, new_new_n55043__,
    new_new_n55044__, new_new_n55045__, new_new_n55046__, new_new_n55047__,
    new_new_n55048__, new_new_n55049__, new_new_n55050__, new_new_n55051__,
    new_new_n55053__, new_new_n55054__, new_new_n55055__, new_new_n55056__,
    new_new_n55057__, new_new_n55058__, new_new_n55059__, new_new_n55060__,
    new_new_n55061__, new_new_n55062__, new_new_n55063__, new_new_n55064__,
    new_new_n55065__, new_new_n55066__, new_new_n55067__, new_new_n55068__,
    new_new_n55069__, new_new_n55070__, new_new_n55071__, new_new_n55072__,
    new_new_n55073__, new_new_n55074__, new_new_n55075__, new_new_n55076__,
    new_new_n55077__, new_new_n55078__, new_new_n55079__, new_new_n55080__,
    new_new_n55081__, new_new_n55082__, new_new_n55083__, new_new_n55084__,
    new_new_n55085__, new_new_n55086__, new_new_n55087__, new_new_n55088__,
    new_new_n55089__, new_new_n55090__, new_new_n55091__, new_new_n55092__,
    new_new_n55093__, new_new_n55094__, new_new_n55095__, new_new_n55096__,
    new_new_n55097__, new_new_n55098__, new_new_n55099__, new_new_n55100__,
    new_new_n55101__, new_new_n55102__, new_new_n55103__, new_new_n55104__,
    new_new_n55105__, new_new_n55106__, new_new_n55107__, new_new_n55108__,
    new_new_n55109__, new_new_n55110__, new_new_n55111__, new_new_n55112__,
    new_new_n55113__, new_new_n55114__, new_new_n55115__, new_new_n55116__,
    new_new_n55117__, new_new_n55118__, new_new_n55119__, new_new_n55120__,
    new_new_n55121__, new_new_n55122__, new_new_n55123__, new_new_n55124__,
    new_new_n55125__, new_new_n55126__, new_new_n55127__, new_new_n55128__,
    new_new_n55129__, new_new_n55130__, new_new_n55131__, new_new_n55132__,
    new_new_n55133__, new_new_n55134__, new_new_n55135__, new_new_n55136__,
    new_new_n55137__, new_new_n55138__, new_new_n55139__, new_new_n55140__,
    new_new_n55141__, new_new_n55142__, new_new_n55143__, new_new_n55144__,
    new_new_n55145__, new_new_n55146__, new_new_n55147__, new_new_n55148__,
    new_new_n55149__, new_new_n55150__, new_new_n55151__, new_new_n55152__,
    new_new_n55153__, new_new_n55154__, new_new_n55155__, new_new_n55156__,
    new_new_n55157__, new_new_n55158__, new_new_n55159__, new_new_n55160__,
    new_new_n55161__, new_new_n55162__, new_new_n55163__, new_new_n55164__,
    new_new_n55165__, new_new_n55166__, new_new_n55167__, new_new_n55168__,
    new_new_n55169__, new_new_n55170__, new_new_n55171__, new_new_n55172__,
    new_new_n55173__, new_new_n55174__, new_new_n55175__, new_new_n55176__,
    new_new_n55177__, new_new_n55178__, new_new_n55179__, new_new_n55180__,
    new_new_n55181__, new_new_n55182__, new_new_n55183__, new_new_n55185__,
    new_new_n55186__, new_new_n55187__, new_new_n55188__, new_new_n55189__,
    new_new_n55190__, new_new_n55191__, new_new_n55192__, new_new_n55193__,
    new_new_n55195__, new_new_n55196__, new_new_n55197__, new_new_n55198__,
    new_new_n55199__, new_new_n55200__, new_new_n55201__, new_new_n55202__,
    new_new_n55203__, new_new_n55204__, new_new_n55205__, new_new_n55206__,
    new_new_n55207__, new_new_n55208__, new_new_n55209__, new_new_n55210__,
    new_new_n55211__, new_new_n55212__, new_new_n55213__, new_new_n55214__,
    new_new_n55215__, new_new_n55216__, new_new_n55217__, new_new_n55218__,
    new_new_n55219__, new_new_n55220__, new_new_n55221__, new_new_n55222__,
    new_new_n55223__, new_new_n55224__, new_new_n55225__, new_new_n55226__,
    new_new_n55227__, new_new_n55228__, new_new_n55229__, new_new_n55230__,
    new_new_n55231__, new_new_n55232__, new_new_n55233__, new_new_n55234__,
    new_new_n55235__, new_new_n55236__, new_new_n55237__, new_new_n55238__,
    new_new_n55239__, new_new_n55240__, new_new_n55241__, new_new_n55242__,
    new_new_n55243__, new_new_n55244__, new_new_n55245__, new_new_n55246__,
    new_new_n55247__, new_new_n55248__, new_new_n55249__, new_new_n55250__,
    new_new_n55251__, new_new_n55252__, new_new_n55253__, new_new_n55254__,
    new_new_n55255__, new_new_n55256__, new_new_n55257__, new_new_n55258__,
    new_new_n55259__, new_new_n55260__, new_new_n55261__, new_new_n55262__,
    new_new_n55263__, new_new_n55264__, new_new_n55265__, new_new_n55266__,
    new_new_n55267__, new_new_n55268__, new_new_n55269__, new_new_n55270__,
    new_new_n55271__, new_new_n55272__, new_new_n55273__, new_new_n55274__,
    new_new_n55275__, new_new_n55276__, new_new_n55277__, new_new_n55278__,
    new_new_n55279__, new_new_n55280__, new_new_n55281__, new_new_n55282__,
    new_new_n55283__, new_new_n55284__, new_new_n55285__, new_new_n55286__,
    new_new_n55287__, new_new_n55288__, new_new_n55289__, new_new_n55290__,
    new_new_n55291__, new_new_n55292__, new_new_n55293__, new_new_n55294__,
    new_new_n55295__, new_new_n55296__, new_new_n55297__, new_new_n55298__,
    new_new_n55299__, new_new_n55300__, new_new_n55301__, new_new_n55302__,
    new_new_n55303__, new_new_n55304__, new_new_n55305__, new_new_n55306__,
    new_new_n55307__, new_new_n55308__, new_new_n55309__, new_new_n55310__,
    new_new_n55311__, new_new_n55312__, new_new_n55313__, new_new_n55314__,
    new_new_n55315__, new_new_n55316__, new_new_n55317__, new_new_n55318__,
    new_new_n55319__, new_new_n55320__, new_new_n55321__, new_new_n55322__,
    new_new_n55323__, new_new_n55324__, new_new_n55325__, new_new_n55327__,
    new_new_n55328__, new_new_n55329__, new_new_n55330__, new_new_n55331__,
    new_new_n55332__, new_new_n55333__, new_new_n55334__, new_new_n55335__,
    new_new_n55337__, new_new_n55338__, new_new_n55339__, new_new_n55340__,
    new_new_n55341__, new_new_n55342__, new_new_n55343__, new_new_n55344__,
    new_new_n55345__, new_new_n55346__, new_new_n55347__, new_new_n55348__,
    new_new_n55349__, new_new_n55350__, new_new_n55351__, new_new_n55352__,
    new_new_n55353__, new_new_n55354__, new_new_n55355__, new_new_n55356__,
    new_new_n55357__, new_new_n55358__, new_new_n55359__, new_new_n55360__,
    new_new_n55361__, new_new_n55362__, new_new_n55363__, new_new_n55364__,
    new_new_n55365__, new_new_n55366__, new_new_n55367__, new_new_n55368__,
    new_new_n55369__, new_new_n55370__, new_new_n55371__, new_new_n55372__,
    new_new_n55373__, new_new_n55374__, new_new_n55375__, new_new_n55376__,
    new_new_n55377__, new_new_n55378__, new_new_n55379__, new_new_n55380__,
    new_new_n55381__, new_new_n55382__, new_new_n55383__, new_new_n55384__,
    new_new_n55385__, new_new_n55386__, new_new_n55387__, new_new_n55388__,
    new_new_n55389__, new_new_n55390__, new_new_n55391__, new_new_n55392__,
    new_new_n55393__, new_new_n55394__, new_new_n55395__, new_new_n55396__,
    new_new_n55397__, new_new_n55398__, new_new_n55399__, new_new_n55400__,
    new_new_n55401__, new_new_n55402__, new_new_n55403__, new_new_n55404__,
    new_new_n55405__, new_new_n55406__, new_new_n55407__, new_new_n55408__,
    new_new_n55409__, new_new_n55410__, new_new_n55411__, new_new_n55412__,
    new_new_n55413__, new_new_n55414__, new_new_n55415__, new_new_n55416__,
    new_new_n55417__, new_new_n55418__, new_new_n55419__, new_new_n55420__,
    new_new_n55421__, new_new_n55422__, new_new_n55423__, new_new_n55424__,
    new_new_n55425__, new_new_n55426__, new_new_n55427__, new_new_n55428__,
    new_new_n55429__, new_new_n55430__, new_new_n55431__, new_new_n55432__,
    new_new_n55433__, new_new_n55434__, new_new_n55435__, new_new_n55436__,
    new_new_n55437__, new_new_n55438__, new_new_n55439__, new_new_n55440__,
    new_new_n55441__, new_new_n55442__, new_new_n55443__, new_new_n55444__,
    new_new_n55445__, new_new_n55446__, new_new_n55447__, new_new_n55448__,
    new_new_n55449__, new_new_n55450__, new_new_n55451__, new_new_n55452__,
    new_new_n55453__, new_new_n55454__, new_new_n55455__, new_new_n55456__,
    new_new_n55457__, new_new_n55458__, new_new_n55459__, new_new_n55460__,
    new_new_n55461__, new_new_n55462__, new_new_n55463__, new_new_n55464__,
    new_new_n55465__, new_new_n55466__, new_new_n55467__, new_new_n55469__,
    new_new_n55470__, new_new_n55471__, new_new_n55472__, new_new_n55473__,
    new_new_n55474__, new_new_n55475__, new_new_n55476__, new_new_n55477__,
    new_new_n55479__, new_new_n55480__, new_new_n55481__, new_new_n55482__,
    new_new_n55483__, new_new_n55484__, new_new_n55485__, new_new_n55486__,
    new_new_n55487__, new_new_n55488__, new_new_n55489__, new_new_n55490__,
    new_new_n55491__, new_new_n55492__, new_new_n55493__, new_new_n55494__,
    new_new_n55495__, new_new_n55496__, new_new_n55497__, new_new_n55498__,
    new_new_n55499__, new_new_n55500__, new_new_n55501__, new_new_n55502__,
    new_new_n55503__, new_new_n55504__, new_new_n55505__, new_new_n55506__,
    new_new_n55507__, new_new_n55508__, new_new_n55509__, new_new_n55510__,
    new_new_n55511__, new_new_n55512__, new_new_n55513__, new_new_n55514__,
    new_new_n55515__, new_new_n55516__, new_new_n55517__, new_new_n55518__,
    new_new_n55519__, new_new_n55520__, new_new_n55521__, new_new_n55522__,
    new_new_n55523__, new_new_n55524__, new_new_n55525__, new_new_n55526__,
    new_new_n55527__, new_new_n55528__, new_new_n55529__, new_new_n55530__,
    new_new_n55531__, new_new_n55532__, new_new_n55533__, new_new_n55534__,
    new_new_n55535__, new_new_n55536__, new_new_n55537__, new_new_n55538__,
    new_new_n55539__, new_new_n55540__, new_new_n55541__, new_new_n55542__,
    new_new_n55543__, new_new_n55544__, new_new_n55545__, new_new_n55546__,
    new_new_n55547__, new_new_n55548__, new_new_n55549__, new_new_n55550__,
    new_new_n55551__, new_new_n55552__, new_new_n55553__, new_new_n55554__,
    new_new_n55555__, new_new_n55556__, new_new_n55557__, new_new_n55558__,
    new_new_n55559__, new_new_n55560__, new_new_n55561__, new_new_n55562__,
    new_new_n55563__, new_new_n55564__, new_new_n55565__, new_new_n55566__,
    new_new_n55567__, new_new_n55568__, new_new_n55569__, new_new_n55570__,
    new_new_n55571__, new_new_n55572__, new_new_n55573__, new_new_n55574__,
    new_new_n55575__, new_new_n55576__, new_new_n55577__, new_new_n55578__,
    new_new_n55579__, new_new_n55580__, new_new_n55581__, new_new_n55582__,
    new_new_n55583__, new_new_n55584__, new_new_n55585__, new_new_n55586__,
    new_new_n55587__, new_new_n55588__, new_new_n55589__, new_new_n55590__,
    new_new_n55591__, new_new_n55592__, new_new_n55593__, new_new_n55594__,
    new_new_n55595__, new_new_n55596__, new_new_n55597__, new_new_n55598__,
    new_new_n55599__, new_new_n55600__, new_new_n55601__, new_new_n55602__,
    new_new_n55603__, new_new_n55604__, new_new_n55605__, new_new_n55606__,
    new_new_n55607__, new_new_n55608__, new_new_n55609__, new_new_n55611__,
    new_new_n55612__, new_new_n55613__, new_new_n55614__, new_new_n55615__,
    new_new_n55616__, new_new_n55617__, new_new_n55618__, new_new_n55619__,
    new_new_n55621__, new_new_n55622__, new_new_n55623__, new_new_n55624__,
    new_new_n55625__, new_new_n55626__, new_new_n55627__, new_new_n55628__,
    new_new_n55629__, new_new_n55630__, new_new_n55631__, new_new_n55632__,
    new_new_n55633__, new_new_n55634__, new_new_n55635__, new_new_n55636__,
    new_new_n55637__, new_new_n55638__, new_new_n55639__, new_new_n55640__,
    new_new_n55641__, new_new_n55642__, new_new_n55643__, new_new_n55644__,
    new_new_n55645__, new_new_n55646__, new_new_n55647__, new_new_n55648__,
    new_new_n55649__, new_new_n55650__, new_new_n55651__, new_new_n55652__,
    new_new_n55653__, new_new_n55654__, new_new_n55655__, new_new_n55656__,
    new_new_n55657__, new_new_n55658__, new_new_n55659__, new_new_n55660__,
    new_new_n55661__, new_new_n55662__, new_new_n55663__, new_new_n55664__,
    new_new_n55665__, new_new_n55666__, new_new_n55667__, new_new_n55668__,
    new_new_n55669__, new_new_n55670__, new_new_n55671__, new_new_n55672__,
    new_new_n55673__, new_new_n55674__, new_new_n55675__, new_new_n55676__,
    new_new_n55677__, new_new_n55678__, new_new_n55679__, new_new_n55680__,
    new_new_n55681__, new_new_n55682__, new_new_n55683__, new_new_n55684__,
    new_new_n55685__, new_new_n55686__, new_new_n55687__, new_new_n55688__,
    new_new_n55689__, new_new_n55690__, new_new_n55691__, new_new_n55692__,
    new_new_n55693__, new_new_n55694__, new_new_n55695__, new_new_n55696__,
    new_new_n55697__, new_new_n55698__, new_new_n55699__, new_new_n55700__,
    new_new_n55701__, new_new_n55702__, new_new_n55703__, new_new_n55704__,
    new_new_n55705__, new_new_n55706__, new_new_n55707__, new_new_n55708__,
    new_new_n55709__, new_new_n55710__, new_new_n55711__, new_new_n55712__,
    new_new_n55713__, new_new_n55714__, new_new_n55715__, new_new_n55716__,
    new_new_n55717__, new_new_n55718__, new_new_n55719__, new_new_n55720__,
    new_new_n55721__, new_new_n55722__, new_new_n55723__, new_new_n55724__,
    new_new_n55725__, new_new_n55726__, new_new_n55727__, new_new_n55728__,
    new_new_n55729__, new_new_n55730__, new_new_n55731__, new_new_n55732__,
    new_new_n55733__, new_new_n55734__, new_new_n55735__, new_new_n55736__,
    new_new_n55737__, new_new_n55738__, new_new_n55739__, new_new_n55740__,
    new_new_n55741__, new_new_n55742__, new_new_n55743__, new_new_n55744__,
    new_new_n55745__, new_new_n55746__, new_new_n55747__, new_new_n55748__,
    new_new_n55749__, new_new_n55750__, new_new_n55751__, new_new_n55753__,
    new_new_n55754__, new_new_n55755__, new_new_n55756__, new_new_n55757__,
    new_new_n55758__, new_new_n55759__, new_new_n55760__, new_new_n55761__,
    new_new_n55763__, new_new_n55764__, new_new_n55765__, new_new_n55766__,
    new_new_n55767__, new_new_n55768__, new_new_n55769__, new_new_n55770__,
    new_new_n55771__, new_new_n55772__, new_new_n55773__, new_new_n55774__,
    new_new_n55775__, new_new_n55776__, new_new_n55777__, new_new_n55778__,
    new_new_n55779__, new_new_n55780__, new_new_n55781__, new_new_n55782__,
    new_new_n55783__, new_new_n55784__, new_new_n55785__, new_new_n55786__,
    new_new_n55787__, new_new_n55788__, new_new_n55789__, new_new_n55790__,
    new_new_n55791__, new_new_n55792__, new_new_n55793__, new_new_n55794__,
    new_new_n55795__, new_new_n55796__, new_new_n55797__, new_new_n55798__,
    new_new_n55799__, new_new_n55800__, new_new_n55801__, new_new_n55802__,
    new_new_n55803__, new_new_n55804__, new_new_n55805__, new_new_n55806__,
    new_new_n55807__, new_new_n55808__, new_new_n55809__, new_new_n55810__,
    new_new_n55811__, new_new_n55812__, new_new_n55813__, new_new_n55814__,
    new_new_n55815__, new_new_n55816__, new_new_n55817__, new_new_n55818__,
    new_new_n55819__, new_new_n55820__, new_new_n55821__, new_new_n55822__,
    new_new_n55823__, new_new_n55824__, new_new_n55825__, new_new_n55826__,
    new_new_n55827__, new_new_n55828__, new_new_n55829__, new_new_n55830__,
    new_new_n55831__, new_new_n55832__, new_new_n55833__, new_new_n55834__,
    new_new_n55835__, new_new_n55836__, new_new_n55837__, new_new_n55838__,
    new_new_n55839__, new_new_n55840__, new_new_n55841__, new_new_n55842__,
    new_new_n55843__, new_new_n55844__, new_new_n55845__, new_new_n55846__,
    new_new_n55847__, new_new_n55848__, new_new_n55849__, new_new_n55850__,
    new_new_n55851__, new_new_n55852__, new_new_n55853__, new_new_n55854__,
    new_new_n55855__, new_new_n55856__, new_new_n55857__, new_new_n55858__,
    new_new_n55859__, new_new_n55860__, new_new_n55861__, new_new_n55862__,
    new_new_n55863__, new_new_n55864__, new_new_n55865__, new_new_n55866__,
    new_new_n55867__, new_new_n55868__, new_new_n55869__, new_new_n55870__,
    new_new_n55871__, new_new_n55872__, new_new_n55873__, new_new_n55874__,
    new_new_n55875__, new_new_n55876__, new_new_n55877__, new_new_n55878__,
    new_new_n55879__, new_new_n55880__, new_new_n55881__, new_new_n55882__,
    new_new_n55883__, new_new_n55884__, new_new_n55885__, new_new_n55886__,
    new_new_n55887__, new_new_n55888__, new_new_n55889__, new_new_n55890__,
    new_new_n55891__, new_new_n55892__, new_new_n55893__, new_new_n55895__,
    new_new_n55896__, new_new_n55897__, new_new_n55898__, new_new_n55899__,
    new_new_n55900__, new_new_n55901__, new_new_n55902__, new_new_n55903__,
    new_new_n55905__, new_new_n55906__, new_new_n55907__, new_new_n55908__,
    new_new_n55909__, new_new_n55910__, new_new_n55911__, new_new_n55912__,
    new_new_n55913__, new_new_n55914__, new_new_n55915__, new_new_n55916__,
    new_new_n55917__, new_new_n55918__, new_new_n55919__, new_new_n55920__,
    new_new_n55921__, new_new_n55922__, new_new_n55923__, new_new_n55924__,
    new_new_n55925__, new_new_n55926__, new_new_n55927__, new_new_n55928__,
    new_new_n55929__, new_new_n55930__, new_new_n55931__, new_new_n55932__,
    new_new_n55933__, new_new_n55934__, new_new_n55935__, new_new_n55936__,
    new_new_n55937__, new_new_n55938__, new_new_n55939__, new_new_n55940__,
    new_new_n55941__, new_new_n55942__, new_new_n55943__, new_new_n55944__,
    new_new_n55945__, new_new_n55946__, new_new_n55947__, new_new_n55948__,
    new_new_n55949__, new_new_n55950__, new_new_n55951__, new_new_n55952__,
    new_new_n55953__, new_new_n55954__, new_new_n55955__, new_new_n55956__,
    new_new_n55957__, new_new_n55958__, new_new_n55959__, new_new_n55960__,
    new_new_n55961__, new_new_n55962__, new_new_n55963__, new_new_n55964__,
    new_new_n55965__, new_new_n55966__, new_new_n55967__, new_new_n55968__,
    new_new_n55969__, new_new_n55970__, new_new_n55971__, new_new_n55972__,
    new_new_n55973__, new_new_n55974__, new_new_n55975__, new_new_n55976__,
    new_new_n55977__, new_new_n55978__, new_new_n55979__, new_new_n55980__,
    new_new_n55981__, new_new_n55982__, new_new_n55983__, new_new_n55984__,
    new_new_n55985__, new_new_n55986__, new_new_n55987__, new_new_n55988__,
    new_new_n55989__, new_new_n55990__, new_new_n55991__, new_new_n55992__,
    new_new_n55993__, new_new_n55994__, new_new_n55995__, new_new_n55996__,
    new_new_n55997__, new_new_n55998__, new_new_n55999__, new_new_n56000__,
    new_new_n56001__, new_new_n56002__, new_new_n56003__, new_new_n56004__,
    new_new_n56005__, new_new_n56006__, new_new_n56007__, new_new_n56008__,
    new_new_n56009__, new_new_n56010__, new_new_n56011__, new_new_n56012__,
    new_new_n56013__, new_new_n56014__, new_new_n56015__, new_new_n56016__,
    new_new_n56017__, new_new_n56018__, new_new_n56019__, new_new_n56020__,
    new_new_n56021__, new_new_n56022__, new_new_n56023__, new_new_n56024__,
    new_new_n56025__, new_new_n56026__, new_new_n56027__, new_new_n56028__,
    new_new_n56029__, new_new_n56030__, new_new_n56031__, new_new_n56032__,
    new_new_n56033__, new_new_n56034__, new_new_n56035__, new_new_n56037__,
    new_new_n56038__, new_new_n56039__, new_new_n56040__, new_new_n56041__,
    new_new_n56042__, new_new_n56043__, new_new_n56044__, new_new_n56045__,
    new_new_n56047__, new_new_n56048__, new_new_n56049__, new_new_n56050__,
    new_new_n56051__, new_new_n56052__, new_new_n56053__, new_new_n56054__,
    new_new_n56055__, new_new_n56056__, new_new_n56057__, new_new_n56058__,
    new_new_n56059__, new_new_n56060__, new_new_n56061__, new_new_n56062__,
    new_new_n56063__, new_new_n56064__, new_new_n56065__, new_new_n56066__,
    new_new_n56067__, new_new_n56068__, new_new_n56069__, new_new_n56070__,
    new_new_n56071__, new_new_n56072__, new_new_n56073__, new_new_n56074__,
    new_new_n56075__, new_new_n56076__, new_new_n56077__, new_new_n56078__,
    new_new_n56079__, new_new_n56080__, new_new_n56081__, new_new_n56082__,
    new_new_n56083__, new_new_n56084__, new_new_n56085__, new_new_n56086__,
    new_new_n56087__, new_new_n56088__, new_new_n56089__, new_new_n56090__,
    new_new_n56091__, new_new_n56092__, new_new_n56093__, new_new_n56094__,
    new_new_n56095__, new_new_n56096__, new_new_n56097__, new_new_n56098__,
    new_new_n56099__, new_new_n56100__, new_new_n56101__, new_new_n56102__,
    new_new_n56103__, new_new_n56104__, new_new_n56105__, new_new_n56106__,
    new_new_n56107__, new_new_n56108__, new_new_n56109__, new_new_n56110__,
    new_new_n56111__, new_new_n56112__, new_new_n56113__, new_new_n56114__,
    new_new_n56115__, new_new_n56116__, new_new_n56117__, new_new_n56118__,
    new_new_n56119__, new_new_n56120__, new_new_n56121__, new_new_n56122__,
    new_new_n56123__, new_new_n56124__, new_new_n56125__, new_new_n56126__,
    new_new_n56127__, new_new_n56128__, new_new_n56129__, new_new_n56130__,
    new_new_n56131__, new_new_n56132__, new_new_n56133__, new_new_n56134__,
    new_new_n56135__, new_new_n56136__, new_new_n56137__, new_new_n56138__,
    new_new_n56139__, new_new_n56140__, new_new_n56141__, new_new_n56142__,
    new_new_n56143__, new_new_n56144__, new_new_n56145__, new_new_n56146__,
    new_new_n56147__, new_new_n56148__, new_new_n56149__, new_new_n56150__,
    new_new_n56151__, new_new_n56152__, new_new_n56153__, new_new_n56154__,
    new_new_n56155__, new_new_n56156__, new_new_n56157__, new_new_n56158__,
    new_new_n56159__, new_new_n56160__, new_new_n56161__, new_new_n56162__,
    new_new_n56163__, new_new_n56164__, new_new_n56165__, new_new_n56166__,
    new_new_n56167__, new_new_n56168__, new_new_n56169__, new_new_n56170__,
    new_new_n56171__, new_new_n56172__, new_new_n56173__, new_new_n56174__,
    new_new_n56175__, new_new_n56176__, new_new_n56177__, new_new_n56179__,
    new_new_n56180__, new_new_n56181__, new_new_n56182__, new_new_n56183__,
    new_new_n56184__, new_new_n56185__, new_new_n56186__, new_new_n56187__,
    new_new_n56189__, new_new_n56190__, new_new_n56191__, new_new_n56192__,
    new_new_n56193__, new_new_n56194__, new_new_n56195__, new_new_n56196__,
    new_new_n56197__, new_new_n56198__, new_new_n56199__, new_new_n56200__,
    new_new_n56201__, new_new_n56202__, new_new_n56203__, new_new_n56204__,
    new_new_n56205__, new_new_n56206__, new_new_n56207__, new_new_n56208__,
    new_new_n56209__, new_new_n56210__, new_new_n56211__, new_new_n56212__,
    new_new_n56213__, new_new_n56214__, new_new_n56215__, new_new_n56216__,
    new_new_n56217__, new_new_n56218__, new_new_n56219__, new_new_n56220__,
    new_new_n56221__, new_new_n56222__, new_new_n56223__, new_new_n56224__,
    new_new_n56225__, new_new_n56226__, new_new_n56227__, new_new_n56228__,
    new_new_n56229__, new_new_n56230__, new_new_n56231__, new_new_n56232__,
    new_new_n56233__, new_new_n56234__, new_new_n56235__, new_new_n56236__,
    new_new_n56237__, new_new_n56238__, new_new_n56239__, new_new_n56240__,
    new_new_n56241__, new_new_n56242__, new_new_n56243__, new_new_n56244__,
    new_new_n56245__, new_new_n56246__, new_new_n56247__, new_new_n56248__,
    new_new_n56249__, new_new_n56250__, new_new_n56251__, new_new_n56252__,
    new_new_n56253__, new_new_n56254__, new_new_n56255__, new_new_n56256__,
    new_new_n56257__, new_new_n56258__, new_new_n56259__, new_new_n56260__,
    new_new_n56261__, new_new_n56262__, new_new_n56263__, new_new_n56264__,
    new_new_n56265__, new_new_n56266__, new_new_n56267__, new_new_n56268__,
    new_new_n56269__, new_new_n56270__, new_new_n56271__, new_new_n56272__,
    new_new_n56273__, new_new_n56274__, new_new_n56275__, new_new_n56276__,
    new_new_n56277__, new_new_n56278__, new_new_n56279__, new_new_n56280__,
    new_new_n56281__, new_new_n56282__, new_new_n56283__, new_new_n56284__,
    new_new_n56285__, new_new_n56286__, new_new_n56287__, new_new_n56288__,
    new_new_n56289__, new_new_n56290__, new_new_n56291__, new_new_n56292__,
    new_new_n56293__, new_new_n56294__, new_new_n56295__, new_new_n56296__,
    new_new_n56297__, new_new_n56298__, new_new_n56299__, new_new_n56300__,
    new_new_n56301__, new_new_n56302__, new_new_n56303__, new_new_n56304__,
    new_new_n56305__, new_new_n56306__, new_new_n56307__, new_new_n56308__,
    new_new_n56309__, new_new_n56310__, new_new_n56311__, new_new_n56312__,
    new_new_n56313__, new_new_n56314__, new_new_n56315__, new_new_n56316__,
    new_new_n56317__, new_new_n56318__, new_new_n56319__, new_new_n56321__,
    new_new_n56322__, new_new_n56323__, new_new_n56324__, new_new_n56325__,
    new_new_n56326__, new_new_n56327__, new_new_n56328__, new_new_n56329__,
    new_new_n56331__, new_new_n56332__, new_new_n56333__, new_new_n56334__,
    new_new_n56335__, new_new_n56336__, new_new_n56337__, new_new_n56338__,
    new_new_n56339__, new_new_n56340__, new_new_n56341__, new_new_n56342__,
    new_new_n56343__, new_new_n56344__, new_new_n56345__, new_new_n56346__,
    new_new_n56347__, new_new_n56348__, new_new_n56349__, new_new_n56350__,
    new_new_n56351__, new_new_n56352__, new_new_n56353__, new_new_n56354__,
    new_new_n56355__, new_new_n56356__, new_new_n56357__, new_new_n56358__,
    new_new_n56359__, new_new_n56360__, new_new_n56361__, new_new_n56362__,
    new_new_n56363__, new_new_n56364__, new_new_n56365__, new_new_n56366__,
    new_new_n56367__, new_new_n56368__, new_new_n56369__, new_new_n56370__,
    new_new_n56371__, new_new_n56372__, new_new_n56373__, new_new_n56374__,
    new_new_n56375__, new_new_n56376__, new_new_n56377__, new_new_n56378__,
    new_new_n56379__, new_new_n56380__, new_new_n56381__, new_new_n56382__,
    new_new_n56383__, new_new_n56384__, new_new_n56385__, new_new_n56386__,
    new_new_n56387__, new_new_n56388__, new_new_n56389__, new_new_n56390__,
    new_new_n56391__, new_new_n56392__, new_new_n56393__, new_new_n56394__,
    new_new_n56395__, new_new_n56396__, new_new_n56397__, new_new_n56398__,
    new_new_n56399__, new_new_n56400__, new_new_n56401__, new_new_n56402__,
    new_new_n56403__, new_new_n56404__, new_new_n56405__, new_new_n56406__,
    new_new_n56407__, new_new_n56408__, new_new_n56409__, new_new_n56410__,
    new_new_n56411__, new_new_n56412__, new_new_n56413__, new_new_n56414__,
    new_new_n56415__, new_new_n56416__, new_new_n56417__, new_new_n56418__,
    new_new_n56419__, new_new_n56420__, new_new_n56421__, new_new_n56422__,
    new_new_n56423__, new_new_n56424__, new_new_n56425__, new_new_n56426__,
    new_new_n56427__, new_new_n56428__, new_new_n56429__, new_new_n56430__,
    new_new_n56431__, new_new_n56432__, new_new_n56433__, new_new_n56434__,
    new_new_n56435__, new_new_n56436__, new_new_n56437__, new_new_n56438__,
    new_new_n56439__, new_new_n56440__, new_new_n56441__, new_new_n56442__,
    new_new_n56443__, new_new_n56444__, new_new_n56445__, new_new_n56446__,
    new_new_n56447__, new_new_n56448__, new_new_n56449__, new_new_n56450__,
    new_new_n56451__, new_new_n56452__, new_new_n56453__, new_new_n56454__,
    new_new_n56455__, new_new_n56456__, new_new_n56457__, new_new_n56459__,
    new_new_n56460__, new_new_n56461__, new_new_n56462__, new_new_n56463__,
    new_new_n56464__, new_new_n56465__, new_new_n56466__, new_new_n56467__,
    new_new_n56469__, new_new_n56470__, new_new_n56471__, new_new_n56472__,
    new_new_n56473__, new_new_n56474__, new_new_n56475__, new_new_n56476__,
    new_new_n56477__, new_new_n56478__, new_new_n56479__, new_new_n56480__,
    new_new_n56481__, new_new_n56482__, new_new_n56483__, new_new_n56484__,
    new_new_n56485__, new_new_n56486__, new_new_n56487__, new_new_n56488__,
    new_new_n56489__, new_new_n56490__, new_new_n56491__, new_new_n56492__,
    new_new_n56493__, new_new_n56494__, new_new_n56495__, new_new_n56496__,
    new_new_n56497__, new_new_n56498__, new_new_n56499__, new_new_n56500__,
    new_new_n56501__, new_new_n56502__, new_new_n56503__, new_new_n56504__,
    new_new_n56505__, new_new_n56506__, new_new_n56507__, new_new_n56508__,
    new_new_n56509__, new_new_n56510__, new_new_n56511__, new_new_n56512__,
    new_new_n56513__, new_new_n56514__, new_new_n56515__, new_new_n56516__,
    new_new_n56517__, new_new_n56518__, new_new_n56519__, new_new_n56520__,
    new_new_n56521__, new_new_n56522__, new_new_n56523__, new_new_n56524__,
    new_new_n56525__, new_new_n56526__, new_new_n56527__, new_new_n56528__,
    new_new_n56529__, new_new_n56530__, new_new_n56531__, new_new_n56532__,
    new_new_n56533__, new_new_n56534__, new_new_n56535__, new_new_n56536__,
    new_new_n56537__, new_new_n56538__, new_new_n56539__, new_new_n56540__,
    new_new_n56541__, new_new_n56542__, new_new_n56543__, new_new_n56544__,
    new_new_n56545__, new_new_n56546__, new_new_n56547__, new_new_n56548__,
    new_new_n56549__, new_new_n56550__, new_new_n56551__, new_new_n56552__,
    new_new_n56553__, new_new_n56554__, new_new_n56555__, new_new_n56556__,
    new_new_n56557__, new_new_n56558__, new_new_n56559__, new_new_n56560__,
    new_new_n56561__, new_new_n56562__, new_new_n56563__, new_new_n56564__,
    new_new_n56565__, new_new_n56566__, new_new_n56567__, new_new_n56568__,
    new_new_n56569__, new_new_n56570__, new_new_n56571__, new_new_n56572__,
    new_new_n56573__, new_new_n56574__, new_new_n56575__, new_new_n56576__,
    new_new_n56577__, new_new_n56578__, new_new_n56579__, new_new_n56580__,
    new_new_n56581__, new_new_n56582__, new_new_n56583__, new_new_n56584__,
    new_new_n56585__, new_new_n56586__, new_new_n56587__, new_new_n56588__,
    new_new_n56590__, new_new_n56591__, new_new_n56592__, new_new_n56593__,
    new_new_n56594__, new_new_n56595__, new_new_n56596__, new_new_n56597__,
    new_new_n56598__, new_new_n56600__, new_new_n56601__, new_new_n56602__,
    new_new_n56603__, new_new_n56604__, new_new_n56605__, new_new_n56606__,
    new_new_n56607__, new_new_n56608__, new_new_n56609__, new_new_n56610__,
    new_new_n56611__, new_new_n56612__, new_new_n56613__, new_new_n56614__,
    new_new_n56615__, new_new_n56616__, new_new_n56617__, new_new_n56618__,
    new_new_n56619__, new_new_n56620__, new_new_n56621__, new_new_n56622__,
    new_new_n56623__, new_new_n56624__, new_new_n56625__, new_new_n56626__,
    new_new_n56627__, new_new_n56628__, new_new_n56629__, new_new_n56630__,
    new_new_n56631__, new_new_n56632__, new_new_n56633__, new_new_n56634__,
    new_new_n56635__, new_new_n56636__, new_new_n56637__, new_new_n56638__,
    new_new_n56639__, new_new_n56640__, new_new_n56641__, new_new_n56642__,
    new_new_n56643__, new_new_n56644__, new_new_n56645__, new_new_n56646__,
    new_new_n56647__, new_new_n56648__, new_new_n56649__, new_new_n56650__,
    new_new_n56651__, new_new_n56652__, new_new_n56653__, new_new_n56654__,
    new_new_n56655__, new_new_n56656__, new_new_n56657__, new_new_n56658__,
    new_new_n56659__, new_new_n56660__, new_new_n56661__, new_new_n56662__,
    new_new_n56663__, new_new_n56664__, new_new_n56665__, new_new_n56666__,
    new_new_n56667__, new_new_n56668__, new_new_n56669__, new_new_n56670__,
    new_new_n56671__, new_new_n56672__, new_new_n56673__, new_new_n56674__,
    new_new_n56675__, new_new_n56676__, new_new_n56677__, new_new_n56678__,
    new_new_n56679__, new_new_n56680__, new_new_n56681__, new_new_n56682__,
    new_new_n56683__, new_new_n56684__, new_new_n56685__, new_new_n56686__,
    new_new_n56687__, new_new_n56688__, new_new_n56689__, new_new_n56690__,
    new_new_n56691__, new_new_n56692__, new_new_n56693__, new_new_n56694__,
    new_new_n56695__, new_new_n56696__, new_new_n56697__, new_new_n56698__,
    new_new_n56699__, new_new_n56700__, new_new_n56701__, new_new_n56702__,
    new_new_n56703__, new_new_n56704__, new_new_n56705__, new_new_n56706__,
    new_new_n56707__, new_new_n56708__, new_new_n56710__, new_new_n56711__,
    new_new_n56712__, new_new_n56713__, new_new_n56714__, new_new_n56715__,
    new_new_n56716__, new_new_n56717__, new_new_n56718__, new_new_n56720__,
    new_new_n56721__, new_new_n56722__, new_new_n56723__, new_new_n56724__,
    new_new_n56725__, new_new_n56726__, new_new_n56727__, new_new_n56728__,
    new_new_n56729__, new_new_n56730__, new_new_n56731__, new_new_n56732__,
    new_new_n56733__, new_new_n56734__, new_new_n56735__, new_new_n56736__,
    new_new_n56737__, new_new_n56738__, new_new_n56739__, new_new_n56740__,
    new_new_n56741__, new_new_n56742__, new_new_n56743__, new_new_n56744__,
    new_new_n56745__, new_new_n56746__, new_new_n56747__, new_new_n56748__,
    new_new_n56749__, new_new_n56750__, new_new_n56751__, new_new_n56752__,
    new_new_n56753__, new_new_n56754__, new_new_n56755__, new_new_n56756__,
    new_new_n56757__, new_new_n56758__, new_new_n56759__, new_new_n56760__,
    new_new_n56761__, new_new_n56762__, new_new_n56763__, new_new_n56764__,
    new_new_n56765__, new_new_n56766__, new_new_n56767__, new_new_n56768__,
    new_new_n56769__, new_new_n56770__, new_new_n56771__, new_new_n56772__,
    new_new_n56773__, new_new_n56774__, new_new_n56775__, new_new_n56776__,
    new_new_n56777__, new_new_n56778__, new_new_n56779__, new_new_n56780__,
    new_new_n56781__, new_new_n56782__, new_new_n56783__, new_new_n56784__,
    new_new_n56785__, new_new_n56786__, new_new_n56787__, new_new_n56788__,
    new_new_n56789__, new_new_n56790__, new_new_n56791__, new_new_n56792__,
    new_new_n56793__, new_new_n56794__, new_new_n56795__, new_new_n56796__,
    new_new_n56797__, new_new_n56798__, new_new_n56799__, new_new_n56800__,
    new_new_n56801__, new_new_n56802__, new_new_n56803__, new_new_n56804__,
    new_new_n56805__, new_new_n56806__, new_new_n56807__, new_new_n56808__,
    new_new_n56809__, new_new_n56810__, new_new_n56811__, new_new_n56812__,
    new_new_n56813__, new_new_n56814__, new_new_n56815__, new_new_n56816__,
    new_new_n56817__, new_new_n56818__, new_new_n56819__, new_new_n56820__,
    new_new_n56821__, new_new_n56822__, new_new_n56823__, new_new_n56824__,
    new_new_n56825__, new_new_n56826__, new_new_n56827__, new_new_n56828__,
    new_new_n56830__, new_new_n56831__, new_new_n56832__, new_new_n56833__,
    new_new_n56834__, new_new_n56835__, new_new_n56836__, new_new_n56837__,
    new_new_n56838__, new_new_n56840__, new_new_n56841__, new_new_n56842__,
    new_new_n56843__, new_new_n56844__, new_new_n56845__, new_new_n56846__,
    new_new_n56847__, new_new_n56848__, new_new_n56849__, new_new_n56850__,
    new_new_n56851__, new_new_n56852__, new_new_n56853__, new_new_n56854__,
    new_new_n56855__, new_new_n56856__, new_new_n56857__, new_new_n56858__,
    new_new_n56859__, new_new_n56860__, new_new_n56861__, new_new_n56862__,
    new_new_n56863__, new_new_n56864__, new_new_n56865__, new_new_n56866__,
    new_new_n56867__, new_new_n56868__, new_new_n56869__, new_new_n56870__,
    new_new_n56871__, new_new_n56872__, new_new_n56873__, new_new_n56874__,
    new_new_n56875__, new_new_n56876__, new_new_n56877__, new_new_n56878__,
    new_new_n56879__, new_new_n56880__, new_new_n56881__, new_new_n56882__,
    new_new_n56883__, new_new_n56884__, new_new_n56885__, new_new_n56886__,
    new_new_n56887__, new_new_n56888__, new_new_n56889__, new_new_n56890__,
    new_new_n56891__, new_new_n56892__, new_new_n56893__, new_new_n56894__,
    new_new_n56895__, new_new_n56896__, new_new_n56897__, new_new_n56898__,
    new_new_n56899__, new_new_n56900__, new_new_n56901__, new_new_n56902__,
    new_new_n56903__, new_new_n56904__, new_new_n56905__, new_new_n56906__,
    new_new_n56907__, new_new_n56908__, new_new_n56909__, new_new_n56910__,
    new_new_n56911__, new_new_n56912__, new_new_n56913__, new_new_n56914__,
    new_new_n56915__, new_new_n56916__, new_new_n56917__, new_new_n56918__,
    new_new_n56919__, new_new_n56920__, new_new_n56921__, new_new_n56922__,
    new_new_n56923__, new_new_n56924__, new_new_n56926__, new_new_n56927__,
    new_new_n56928__, new_new_n56929__, new_new_n56930__, new_new_n56931__,
    new_new_n56932__, new_new_n56933__, new_new_n56934__, new_new_n56936__,
    new_new_n56937__, new_new_n56938__, new_new_n56939__, new_new_n56940__,
    new_new_n56941__, new_new_n56942__, new_new_n56943__, new_new_n56944__,
    new_new_n56945__, new_new_n56946__, new_new_n56947__, new_new_n56948__,
    new_new_n56949__, new_new_n56950__, new_new_n56951__, new_new_n56952__,
    new_new_n56953__, new_new_n56954__, new_new_n56955__, new_new_n56956__,
    new_new_n56957__, new_new_n56958__, new_new_n56959__, new_new_n56960__,
    new_new_n56961__, new_new_n56962__, new_new_n56963__, new_new_n56964__,
    new_new_n56965__, new_new_n56966__, new_new_n56967__, new_new_n56968__,
    new_new_n56969__, new_new_n56970__, new_new_n56971__, new_new_n56972__,
    new_new_n56973__, new_new_n56974__, new_new_n56975__, new_new_n56976__,
    new_new_n56977__, new_new_n56978__, new_new_n56979__, new_new_n56980__,
    new_new_n56981__, new_new_n56982__, new_new_n56983__, new_new_n56984__,
    new_new_n56985__, new_new_n56986__, new_new_n56987__, new_new_n56988__,
    new_new_n56989__, new_new_n56990__, new_new_n56991__, new_new_n56992__,
    new_new_n56993__, new_new_n56994__, new_new_n56995__, new_new_n56996__,
    new_new_n56997__, new_new_n56998__, new_new_n56999__, new_new_n57000__,
    new_new_n57001__, new_new_n57002__, new_new_n57003__, new_new_n57004__,
    new_new_n57005__, new_new_n57006__, new_new_n57007__, new_new_n57008__,
    new_new_n57009__, new_new_n57010__, new_new_n57011__, new_new_n57012__,
    new_new_n57013__, new_new_n57014__, new_new_n57015__, new_new_n57016__,
    new_new_n57017__, new_new_n57018__, new_new_n57020__, new_new_n57021__,
    new_new_n57022__, new_new_n57023__, new_new_n57024__, new_new_n57025__,
    new_new_n57026__, new_new_n57027__, new_new_n57028__, new_new_n57030__,
    new_new_n57031__, new_new_n57032__, new_new_n57033__, new_new_n57034__,
    new_new_n57035__, new_new_n57036__, new_new_n57037__, new_new_n57038__,
    new_new_n57039__, new_new_n57040__, new_new_n57041__, new_new_n57042__,
    new_new_n57043__, new_new_n57044__, new_new_n57045__, new_new_n57046__,
    new_new_n57047__, new_new_n57048__, new_new_n57049__, new_new_n57050__,
    new_new_n57051__, new_new_n57052__, new_new_n57053__, new_new_n57054__,
    new_new_n57055__, new_new_n57056__, new_new_n57057__, new_new_n57058__,
    new_new_n57059__, new_new_n57060__, new_new_n57061__, new_new_n57062__,
    new_new_n57063__, new_new_n57064__, new_new_n57065__, new_new_n57066__,
    new_new_n57067__, new_new_n57068__, new_new_n57069__, new_new_n57070__,
    new_new_n57071__, new_new_n57072__, new_new_n57073__, new_new_n57074__,
    new_new_n57075__, new_new_n57076__, new_new_n57077__, new_new_n57078__,
    new_new_n57079__, new_new_n57080__, new_new_n57081__, new_new_n57082__,
    new_new_n57083__, new_new_n57084__, new_new_n57085__, new_new_n57086__,
    new_new_n57087__, new_new_n57088__, new_new_n57089__, new_new_n57090__,
    new_new_n57091__, new_new_n57092__, new_new_n57093__, new_new_n57094__,
    new_new_n57095__, new_new_n57096__, new_new_n57097__, new_new_n57098__,
    new_new_n57099__, new_new_n57100__, new_new_n57101__, new_new_n57102__,
    new_new_n57103__, new_new_n57104__, new_new_n57105__, new_new_n57106__,
    new_new_n57107__, new_new_n57108__, new_new_n57109__, new_new_n57110__,
    new_new_n57111__, new_new_n57112__, new_new_n57113__, new_new_n57114__,
    new_new_n57115__, new_new_n57116__, new_new_n57117__, new_new_n57118__,
    new_new_n57119__, new_new_n57120__, new_new_n57122__, new_new_n57123__,
    new_new_n57124__, new_new_n57125__, new_new_n57126__, new_new_n57127__,
    new_new_n57128__, new_new_n57129__, new_new_n57130__, new_new_n57132__,
    new_new_n57133__, new_new_n57134__, new_new_n57135__, new_new_n57136__,
    new_new_n57137__, new_new_n57138__, new_new_n57139__, new_new_n57140__,
    new_new_n57141__, new_new_n57142__, new_new_n57143__, new_new_n57144__,
    new_new_n57145__, new_new_n57146__, new_new_n57147__, new_new_n57148__,
    new_new_n57149__, new_new_n57150__, new_new_n57151__, new_new_n57152__,
    new_new_n57153__, new_new_n57154__, new_new_n57155__, new_new_n57156__,
    new_new_n57157__, new_new_n57158__, new_new_n57159__, new_new_n57160__,
    new_new_n57161__, new_new_n57162__, new_new_n57163__, new_new_n57164__,
    new_new_n57165__, new_new_n57166__, new_new_n57167__, new_new_n57168__,
    new_new_n57169__, new_new_n57170__, new_new_n57171__, new_new_n57172__,
    new_new_n57173__, new_new_n57174__, new_new_n57175__, new_new_n57176__,
    new_new_n57177__, new_new_n57178__, new_new_n57179__, new_new_n57180__,
    new_new_n57181__, new_new_n57182__, new_new_n57183__, new_new_n57184__,
    new_new_n57185__, new_new_n57186__, new_new_n57187__, new_new_n57188__,
    new_new_n57189__, new_new_n57190__, new_new_n57191__, new_new_n57192__,
    new_new_n57193__, new_new_n57194__, new_new_n57195__, new_new_n57196__,
    new_new_n57197__, new_new_n57198__, new_new_n57199__, new_new_n57200__,
    new_new_n57201__, new_new_n57202__, new_new_n57203__, new_new_n57204__,
    new_new_n57205__, new_new_n57206__, new_new_n57207__, new_new_n57208__,
    new_new_n57209__, new_new_n57211__, new_new_n57212__, new_new_n57213__,
    new_new_n57214__, new_new_n57215__, new_new_n57216__, new_new_n57217__,
    new_new_n57218__, new_new_n57219__, new_new_n57221__, new_new_n57222__,
    new_new_n57223__, new_new_n57224__, new_new_n57225__, new_new_n57226__,
    new_new_n57227__, new_new_n57228__, new_new_n57229__, new_new_n57230__,
    new_new_n57231__, new_new_n57232__, new_new_n57233__, new_new_n57235__,
    new_new_n57236__, new_new_n57238__, new_new_n57239__, new_new_n57240__,
    new_new_n57241__, new_new_n57242__, new_new_n57243__, new_new_n57244__,
    new_new_n57245__, new_new_n57246__, new_new_n57247__, new_new_n57248__,
    new_new_n57249__, new_new_n57250__, new_new_n57251__, new_new_n57252__,
    new_new_n57253__, new_new_n57254__, new_new_n57255__, new_new_n57256__,
    new_new_n57257__, new_new_n57258__, new_new_n57259__, new_new_n57260__,
    new_new_n57261__, new_new_n57262__, new_new_n57263__, new_new_n57264__,
    new_new_n57265__, new_new_n57266__, new_new_n57267__, new_new_n57268__,
    new_new_n57269__, new_new_n57270__, new_new_n57271__, new_new_n57272__,
    new_new_n57273__, new_new_n57274__, new_new_n57275__, new_new_n57276__,
    new_new_n57277__, new_new_n57278__, new_new_n57279__, new_new_n57280__,
    new_new_n57281__, new_new_n57282__, new_new_n57283__, new_new_n57284__,
    new_new_n57285__, new_new_n57286__, new_new_n57287__, new_new_n57288__,
    new_new_n57289__, new_new_n57290__, new_new_n57291__, new_new_n57292__,
    new_new_n57293__, new_new_n57295__, new_new_n57296__, new_new_n57298__,
    new_new_n57299__, new_new_n57300__, new_new_n57301__, new_new_n57302__,
    new_new_n57303__, new_new_n57304__, new_new_n57305__, new_new_n57306__,
    new_new_n57307__, new_new_n57308__, new_new_n57309__, new_new_n57310__,
    new_new_n57311__, new_new_n57312__, new_new_n57313__, new_new_n57314__,
    new_new_n57315__, new_new_n57316__, new_new_n57317__, new_new_n57318__,
    new_new_n57319__, new_new_n57320__, new_new_n57321__, new_new_n57322__,
    new_new_n57323__, new_new_n57324__, new_new_n57325__, new_new_n57326__,
    new_new_n57327__, new_new_n57328__, new_new_n57329__, new_new_n57330__,
    new_new_n57331__, new_new_n57332__, new_new_n57333__, new_new_n57334__,
    new_new_n57335__, new_new_n57336__, new_new_n57337__, new_new_n57338__,
    new_new_n57339__, new_new_n57340__, new_new_n57341__, new_new_n57342__,
    new_new_n57343__, new_new_n57344__, new_new_n57345__, new_new_n57346__,
    new_new_n57347__, new_new_n57348__, new_new_n57349__, new_new_n57350__,
    new_new_n57351__, new_new_n57352__, new_new_n57353__, new_new_n57354__,
    new_new_n57355__, new_new_n57356__, new_new_n57357__, new_new_n57358__,
    new_new_n57359__, new_new_n57360__, new_new_n57361__, new_new_n57362__,
    new_new_n57363__, new_new_n57364__, new_new_n57365__, new_new_n57366__,
    new_new_n57367__, new_new_n57368__, new_new_n57369__, new_new_n57370__,
    new_new_n57371__, new_new_n57372__, new_new_n57373__, new_new_n57374__,
    new_new_n57375__, new_new_n57376__, new_new_n57377__, new_new_n57378__,
    new_new_n57379__, new_new_n57380__, new_new_n57381__, new_new_n57382__,
    new_new_n57383__, new_new_n57384__, new_new_n57385__, new_new_n57387__,
    new_new_n57388__, new_new_n57389__, new_new_n57390__, new_new_n57391__,
    new_new_n57392__, new_new_n57393__, new_new_n57394__, new_new_n57395__,
    new_new_n57397__, new_new_n57398__, new_new_n57399__, new_new_n57400__,
    new_new_n57401__, new_new_n57402__, new_new_n57403__, new_new_n57404__,
    new_new_n57405__, new_new_n57406__, new_new_n57407__, new_new_n57408__,
    new_new_n57409__, new_new_n57411__, new_new_n57412__, new_new_n57414__,
    new_new_n57415__, new_new_n57416__, new_new_n57417__, new_new_n57418__,
    new_new_n57419__, new_new_n57420__, new_new_n57421__, new_new_n57422__,
    new_new_n57423__, new_new_n57424__, new_new_n57425__, new_new_n57426__,
    new_new_n57427__, new_new_n57428__, new_new_n57429__, new_new_n57430__,
    new_new_n57431__, new_new_n57432__, new_new_n57433__, new_new_n57434__,
    new_new_n57435__, new_new_n57436__, new_new_n57437__, new_new_n57438__,
    new_new_n57439__, new_new_n57440__, new_new_n57441__, new_new_n57442__,
    new_new_n57443__, new_new_n57445__, new_new_n57446__, new_new_n57448__,
    new_new_n57449__, new_new_n57450__, new_new_n57451__, new_new_n57452__,
    new_new_n57453__, new_new_n57454__, new_new_n57455__, new_new_n57456__,
    new_new_n57457__, new_new_n57458__, new_new_n57459__, new_new_n57460__,
    new_new_n57461__, new_new_n57462__, new_new_n57463__, new_new_n57464__,
    new_new_n57465__, new_new_n57466__, new_new_n57467__, new_new_n57468__,
    new_new_n57469__, new_new_n57470__, new_new_n57471__, new_new_n57472__,
    new_new_n57473__, new_new_n57474__, new_new_n57475__, new_new_n57476__,
    new_new_n57477__, new_new_n57479__, new_new_n57480__, new_new_n57482__,
    new_new_n57483__, new_new_n57484__, new_new_n57485__, new_new_n57486__,
    new_new_n57487__, new_new_n57488__, new_new_n57489__, new_new_n57490__,
    new_new_n57492__, new_new_n57493__, new_new_n57494__, new_new_n57495__,
    new_new_n57496__, new_new_n57497__, new_new_n57498__, new_new_n57499__,
    new_new_n57500__, new_new_n57501__, new_new_n57502__, new_new_n57503__,
    new_new_n57504__, new_new_n57505__, new_new_n57506__, new_new_n57507__,
    new_new_n57508__, new_new_n57509__, new_new_n57510__, new_new_n57512__,
    new_new_n57513__, new_new_n57515__, new_new_n57516__, new_new_n57518__,
    new_new_n57519__, new_new_n57523__, new_new_n57524__, new_new_n57525__,
    new_new_n57526__, new_new_n57527__, new_new_n57530__, new_new_n57531__,
    new_new_n57532__, new_new_n57533__, new_new_n57534__, new_new_n57535__,
    new_new_n57536__, new_new_n57537__, new_new_n57538__, new_new_n57542__,
    new_new_n57543__, new_new_n57544__, new_new_n57545__, new_new_n57546__,
    new_new_n57547__, new_new_n57548__, new_new_n57549__, new_new_n57550__,
    new_new_n57551__, new_new_n57552__, new_new_n57553__, new_new_n57555__,
    new_new_n57556__, new_new_n57559__, new_new_n57560__, new_new_n57561__,
    new_new_n57562__, new_new_n57563__, new_new_n57565__, new_new_n57567__,
    new_new_n57568__, new_new_n57569__, new_new_n57570__, new_new_n57571__,
    new_new_n57572__, new_new_n57573__, new_new_n57574__, new_new_n57575__,
    new_new_n57576__, new_new_n57577__, new_new_n57578__, new_new_n57579__,
    new_new_n57580__, new_new_n57581__, new_new_n57582__, new_new_n57583__,
    new_new_n57584__, new_new_n57585__, new_new_n57586__, new_new_n57587__,
    new_new_n57588__, new_new_n57589__, new_new_n57590__, new_new_n57591__,
    new_new_n57592__, new_new_n57593__, new_new_n57594__, new_new_n57595__,
    new_new_n57596__, new_new_n57597__, new_new_n57598__, new_new_n57599__,
    new_new_n57600__, new_new_n57601__, new_new_n57602__, new_new_n57603__,
    new_new_n57604__, new_new_n57605__, new_new_n57606__, new_new_n57607__,
    new_new_n57608__, new_new_n57609__, new_new_n57610__, new_new_n57611__,
    new_new_n57612__, new_new_n57613__, new_new_n57614__, new_new_n57615__,
    new_new_n57616__, new_new_n57617__, new_new_n57618__, new_new_n57619__,
    new_new_n57620__, new_new_n57621__, new_new_n57622__, new_new_n57623__,
    new_new_n57624__, new_new_n57625__, new_new_n57626__, new_new_n57627__,
    new_new_n57628__, new_new_n57629__, new_new_n57630__, new_new_n57631__,
    new_new_n57632__, new_new_n57633__, new_new_n57634__, new_new_n57635__,
    new_new_n57636__, new_new_n57637__, new_new_n57638__, new_new_n57639__,
    new_new_n57640__, new_new_n57641__, new_new_n57642__, new_new_n57643__,
    new_new_n57644__, new_new_n57645__, new_new_n57646__, new_new_n57647__,
    new_new_n57648__, new_new_n57649__, new_new_n57650__, new_new_n57651__,
    new_new_n57652__, new_new_n57653__, new_new_n57654__, new_new_n57655__,
    new_new_n57656__, new_new_n57657__, new_new_n57658__, new_new_n57659__,
    new_new_n57660__, new_new_n57661__, new_new_n57665__, new_new_n57666__,
    new_new_n57667__, new_new_n57668__, new_new_n57669__, new_new_n57670__,
    new_new_n57672__, new_new_n57674__, new_new_n57675__, new_new_n57677__,
    new_new_n57679__, new_new_n57681__, new_new_n57683__, new_new_n57685__,
    new_new_n57686__, new_new_n57687__, new_new_n57688__, new_new_n57689__,
    new_new_n57691__, new_new_n57692__, new_new_n57693__, new_new_n57695__,
    new_new_n57697__, new_new_n57698__, new_new_n57699__, new_new_n57700__,
    new_new_n57701__, new_new_n57703__, new_new_n57704__, new_new_n57705__,
    new_new_n57706__, new_new_n57707__, new_new_n57709__, new_new_n57711__,
    new_new_n57712__, new_new_n57714__, new_new_n57715__, new_new_n57717__,
    new_new_n57718__, new_new_n57719__, new_new_n57720__, new_new_n57721__,
    new_new_n57723__, new_new_n57724__, new_new_n57725__, new_new_n57726__,
    new_new_n57728__, new_new_n57729__, new_new_n57731__, new_new_n57732__,
    new_new_n57734__, new_new_n57735__, new_new_n57736__, new_new_n57737__,
    new_new_n57738__, new_new_n57740__, new_new_n57741__, new_new_n57742__,
    new_new_n57743__, new_new_n57744__, new_new_n57746__, new_new_n57747__,
    new_new_n57749__, new_new_n57750__, new_new_n57752__, new_new_n57753__,
    new_new_n57754__, new_new_n57755__, new_new_n57756__, new_new_n57758__,
    new_new_n57759__, new_new_n57760__, new_new_n57761__, new_new_n57762__,
    new_new_n57764__, new_new_n57765__, new_new_n57767__, new_new_n57768__,
    new_new_n57770__, new_new_n57771__, new_new_n57772__, new_new_n57773__,
    new_new_n57774__, new_new_n57776__, new_new_n57777__, new_new_n57778__,
    new_new_n57779__, new_new_n57780__, new_new_n57782__, new_new_n57783__,
    new_new_n57785__, new_new_n57786__, new_new_n57789__, new_new_n57791__,
    new_new_n57792__, new_new_n57794__, new_new_n57795__, new_new_n57797__,
    new_new_n57798__, new_new_n57799__, new_new_n57801__, new_new_n57802__,
    new_new_n57804__, new_new_n57805__, new_new_n57806__, new_new_n57808__,
    new_new_n57809__, new_new_n57810__, new_new_n57812__, new_new_n57813__,
    new_new_n57815__, new_new_n57816__, new_new_n57817__, new_new_n57818__,
    new_new_n57820__, new_new_n57821__, new_new_n57823__, new_new_n57824__,
    new_new_n57825__, new_new_n57826__, new_new_n57828__, new_new_n57829__,
    new_new_n57830__, new_new_n57831__, new_new_n57833__, new_new_n57834__,
    new_new_n57835__, new_new_n57836__, new_new_n57838__, new_new_n57839__,
    new_new_n57841__, new_new_n57842__, new_new_n57843__, new_new_n57844__,
    new_new_n57846__, new_new_n57847__, new_new_n57848__, new_new_n57849__,
    new_new_n57851__, new_new_n57852__, new_new_n57853__, new_new_n57854__,
    new_new_n57856__, new_new_n57857__, new_new_n57858__, new_new_n57859__,
    new_new_n57861__, new_new_n57862__, new_new_n57863__, new_new_n57864__,
    new_new_n57866__, new_new_n57867__, new_new_n57868__, new_new_n57869__,
    new_new_n57871__, new_new_n57872__, new_new_n57873__, new_new_n57874__,
    new_new_n98_9_, new_new_n99_9_, new_new_n101_9_, new_new_n102_9_,
    new_new_n104_9_, new_new_n105_9_, new_new_n107_9_, new_new_n108_9_,
    new_new_n110_9_, new_new_n111_9_, new_new_n113_9_, new_new_n114_9_,
    new_new_n116_9_, new_new_n117_9_, new_new_n119_9_, new_new_n120_9_,
    new_new_n122_9_, new_new_n123_9_, new_new_n125_9_, new_new_n126_9_,
    new_new_n128_9_, new_new_n129_9_, new_new_n131_9_, new_new_n132_9_,
    new_new_n134_9_, new_new_n135_9_, new_new_n137_9_, new_new_n138_9_,
    new_new_n140_9_, new_new_n141_9_, new_new_n143_9_, new_new_n144_9_,
    new_new_n146_9_, new_new_n147_9_, new_new_n149_9_, new_new_n150_9_,
    new_new_n152_9_, new_new_n153_9_, new_new_n155_9_, new_new_n156_9_,
    new_new_n158_9_, new_new_n159_9_, new_new_n161_9_, new_new_n162_9_,
    new_new_n164_9_, new_new_n165_9_, new_new_n167_9_, new_new_n168_9_,
    new_new_n170_9_, new_new_n171_9_, new_new_n173_9_, new_new_n174_9_,
    new_new_n176_9_, new_new_n177_9_, new_new_n179_9_, new_new_n180_9_,
    new_new_n182_9_, new_new_n183_9_, new_new_n185_9_, new_new_n186_9_,
    new_new_n188_9_, new_new_n189_9_, new_new_n191_9_, new_new_n192_9_;
  assign ys__n33337 = ~ys__n33336;
  assign new_new_n98__ = ys__n29119 & ~ys__n29121;
  assign new_new_n99__ = ys__n29120 & ys__n29121;
  assign ys__n29122 = new_new_n98__ | new_new_n99__;
  assign new_new_n101__ = ~ys__n29121 & ys__n29123;
  assign new_new_n102__ = ys__n29121 & ys__n29124;
  assign ys__n29125 = new_new_n101__ | new_new_n102__;
  assign new_new_n104__ = ~ys__n29121 & ys__n29126;
  assign new_new_n105__ = ys__n29121 & ys__n29127;
  assign ys__n29128 = new_new_n104__ | new_new_n105__;
  assign new_new_n107__ = ~ys__n29121 & ys__n29129;
  assign new_new_n108__ = ys__n29121 & ys__n29130;
  assign ys__n29131 = new_new_n107__ | new_new_n108__;
  assign new_new_n110__ = ~ys__n29121 & ys__n29132;
  assign new_new_n111__ = ys__n29121 & ys__n29133;
  assign ys__n29134 = new_new_n110__ | new_new_n111__;
  assign new_new_n113__ = ~ys__n29121 & ys__n29135;
  assign new_new_n114__ = ys__n29121 & ys__n29136;
  assign ys__n29137 = new_new_n113__ | new_new_n114__;
  assign new_new_n116__ = ~ys__n29121 & ys__n29138;
  assign new_new_n117__ = ys__n29121 & ys__n29139;
  assign ys__n29140 = new_new_n116__ | new_new_n117__;
  assign new_new_n119__ = ~ys__n29121 & ys__n29141;
  assign new_new_n120__ = ys__n29121 & ys__n29142;
  assign ys__n29143 = new_new_n119__ | new_new_n120__;
  assign new_new_n122__ = ~ys__n29121 & ys__n29144;
  assign new_new_n123__ = ys__n29121 & ys__n29145;
  assign ys__n29146 = new_new_n122__ | new_new_n123__;
  assign new_new_n125__ = ~ys__n29121 & ys__n29147;
  assign new_new_n126__ = ys__n29121 & ys__n29148;
  assign ys__n29149 = new_new_n125__ | new_new_n126__;
  assign new_new_n128__ = ~ys__n29121 & ys__n29150;
  assign new_new_n129__ = ys__n29121 & ys__n29151;
  assign ys__n29152 = new_new_n128__ | new_new_n129__;
  assign new_new_n131__ = ~ys__n29121 & ys__n29153;
  assign new_new_n132__ = ys__n29121 & ys__n29154;
  assign ys__n29155 = new_new_n131__ | new_new_n132__;
  assign new_new_n134__ = ~ys__n29121 & ys__n29156;
  assign new_new_n135__ = ys__n29121 & ys__n29157;
  assign ys__n29158 = new_new_n134__ | new_new_n135__;
  assign new_new_n137__ = ~ys__n29121 & ys__n29159;
  assign new_new_n138__ = ys__n29121 & ys__n29160;
  assign ys__n29161 = new_new_n137__ | new_new_n138__;
  assign new_new_n140__ = ~ys__n29121 & ys__n29162;
  assign new_new_n141__ = ys__n29121 & ys__n29163;
  assign ys__n29164 = new_new_n140__ | new_new_n141__;
  assign new_new_n143__ = ~ys__n29121 & ys__n29165;
  assign new_new_n144__ = ys__n29121 & ys__n29166;
  assign ys__n29167 = new_new_n143__ | new_new_n144__;
  assign new_new_n146__ = ~ys__n29121 & ys__n29168;
  assign new_new_n147__ = ys__n29121 & ys__n29169;
  assign ys__n29170 = new_new_n146__ | new_new_n147__;
  assign new_new_n149__ = ~ys__n29121 & ys__n29171;
  assign new_new_n150__ = ys__n29121 & ys__n29172;
  assign ys__n29173 = new_new_n149__ | new_new_n150__;
  assign new_new_n152__ = ~ys__n29121 & ys__n29174;
  assign new_new_n153__ = ys__n29121 & ys__n29175;
  assign ys__n29176 = new_new_n152__ | new_new_n153__;
  assign new_new_n155__ = ~ys__n29121 & ys__n29177;
  assign new_new_n156__ = ys__n29121 & ys__n29178;
  assign ys__n29179 = new_new_n155__ | new_new_n156__;
  assign new_new_n158__ = ~ys__n29121 & ys__n29180;
  assign new_new_n159__ = ys__n29121 & ys__n29181;
  assign ys__n29182 = new_new_n158__ | new_new_n159__;
  assign new_new_n161__ = ~ys__n29121 & ys__n29183;
  assign new_new_n162__ = ys__n29121 & ys__n29184;
  assign ys__n29185 = new_new_n161__ | new_new_n162__;
  assign new_new_n164__ = ~ys__n29121 & ys__n29186;
  assign new_new_n165__ = ys__n29121 & ys__n29187;
  assign ys__n29188 = new_new_n164__ | new_new_n165__;
  assign new_new_n167__ = ~ys__n29121 & ys__n29189;
  assign new_new_n168__ = ys__n29121 & ys__n29190;
  assign ys__n29191 = new_new_n167__ | new_new_n168__;
  assign new_new_n170__ = ~ys__n29121 & ys__n29192;
  assign new_new_n171__ = ys__n29121 & ys__n29193;
  assign ys__n29194 = new_new_n170__ | new_new_n171__;
  assign new_new_n173__ = ~ys__n29121 & ys__n29195;
  assign new_new_n174__ = ys__n29121 & ys__n29196;
  assign ys__n29197 = new_new_n173__ | new_new_n174__;
  assign new_new_n176__ = ~ys__n29121 & ys__n29198;
  assign new_new_n177__ = ys__n29121 & ys__n29199;
  assign ys__n29200 = new_new_n176__ | new_new_n177__;
  assign new_new_n179__ = ~ys__n29121 & ys__n29201;
  assign new_new_n180__ = ys__n29121 & ys__n29202;
  assign ys__n29203 = new_new_n179__ | new_new_n180__;
  assign new_new_n182__ = ~ys__n29121 & ys__n29204;
  assign new_new_n183__ = ys__n29121 & ys__n29205;
  assign ys__n29206 = new_new_n182__ | new_new_n183__;
  assign new_new_n185__ = ~ys__n29121 & ys__n29207;
  assign new_new_n186__ = ys__n29121 & ys__n29208;
  assign ys__n29209 = new_new_n185__ | new_new_n186__;
  assign new_new_n188__ = ~ys__n29121 & ys__n29210;
  assign new_new_n189__ = ys__n29121 & ys__n29211;
  assign ys__n29212 = new_new_n188__ | new_new_n189__;
  assign new_new_n191__ = ~ys__n29121 & ys__n29213;
  assign new_new_n192__ = ys__n29121 & ys__n29214;
  assign ys__n29215 = new_new_n191__ | new_new_n192__;
  assign ys__n33335 = ~ys__n33334;
  assign ys__n33329 = ~ys__n33328;
  assign ys__n33331 = ~ys__n33330;
  assign new_new_n98_5_ = ys__n29432 & ~ys__n29434;
  assign new_new_n99_5_ = ys__n29433 & ys__n29434;
  assign ys__n29435 = new_new_n98_5_ | new_new_n99_5_;
  assign new_new_n101_5_ = ~ys__n29434 & ys__n29436;
  assign new_new_n102_5_ = ys__n29434 & ys__n29437;
  assign ys__n29438 = new_new_n101_5_ | new_new_n102_5_;
  assign new_new_n104_5_ = ~ys__n29434 & ys__n29439;
  assign new_new_n105_5_ = ys__n29434 & ys__n29440;
  assign ys__n29441 = new_new_n104_5_ | new_new_n105_5_;
  assign new_new_n107_5_ = ~ys__n29434 & ys__n29442;
  assign new_new_n108_5_ = ys__n29434 & ys__n29443;
  assign ys__n29444 = new_new_n107_5_ | new_new_n108_5_;
  assign new_new_n110_5_ = ~ys__n29434 & ys__n29445;
  assign new_new_n111_5_ = ys__n29434 & ys__n29446;
  assign ys__n29447 = new_new_n110_5_ | new_new_n111_5_;
  assign new_new_n113_5_ = ~ys__n29434 & ys__n29448;
  assign new_new_n114_5_ = ys__n29434 & ys__n29449;
  assign ys__n29450 = new_new_n113_5_ | new_new_n114_5_;
  assign new_new_n116_5_ = ~ys__n29434 & ys__n29451;
  assign new_new_n117_5_ = ys__n29434 & ys__n29452;
  assign ys__n29453 = new_new_n116_5_ | new_new_n117_5_;
  assign new_new_n119_5_ = ~ys__n29434 & ys__n29454;
  assign new_new_n120_5_ = ys__n29434 & ys__n29455;
  assign ys__n29456 = new_new_n119_5_ | new_new_n120_5_;
  assign new_new_n122_5_ = ~ys__n29434 & ys__n29457;
  assign new_new_n123_5_ = ys__n29434 & ys__n29458;
  assign ys__n29459 = new_new_n122_5_ | new_new_n123_5_;
  assign new_new_n125_5_ = ~ys__n29434 & ys__n29460;
  assign new_new_n126_5_ = ys__n29434 & ys__n29461;
  assign ys__n29462 = new_new_n125_5_ | new_new_n126_5_;
  assign new_new_n128_5_ = ~ys__n29434 & ys__n29463;
  assign new_new_n129_5_ = ys__n29434 & ys__n29464;
  assign ys__n29465 = new_new_n128_5_ | new_new_n129_5_;
  assign new_new_n131_5_ = ~ys__n29434 & ys__n29466;
  assign new_new_n132_5_ = ys__n29434 & ys__n29467;
  assign ys__n29468 = new_new_n131_5_ | new_new_n132_5_;
  assign new_new_n134_5_ = ~ys__n29434 & ys__n29469;
  assign new_new_n135_5_ = ys__n29434 & ys__n29470;
  assign ys__n29471 = new_new_n134_5_ | new_new_n135_5_;
  assign new_new_n137_5_ = ~ys__n29434 & ys__n29472;
  assign new_new_n138_5_ = ys__n29434 & ys__n29473;
  assign ys__n29474 = new_new_n137_5_ | new_new_n138_5_;
  assign new_new_n140_5_ = ~ys__n29434 & ys__n29475;
  assign new_new_n141_5_ = ys__n29434 & ys__n29476;
  assign ys__n29477 = new_new_n140_5_ | new_new_n141_5_;
  assign new_new_n143_5_ = ~ys__n29434 & ys__n29478;
  assign new_new_n144_5_ = ys__n29434 & ys__n29479;
  assign ys__n29480 = new_new_n143_5_ | new_new_n144_5_;
  assign new_new_n146_5_ = ~ys__n29434 & ys__n29481;
  assign new_new_n147_5_ = ys__n29434 & ys__n29482;
  assign ys__n29483 = new_new_n146_5_ | new_new_n147_5_;
  assign new_new_n149_5_ = ~ys__n29434 & ys__n29484;
  assign new_new_n150_5_ = ys__n29434 & ys__n29485;
  assign ys__n29486 = new_new_n149_5_ | new_new_n150_5_;
  assign new_new_n152_5_ = ~ys__n29434 & ys__n29487;
  assign new_new_n153_5_ = ys__n29434 & ys__n29488;
  assign ys__n29489 = new_new_n152_5_ | new_new_n153_5_;
  assign new_new_n155_5_ = ~ys__n29434 & ys__n29490;
  assign new_new_n156_5_ = ys__n29434 & ys__n29491;
  assign ys__n29492 = new_new_n155_5_ | new_new_n156_5_;
  assign new_new_n158_5_ = ~ys__n29434 & ys__n29493;
  assign new_new_n159_5_ = ys__n29434 & ys__n29494;
  assign ys__n29495 = new_new_n158_5_ | new_new_n159_5_;
  assign new_new_n161_5_ = ~ys__n29434 & ys__n29496;
  assign new_new_n162_5_ = ys__n29434 & ys__n29497;
  assign ys__n29498 = new_new_n161_5_ | new_new_n162_5_;
  assign new_new_n164_5_ = ~ys__n29434 & ys__n29499;
  assign new_new_n165_5_ = ys__n29434 & ys__n29500;
  assign ys__n29501 = new_new_n164_5_ | new_new_n165_5_;
  assign new_new_n167_5_ = ~ys__n29434 & ys__n29502;
  assign new_new_n168_5_ = ys__n29434 & ys__n29503;
  assign ys__n29504 = new_new_n167_5_ | new_new_n168_5_;
  assign new_new_n170_5_ = ~ys__n29434 & ys__n29505;
  assign new_new_n171_5_ = ys__n29434 & ys__n29506;
  assign ys__n29507 = new_new_n170_5_ | new_new_n171_5_;
  assign new_new_n173_5_ = ~ys__n29434 & ys__n29508;
  assign new_new_n174_5_ = ys__n29434 & ys__n29509;
  assign ys__n29510 = new_new_n173_5_ | new_new_n174_5_;
  assign new_new_n176_5_ = ~ys__n29434 & ys__n29511;
  assign new_new_n177_5_ = ys__n29434 & ys__n29512;
  assign ys__n29513 = new_new_n176_5_ | new_new_n177_5_;
  assign new_new_n179_5_ = ~ys__n29434 & ys__n29514;
  assign new_new_n180_5_ = ys__n29434 & ys__n29515;
  assign ys__n29516 = new_new_n179_5_ | new_new_n180_5_;
  assign new_new_n182_5_ = ~ys__n29434 & ys__n29517;
  assign new_new_n183_5_ = ys__n29434 & ys__n29518;
  assign ys__n29519 = new_new_n182_5_ | new_new_n183_5_;
  assign new_new_n185_5_ = ~ys__n29434 & ys__n29520;
  assign new_new_n186_5_ = ys__n29434 & ys__n29521;
  assign ys__n29522 = new_new_n185_5_ | new_new_n186_5_;
  assign new_new_n188_5_ = ~ys__n29434 & ys__n29523;
  assign new_new_n189_5_ = ys__n29434 & ys__n29524;
  assign ys__n29525 = new_new_n188_5_ | new_new_n189_5_;
  assign new_new_n191_5_ = ~ys__n29434 & ys__n29526;
  assign new_new_n192_5_ = ys__n29434 & ys__n29527;
  assign ys__n29528 = new_new_n191_5_ | new_new_n192_5_;
  assign new_new_n10398__ = ~ys__n35124 & ~ys__n35727;
  assign new_new_n10399__ = ys__n35124 & ys__n35727;
  assign new_new_n10400__ = ~new_new_n10398__ & ~new_new_n10399__;
  assign new_new_n10401__ = ~ys__n35122 & ~ys__n35725;
  assign new_new_n10402__ = ys__n35122 & ys__n35725;
  assign new_new_n10403__ = ~new_new_n10401__ & ~new_new_n10402__;
  assign new_new_n10404__ = ~new_new_n10400__ & ~new_new_n10403__;
  assign new_new_n10405__ = ~ys__n35120 & ~ys__n35723;
  assign new_new_n10406__ = ys__n35120 & ys__n35723;
  assign new_new_n10407__ = ~new_new_n10405__ & ~new_new_n10406__;
  assign new_new_n10408__ = ~ys__n35118 & ~ys__n35721;
  assign new_new_n10409__ = ys__n35118 & ys__n35721;
  assign new_new_n10410__ = ~new_new_n10408__ & ~new_new_n10409__;
  assign new_new_n10411__ = ~new_new_n10407__ & ~new_new_n10410__;
  assign new_new_n10412__ = new_new_n10404__ & new_new_n10411__;
  assign new_new_n10413__ = ~ys__n35116 & ~ys__n35719;
  assign new_new_n10414__ = ys__n35116 & ys__n35719;
  assign new_new_n10415__ = ~new_new_n10413__ & ~new_new_n10414__;
  assign new_new_n10416__ = ~ys__n35114 & ~ys__n35717;
  assign new_new_n10417__ = ys__n35114 & ys__n35717;
  assign new_new_n10418__ = ~new_new_n10416__ & ~new_new_n10417__;
  assign new_new_n10419__ = ~new_new_n10415__ & ~new_new_n10418__;
  assign new_new_n10420__ = ~ys__n24207 & ~ys__n35112;
  assign new_new_n10421__ = ys__n24207 & ys__n35112;
  assign new_new_n10422__ = ~new_new_n10420__ & ~new_new_n10421__;
  assign new_new_n10423__ = ~ys__n24205 & ~ys__n35110;
  assign new_new_n10424__ = ys__n24205 & ys__n35110;
  assign new_new_n10425__ = ~new_new_n10423__ & ~new_new_n10424__;
  assign new_new_n10426__ = ~new_new_n10422__ & ~new_new_n10425__;
  assign new_new_n10427__ = new_new_n10419__ & new_new_n10426__;
  assign new_new_n10428__ = ~ys__n24203 & ~ys__n35108;
  assign new_new_n10429__ = ys__n24203 & ys__n35108;
  assign new_new_n10430__ = ~new_new_n10428__ & ~new_new_n10429__;
  assign new_new_n10431__ = ~ys__n24201 & ~ys__n35106;
  assign new_new_n10432__ = ys__n24201 & ys__n35106;
  assign new_new_n10433__ = ~new_new_n10431__ & ~new_new_n10432__;
  assign new_new_n10434__ = ~new_new_n10430__ & ~new_new_n10433__;
  assign new_new_n10435__ = ys__n24199 & ~ys__n35104;
  assign new_new_n10436__ = ~ys__n24199 & ~ys__n35104;
  assign new_new_n10437__ = ys__n24199 & ys__n35104;
  assign new_new_n10438__ = ~new_new_n10436__ & ~new_new_n10437__;
  assign new_new_n10439__ = ys__n24197 & ~ys__n35102;
  assign new_new_n10440__ = ~ys__n24197 & ~ys__n35102;
  assign new_new_n10441__ = ys__n24197 & ys__n35102;
  assign new_new_n10442__ = ~new_new_n10440__ & ~new_new_n10441__;
  assign new_new_n10443__ = ~new_new_n10439__ & new_new_n10442__;
  assign new_new_n10444__ = ~new_new_n10438__ & ~new_new_n10443__;
  assign new_new_n10445__ = ~new_new_n10435__ & ~new_new_n10444__;
  assign new_new_n10446__ = new_new_n10434__ & ~new_new_n10445__;
  assign new_new_n10447__ = ys__n24203 & ~ys__n35108;
  assign new_new_n10448__ = ys__n24201 & ~ys__n35106;
  assign new_new_n10449__ = ~new_new_n10430__ & new_new_n10448__;
  assign new_new_n10450__ = ~new_new_n10447__ & ~new_new_n10449__;
  assign new_new_n10451__ = ~new_new_n10446__ & new_new_n10450__;
  assign new_new_n10452__ = new_new_n10427__ & ~new_new_n10451__;
  assign new_new_n10453__ = ys__n24207 & ~ys__n35112;
  assign new_new_n10454__ = ys__n24205 & ~ys__n35110;
  assign new_new_n10455__ = ~new_new_n10422__ & new_new_n10454__;
  assign new_new_n10456__ = ~new_new_n10453__ & ~new_new_n10455__;
  assign new_new_n10457__ = new_new_n10419__ & ~new_new_n10456__;
  assign new_new_n10458__ = ~ys__n35116 & ys__n35719;
  assign new_new_n10459__ = ~ys__n35114 & ys__n35717;
  assign new_new_n10460__ = ~new_new_n10415__ & new_new_n10459__;
  assign new_new_n10461__ = ~new_new_n10458__ & ~new_new_n10460__;
  assign new_new_n10462__ = ~new_new_n10457__ & new_new_n10461__;
  assign new_new_n10463__ = ~new_new_n10452__ & new_new_n10462__;
  assign new_new_n10464__ = new_new_n10412__ & ~new_new_n10463__;
  assign new_new_n10465__ = ~ys__n35120 & ys__n35723;
  assign new_new_n10466__ = ~ys__n35118 & ys__n35721;
  assign new_new_n10467__ = ~new_new_n10407__ & new_new_n10466__;
  assign new_new_n10468__ = ~new_new_n10465__ & ~new_new_n10467__;
  assign new_new_n10469__ = new_new_n10404__ & ~new_new_n10468__;
  assign new_new_n10470__ = ~ys__n35124 & ys__n35727;
  assign new_new_n10471__ = ~ys__n35122 & ys__n35725;
  assign new_new_n10472__ = ~new_new_n10400__ & new_new_n10471__;
  assign new_new_n10473__ = ~new_new_n10470__ & ~new_new_n10472__;
  assign new_new_n10474__ = ~new_new_n10469__ & new_new_n10473__;
  assign new_new_n10475__ = ~new_new_n10464__ & new_new_n10474__;
  assign new_new_n10476__ = ~new_new_n10438__ & ~new_new_n10442__;
  assign new_new_n10477__ = new_new_n10434__ & new_new_n10476__;
  assign new_new_n10478__ = new_new_n10412__ & new_new_n10477__;
  assign new_new_n10479__ = new_new_n10427__ & new_new_n10478__;
  assign new_new_n10480__ = ~new_new_n10475__ & ~new_new_n10479__;
  assign new_new_n10481__ = ~ys__n33265 & ~ys__n35723;
  assign new_new_n10482__ = ys__n33265 & ys__n35723;
  assign new_new_n10483__ = ~new_new_n10481__ & ~new_new_n10482__;
  assign new_new_n10484__ = ~ys__n33263 & ~ys__n35721;
  assign new_new_n10485__ = ys__n33263 & ys__n35721;
  assign new_new_n10486__ = ~new_new_n10484__ & ~new_new_n10485__;
  assign new_new_n10487__ = ~new_new_n10483__ & ~new_new_n10486__;
  assign new_new_n10488__ = ~ys__n33269 & ~ys__n35727;
  assign new_new_n10489__ = ys__n33269 & ys__n35727;
  assign new_new_n10490__ = ~new_new_n10488__ & ~new_new_n10489__;
  assign new_new_n10491__ = ~ys__n33267 & ~ys__n35725;
  assign new_new_n10492__ = ys__n33267 & ys__n35725;
  assign new_new_n10493__ = ~new_new_n10491__ & ~new_new_n10492__;
  assign new_new_n10494__ = ~new_new_n10490__ & ~new_new_n10493__;
  assign new_new_n10495__ = ~ys__n33261 & ~ys__n35719;
  assign new_new_n10496__ = ys__n33261 & ys__n35719;
  assign new_new_n10497__ = ~new_new_n10495__ & ~new_new_n10496__;
  assign new_new_n10498__ = ~ys__n33259 & ~ys__n35717;
  assign new_new_n10499__ = ys__n33259 & ys__n35717;
  assign new_new_n10500__ = ~new_new_n10498__ & ~new_new_n10499__;
  assign new_new_n10501__ = ~new_new_n10497__ & ~new_new_n10500__;
  assign new_new_n10502__ = new_new_n10494__ & new_new_n10501__;
  assign new_new_n10503__ = new_new_n10487__ & new_new_n10502__;
  assign new_new_n10504__ = ~ys__n33261 & ys__n35719;
  assign new_new_n10505__ = ~ys__n33259 & ys__n35717;
  assign new_new_n10506__ = new_new_n10500__ & ~new_new_n10505__;
  assign new_new_n10507__ = ~new_new_n10497__ & ~new_new_n10506__;
  assign new_new_n10508__ = ~new_new_n10504__ & ~new_new_n10507__;
  assign new_new_n10509__ = new_new_n10487__ & ~new_new_n10508__;
  assign new_new_n10510__ = ~ys__n33265 & ys__n35723;
  assign new_new_n10511__ = ~ys__n33263 & ys__n35721;
  assign new_new_n10512__ = ~new_new_n10483__ & new_new_n10511__;
  assign new_new_n10513__ = ~new_new_n10510__ & ~new_new_n10512__;
  assign new_new_n10514__ = ~new_new_n10509__ & new_new_n10513__;
  assign new_new_n10515__ = new_new_n10494__ & ~new_new_n10514__;
  assign new_new_n10516__ = ~ys__n33269 & ys__n35727;
  assign new_new_n10517__ = ~ys__n33267 & ys__n35725;
  assign new_new_n10518__ = ~new_new_n10490__ & new_new_n10517__;
  assign new_new_n10519__ = ~new_new_n10516__ & ~new_new_n10518__;
  assign new_new_n10520__ = ~new_new_n10515__ & new_new_n10519__;
  assign new_new_n10521__ = ~new_new_n10503__ & ~new_new_n10520__;
  assign new_new_n10522__ = ~new_new_n10503__ & ~new_new_n10521__;
  assign new_new_n10523__ = ys__n128 & ~ys__n38605;
  assign new_new_n10524__ = ~ys__n38606 & ys__n38607;
  assign new_new_n10525__ = ~new_new_n10523__ & ~new_new_n10524__;
  assign new_new_n10526__ = ys__n38606 & ~ys__n38607;
  assign new_new_n10527__ = ~ys__n38608 & ys__n38609;
  assign new_new_n10528__ = ~new_new_n10526__ & ~new_new_n10527__;
  assign new_new_n10529__ = new_new_n10525__ & new_new_n10528__;
  assign new_new_n10530__ = ys__n132 & ~ys__n38603;
  assign new_new_n10531__ = ~ys__n130 & ys__n38604;
  assign new_new_n10532__ = ~new_new_n10530__ & ~new_new_n10531__;
  assign new_new_n10533__ = ys__n130 & ~ys__n38604;
  assign new_new_n10534__ = ~ys__n128 & ys__n38605;
  assign new_new_n10535__ = ~new_new_n10533__ & ~new_new_n10534__;
  assign new_new_n10536__ = new_new_n10532__ & new_new_n10535__;
  assign new_new_n10537__ = new_new_n10529__ & new_new_n10536__;
  assign new_new_n10538__ = ys__n130 & ys__n132;
  assign new_new_n10539__ = ys__n134 & ys__n136;
  assign new_new_n10540__ = new_new_n10538__ & new_new_n10539__;
  assign new_new_n10541__ = ys__n122 & ys__n124;
  assign new_new_n10542__ = ys__n126 & ys__n128;
  assign new_new_n10543__ = new_new_n10541__ & new_new_n10542__;
  assign new_new_n10544__ = new_new_n10540__ & new_new_n10543__;
  assign new_new_n10545__ = ys__n38610 & ~ys__n38611;
  assign new_new_n10546__ = ys__n38608 & ~ys__n38609;
  assign new_new_n10547__ = ~ys__n38610 & ys__n38611;
  assign new_new_n10548__ = ~new_new_n10546__ & ~new_new_n10547__;
  assign new_new_n10549__ = ~new_new_n10545__ & new_new_n10548__;
  assign new_new_n10550__ = ~new_new_n10544__ & new_new_n10549__;
  assign new_new_n10551__ = new_new_n10537__ & new_new_n10550__;
  assign new_new_n10552__ = ~ys__n38585 & ys__n38586;
  assign new_new_n10553__ = ~ys__n38557 & ~new_new_n10552__;
  assign new_new_n10554__ = ys__n38585 & ~ys__n38586;
  assign new_new_n10555__ = ~ys__n38587 & ys__n38588;
  assign new_new_n10556__ = ~new_new_n10554__ & ~new_new_n10555__;
  assign new_new_n10557__ = ys__n38587 & ~ys__n38588;
  assign new_new_n10558__ = ~ys__n38589 & ys__n38590;
  assign new_new_n10559__ = ~new_new_n10557__ & ~new_new_n10558__;
  assign new_new_n10560__ = new_new_n10556__ & new_new_n10559__;
  assign new_new_n10561__ = new_new_n10553__ & new_new_n10560__;
  assign new_new_n10562__ = ys__n38593 & ~ys__n38594;
  assign new_new_n10563__ = ~ys__n38595 & ys__n38596;
  assign new_new_n10564__ = ~new_new_n10562__ & ~new_new_n10563__;
  assign new_new_n10565__ = ys__n38595 & ~ys__n38596;
  assign new_new_n10566__ = ~ys__n38597 & ys__n38598;
  assign new_new_n10567__ = ~new_new_n10565__ & ~new_new_n10566__;
  assign new_new_n10568__ = new_new_n10564__ & new_new_n10567__;
  assign new_new_n10569__ = ys__n38589 & ~ys__n38590;
  assign new_new_n10570__ = ~ys__n38591 & ys__n38592;
  assign new_new_n10571__ = ~new_new_n10569__ & ~new_new_n10570__;
  assign new_new_n10572__ = ys__n38591 & ~ys__n38592;
  assign new_new_n10573__ = ~ys__n38593 & ys__n38594;
  assign new_new_n10574__ = ~new_new_n10572__ & ~new_new_n10573__;
  assign new_new_n10575__ = new_new_n10571__ & new_new_n10574__;
  assign new_new_n10576__ = new_new_n10568__ & new_new_n10575__;
  assign new_new_n10577__ = ys__n136 & ~ys__n38601;
  assign new_new_n10578__ = ~ys__n134 & ys__n38602;
  assign new_new_n10579__ = ~new_new_n10577__ & ~new_new_n10578__;
  assign new_new_n10580__ = ys__n134 & ~ys__n38602;
  assign new_new_n10581__ = ~ys__n132 & ys__n38603;
  assign new_new_n10582__ = ~new_new_n10580__ & ~new_new_n10581__;
  assign new_new_n10583__ = new_new_n10579__ & new_new_n10582__;
  assign new_new_n10584__ = ys__n38597 & ~ys__n38598;
  assign new_new_n10585__ = ~ys__n38599 & ys__n38600;
  assign new_new_n10586__ = ~new_new_n10584__ & ~new_new_n10585__;
  assign new_new_n10587__ = ys__n38599 & ~ys__n38600;
  assign new_new_n10588__ = ~ys__n136 & ys__n38601;
  assign new_new_n10589__ = ~new_new_n10587__ & ~new_new_n10588__;
  assign new_new_n10590__ = new_new_n10586__ & new_new_n10589__;
  assign new_new_n10591__ = new_new_n10583__ & new_new_n10590__;
  assign new_new_n10592__ = new_new_n10576__ & new_new_n10591__;
  assign new_new_n10593__ = new_new_n10561__ & new_new_n10592__;
  assign new_new_n10594__ = new_new_n10551__ & new_new_n10593__;
  assign new_new_n10595__ = ~new_new_n10522__ & new_new_n10594__;
  assign new_new_n10596__ = ~new_new_n10480__ & new_new_n10595__;
  assign new_new_n10597__ = ys__n1072 & new_new_n10596__;
  assign new_new_n10598__ = ~ys__n4613 & ~new_new_n10597__;
  assign new_new_n10599__ = ~ys__n4185 & ~new_new_n10598__;
  assign new_new_n10600__ = ys__n1029 & ~ys__n24131;
  assign new_new_n10601__ = ~new_new_n10599__ & new_new_n10600__;
  assign new_new_n10602__ = ys__n1072 & ~ys__n4185;
  assign new_new_n10603__ = new_new_n10596__ & new_new_n10602__;
  assign new_new_n10604__ = ys__n29897 & ~new_new_n10603__;
  assign new_new_n10605__ = ~new_new_n10601__ & new_new_n10604__;
  assign ys__n4192 = ys__n4185 | ys__n4613;
  assign new_new_n10607__ = ~ys__n4184 & ~ys__n4190;
  assign new_new_n10608__ = ~ys__n4192 & new_new_n10607__;
  assign new_new_n10609__ = ~ys__n4625 & ~ys__n4627;
  assign new_new_n10610__ = ~ys__n4176 & ~ys__n4698;
  assign new_new_n10611__ = new_new_n10609__ & new_new_n10610__;
  assign new_new_n10612__ = new_new_n10608__ & new_new_n10611__;
  assign new_new_n10613__ = ~ys__n846 & ~ys__n4177;
  assign ys__n738 = ~new_new_n10612__ | ~new_new_n10613__;
  assign new_new_n10615__ = ys__n23339 & ~ys__n738;
  assign new_new_n10616__ = ys__n23763 & ys__n738;
  assign ys__n23764 = new_new_n10615__ | new_new_n10616__;
  assign new_new_n10618__ = new_new_n10605__ & ~ys__n23764;
  assign new_new_n10619__ = ys__n29913 & ~new_new_n10603__;
  assign new_new_n10620__ = ~new_new_n10601__ & new_new_n10619__;
  assign new_new_n10621__ = ys__n22464 & ~ys__n738;
  assign new_new_n10622__ = ys__n22465 & ys__n738;
  assign ys__n22466 = new_new_n10621__ | new_new_n10622__;
  assign new_new_n10624__ = new_new_n10620__ & ~ys__n22466;
  assign new_new_n10625__ = new_new_n10605__ & ys__n22466;
  assign new_new_n10626__ = ~new_new_n10624__ & ~new_new_n10625__;
  assign new_new_n10627__ = ys__n23764 & ~new_new_n10626__;
  assign new_new_n10628__ = ~new_new_n10618__ & ~new_new_n10627__;
  assign new_new_n10629__ = ~ys__n532 & ~ys__n746;
  assign new_new_n10630__ = ys__n742 & ys__n744;
  assign new_new_n10631__ = new_new_n10629__ & new_new_n10630__;
  assign new_new_n10632__ = ~ys__n748 & ~ys__n750;
  assign new_new_n10633__ = new_new_n10631__ & new_new_n10632__;
  assign new_new_n10634__ = ys__n518 & ~ys__n548;
  assign new_new_n10635__ = ~ys__n550 & new_new_n10634__;
  assign new_new_n10636__ = ~ys__n518 & ~ys__n548;
  assign new_new_n10637__ = ~ys__n550 & new_new_n10636__;
  assign new_new_n10638__ = ~new_new_n10635__ & ~new_new_n10637__;
  assign new_new_n10639__ = ~ys__n23730 & ~new_new_n10638__;
  assign new_new_n10640__ = new_new_n10633__ & new_new_n10639__;
  assign new_new_n10641__ = ~ys__n742 & ys__n744;
  assign new_new_n10642__ = new_new_n10629__ & new_new_n10641__;
  assign new_new_n10643__ = new_new_n10632__ & new_new_n10642__;
  assign new_new_n10644__ = ys__n532 & ~ys__n746;
  assign new_new_n10645__ = new_new_n10641__ & new_new_n10644__;
  assign new_new_n10646__ = new_new_n10632__ & new_new_n10645__;
  assign new_new_n10647__ = ~new_new_n10643__ & ~new_new_n10646__;
  assign new_new_n10648__ = ~ys__n532 & ys__n746;
  assign new_new_n10649__ = ~ys__n742 & ~ys__n744;
  assign new_new_n10650__ = new_new_n10648__ & new_new_n10649__;
  assign new_new_n10651__ = new_new_n10632__ & new_new_n10650__;
  assign new_new_n10652__ = new_new_n10647__ & ~new_new_n10651__;
  assign new_new_n10653__ = ~ys__n23730 & ~new_new_n10652__;
  assign new_new_n10654__ = ~new_new_n10640__ & ~new_new_n10653__;
  assign new_new_n10655__ = ~new_new_n10633__ & new_new_n10652__;
  assign new_new_n10656__ = ~new_new_n10654__ & ~new_new_n10655__;
  assign new_new_n10657__ = new_new_n10629__ & new_new_n10649__;
  assign new_new_n10658__ = ys__n748 & ~ys__n750;
  assign new_new_n10659__ = new_new_n10657__ & new_new_n10658__;
  assign new_new_n10660__ = new_new_n10642__ & new_new_n10658__;
  assign new_new_n10661__ = ~new_new_n10659__ & ~new_new_n10660__;
  assign new_new_n10662__ = new_new_n10644__ & new_new_n10649__;
  assign new_new_n10663__ = new_new_n10658__ & new_new_n10662__;
  assign new_new_n10664__ = new_new_n10645__ & new_new_n10658__;
  assign new_new_n10665__ = ~new_new_n10663__ & ~new_new_n10664__;
  assign new_new_n10666__ = new_new_n10661__ & new_new_n10665__;
  assign new_new_n10667__ = ys__n532 & ys__n746;
  assign new_new_n10668__ = new_new_n10649__ & new_new_n10667__;
  assign new_new_n10669__ = new_new_n10658__ & new_new_n10668__;
  assign new_new_n10670__ = new_new_n10650__ & new_new_n10658__;
  assign new_new_n10671__ = ~new_new_n10669__ & ~new_new_n10670__;
  assign new_new_n10672__ = new_new_n10641__ & new_new_n10648__;
  assign new_new_n10673__ = new_new_n10658__ & new_new_n10672__;
  assign new_new_n10674__ = new_new_n10671__ & ~new_new_n10673__;
  assign new_new_n10675__ = new_new_n10666__ & new_new_n10674__;
  assign new_new_n10676__ = ~ys__n23730 & ~new_new_n10675__;
  assign new_new_n10677__ = ~new_new_n10656__ & ~new_new_n10676__;
  assign new_new_n10678__ = ys__n28243 & ~new_new_n10677__;
  assign new_new_n10679__ = ys__n23332 & ys__n38438;
  assign new_new_n10680__ = ~ys__n23332 & ys__n38449;
  assign new_new_n10681__ = ys__n23332 & ys__n38448;
  assign new_new_n10682__ = ~new_new_n10680__ & ~new_new_n10681__;
  assign new_new_n10683__ = ~new_new_n10679__ & new_new_n10682__;
  assign new_new_n10684__ = ~ys__n38437 & ~ys__n38438;
  assign new_new_n10685__ = new_new_n10683__ & new_new_n10684__;
  assign new_new_n10686__ = ys__n23627 & ~new_new_n10685__;
  assign new_new_n10687__ = ~ys__n23310 & ys__n28019;
  assign new_new_n10688__ = ys__n23310 & ~ys__n28019;
  assign new_new_n10689__ = ~new_new_n10687__ & ~new_new_n10688__;
  assign new_new_n10690__ = ~ys__n23312 & ys__n28020;
  assign new_new_n10691__ = ys__n23312 & ~ys__n28020;
  assign new_new_n10692__ = ~new_new_n10690__ & ~new_new_n10691__;
  assign new_new_n10693__ = new_new_n10689__ & new_new_n10692__;
  assign new_new_n10694__ = ~ys__n23314 & ys__n28021;
  assign new_new_n10695__ = ys__n23314 & ~ys__n28021;
  assign new_new_n10696__ = ~new_new_n10694__ & ~new_new_n10695__;
  assign new_new_n10697__ = ~ys__n23316 & ys__n28022;
  assign new_new_n10698__ = ys__n23316 & ~ys__n28022;
  assign new_new_n10699__ = ~new_new_n10697__ & ~new_new_n10698__;
  assign new_new_n10700__ = new_new_n10696__ & new_new_n10699__;
  assign new_new_n10701__ = new_new_n10693__ & new_new_n10700__;
  assign new_new_n10702__ = ~ys__n23302 & ys__n28015;
  assign new_new_n10703__ = ys__n23302 & ~ys__n28015;
  assign new_new_n10704__ = ~new_new_n10702__ & ~new_new_n10703__;
  assign new_new_n10705__ = ~ys__n23304 & ys__n28016;
  assign new_new_n10706__ = ys__n23304 & ~ys__n28016;
  assign new_new_n10707__ = ~new_new_n10705__ & ~new_new_n10706__;
  assign new_new_n10708__ = new_new_n10704__ & new_new_n10707__;
  assign new_new_n10709__ = ~ys__n23306 & ys__n28017;
  assign new_new_n10710__ = ys__n23306 & ~ys__n28017;
  assign new_new_n10711__ = ~new_new_n10709__ & ~new_new_n10710__;
  assign new_new_n10712__ = ~ys__n23308 & ys__n28018;
  assign new_new_n10713__ = ys__n23308 & ~ys__n28018;
  assign new_new_n10714__ = ~new_new_n10712__ & ~new_new_n10713__;
  assign new_new_n10715__ = new_new_n10711__ & new_new_n10714__;
  assign new_new_n10716__ = new_new_n10708__ & new_new_n10715__;
  assign new_new_n10717__ = new_new_n10701__ & new_new_n10716__;
  assign new_new_n10718__ = ~ys__n23326 & ys__n28027;
  assign new_new_n10719__ = ys__n23326 & ~ys__n28027;
  assign new_new_n10720__ = ~new_new_n10718__ & ~new_new_n10719__;
  assign new_new_n10721__ = ~ys__n23328 & ys__n28028;
  assign new_new_n10722__ = ys__n23328 & ~ys__n28028;
  assign new_new_n10723__ = ~new_new_n10721__ & ~new_new_n10722__;
  assign new_new_n10724__ = new_new_n10720__ & new_new_n10723__;
  assign new_new_n10725__ = ~ys__n23330 & ys__n28029;
  assign new_new_n10726__ = ys__n23330 & ~ys__n28029;
  assign new_new_n10727__ = ~new_new_n10725__ & ~new_new_n10726__;
  assign new_new_n10728__ = ~ys__n23332 & ys__n28030;
  assign new_new_n10729__ = ys__n23332 & ~ys__n28030;
  assign new_new_n10730__ = ~new_new_n10728__ & ~new_new_n10729__;
  assign new_new_n10731__ = new_new_n10727__ & new_new_n10730__;
  assign new_new_n10732__ = new_new_n10724__ & new_new_n10731__;
  assign new_new_n10733__ = ~ys__n23318 & ys__n28023;
  assign new_new_n10734__ = ys__n23318 & ~ys__n28023;
  assign new_new_n10735__ = ~new_new_n10733__ & ~new_new_n10734__;
  assign new_new_n10736__ = ~ys__n23320 & ys__n28024;
  assign new_new_n10737__ = ys__n23320 & ~ys__n28024;
  assign new_new_n10738__ = ~new_new_n10736__ & ~new_new_n10737__;
  assign new_new_n10739__ = new_new_n10735__ & new_new_n10738__;
  assign new_new_n10740__ = ~ys__n23322 & ys__n28025;
  assign new_new_n10741__ = ys__n23322 & ~ys__n28025;
  assign new_new_n10742__ = ~new_new_n10740__ & ~new_new_n10741__;
  assign new_new_n10743__ = ~ys__n23324 & ys__n28026;
  assign new_new_n10744__ = ys__n23324 & ~ys__n28026;
  assign new_new_n10745__ = ~new_new_n10743__ & ~new_new_n10744__;
  assign new_new_n10746__ = new_new_n10742__ & new_new_n10745__;
  assign new_new_n10747__ = new_new_n10739__ & new_new_n10746__;
  assign new_new_n10748__ = new_new_n10732__ & new_new_n10747__;
  assign new_new_n10749__ = new_new_n10717__ & new_new_n10748__;
  assign new_new_n10750__ = ~ys__n23278 & ys__n27863;
  assign new_new_n10751__ = ys__n23278 & ~ys__n27863;
  assign new_new_n10752__ = ~new_new_n10750__ & ~new_new_n10751__;
  assign new_new_n10753__ = ~ys__n23280 & ys__n27865;
  assign new_new_n10754__ = ys__n23280 & ~ys__n27865;
  assign new_new_n10755__ = ~new_new_n10753__ & ~new_new_n10754__;
  assign new_new_n10756__ = new_new_n10752__ & new_new_n10755__;
  assign new_new_n10757__ = ~ys__n23282 & ys__n27867;
  assign new_new_n10758__ = ys__n23282 & ~ys__n27867;
  assign new_new_n10759__ = ~new_new_n10757__ & ~new_new_n10758__;
  assign new_new_n10760__ = ~ys__n23284 & ys__n27869;
  assign new_new_n10761__ = ys__n23284 & ~ys__n27869;
  assign new_new_n10762__ = ~new_new_n10760__ & ~new_new_n10761__;
  assign new_new_n10763__ = new_new_n10759__ & new_new_n10762__;
  assign new_new_n10764__ = new_new_n10756__ & new_new_n10763__;
  assign new_new_n10765__ = ~ys__n23335 & ys__n27855;
  assign new_new_n10766__ = ys__n23335 & ~ys__n27855;
  assign new_new_n10767__ = ~new_new_n10765__ & ~new_new_n10766__;
  assign new_new_n10768__ = ~ys__n23272 & ys__n27857;
  assign new_new_n10769__ = ys__n23272 & ~ys__n27857;
  assign new_new_n10770__ = ~new_new_n10768__ & ~new_new_n10769__;
  assign new_new_n10771__ = new_new_n10767__ & new_new_n10770__;
  assign new_new_n10772__ = ~ys__n23274 & ys__n27859;
  assign new_new_n10773__ = ys__n23274 & ~ys__n27859;
  assign new_new_n10774__ = ~new_new_n10772__ & ~new_new_n10773__;
  assign new_new_n10775__ = ~ys__n23276 & ys__n27861;
  assign new_new_n10776__ = ys__n23276 & ~ys__n27861;
  assign new_new_n10777__ = ~new_new_n10775__ & ~new_new_n10776__;
  assign new_new_n10778__ = new_new_n10774__ & new_new_n10777__;
  assign new_new_n10779__ = new_new_n10771__ & new_new_n10778__;
  assign new_new_n10780__ = new_new_n10764__ & new_new_n10779__;
  assign new_new_n10781__ = ~ys__n23294 & ys__n27879;
  assign new_new_n10782__ = ys__n23294 & ~ys__n27879;
  assign new_new_n10783__ = ~new_new_n10781__ & ~new_new_n10782__;
  assign new_new_n10784__ = ~ys__n23296 & ys__n27881;
  assign new_new_n10785__ = ys__n23296 & ~ys__n27881;
  assign new_new_n10786__ = ~new_new_n10784__ & ~new_new_n10785__;
  assign new_new_n10787__ = new_new_n10783__ & new_new_n10786__;
  assign new_new_n10788__ = ~ys__n23298 & ys__n27883;
  assign new_new_n10789__ = ys__n23298 & ~ys__n27883;
  assign new_new_n10790__ = ~new_new_n10788__ & ~new_new_n10789__;
  assign new_new_n10791__ = ~ys__n23300 & ys__n27885;
  assign new_new_n10792__ = ys__n23300 & ~ys__n27885;
  assign new_new_n10793__ = ~new_new_n10791__ & ~new_new_n10792__;
  assign new_new_n10794__ = new_new_n10790__ & new_new_n10793__;
  assign new_new_n10795__ = new_new_n10787__ & new_new_n10794__;
  assign new_new_n10796__ = ~ys__n23286 & ys__n27871;
  assign new_new_n10797__ = ys__n23286 & ~ys__n27871;
  assign new_new_n10798__ = ~new_new_n10796__ & ~new_new_n10797__;
  assign new_new_n10799__ = ~ys__n23288 & ys__n27873;
  assign new_new_n10800__ = ys__n23288 & ~ys__n27873;
  assign new_new_n10801__ = ~new_new_n10799__ & ~new_new_n10800__;
  assign new_new_n10802__ = new_new_n10798__ & new_new_n10801__;
  assign new_new_n10803__ = ~ys__n23290 & ys__n27875;
  assign new_new_n10804__ = ys__n23290 & ~ys__n27875;
  assign new_new_n10805__ = ~new_new_n10803__ & ~new_new_n10804__;
  assign new_new_n10806__ = ~ys__n23292 & ys__n27877;
  assign new_new_n10807__ = ys__n23292 & ~ys__n27877;
  assign new_new_n10808__ = ~new_new_n10806__ & ~new_new_n10807__;
  assign new_new_n10809__ = new_new_n10805__ & new_new_n10808__;
  assign new_new_n10810__ = new_new_n10802__ & new_new_n10809__;
  assign new_new_n10811__ = new_new_n10795__ & new_new_n10810__;
  assign new_new_n10812__ = new_new_n10780__ & new_new_n10811__;
  assign new_new_n10813__ = new_new_n10749__ & new_new_n10812__;
  assign new_new_n10814__ = new_new_n10686__ & new_new_n10813__;
  assign new_new_n10815__ = ~ys__n23332 & ys__n38443;
  assign new_new_n10816__ = ~ys__n38441 & ~new_new_n10815__;
  assign new_new_n10817__ = new_new_n10683__ & new_new_n10816__;
  assign new_new_n10818__ = ys__n23627 & ~new_new_n10817__;
  assign new_new_n10819__ = ~new_new_n10813__ & new_new_n10818__;
  assign new_new_n10820__ = ~new_new_n10814__ & ~new_new_n10819__;
  assign new_new_n10821__ = ~ys__n23641 & ~ys__n23645;
  assign new_new_n10822__ = ~ys__n23652 & ~ys__n38413;
  assign new_new_n10823__ = new_new_n10821__ & new_new_n10822__;
  assign new_new_n10824__ = ys__n935 & ys__n33340;
  assign new_new_n10825__ = ~ys__n33380 & ~ys__n33384;
  assign new_new_n10826__ = ~ys__n33386 & new_new_n10825__;
  assign new_new_n10827__ = ~new_new_n10824__ & new_new_n10826__;
  assign ys__n478 = ~new_new_n10823__ & new_new_n10827__;
  assign ys__n4566 = ys__n935 | ys__n478;
  assign new_new_n10830__ = ys__n23627 & ~ys__n23717;
  assign new_new_n10831__ = ~ys__n4566 & new_new_n10830__;
  assign new_new_n10832__ = new_new_n10820__ & new_new_n10831__;
  assign ys__n18120 = new_new_n10678__ | ~new_new_n10832__;
  assign new_new_n10834__ = ys__n19245 & ~ys__n19253;
  assign new_new_n10835__ = ~ys__n738 & new_new_n10834__;
  assign new_new_n10836__ = ~ys__n18120 & new_new_n10835__;
  assign new_new_n10837__ = ~ys__n306 & ys__n38567;
  assign new_new_n10838__ = ys__n306 & ~ys__n38567;
  assign new_new_n10839__ = ~new_new_n10837__ & ~new_new_n10838__;
  assign new_new_n10840__ = ~ys__n38568 & ys__n38569;
  assign new_new_n10841__ = ys__n38568 & ~ys__n38569;
  assign new_new_n10842__ = ~new_new_n10840__ & ~new_new_n10841__;
  assign new_new_n10843__ = new_new_n10839__ & new_new_n10842__;
  assign ys__n1073 = ys__n18124 & ys__n24177;
  assign new_new_n10845__ = new_new_n10843__ & ys__n1073;
  assign new_new_n10846__ = ~ys__n418 & ys__n38528;
  assign new_new_n10847__ = ys__n18121 & ys__n18124;
  assign new_new_n10848__ = ~new_new_n10846__ & new_new_n10847__;
  assign new_new_n10849__ = ys__n35704 & ~ys__n38529;
  assign new_new_n10850__ = ys__n418 & ~ys__n38528;
  assign new_new_n10851__ = ~ys__n35704 & ys__n38529;
  assign new_new_n10852__ = ~new_new_n10850__ & ~new_new_n10851__;
  assign new_new_n10853__ = ~new_new_n10849__ & new_new_n10852__;
  assign new_new_n10854__ = new_new_n10848__ & new_new_n10853__;
  assign new_new_n10855__ = ys__n18122 & ys__n18124;
  assign new_new_n10856__ = ~new_new_n10854__ & ~new_new_n10855__;
  assign ys__n30223 = new_new_n10845__ | ~new_new_n10856__;
  assign new_new_n10858__ = ys__n19253 & ys__n30223;
  assign new_new_n10859__ = ~new_new_n10836__ & ~new_new_n10858__;
  assign new_new_n10860__ = ys__n140 & ~ys__n19245;
  assign new_new_n10861__ = ~ys__n738 & new_new_n10860__;
  assign new_new_n10862__ = ys__n19245 & ~ys__n738;
  assign new_new_n10863__ = ys__n18120 & new_new_n10862__;
  assign new_new_n10864__ = ~new_new_n10861__ & ~new_new_n10863__;
  assign new_new_n10865__ = new_new_n10859__ & new_new_n10864__;
  assign new_new_n10866__ = ~new_new_n10859__ & ~new_new_n10865__;
  assign ys__n25436 = ~new_new_n10628__ & new_new_n10866__;
  assign new_new_n10868__ = ys__n738 & new_new_n10860__;
  assign new_new_n10869__ = ys__n19245 & ys__n738;
  assign new_new_n10870__ = ~new_new_n10868__ & ~new_new_n10869__;
  assign new_new_n10871__ = ~ys__n19253 & ~new_new_n10870__;
  assign new_new_n10872__ = ys__n19253 & ~ys__n30223;
  assign ys__n19256 = new_new_n10871__ | new_new_n10872__;
  assign new_new_n10874__ = ys__n25436 & ~ys__n19256;
  assign new_new_n10875__ = ys__n642 & ys__n19256;
  assign new_new_n10876__ = ~new_new_n10874__ & ~new_new_n10875__;
  assign ys__n2 = ys__n874 & ~new_new_n10876__;
  assign new_new_n10878__ = ~ys__n4299 & ~ys__n4300;
  assign new_new_n10879__ = ~ys__n4305 & ys__n19263;
  assign new_new_n10880__ = new_new_n10878__ & new_new_n10879__;
  assign new_new_n10881__ = ys__n244 & ~ys__n4291;
  assign new_new_n10882__ = ~ys__n4292 & ~ys__n4294;
  assign new_new_n10883__ = ~ys__n4296 & ~ys__n4297;
  assign new_new_n10884__ = new_new_n10882__ & new_new_n10883__;
  assign new_new_n10885__ = new_new_n10881__ & new_new_n10884__;
  assign new_new_n10886__ = new_new_n10880__ & new_new_n10885__;
  assign new_new_n10887__ = ys__n20273 & ~ys__n28243;
  assign new_new_n10888__ = ~ys__n738 & new_new_n10887__;
  assign ys__n246 = ~new_new_n10886__ & new_new_n10888__;
  assign new_new_n10890__ = ys__n28243 & ~ys__n38203;
  assign new_new_n10891__ = ys__n28243 & ~ys__n38202;
  assign new_new_n10892__ = ~ys__n28243 & ys__n38203;
  assign new_new_n10893__ = ~new_new_n10891__ & ~new_new_n10892__;
  assign new_new_n10894__ = ~new_new_n10890__ & new_new_n10893__;
  assign new_new_n10895__ = ~ys__n28243 & ys__n38199;
  assign new_new_n10896__ = ys__n38183 & ~ys__n38200;
  assign new_new_n10897__ = ~new_new_n10895__ & new_new_n10896__;
  assign new_new_n10898__ = ys__n28243 & ~ys__n38199;
  assign new_new_n10899__ = ~ys__n28243 & ys__n38201;
  assign new_new_n10900__ = ~new_new_n10898__ & ~new_new_n10899__;
  assign new_new_n10901__ = ys__n28243 & ~ys__n38201;
  assign new_new_n10902__ = ~ys__n28243 & ys__n38202;
  assign new_new_n10903__ = ~new_new_n10901__ & ~new_new_n10902__;
  assign new_new_n10904__ = new_new_n10900__ & new_new_n10903__;
  assign new_new_n10905__ = new_new_n10897__ & new_new_n10904__;
  assign new_new_n10906__ = new_new_n10894__ & new_new_n10905__;
  assign new_new_n10907__ = ys__n20273 & ys__n28243;
  assign new_new_n10908__ = ~ys__n738 & new_new_n10907__;
  assign new_new_n10909__ = ~new_new_n10886__ & new_new_n10908__;
  assign ys__n250 = new_new_n10906__ & new_new_n10909__;
  assign new_new_n10911__ = ~ys__n19263 & ys__n20279;
  assign new_new_n10912__ = ~ys__n738 & new_new_n10911__;
  assign new_new_n10913__ = ~ys__n19263 & ~new_new_n10912__;
  assign new_new_n10914__ = ~ys__n19263 & ys__n20273;
  assign new_new_n10915__ = ys__n20280 & new_new_n10914__;
  assign new_new_n10916__ = ~ys__n738 & new_new_n10915__;
  assign new_new_n10917__ = ys__n738 & new_new_n10914__;
  assign new_new_n10918__ = ys__n20273 & ~new_new_n10917__;
  assign new_new_n10919__ = ~new_new_n10916__ & new_new_n10918__;
  assign new_new_n10920__ = ~new_new_n10913__ & new_new_n10919__;
  assign new_new_n10921__ = ~ys__n766 & ys__n28243;
  assign new_new_n10922__ = ~ys__n764 & ys__n28243;
  assign new_new_n10923__ = ys__n766 & ~ys__n28243;
  assign new_new_n10924__ = ~new_new_n10922__ & ~new_new_n10923__;
  assign new_new_n10925__ = ~new_new_n10921__ & new_new_n10924__;
  assign new_new_n10926__ = ys__n758 & ~ys__n28243;
  assign new_new_n10927__ = ~ys__n760 & ys__n38198;
  assign new_new_n10928__ = ~new_new_n10926__ & new_new_n10927__;
  assign new_new_n10929__ = ~ys__n758 & ys__n28243;
  assign new_new_n10930__ = ys__n762 & ~ys__n28243;
  assign new_new_n10931__ = ~new_new_n10929__ & ~new_new_n10930__;
  assign new_new_n10932__ = ~ys__n762 & ys__n28243;
  assign new_new_n10933__ = ys__n764 & ~ys__n28243;
  assign new_new_n10934__ = ~new_new_n10932__ & ~new_new_n10933__;
  assign new_new_n10935__ = new_new_n10931__ & new_new_n10934__;
  assign new_new_n10936__ = new_new_n10928__ & new_new_n10935__;
  assign new_new_n10937__ = new_new_n10925__ & new_new_n10936__;
  assign new_new_n10938__ = ~new_new_n10906__ & new_new_n10937__;
  assign new_new_n10939__ = new_new_n10909__ & new_new_n10938__;
  assign ys__n252 = ~new_new_n10920__ & new_new_n10939__;
  assign new_new_n10941__ = ys__n28243 & ~ys__n738;
  assign new_new_n10942__ = ~new_new_n10886__ & new_new_n10941__;
  assign new_new_n10943__ = new_new_n10938__ & new_new_n10942__;
  assign new_new_n10944__ = new_new_n10920__ & new_new_n10943__;
  assign new_new_n10945__ = ~new_new_n10886__ & ~new_new_n10944__;
  assign ys__n254 = ys__n20273 & ~new_new_n10945__;
  assign new_new_n10947__ = ys__n28243 & ~ys__n38197;
  assign new_new_n10948__ = ys__n28243 & ~ys__n38196;
  assign new_new_n10949__ = ~ys__n28243 & ys__n38197;
  assign new_new_n10950__ = ~new_new_n10948__ & ~new_new_n10949__;
  assign new_new_n10951__ = ~new_new_n10947__ & new_new_n10950__;
  assign new_new_n10952__ = ~ys__n28243 & ys__n38193;
  assign new_new_n10953__ = ys__n38192 & ~ys__n38194;
  assign new_new_n10954__ = ~new_new_n10952__ & new_new_n10953__;
  assign new_new_n10955__ = ys__n28243 & ~ys__n38193;
  assign new_new_n10956__ = ~ys__n28243 & ys__n38195;
  assign new_new_n10957__ = ~new_new_n10955__ & ~new_new_n10956__;
  assign new_new_n10958__ = ys__n28243 & ~ys__n38195;
  assign new_new_n10959__ = ~ys__n28243 & ys__n38196;
  assign new_new_n10960__ = ~new_new_n10958__ & ~new_new_n10959__;
  assign new_new_n10961__ = new_new_n10957__ & new_new_n10960__;
  assign new_new_n10962__ = new_new_n10954__ & new_new_n10961__;
  assign new_new_n10963__ = new_new_n10951__ & new_new_n10962__;
  assign new_new_n10964__ = ~new_new_n10906__ & ~new_new_n10937__;
  assign new_new_n10965__ = new_new_n10963__ & new_new_n10964__;
  assign ys__n270 = new_new_n10909__ & new_new_n10965__;
  assign new_new_n10967__ = ~new_new_n10963__ & new_new_n10964__;
  assign ys__n278 = new_new_n10909__ & new_new_n10967__;
  assign ys__n404 = ys__n17849 & ~ys__n18156;
  assign new_new_n10970__ = ~ys__n33384 & ys__n38315;
  assign new_new_n10971__ = ys__n38323 & new_new_n10970__;
  assign new_new_n10972__ = ~ys__n38320 & ~new_new_n10971__;
  assign new_new_n10973__ = ys__n38217 & ~new_new_n10972__;
  assign new_new_n10974__ = ys__n38215 & ~new_new_n10972__;
  assign new_new_n10975__ = ~new_new_n10973__ & new_new_n10974__;
  assign new_new_n10976__ = ~new_new_n10973__ & ~new_new_n10975__;
  assign new_new_n10977__ = ~ys__n23641 & ~new_new_n10976__;
  assign new_new_n10978__ = ~ys__n23641 & ~new_new_n10977__;
  assign new_new_n10979__ = ~ys__n23645 & ~ys__n23652;
  assign new_new_n10980__ = ~new_new_n10978__ & new_new_n10979__;
  assign ys__n480 = ys__n23652 | new_new_n10980__;
  assign new_new_n10982__ = new_new_n10821__ & new_new_n10975__;
  assign new_new_n10983__ = ys__n23644 & ys__n23645;
  assign new_new_n10984__ = ~new_new_n10982__ & ~new_new_n10983__;
  assign ys__n482 = ~ys__n23652 & ~new_new_n10984__;
  assign new_new_n10986__ = ~ys__n206 & ~ys__n208;
  assign new_new_n10987__ = ~ys__n190 & ~ys__n192;
  assign new_new_n10988__ = ~ys__n204 & ~ys__n860;
  assign new_new_n10989__ = new_new_n10987__ & new_new_n10988__;
  assign new_new_n10990__ = new_new_n10986__ & new_new_n10989__;
  assign new_new_n10991__ = ys__n33403 & ~new_new_n10990__;
  assign new_new_n10992__ = ys__n30863 & ~ys__n33384;
  assign new_new_n10993__ = ys__n176 & ~ys__n178;
  assign new_new_n10994__ = new_new_n10992__ & new_new_n10993__;
  assign new_new_n10995__ = ~new_new_n10991__ & new_new_n10994__;
  assign new_new_n10996__ = ~ys__n176 & ys__n178;
  assign new_new_n10997__ = new_new_n10992__ & new_new_n10996__;
  assign new_new_n10998__ = new_new_n10990__ & new_new_n10997__;
  assign new_new_n10999__ = ~new_new_n10995__ & ~new_new_n10998__;
  assign new_new_n11000__ = ~ys__n176 & ~ys__n178;
  assign new_new_n11001__ = ys__n176 & ys__n178;
  assign new_new_n11002__ = ~new_new_n11000__ & ~new_new_n11001__;
  assign new_new_n11003__ = ~new_new_n10993__ & ~new_new_n10996__;
  assign new_new_n11004__ = new_new_n11002__ & new_new_n11003__;
  assign new_new_n11005__ = ~new_new_n10999__ & ~new_new_n11004__;
  assign new_new_n11006__ = ~ys__n738 & ~ys__n4566;
  assign ys__n502 = new_new_n11005__ & new_new_n11006__;
  assign new_new_n11008__ = ys__n568 & ~ys__n572;
  assign new_new_n11009__ = ~ys__n566 & ys__n570;
  assign new_new_n11010__ = new_new_n11008__ & new_new_n11009__;
  assign new_new_n11011__ = ~ys__n568 & ~ys__n572;
  assign new_new_n11012__ = new_new_n11009__ & new_new_n11011__;
  assign new_new_n11013__ = ys__n568 & ys__n572;
  assign new_new_n11014__ = ys__n566 & ~ys__n570;
  assign new_new_n11015__ = new_new_n11013__ & new_new_n11014__;
  assign new_new_n11016__ = ~new_new_n11012__ & ~new_new_n11015__;
  assign new_new_n11017__ = ~new_new_n11010__ & new_new_n11016__;
  assign new_new_n11018__ = ~ys__n568 & ys__n572;
  assign new_new_n11019__ = new_new_n11014__ & new_new_n11018__;
  assign new_new_n11020__ = new_new_n11008__ & new_new_n11014__;
  assign new_new_n11021__ = ~new_new_n11019__ & ~new_new_n11020__;
  assign new_new_n11022__ = new_new_n11011__ & new_new_n11014__;
  assign new_new_n11023__ = ~ys__n566 & ~ys__n570;
  assign new_new_n11024__ = new_new_n11013__ & new_new_n11023__;
  assign new_new_n11025__ = ~new_new_n11022__ & ~new_new_n11024__;
  assign new_new_n11026__ = new_new_n11021__ & new_new_n11025__;
  assign ys__n17780 = ~new_new_n11011__ | ~new_new_n11023__;
  assign new_new_n11028__ = new_new_n11009__ & new_new_n11018__;
  assign new_new_n11029__ = ~new_new_n11010__ & ~new_new_n11028__;
  assign new_new_n11030__ = ys__n17780 & new_new_n11029__;
  assign new_new_n11031__ = new_new_n11018__ & new_new_n11023__;
  assign new_new_n11032__ = new_new_n11008__ & new_new_n11023__;
  assign new_new_n11033__ = ~new_new_n11031__ & ~new_new_n11032__;
  assign new_new_n11034__ = new_new_n11016__ & new_new_n11033__;
  assign new_new_n11035__ = new_new_n11030__ & new_new_n11034__;
  assign new_new_n11036__ = new_new_n11026__ & new_new_n11035__;
  assign ys__n574 = ~new_new_n11017__ & ~new_new_n11036__;
  assign new_new_n11038__ = ~ys__n33563 & ~ys__n38922;
  assign new_new_n11039__ = ys__n38919 & new_new_n10613__;
  assign new_new_n11040__ = ~new_new_n11038__ & new_new_n11039__;
  assign new_new_n11041__ = ~ys__n4184 & ~ys__n4810;
  assign new_new_n11042__ = ~ys__n4192 & new_new_n11041__;
  assign new_new_n11043__ = new_new_n10611__ & ~ys__n17780;
  assign new_new_n11044__ = new_new_n11042__ & new_new_n11043__;
  assign new_new_n11045__ = new_new_n11040__ & new_new_n11044__;
  assign new_new_n11046__ = new_new_n10610__ & new_new_n10613__;
  assign new_new_n11047__ = ~ys__n4613 & ~ys__n4625;
  assign new_new_n11048__ = ~ys__n4185 & ~ys__n4810;
  assign new_new_n11049__ = new_new_n11047__ & new_new_n11048__;
  assign new_new_n11050__ = new_new_n11031__ & new_new_n11049__;
  assign new_new_n11051__ = new_new_n11046__ & new_new_n11050__;
  assign new_new_n11052__ = ys__n47107 & new_new_n11012__;
  assign new_new_n11053__ = ys__n30230 & ~ys__n30232;
  assign new_new_n11054__ = ys__n30232 & ~ys__n33563;
  assign new_new_n11055__ = ~new_new_n11053__ & ~new_new_n11054__;
  assign new_new_n11056__ = new_new_n11010__ & new_new_n11055__;
  assign new_new_n11057__ = ~new_new_n11019__ & ~new_new_n11022__;
  assign new_new_n11058__ = ~new_new_n11056__ & new_new_n11057__;
  assign new_new_n11059__ = ~new_new_n11052__ & new_new_n11058__;
  assign new_new_n11060__ = ~new_new_n11051__ & new_new_n11059__;
  assign new_new_n11061__ = ~new_new_n11045__ & new_new_n11060__;
  assign ys__n576 = ~new_new_n11036__ & ~new_new_n11061__;
  assign new_new_n11063__ = ~ys__n108 & ~ys__n290;
  assign new_new_n11064__ = ~ys__n110 & ys__n112;
  assign new_new_n11065__ = ~ys__n1309 & new_new_n11064__;
  assign new_new_n11066__ = new_new_n11063__ & new_new_n11065__;
  assign new_new_n11067__ = ~ys__n108 & ~ys__n1309;
  assign new_new_n11068__ = ~ys__n110 & ~ys__n112;
  assign new_new_n11069__ = ys__n114 & ~ys__n290;
  assign new_new_n11070__ = new_new_n11068__ & new_new_n11069__;
  assign new_new_n11071__ = new_new_n11067__ & new_new_n11070__;
  assign new_new_n11072__ = ~new_new_n11066__ & ~new_new_n11071__;
  assign new_new_n11073__ = ~ys__n114 & ys__n118;
  assign new_new_n11074__ = ~ys__n1309 & new_new_n11073__;
  assign new_new_n11075__ = new_new_n11063__ & new_new_n11068__;
  assign new_new_n11076__ = new_new_n11074__ & new_new_n11075__;
  assign new_new_n11077__ = ys__n110 & ~ys__n290;
  assign new_new_n11078__ = new_new_n11067__ & new_new_n11077__;
  assign new_new_n11079__ = ~ys__n108 & ys__n290;
  assign new_new_n11080__ = ~ys__n1309 & new_new_n11079__;
  assign new_new_n11081__ = ys__n108 & ~ys__n1309;
  assign new_new_n11082__ = ~ys__n1309 & ~new_new_n11081__;
  assign new_new_n11083__ = ~new_new_n11080__ & new_new_n11082__;
  assign new_new_n11084__ = ~new_new_n11078__ & new_new_n11083__;
  assign new_new_n11085__ = ~new_new_n11076__ & new_new_n11084__;
  assign new_new_n11086__ = new_new_n11072__ & new_new_n11085__;
  assign new_new_n11087__ = ys__n112 & new_new_n11086__;
  assign new_new_n11088__ = ~ys__n37672 & ys__n37673;
  assign new_new_n11089__ = ys__n37672 & ~ys__n37673;
  assign new_new_n11090__ = ~new_new_n11088__ & ~new_new_n11089__;
  assign new_new_n11091__ = ~ys__n18393 & ~new_new_n11090__;
  assign new_new_n11092__ = ys__n38861 & ys__n38862;
  assign new_new_n11093__ = ys__n38863 & ~new_new_n11092__;
  assign new_new_n11094__ = ~ys__n33541 & ~ys__n33552;
  assign new_new_n11095__ = ~ys__n38865 & ~new_new_n11094__;
  assign new_new_n11096__ = new_new_n11093__ & ~new_new_n11095__;
  assign new_new_n11097__ = ys__n38864 & ys__n38865;
  assign new_new_n11098__ = ~ys__n33541 & ys__n38863;
  assign new_new_n11099__ = ~new_new_n11093__ & new_new_n11098__;
  assign new_new_n11100__ = ~new_new_n11097__ & ~new_new_n11099__;
  assign new_new_n11101__ = ~new_new_n11096__ & new_new_n11100__;
  assign new_new_n11102__ = ~ys__n4750 & ~ys__n4751;
  assign new_new_n11103__ = ~ys__n4753 & ~ys__n4754;
  assign new_new_n11104__ = ~ys__n4759 & ~ys__n4761;
  assign new_new_n11105__ = new_new_n11103__ & new_new_n11104__;
  assign new_new_n11106__ = new_new_n11102__ & new_new_n11105__;
  assign new_new_n11107__ = ~ys__n4756 & ~ys__n4757;
  assign new_new_n11108__ = ~ys__n4744 & ~ys__n4746;
  assign new_new_n11109__ = new_new_n11107__ & new_new_n11108__;
  assign ys__n4764 = ~new_new_n11106__ | ~new_new_n11109__;
  assign new_new_n11111__ = ~ys__n29117 & ~ys__n4764;
  assign new_new_n11112__ = ~new_new_n11101__ & new_new_n11111__;
  assign ys__n37703 = ys__n24675 | new_new_n11112__;
  assign new_new_n11114__ = ys__n33552 & ys__n38865;
  assign new_new_n11115__ = new_new_n11093__ & new_new_n11114__;
  assign new_new_n11116__ = ~ys__n24675 & ys__n24711;
  assign new_new_n11117__ = ys__n24675 & ys__n24712;
  assign ys__n18759 = new_new_n11116__ | new_new_n11117__;
  assign new_new_n11119__ = new_new_n11115__ & ~ys__n18759;
  assign new_new_n11120__ = ~ys__n38864 & ~new_new_n11119__;
  assign new_new_n11121__ = ~ys__n24675 & ~new_new_n11120__;
  assign new_new_n11122__ = ys__n37703 & new_new_n11121__;
  assign ys__n1020 = ys__n4783 | ys__n4784;
  assign new_new_n11124__ = ~ys__n33545 & ys__n1020;
  assign new_new_n11125__ = ~ys__n4764 & new_new_n11124__;
  assign new_new_n11126__ = ~ys__n844 & ~ys__n3214;
  assign new_new_n11127__ = ~ys__n18070 & ~ys__n18071;
  assign new_new_n11128__ = new_new_n11126__ & new_new_n11127__;
  assign new_new_n11129__ = ~new_new_n11125__ & new_new_n11128__;
  assign new_new_n11130__ = ~new_new_n11122__ & new_new_n11129__;
  assign new_new_n11131__ = ys__n18270 & new_new_n11130__;
  assign new_new_n11132__ = ~ys__n18270 & ~new_new_n11130__;
  assign new_new_n11133__ = ~new_new_n11131__ & ~new_new_n11132__;
  assign new_new_n11134__ = ~ys__n18271 & ~new_new_n11133__;
  assign new_new_n11135__ = ys__n18270 & ys__n18271;
  assign ys__n18272 = new_new_n11134__ | new_new_n11135__;
  assign new_new_n11137__ = ~ys__n18393 & ys__n18272;
  assign new_new_n11138__ = ys__n18271 & ys__n18393;
  assign ys__n27603 = new_new_n11137__ | new_new_n11138__;
  assign new_new_n11140__ = ys__n18393 & ys__n27603;
  assign new_new_n11141__ = ~new_new_n11091__ & ~new_new_n11140__;
  assign new_new_n11142__ = ~ys__n18208 & ~new_new_n11141__;
  assign new_new_n11143__ = ys__n18090 & new_new_n11142__;
  assign new_new_n11144__ = ys__n19203 & ~ys__n19215;
  assign new_new_n11145__ = new_new_n11081__ & new_new_n11144__;
  assign new_new_n11146__ = new_new_n11143__ & new_new_n11145__;
  assign new_new_n11147__ = ys__n18317 & ~new_new_n11141__;
  assign new_new_n11148__ = ~ys__n17941 & ~ys__n17943;
  assign new_new_n11149__ = ys__n18090 & new_new_n11148__;
  assign new_new_n11150__ = new_new_n11076__ & new_new_n11149__;
  assign new_new_n11151__ = ~new_new_n11141__ & new_new_n11150__;
  assign new_new_n11152__ = new_new_n11142__ & new_new_n11151__;
  assign new_new_n11153__ = ~new_new_n11147__ & new_new_n11152__;
  assign new_new_n11154__ = ~new_new_n11146__ & ~new_new_n11153__;
  assign new_new_n11155__ = ~new_new_n11086__ & ~new_new_n11154__;
  assign ys__n628 = new_new_n11087__ | new_new_n11155__;
  assign new_new_n11157__ = ys__n114 & new_new_n11086__;
  assign new_new_n11158__ = ~new_new_n11086__ & new_new_n11150__;
  assign new_new_n11159__ = ~new_new_n11141__ & new_new_n11158__;
  assign new_new_n11160__ = ~new_new_n11142__ & new_new_n11159__;
  assign new_new_n11161__ = ~new_new_n11147__ & new_new_n11160__;
  assign ys__n630 = new_new_n11157__ | new_new_n11161__;
  assign new_new_n11163__ = ~ys__n748 & ys__n750;
  assign new_new_n11164__ = new_new_n10657__ & new_new_n11163__;
  assign new_new_n11165__ = ys__n522 & ys__n524;
  assign new_new_n11166__ = ys__n526 & ys__n528;
  assign new_new_n11167__ = new_new_n11165__ & new_new_n11166__;
  assign new_new_n11168__ = ~ys__n512 & ys__n520;
  assign new_new_n11169__ = ys__n530 & ~ys__n752;
  assign new_new_n11170__ = new_new_n11168__ & new_new_n11169__;
  assign new_new_n11171__ = new_new_n11167__ & new_new_n11170__;
  assign new_new_n11172__ = ~ys__n23730 & ~ys__n28243;
  assign new_new_n11173__ = new_new_n10830__ & new_new_n11172__;
  assign new_new_n11174__ = new_new_n11171__ & new_new_n11173__;
  assign new_new_n11175__ = new_new_n11164__ & new_new_n11174__;
  assign new_new_n11176__ = ~ys__n23627 & ~new_new_n11175__;
  assign new_new_n11177__ = ys__n22880 & new_new_n11175__;
  assign new_new_n11178__ = ~new_new_n11176__ & ~new_new_n11177__;
  assign new_new_n11179__ = ys__n23627 & ys__n23717;
  assign new_new_n11180__ = ~ys__n23730 & new_new_n11179__;
  assign new_new_n11181__ = ~new_new_n11178__ & ~new_new_n11180__;
  assign new_new_n11182__ = ys__n23328 & new_new_n11180__;
  assign new_new_n11183__ = ~new_new_n11181__ & ~new_new_n11182__;
  assign new_new_n11184__ = ~ys__n23730 & ys__n28243;
  assign new_new_n11185__ = new_new_n10830__ & new_new_n11184__;
  assign new_new_n11186__ = new_new_n10676__ & new_new_n11185__;
  assign new_new_n11187__ = ~new_new_n11183__ & ~new_new_n11186__;
  assign new_new_n11188__ = ys__n450 & new_new_n11186__;
  assign new_new_n11189__ = ~new_new_n11187__ & ~new_new_n11188__;
  assign new_new_n11190__ = new_new_n10668__ & new_new_n11163__;
  assign new_new_n11191__ = new_new_n10650__ & new_new_n11163__;
  assign new_new_n11192__ = ~new_new_n11190__ & ~new_new_n11191__;
  assign new_new_n11193__ = new_new_n10632__ & new_new_n10662__;
  assign new_new_n11194__ = new_new_n10662__ & new_new_n11163__;
  assign new_new_n11195__ = ~new_new_n11164__ & ~new_new_n11194__;
  assign new_new_n11196__ = ~new_new_n11193__ & new_new_n11195__;
  assign new_new_n11197__ = new_new_n11192__ & new_new_n11196__;
  assign new_new_n11198__ = new_new_n10632__ & new_new_n10672__;
  assign new_new_n11199__ = new_new_n10641__ & new_new_n10667__;
  assign new_new_n11200__ = new_new_n10632__ & new_new_n11199__;
  assign new_new_n11201__ = ~new_new_n11198__ & ~new_new_n11200__;
  assign new_new_n11202__ = new_new_n10647__ & new_new_n11201__;
  assign new_new_n11203__ = new_new_n10632__ & new_new_n10668__;
  assign new_new_n11204__ = new_new_n10630__ & new_new_n10644__;
  assign new_new_n11205__ = new_new_n11163__ & new_new_n11204__;
  assign new_new_n11206__ = ~new_new_n10651__ & ~new_new_n11205__;
  assign new_new_n11207__ = ~new_new_n11203__ & new_new_n11206__;
  assign new_new_n11208__ = new_new_n11202__ & new_new_n11207__;
  assign new_new_n11209__ = new_new_n11197__ & new_new_n11208__;
  assign new_new_n11210__ = ~ys__n4494 & ~ys__n4496;
  assign new_new_n11211__ = ys__n512 & ~ys__n632;
  assign new_new_n11212__ = new_new_n11210__ & new_new_n11211__;
  assign new_new_n11213__ = ~ys__n520 & new_new_n11212__;
  assign new_new_n11214__ = ~ys__n4478 & ~ys__n4480;
  assign new_new_n11215__ = ~ys__n514 & ~ys__n2024;
  assign new_new_n11216__ = new_new_n11214__ & new_new_n11215__;
  assign new_new_n11217__ = ~ys__n516 & new_new_n11216__;
  assign new_new_n11218__ = new_new_n11213__ & new_new_n11217__;
  assign new_new_n11219__ = ~ys__n28720 & new_new_n11218__;
  assign new_new_n11220__ = ys__n514 & ~ys__n2024;
  assign new_new_n11221__ = new_new_n11214__ & new_new_n11220__;
  assign new_new_n11222__ = ~ys__n516 & new_new_n11221__;
  assign new_new_n11223__ = new_new_n11213__ & new_new_n11222__;
  assign new_new_n11224__ = ys__n28720 & new_new_n11223__;
  assign new_new_n11225__ = ~new_new_n11219__ & ~new_new_n11224__;
  assign new_new_n11226__ = new_new_n11190__ & new_new_n11225__;
  assign new_new_n11227__ = new_new_n11164__ & ~new_new_n11171__;
  assign new_new_n11228__ = ys__n516 & new_new_n11216__;
  assign new_new_n11229__ = ys__n516 & new_new_n11221__;
  assign new_new_n11230__ = ~new_new_n11228__ & ~new_new_n11229__;
  assign new_new_n11231__ = ~new_new_n11217__ & ~new_new_n11222__;
  assign new_new_n11232__ = new_new_n11230__ & new_new_n11231__;
  assign new_new_n11233__ = new_new_n11193__ & new_new_n11232__;
  assign new_new_n11234__ = ~new_new_n11227__ & ~new_new_n11233__;
  assign new_new_n11235__ = ~new_new_n11226__ & new_new_n11234__;
  assign new_new_n11236__ = ~ys__n28719 & new_new_n11218__;
  assign new_new_n11237__ = ys__n28719 & new_new_n11223__;
  assign new_new_n11238__ = ~new_new_n11236__ & ~new_new_n11237__;
  assign new_new_n11239__ = new_new_n11191__ & new_new_n11238__;
  assign new_new_n11240__ = ~ys__n28718 & new_new_n11218__;
  assign new_new_n11241__ = ys__n28718 & new_new_n11223__;
  assign new_new_n11242__ = ~new_new_n11240__ & ~new_new_n11241__;
  assign new_new_n11243__ = new_new_n11194__ & new_new_n11242__;
  assign new_new_n11244__ = ~new_new_n11239__ & ~new_new_n11243__;
  assign new_new_n11245__ = new_new_n11235__ & new_new_n11244__;
  assign new_new_n11246__ = ~new_new_n11209__ & ~new_new_n11245__;
  assign new_new_n11247__ = ~new_new_n11209__ & ~new_new_n11246__;
  assign new_new_n11248__ = ~ys__n28243 & ~new_new_n11247__;
  assign new_new_n11249__ = ~new_new_n10633__ & ~new_new_n10651__;
  assign new_new_n11250__ = new_new_n10658__ & new_new_n11204__;
  assign new_new_n11251__ = ~new_new_n10673__ & ~new_new_n11250__;
  assign new_new_n11252__ = new_new_n11249__ & new_new_n11251__;
  assign new_new_n11253__ = new_new_n10647__ & new_new_n10671__;
  assign new_new_n11254__ = new_new_n11252__ & new_new_n11253__;
  assign new_new_n11255__ = new_new_n10666__ & new_new_n11254__;
  assign new_new_n11256__ = new_new_n10633__ & new_new_n10638__;
  assign new_new_n11257__ = ~ys__n526 & ~ys__n528;
  assign new_new_n11258__ = ~ys__n522 & ~ys__n524;
  assign new_new_n11259__ = new_new_n11257__ & new_new_n11258__;
  assign new_new_n11260__ = ~ys__n530 & new_new_n11259__;
  assign new_new_n11261__ = ~ys__n23730 & new_new_n11260__;
  assign new_new_n11262__ = new_new_n11260__ & ~new_new_n11261__;
  assign new_new_n11263__ = new_new_n11250__ & ~new_new_n11262__;
  assign new_new_n11264__ = ~new_new_n11256__ & ~new_new_n11263__;
  assign new_new_n11265__ = ~new_new_n11255__ & ~new_new_n11264__;
  assign new_new_n11266__ = ~new_new_n11255__ & ~new_new_n11265__;
  assign new_new_n11267__ = ys__n28243 & ~new_new_n11266__;
  assign new_new_n11268__ = ~new_new_n11248__ & ~new_new_n11267__;
  assign new_new_n11269__ = ~ys__n23730 & new_new_n10830__;
  assign new_new_n11270__ = ~new_new_n11268__ & new_new_n11269__;
  assign new_new_n11271__ = ~new_new_n11189__ & ~new_new_n11270__;
  assign new_new_n11272__ = ~ys__n23339 & ys__n23548;
  assign new_new_n11273__ = ys__n23550 & new_new_n11272__;
  assign new_new_n11274__ = ~ys__n23339 & ~ys__n23548;
  assign new_new_n11275__ = ys__n23339 & ys__n23548;
  assign new_new_n11276__ = ~new_new_n11274__ & ~new_new_n11275__;
  assign new_new_n11277__ = ys__n22464 & ys__n23339;
  assign new_new_n11278__ = ys__n23550 & new_new_n11277__;
  assign new_new_n11279__ = ~new_new_n11276__ & new_new_n11278__;
  assign new_new_n11280__ = ~new_new_n11273__ & ~new_new_n11279__;
  assign new_new_n11281__ = ys__n23552 & ys__n23554;
  assign new_new_n11282__ = ys__n23556 & ys__n23558;
  assign new_new_n11283__ = new_new_n11281__ & new_new_n11282__;
  assign new_new_n11284__ = ~new_new_n11280__ & new_new_n11283__;
  assign new_new_n11285__ = ys__n23560 & ys__n23562;
  assign new_new_n11286__ = ys__n23564 & ys__n23566;
  assign new_new_n11287__ = new_new_n11285__ & new_new_n11286__;
  assign new_new_n11288__ = ys__n23568 & ys__n23570;
  assign new_new_n11289__ = ys__n23572 & ys__n23574;
  assign new_new_n11290__ = new_new_n11288__ & new_new_n11289__;
  assign new_new_n11291__ = new_new_n11287__ & new_new_n11290__;
  assign new_new_n11292__ = new_new_n11284__ & new_new_n11291__;
  assign new_new_n11293__ = ys__n450 & ~new_new_n11292__;
  assign new_new_n11294__ = ys__n420 & ys__n442;
  assign new_new_n11295__ = ys__n440 & ys__n444;
  assign new_new_n11296__ = new_new_n11294__ & new_new_n11295__;
  assign new_new_n11297__ = ys__n438 & ys__n446;
  assign new_new_n11298__ = ys__n434 & ys__n436;
  assign new_new_n11299__ = new_new_n11297__ & new_new_n11298__;
  assign new_new_n11300__ = new_new_n11296__ & new_new_n11299__;
  assign new_new_n11301__ = ys__n432 & ys__n448;
  assign new_new_n11302__ = ys__n428 & ys__n430;
  assign new_new_n11303__ = new_new_n11301__ & new_new_n11302__;
  assign new_new_n11304__ = new_new_n11300__ & new_new_n11303__;
  assign new_new_n11305__ = ys__n426 & new_new_n11304__;
  assign new_new_n11306__ = ~ys__n450 & new_new_n11305__;
  assign new_new_n11307__ = ys__n450 & ~new_new_n11305__;
  assign new_new_n11308__ = ~new_new_n11306__ & ~new_new_n11307__;
  assign new_new_n11309__ = new_new_n11292__ & ~new_new_n11308__;
  assign ys__n23539 = new_new_n11293__ | new_new_n11309__;
  assign new_new_n11311__ = new_new_n11270__ & ys__n23539;
  assign new_new_n11312__ = ~new_new_n11271__ & ~new_new_n11311__;
  assign new_new_n11313__ = ~new_new_n10651__ & ~new_new_n11203__;
  assign new_new_n11314__ = ~ys__n23717 & ~ys__n23730;
  assign new_new_n11315__ = ~ys__n28243 & new_new_n11314__;
  assign new_new_n11316__ = ~new_new_n11313__ & new_new_n11315__;
  assign new_new_n11317__ = ~ys__n23729 & ys__n23730;
  assign new_new_n11318__ = ~new_new_n11316__ & ~new_new_n11317__;
  assign new_new_n11319__ = ys__n23627 & ~new_new_n11318__;
  assign new_new_n11320__ = new_new_n11205__ & new_new_n11315__;
  assign new_new_n11321__ = ys__n23729 & ys__n23730;
  assign new_new_n11322__ = ~new_new_n11320__ & ~new_new_n11321__;
  assign new_new_n11323__ = ys__n23627 & ~new_new_n11322__;
  assign new_new_n11324__ = ~new_new_n11319__ & ~new_new_n11323__;
  assign new_new_n11325__ = ~new_new_n11312__ & new_new_n11324__;
  assign new_new_n11326__ = ys__n450 & ~new_new_n11324__;
  assign new_new_n11327__ = ~new_new_n11325__ & ~new_new_n11326__;
  assign new_new_n11328__ = new_new_n11190__ & ~new_new_n11225__;
  assign new_new_n11329__ = new_new_n11193__ & ~new_new_n11232__;
  assign new_new_n11330__ = new_new_n11202__ & ~new_new_n11329__;
  assign new_new_n11331__ = ~new_new_n11328__ & new_new_n11330__;
  assign new_new_n11332__ = new_new_n11191__ & ~new_new_n11238__;
  assign new_new_n11333__ = new_new_n11194__ & ~new_new_n11242__;
  assign new_new_n11334__ = ~new_new_n11332__ & ~new_new_n11333__;
  assign new_new_n11335__ = new_new_n11331__ & new_new_n11334__;
  assign new_new_n11336__ = ~new_new_n11193__ & ~new_new_n11194__;
  assign new_new_n11337__ = new_new_n11192__ & new_new_n11336__;
  assign new_new_n11338__ = new_new_n11202__ & new_new_n11337__;
  assign new_new_n11339__ = ~ys__n28243 & ~new_new_n11338__;
  assign new_new_n11340__ = ~new_new_n11335__ & new_new_n11339__;
  assign new_new_n11341__ = ys__n28243 & new_new_n10656__;
  assign new_new_n11342__ = ~new_new_n11340__ & ~new_new_n11341__;
  assign new_new_n11343__ = new_new_n11269__ & ~new_new_n11342__;
  assign new_new_n11344__ = ~new_new_n11327__ & ~new_new_n11343__;
  assign new_new_n11345__ = ys__n634 & ~ys__n28243;
  assign new_new_n11346__ = ~ys__n256 & ~ys__n744;
  assign new_new_n11347__ = ys__n550 & new_new_n11346__;
  assign new_new_n11348__ = ys__n256 & ys__n28641;
  assign new_new_n11349__ = ~ys__n256 & ys__n744;
  assign new_new_n11350__ = ys__n4488 & new_new_n11349__;
  assign new_new_n11351__ = ~new_new_n11348__ & ~new_new_n11350__;
  assign new_new_n11352__ = ~new_new_n11347__ & new_new_n11351__;
  assign new_new_n11353__ = ~ys__n256 & ~new_new_n11349__;
  assign new_new_n11354__ = ~new_new_n11346__ & new_new_n11353__;
  assign new_new_n11355__ = ys__n28243 & ~new_new_n11354__;
  assign new_new_n11356__ = ~new_new_n11352__ & new_new_n11355__;
  assign new_new_n11357__ = ~new_new_n11345__ & ~new_new_n11356__;
  assign new_new_n11358__ = ys__n420 & ~new_new_n11357__;
  assign new_new_n11359__ = ~ys__n420 & ~new_new_n11357__;
  assign new_new_n11360__ = ys__n420 & new_new_n11357__;
  assign new_new_n11361__ = ~new_new_n11359__ & ~new_new_n11360__;
  assign new_new_n11362__ = ys__n528 & ~ys__n28243;
  assign new_new_n11363__ = ys__n526 & new_new_n11346__;
  assign new_new_n11364__ = ys__n256 & ys__n526;
  assign new_new_n11365__ = ys__n526 & new_new_n11349__;
  assign new_new_n11366__ = ~new_new_n11364__ & ~new_new_n11365__;
  assign new_new_n11367__ = ~new_new_n11363__ & new_new_n11366__;
  assign new_new_n11368__ = new_new_n11355__ & ~new_new_n11367__;
  assign new_new_n11369__ = ~new_new_n11362__ & ~new_new_n11368__;
  assign new_new_n11370__ = ~ys__n23548 & ~new_new_n11369__;
  assign new_new_n11371__ = ys__n23548 & new_new_n11369__;
  assign new_new_n11372__ = ~new_new_n11370__ & ~new_new_n11371__;
  assign new_new_n11373__ = ys__n526 & ~ys__n28243;
  assign new_new_n11374__ = ys__n524 & new_new_n11346__;
  assign new_new_n11375__ = ys__n256 & ys__n524;
  assign new_new_n11376__ = ys__n524 & new_new_n11349__;
  assign new_new_n11377__ = ~new_new_n11375__ & ~new_new_n11376__;
  assign new_new_n11378__ = ~new_new_n11374__ & new_new_n11377__;
  assign new_new_n11379__ = new_new_n11355__ & ~new_new_n11378__;
  assign new_new_n11380__ = ~new_new_n11373__ & ~new_new_n11379__;
  assign new_new_n11381__ = ~ys__n23550 & ~new_new_n11380__;
  assign new_new_n11382__ = ys__n23550 & new_new_n11380__;
  assign new_new_n11383__ = ~new_new_n11381__ & ~new_new_n11382__;
  assign new_new_n11384__ = ys__n528 & new_new_n11346__;
  assign new_new_n11385__ = ys__n256 & ys__n528;
  assign new_new_n11386__ = ys__n528 & new_new_n11349__;
  assign new_new_n11387__ = ~new_new_n11385__ & ~new_new_n11386__;
  assign new_new_n11388__ = ~new_new_n11384__ & new_new_n11387__;
  assign new_new_n11389__ = new_new_n11355__ & ~new_new_n11388__;
  assign new_new_n11390__ = ys__n22464 & new_new_n11389__;
  assign new_new_n11391__ = ~new_new_n11383__ & new_new_n11390__;
  assign new_new_n11392__ = ~new_new_n11372__ & new_new_n11391__;
  assign new_new_n11393__ = ys__n23550 & ~new_new_n11380__;
  assign new_new_n11394__ = ys__n23548 & ~new_new_n11369__;
  assign new_new_n11395__ = ~new_new_n11383__ & new_new_n11394__;
  assign new_new_n11396__ = ~new_new_n11393__ & ~new_new_n11395__;
  assign new_new_n11397__ = ~new_new_n11392__ & new_new_n11396__;
  assign new_new_n11398__ = ys__n752 & ~ys__n28243;
  assign new_new_n11399__ = ys__n736 & new_new_n11346__;
  assign new_new_n11400__ = ys__n256 & ys__n28633;
  assign new_new_n11401__ = ys__n736 & new_new_n11349__;
  assign new_new_n11402__ = ~new_new_n11400__ & ~new_new_n11401__;
  assign new_new_n11403__ = ~new_new_n11399__ & new_new_n11402__;
  assign new_new_n11404__ = new_new_n11355__ & ~new_new_n11403__;
  assign new_new_n11405__ = ~new_new_n11398__ & ~new_new_n11404__;
  assign new_new_n11406__ = ~ys__n23558 & ~new_new_n11405__;
  assign new_new_n11407__ = ys__n23558 & new_new_n11405__;
  assign new_new_n11408__ = ~new_new_n11406__ & ~new_new_n11407__;
  assign new_new_n11409__ = ys__n530 & ~ys__n28243;
  assign new_new_n11410__ = ys__n752 & new_new_n11346__;
  assign new_new_n11411__ = ys__n256 & ys__n28632;
  assign new_new_n11412__ = ys__n752 & new_new_n11349__;
  assign new_new_n11413__ = ~new_new_n11411__ & ~new_new_n11412__;
  assign new_new_n11414__ = ~new_new_n11410__ & new_new_n11413__;
  assign new_new_n11415__ = new_new_n11355__ & ~new_new_n11414__;
  assign new_new_n11416__ = ~new_new_n11409__ & ~new_new_n11415__;
  assign new_new_n11417__ = ~ys__n23556 & ~new_new_n11416__;
  assign new_new_n11418__ = ys__n23556 & new_new_n11416__;
  assign new_new_n11419__ = ~new_new_n11417__ & ~new_new_n11418__;
  assign new_new_n11420__ = ~new_new_n11408__ & ~new_new_n11419__;
  assign new_new_n11421__ = ys__n522 & ~ys__n28243;
  assign new_new_n11422__ = ys__n530 & new_new_n11346__;
  assign new_new_n11423__ = ys__n256 & ys__n530;
  assign new_new_n11424__ = ys__n530 & new_new_n11349__;
  assign new_new_n11425__ = ~new_new_n11423__ & ~new_new_n11424__;
  assign new_new_n11426__ = ~new_new_n11422__ & new_new_n11425__;
  assign new_new_n11427__ = new_new_n11355__ & ~new_new_n11426__;
  assign new_new_n11428__ = ~new_new_n11421__ & ~new_new_n11427__;
  assign new_new_n11429__ = ~ys__n23554 & ~new_new_n11428__;
  assign new_new_n11430__ = ys__n23554 & new_new_n11428__;
  assign new_new_n11431__ = ~new_new_n11429__ & ~new_new_n11430__;
  assign new_new_n11432__ = ys__n524 & ~ys__n28243;
  assign new_new_n11433__ = ys__n522 & new_new_n11346__;
  assign new_new_n11434__ = ys__n256 & ys__n522;
  assign new_new_n11435__ = ys__n522 & new_new_n11349__;
  assign new_new_n11436__ = ~new_new_n11434__ & ~new_new_n11435__;
  assign new_new_n11437__ = ~new_new_n11433__ & new_new_n11436__;
  assign new_new_n11438__ = new_new_n11355__ & ~new_new_n11437__;
  assign new_new_n11439__ = ~new_new_n11432__ & ~new_new_n11438__;
  assign new_new_n11440__ = ~ys__n23552 & ~new_new_n11439__;
  assign new_new_n11441__ = ys__n23552 & new_new_n11439__;
  assign new_new_n11442__ = ~new_new_n11440__ & ~new_new_n11441__;
  assign new_new_n11443__ = ~new_new_n11431__ & ~new_new_n11442__;
  assign new_new_n11444__ = new_new_n11420__ & new_new_n11443__;
  assign new_new_n11445__ = ~new_new_n11397__ & new_new_n11444__;
  assign new_new_n11446__ = ys__n23554 & ~new_new_n11428__;
  assign new_new_n11447__ = ys__n23552 & ~new_new_n11439__;
  assign new_new_n11448__ = ~new_new_n11431__ & new_new_n11447__;
  assign new_new_n11449__ = ~new_new_n11446__ & ~new_new_n11448__;
  assign new_new_n11450__ = new_new_n11420__ & ~new_new_n11449__;
  assign new_new_n11451__ = ys__n23558 & ~new_new_n11405__;
  assign new_new_n11452__ = ys__n23556 & ~new_new_n11416__;
  assign new_new_n11453__ = ~new_new_n11408__ & new_new_n11452__;
  assign new_new_n11454__ = ~new_new_n11451__ & ~new_new_n11453__;
  assign new_new_n11455__ = ~new_new_n11450__ & new_new_n11454__;
  assign new_new_n11456__ = ~new_new_n11445__ & new_new_n11455__;
  assign new_new_n11457__ = ys__n636 & ~ys__n28243;
  assign new_new_n11458__ = ys__n256 & ys__n28640;
  assign new_new_n11459__ = ~new_new_n11350__ & ~new_new_n11458__;
  assign new_new_n11460__ = ~new_new_n11347__ & new_new_n11459__;
  assign new_new_n11461__ = new_new_n11355__ & ~new_new_n11460__;
  assign new_new_n11462__ = ~new_new_n11457__ & ~new_new_n11461__;
  assign new_new_n11463__ = ~ys__n23574 & ~new_new_n11462__;
  assign new_new_n11464__ = ys__n23574 & new_new_n11462__;
  assign new_new_n11465__ = ~new_new_n11463__ & ~new_new_n11464__;
  assign new_new_n11466__ = ys__n638 & ~ys__n28243;
  assign new_new_n11467__ = ys__n256 & ys__n28639;
  assign new_new_n11468__ = ~new_new_n11350__ & ~new_new_n11467__;
  assign new_new_n11469__ = ~new_new_n11347__ & new_new_n11468__;
  assign new_new_n11470__ = new_new_n11355__ & ~new_new_n11469__;
  assign new_new_n11471__ = ~new_new_n11466__ & ~new_new_n11470__;
  assign new_new_n11472__ = ~ys__n23572 & ~new_new_n11471__;
  assign new_new_n11473__ = ys__n23572 & new_new_n11471__;
  assign new_new_n11474__ = ~new_new_n11472__ & ~new_new_n11473__;
  assign new_new_n11475__ = ~new_new_n11465__ & ~new_new_n11474__;
  assign new_new_n11476__ = ys__n640 & ~ys__n28243;
  assign new_new_n11477__ = ys__n256 & ys__n28638;
  assign new_new_n11478__ = ~new_new_n11350__ & ~new_new_n11477__;
  assign new_new_n11479__ = ~new_new_n11347__ & new_new_n11478__;
  assign new_new_n11480__ = new_new_n11355__ & ~new_new_n11479__;
  assign new_new_n11481__ = ~new_new_n11476__ & ~new_new_n11480__;
  assign new_new_n11482__ = ~ys__n23570 & ~new_new_n11481__;
  assign new_new_n11483__ = ys__n23570 & new_new_n11481__;
  assign new_new_n11484__ = ~new_new_n11482__ & ~new_new_n11483__;
  assign new_new_n11485__ = ys__n550 & ~ys__n28243;
  assign new_new_n11486__ = ys__n256 & ys__n28637;
  assign new_new_n11487__ = ~new_new_n11350__ & ~new_new_n11486__;
  assign new_new_n11488__ = ~new_new_n11347__ & new_new_n11487__;
  assign new_new_n11489__ = new_new_n11355__ & ~new_new_n11488__;
  assign new_new_n11490__ = ~new_new_n11485__ & ~new_new_n11489__;
  assign new_new_n11491__ = ~ys__n23568 & ~new_new_n11490__;
  assign new_new_n11492__ = ys__n23568 & new_new_n11490__;
  assign new_new_n11493__ = ~new_new_n11491__ & ~new_new_n11492__;
  assign new_new_n11494__ = ~new_new_n11484__ & ~new_new_n11493__;
  assign new_new_n11495__ = new_new_n11475__ & new_new_n11494__;
  assign new_new_n11496__ = ys__n548 & ~ys__n28243;
  assign new_new_n11497__ = ys__n256 & ys__n47660;
  assign new_new_n11498__ = ~new_new_n11350__ & ~new_new_n11497__;
  assign new_new_n11499__ = ~new_new_n11347__ & new_new_n11498__;
  assign new_new_n11500__ = new_new_n11355__ & ~new_new_n11499__;
  assign new_new_n11501__ = ~new_new_n11496__ & ~new_new_n11500__;
  assign new_new_n11502__ = ~ys__n23566 & ~new_new_n11501__;
  assign new_new_n11503__ = ys__n23566 & new_new_n11501__;
  assign new_new_n11504__ = ~new_new_n11502__ & ~new_new_n11503__;
  assign new_new_n11505__ = ys__n518 & ~ys__n28243;
  assign new_new_n11506__ = ys__n548 & new_new_n11346__;
  assign new_new_n11507__ = ys__n256 & ys__n28636;
  assign new_new_n11508__ = ~new_new_n11350__ & ~new_new_n11507__;
  assign new_new_n11509__ = ~new_new_n11506__ & new_new_n11508__;
  assign new_new_n11510__ = new_new_n11355__ & ~new_new_n11509__;
  assign new_new_n11511__ = ~new_new_n11505__ & ~new_new_n11510__;
  assign new_new_n11512__ = ~ys__n23564 & ~new_new_n11511__;
  assign new_new_n11513__ = ys__n23564 & new_new_n11511__;
  assign new_new_n11514__ = ~new_new_n11512__ & ~new_new_n11513__;
  assign new_new_n11515__ = ~new_new_n11504__ & ~new_new_n11514__;
  assign new_new_n11516__ = ys__n4488 & ~ys__n28243;
  assign new_new_n11517__ = ys__n518 & new_new_n11346__;
  assign new_new_n11518__ = ys__n256 & ys__n28635;
  assign new_new_n11519__ = ~new_new_n11350__ & ~new_new_n11518__;
  assign new_new_n11520__ = ~new_new_n11517__ & new_new_n11519__;
  assign new_new_n11521__ = new_new_n11355__ & ~new_new_n11520__;
  assign new_new_n11522__ = ~new_new_n11516__ & ~new_new_n11521__;
  assign new_new_n11523__ = ~ys__n23562 & ~new_new_n11522__;
  assign new_new_n11524__ = ys__n23562 & new_new_n11522__;
  assign new_new_n11525__ = ~new_new_n11523__ & ~new_new_n11524__;
  assign new_new_n11526__ = ys__n736 & ~ys__n28243;
  assign new_new_n11527__ = ys__n4488 & new_new_n11346__;
  assign new_new_n11528__ = ys__n256 & ys__n28634;
  assign new_new_n11529__ = ~new_new_n11350__ & ~new_new_n11528__;
  assign new_new_n11530__ = ~new_new_n11527__ & new_new_n11529__;
  assign new_new_n11531__ = new_new_n11355__ & ~new_new_n11530__;
  assign new_new_n11532__ = ~new_new_n11526__ & ~new_new_n11531__;
  assign new_new_n11533__ = ~ys__n23560 & ~new_new_n11532__;
  assign new_new_n11534__ = ys__n23560 & new_new_n11532__;
  assign new_new_n11535__ = ~new_new_n11533__ & ~new_new_n11534__;
  assign new_new_n11536__ = ~new_new_n11525__ & ~new_new_n11535__;
  assign new_new_n11537__ = new_new_n11515__ & new_new_n11536__;
  assign new_new_n11538__ = new_new_n11495__ & new_new_n11537__;
  assign new_new_n11539__ = ~new_new_n11456__ & new_new_n11538__;
  assign new_new_n11540__ = ys__n23562 & ~new_new_n11522__;
  assign new_new_n11541__ = ys__n23560 & ~new_new_n11532__;
  assign new_new_n11542__ = ~new_new_n11525__ & new_new_n11541__;
  assign new_new_n11543__ = ~new_new_n11540__ & ~new_new_n11542__;
  assign new_new_n11544__ = new_new_n11515__ & ~new_new_n11543__;
  assign new_new_n11545__ = ys__n23566 & ~new_new_n11501__;
  assign new_new_n11546__ = ys__n23564 & ~new_new_n11511__;
  assign new_new_n11547__ = ~new_new_n11504__ & new_new_n11546__;
  assign new_new_n11548__ = ~new_new_n11545__ & ~new_new_n11547__;
  assign new_new_n11549__ = ~new_new_n11544__ & new_new_n11548__;
  assign new_new_n11550__ = new_new_n11495__ & ~new_new_n11549__;
  assign new_new_n11551__ = ys__n23570 & ~new_new_n11481__;
  assign new_new_n11552__ = ys__n23568 & ~new_new_n11490__;
  assign new_new_n11553__ = ~new_new_n11484__ & new_new_n11552__;
  assign new_new_n11554__ = ~new_new_n11551__ & ~new_new_n11553__;
  assign new_new_n11555__ = new_new_n11475__ & ~new_new_n11554__;
  assign new_new_n11556__ = ys__n23574 & ~new_new_n11462__;
  assign new_new_n11557__ = ys__n23572 & ~new_new_n11471__;
  assign new_new_n11558__ = ~new_new_n11465__ & new_new_n11557__;
  assign new_new_n11559__ = ~new_new_n11556__ & ~new_new_n11558__;
  assign new_new_n11560__ = ~new_new_n11555__ & new_new_n11559__;
  assign new_new_n11561__ = ~new_new_n11550__ & new_new_n11560__;
  assign new_new_n11562__ = ~new_new_n11539__ & new_new_n11561__;
  assign new_new_n11563__ = ~new_new_n11361__ & ~new_new_n11562__;
  assign new_new_n11564__ = ~new_new_n11358__ & ~new_new_n11563__;
  assign new_new_n11565__ = ys__n642 & ~ys__n28243;
  assign new_new_n11566__ = ~new_new_n11356__ & ~new_new_n11565__;
  assign new_new_n11567__ = new_new_n11564__ & new_new_n11566__;
  assign new_new_n11568__ = ~new_new_n11564__ & ~new_new_n11566__;
  assign new_new_n11569__ = ~new_new_n11567__ & ~new_new_n11568__;
  assign new_new_n11570__ = ys__n450 & ~new_new_n11569__;
  assign new_new_n11571__ = ~ys__n440 & ys__n442;
  assign new_new_n11572__ = ~ys__n440 & ~new_new_n11571__;
  assign new_new_n11573__ = ~ys__n438 & ~ys__n444;
  assign new_new_n11574__ = ~new_new_n11572__ & new_new_n11573__;
  assign new_new_n11575__ = ~ys__n438 & ys__n444;
  assign new_new_n11576__ = ~ys__n438 & ~new_new_n11575__;
  assign new_new_n11577__ = ~new_new_n11574__ & new_new_n11576__;
  assign new_new_n11578__ = ~ys__n432 & ~ys__n436;
  assign new_new_n11579__ = ~ys__n434 & ~ys__n446;
  assign new_new_n11580__ = new_new_n11578__ & new_new_n11579__;
  assign new_new_n11581__ = ~new_new_n11577__ & new_new_n11580__;
  assign new_new_n11582__ = ~ys__n434 & ys__n446;
  assign new_new_n11583__ = ~ys__n434 & ~new_new_n11582__;
  assign new_new_n11584__ = new_new_n11578__ & ~new_new_n11583__;
  assign new_new_n11585__ = ~ys__n432 & ys__n436;
  assign new_new_n11586__ = ~ys__n432 & ~new_new_n11585__;
  assign new_new_n11587__ = ~new_new_n11584__ & new_new_n11586__;
  assign new_new_n11588__ = ~new_new_n11581__ & new_new_n11587__;
  assign new_new_n11589__ = ~ys__n426 & ~ys__n430;
  assign new_new_n11590__ = ~ys__n428 & ~ys__n448;
  assign new_new_n11591__ = new_new_n11589__ & new_new_n11590__;
  assign new_new_n11592__ = ~new_new_n11588__ & new_new_n11591__;
  assign new_new_n11593__ = ~ys__n428 & ys__n448;
  assign new_new_n11594__ = ~ys__n428 & ~new_new_n11593__;
  assign new_new_n11595__ = new_new_n11589__ & ~new_new_n11594__;
  assign new_new_n11596__ = ~ys__n426 & ys__n430;
  assign new_new_n11597__ = ~ys__n426 & ~new_new_n11596__;
  assign new_new_n11598__ = ~new_new_n11595__ & new_new_n11597__;
  assign new_new_n11599__ = ~new_new_n11592__ & new_new_n11598__;
  assign new_new_n11600__ = ys__n450 & ~new_new_n11599__;
  assign new_new_n11601__ = ~ys__n450 & new_new_n11599__;
  assign new_new_n11602__ = ~new_new_n11600__ & ~new_new_n11601__;
  assign new_new_n11603__ = new_new_n11564__ & ~new_new_n11566__;
  assign new_new_n11604__ = ~new_new_n11602__ & new_new_n11603__;
  assign new_new_n11605__ = ys__n428 & ys__n448;
  assign new_new_n11606__ = ys__n426 & ys__n430;
  assign new_new_n11607__ = new_new_n11605__ & new_new_n11606__;
  assign new_new_n11608__ = ys__n440 & ys__n442;
  assign new_new_n11609__ = ys__n438 & ys__n444;
  assign new_new_n11610__ = new_new_n11608__ & new_new_n11609__;
  assign new_new_n11611__ = ys__n434 & ys__n446;
  assign new_new_n11612__ = ys__n432 & ys__n436;
  assign new_new_n11613__ = new_new_n11611__ & new_new_n11612__;
  assign new_new_n11614__ = new_new_n11610__ & new_new_n11613__;
  assign new_new_n11615__ = new_new_n11607__ & new_new_n11614__;
  assign new_new_n11616__ = ~ys__n450 & new_new_n11615__;
  assign new_new_n11617__ = ys__n450 & ~new_new_n11615__;
  assign new_new_n11618__ = ~new_new_n11616__ & ~new_new_n11617__;
  assign new_new_n11619__ = ~new_new_n11564__ & new_new_n11566__;
  assign new_new_n11620__ = ~new_new_n11618__ & new_new_n11619__;
  assign new_new_n11621__ = ~new_new_n11604__ & ~new_new_n11620__;
  assign new_new_n11622__ = ~new_new_n11570__ & new_new_n11621__;
  assign new_new_n11623__ = ~new_new_n11603__ & ~new_new_n11619__;
  assign new_new_n11624__ = new_new_n11569__ & new_new_n11623__;
  assign new_new_n11625__ = new_new_n11343__ & ~new_new_n11624__;
  assign new_new_n11626__ = ~new_new_n11622__ & new_new_n11625__;
  assign new_new_n11627__ = ~new_new_n11344__ & ~new_new_n11626__;
  assign new_new_n11628__ = ys__n23627 & ys__n4566;
  assign new_new_n11629__ = ~new_new_n10686__ & ~new_new_n11628__;
  assign new_new_n11630__ = ~new_new_n11627__ & new_new_n11629__;
  assign new_new_n11631__ = ~ys__n935 & ys__n28446;
  assign new_new_n11632__ = ~ys__n935 & ~new_new_n11631__;
  assign new_new_n11633__ = new_new_n11628__ & ~new_new_n11632__;
  assign new_new_n11634__ = new_new_n10686__ & ~new_new_n11628__;
  assign new_new_n11635__ = ys__n47690 & new_new_n11634__;
  assign new_new_n11636__ = ~new_new_n11633__ & ~new_new_n11635__;
  assign new_new_n11637__ = ~new_new_n11630__ & new_new_n11636__;
  assign new_new_n11638__ = ~new_new_n11628__ & ~new_new_n11634__;
  assign new_new_n11639__ = ~new_new_n11629__ & new_new_n11638__;
  assign new_new_n11640__ = new_new_n10813__ & ~new_new_n11639__;
  assign new_new_n11641__ = ~new_new_n11637__ & new_new_n11640__;
  assign new_new_n11642__ = ~new_new_n10818__ & ~new_new_n11628__;
  assign new_new_n11643__ = ~new_new_n11627__ & new_new_n11642__;
  assign new_new_n11644__ = new_new_n10818__ & ~new_new_n11628__;
  assign new_new_n11645__ = ys__n47690 & new_new_n11644__;
  assign new_new_n11646__ = ~new_new_n11633__ & ~new_new_n11645__;
  assign new_new_n11647__ = ~new_new_n11643__ & new_new_n11646__;
  assign new_new_n11648__ = ~new_new_n11628__ & ~new_new_n11644__;
  assign new_new_n11649__ = ~new_new_n11642__ & new_new_n11648__;
  assign new_new_n11650__ = ~new_new_n10813__ & ~new_new_n11649__;
  assign new_new_n11651__ = ~new_new_n11647__ & new_new_n11650__;
  assign ys__n714 = new_new_n11641__ | new_new_n11651__;
  assign new_new_n11653__ = ys__n22884 & new_new_n11175__;
  assign new_new_n11654__ = ~new_new_n11176__ & ~new_new_n11653__;
  assign new_new_n11655__ = ~new_new_n11180__ & ~new_new_n11654__;
  assign new_new_n11656__ = ys__n23332 & new_new_n11180__;
  assign new_new_n11657__ = ~new_new_n11655__ & ~new_new_n11656__;
  assign new_new_n11658__ = ~new_new_n11186__ & ~new_new_n11657__;
  assign new_new_n11659__ = ys__n422 & new_new_n11186__;
  assign new_new_n11660__ = ~new_new_n11658__ & ~new_new_n11659__;
  assign new_new_n11661__ = ~new_new_n11270__ & ~new_new_n11660__;
  assign new_new_n11662__ = ys__n422 & ~new_new_n11292__;
  assign new_new_n11663__ = ys__n426 & ys__n450;
  assign new_new_n11664__ = new_new_n11304__ & new_new_n11663__;
  assign new_new_n11665__ = ys__n424 & new_new_n11664__;
  assign new_new_n11666__ = ~ys__n422 & new_new_n11665__;
  assign new_new_n11667__ = ys__n422 & ~new_new_n11665__;
  assign new_new_n11668__ = ~new_new_n11666__ & ~new_new_n11667__;
  assign new_new_n11669__ = new_new_n11292__ & ~new_new_n11668__;
  assign ys__n23543 = new_new_n11662__ | new_new_n11669__;
  assign new_new_n11671__ = new_new_n11270__ & ys__n23543;
  assign new_new_n11672__ = ~new_new_n11661__ & ~new_new_n11671__;
  assign new_new_n11673__ = new_new_n11324__ & ~new_new_n11672__;
  assign new_new_n11674__ = ys__n422 & ~new_new_n11324__;
  assign new_new_n11675__ = ~new_new_n11673__ & ~new_new_n11674__;
  assign new_new_n11676__ = ~new_new_n11343__ & ~new_new_n11675__;
  assign new_new_n11677__ = ys__n422 & ~new_new_n11569__;
  assign new_new_n11678__ = ~ys__n424 & ~ys__n450;
  assign new_new_n11679__ = ~new_new_n11599__ & new_new_n11678__;
  assign new_new_n11680__ = ~ys__n424 & ys__n450;
  assign new_new_n11681__ = ~ys__n424 & ~new_new_n11680__;
  assign new_new_n11682__ = ~new_new_n11679__ & new_new_n11681__;
  assign new_new_n11683__ = ys__n422 & ~new_new_n11682__;
  assign new_new_n11684__ = ~ys__n422 & new_new_n11682__;
  assign new_new_n11685__ = ~new_new_n11683__ & ~new_new_n11684__;
  assign new_new_n11686__ = new_new_n11603__ & ~new_new_n11685__;
  assign new_new_n11687__ = ys__n424 & ys__n450;
  assign new_new_n11688__ = new_new_n11615__ & new_new_n11687__;
  assign new_new_n11689__ = ~ys__n422 & new_new_n11688__;
  assign new_new_n11690__ = ys__n422 & ~new_new_n11688__;
  assign new_new_n11691__ = ~new_new_n11689__ & ~new_new_n11690__;
  assign new_new_n11692__ = new_new_n11619__ & ~new_new_n11691__;
  assign new_new_n11693__ = ~new_new_n11686__ & ~new_new_n11692__;
  assign new_new_n11694__ = ~new_new_n11677__ & new_new_n11693__;
  assign new_new_n11695__ = new_new_n11625__ & ~new_new_n11694__;
  assign new_new_n11696__ = ~new_new_n11676__ & ~new_new_n11695__;
  assign new_new_n11697__ = new_new_n11629__ & ~new_new_n11696__;
  assign new_new_n11698__ = ys__n38311 & new_new_n11634__;
  assign new_new_n11699__ = ~new_new_n11628__ & ~new_new_n11698__;
  assign new_new_n11700__ = ~new_new_n11697__ & new_new_n11699__;
  assign new_new_n11701__ = new_new_n11640__ & ~new_new_n11700__;
  assign new_new_n11702__ = new_new_n11642__ & ~new_new_n11696__;
  assign new_new_n11703__ = ys__n38311 & new_new_n11644__;
  assign new_new_n11704__ = ~new_new_n11628__ & ~new_new_n11703__;
  assign new_new_n11705__ = ~new_new_n11702__ & new_new_n11704__;
  assign new_new_n11706__ = new_new_n11650__ & ~new_new_n11705__;
  assign ys__n716 = new_new_n11701__ | new_new_n11706__;
  assign new_new_n11708__ = ys__n19203 & ys__n38178;
  assign new_new_n11709__ = ~new_new_n11078__ & ~new_new_n11080__;
  assign new_new_n11710__ = new_new_n11708__ & ~new_new_n11709__;
  assign new_new_n11711__ = ~ys__n1301 & ys__n1309;
  assign new_new_n11712__ = ~ys__n1301 & ys__n19215;
  assign new_new_n11713__ = ys__n19203 & new_new_n11081__;
  assign new_new_n11714__ = new_new_n11712__ & new_new_n11713__;
  assign new_new_n11715__ = ~new_new_n11711__ & ~new_new_n11714__;
  assign new_new_n11716__ = ~new_new_n11710__ & new_new_n11715__;
  assign new_new_n11717__ = new_new_n11082__ & new_new_n11709__;
  assign ys__n732 = ~new_new_n11716__ & ~new_new_n11717__;
  assign new_new_n11719__ = ~ys__n37670 & ys__n37671;
  assign new_new_n11720__ = ys__n37670 & ~ys__n37671;
  assign new_new_n11721__ = ~new_new_n11719__ & ~new_new_n11720__;
  assign new_new_n11722__ = ~ys__n18393 & ~new_new_n11721__;
  assign new_new_n11723__ = ~ys__n18393 & ~new_new_n11722__;
  assign new_new_n11724__ = ~ys__n18393 & ~new_new_n11723__;
  assign new_new_n11725__ = ys__n18393 & ys__n27738;
  assign new_new_n11726__ = ~new_new_n11724__ & ~new_new_n11725__;
  assign new_new_n11727__ = ys__n732 & new_new_n11726__;
  assign new_new_n11728__ = ys__n826 & ~new_new_n11727__;
  assign new_new_n11729__ = ys__n828 & new_new_n11727__;
  assign new_new_n11730__ = ~new_new_n11728__ & ~new_new_n11729__;
  assign new_new_n11731__ = ~ys__n732 & ~new_new_n11726__;
  assign new_new_n11732__ = ~new_new_n11730__ & ~new_new_n11731__;
  assign new_new_n11733__ = ys__n824 & new_new_n11731__;
  assign ys__n730 = new_new_n11732__ | new_new_n11733__;
  assign new_new_n11735__ = ~ys__n889 & ~ys__n4184;
  assign new_new_n11736__ = ~ys__n4192 & new_new_n11735__;
  assign new_new_n11737__ = new_new_n10613__ & new_new_n11736__;
  assign ys__n740 = ~new_new_n10611__ | ~new_new_n11737__;
  assign new_new_n11739__ = ys__n23641 & ~ys__n23645;
  assign new_new_n11740__ = ys__n23645 & ys__n23650;
  assign new_new_n11741__ = ~new_new_n11739__ & ~new_new_n11740__;
  assign ys__n754 = ~ys__n23652 & ~new_new_n11741__;
  assign new_new_n11743__ = ys__n23645 & ys__n23647;
  assign ys__n756 = ~ys__n23652 & new_new_n11743__;
  assign new_new_n11745__ = ys__n108 & new_new_n11086__;
  assign new_new_n11746__ = ~ys__n19203 & new_new_n11081__;
  assign new_new_n11747__ = ~new_new_n11066__ & ~new_new_n11746__;
  assign new_new_n11748__ = ~new_new_n11086__ & ~new_new_n11747__;
  assign ys__n786 = new_new_n11745__ | new_new_n11748__;
  assign new_new_n11750__ = ys__n1301 & ys__n1309;
  assign new_new_n11751__ = ys__n1301 & ys__n19203;
  assign new_new_n11752__ = ys__n19215 & new_new_n11751__;
  assign new_new_n11753__ = new_new_n11081__ & new_new_n11752__;
  assign new_new_n11754__ = ~new_new_n11750__ & ~new_new_n11753__;
  assign ys__n788 = ~new_new_n11086__ & ~new_new_n11754__;
  assign new_new_n11756__ = ys__n118 & new_new_n11086__;
  assign new_new_n11757__ = ~new_new_n11147__ & ~new_new_n11149__;
  assign new_new_n11758__ = ~new_new_n11147__ & ~new_new_n11757__;
  assign new_new_n11759__ = ~new_new_n11141__ & ~new_new_n11758__;
  assign new_new_n11760__ = ~new_new_n11141__ & ~new_new_n11759__;
  assign new_new_n11761__ = new_new_n11076__ & ~new_new_n11760__;
  assign new_new_n11762__ = ~ys__n19215 & ~new_new_n11143__;
  assign new_new_n11763__ = ~new_new_n11712__ & ~new_new_n11762__;
  assign new_new_n11764__ = new_new_n11713__ & ~new_new_n11763__;
  assign new_new_n11765__ = new_new_n11080__ & new_new_n11708__;
  assign new_new_n11766__ = ~new_new_n11711__ & ~new_new_n11765__;
  assign new_new_n11767__ = ~new_new_n11764__ & new_new_n11766__;
  assign new_new_n11768__ = ~new_new_n11761__ & new_new_n11767__;
  assign new_new_n11769__ = ~new_new_n11086__ & ~new_new_n11768__;
  assign ys__n790 = new_new_n11756__ | new_new_n11769__;
  assign new_new_n11771__ = ys__n290 & new_new_n11086__;
  assign new_new_n11772__ = ~ys__n18389 & new_new_n11071__;
  assign new_new_n11773__ = new_new_n11080__ & ~new_new_n11708__;
  assign new_new_n11774__ = ~ys__n308 & ~ys__n310;
  assign new_new_n11775__ = new_new_n11708__ & new_new_n11774__;
  assign new_new_n11776__ = new_new_n11078__ & new_new_n11775__;
  assign new_new_n11777__ = ~new_new_n11773__ & ~new_new_n11776__;
  assign new_new_n11778__ = ~new_new_n11772__ & new_new_n11777__;
  assign new_new_n11779__ = ~new_new_n11086__ & ~new_new_n11778__;
  assign ys__n792 = new_new_n11771__ | new_new_n11779__;
  assign new_new_n11781__ = ys__n110 & new_new_n11086__;
  assign new_new_n11782__ = new_new_n11708__ & ~new_new_n11774__;
  assign new_new_n11783__ = new_new_n11708__ & ~new_new_n11782__;
  assign new_new_n11784__ = new_new_n11078__ & ~new_new_n11783__;
  assign new_new_n11785__ = ys__n18389 & new_new_n11071__;
  assign new_new_n11786__ = ~new_new_n11784__ & ~new_new_n11785__;
  assign new_new_n11787__ = ~new_new_n11086__ & ~new_new_n11786__;
  assign ys__n794 = new_new_n11781__ | new_new_n11787__;
  assign new_new_n11789__ = ys__n18283 & new_new_n11130__;
  assign ys__n37676 = ys__n18070 | new_new_n11125__;
  assign new_new_n11791__ = ~ys__n3214 & ys__n37676;
  assign new_new_n11792__ = ~ys__n3214 & ~new_new_n11791__;
  assign new_new_n11793__ = ~ys__n844 & new_new_n11122__;
  assign new_new_n11794__ = ~ys__n37678 & ~ys__n37679;
  assign new_new_n11795__ = ys__n844 & ~new_new_n11794__;
  assign new_new_n11796__ = ys__n844 & ys__n37682;
  assign new_new_n11797__ = ys__n18071 & ~new_new_n11796__;
  assign new_new_n11798__ = ~new_new_n11795__ & new_new_n11797__;
  assign new_new_n11799__ = ~new_new_n11793__ & ~new_new_n11798__;
  assign new_new_n11800__ = new_new_n11792__ & ~new_new_n11799__;
  assign new_new_n11801__ = ~new_new_n11130__ & new_new_n11800__;
  assign new_new_n11802__ = ~new_new_n11789__ & ~new_new_n11801__;
  assign new_new_n11803__ = ~ys__n18271 & ~new_new_n11802__;
  assign new_new_n11804__ = ys__n18271 & ys__n18283;
  assign ys__n18284 = new_new_n11803__ | new_new_n11804__;
  assign new_new_n11806__ = ys__n18286 & new_new_n11130__;
  assign new_new_n11807__ = ys__n844 & new_new_n11792__;
  assign new_new_n11808__ = ~new_new_n11130__ & new_new_n11807__;
  assign new_new_n11809__ = ~new_new_n11800__ & new_new_n11808__;
  assign new_new_n11810__ = ~new_new_n11806__ & ~new_new_n11809__;
  assign new_new_n11811__ = ~ys__n18271 & ~new_new_n11810__;
  assign new_new_n11812__ = ys__n18271 & ys__n18286;
  assign ys__n18287 = new_new_n11811__ | new_new_n11812__;
  assign new_new_n11814__ = ys__n18984 & ys__n18287;
  assign new_new_n11815__ = ~ys__n18284 & new_new_n11814__;
  assign new_new_n11816__ = ys__n54 & ~ys__n4764;
  assign new_new_n11817__ = ys__n24667 & ys__n4764;
  assign ys__n18820 = new_new_n11816__ | new_new_n11817__;
  assign new_new_n11819__ = ~ys__n18071 & ys__n18820;
  assign new_new_n11820__ = ys__n18071 & ys__n18821;
  assign new_new_n11821__ = ~new_new_n11819__ & ~new_new_n11820__;
  assign new_new_n11822__ = ~new_new_n11122__ & ~new_new_n11821__;
  assign new_new_n11823__ = ys__n24667 & ~ys__n24675;
  assign new_new_n11824__ = ys__n24675 & ys__n24707;
  assign ys__n18738 = new_new_n11823__ | new_new_n11824__;
  assign new_new_n11826__ = new_new_n11122__ & ys__n18738;
  assign ys__n18739 = new_new_n11822__ | new_new_n11826__;
  assign new_new_n11828__ = ys__n18284 & ys__n18739;
  assign new_new_n11829__ = ~new_new_n11815__ & ~new_new_n11828__;
  assign new_new_n11830__ = ys__n18280 & new_new_n11130__;
  assign new_new_n11831__ = ~new_new_n11130__ & new_new_n11791__;
  assign new_new_n11832__ = ~new_new_n11830__ & ~new_new_n11831__;
  assign new_new_n11833__ = ~ys__n18271 & ~new_new_n11832__;
  assign new_new_n11834__ = ys__n18271 & ys__n18280;
  assign ys__n18281 = new_new_n11833__ | new_new_n11834__;
  assign new_new_n11836__ = ~new_new_n11829__ & ~ys__n18281;
  assign new_new_n11837__ = ys__n18636 & ~new_new_n11125__;
  assign new_new_n11838__ = ys__n74 & new_new_n11125__;
  assign ys__n18637 = new_new_n11837__ | new_new_n11838__;
  assign new_new_n11840__ = ys__n18281 & ys__n18637;
  assign new_new_n11841__ = ~new_new_n11836__ & ~new_new_n11840__;
  assign new_new_n11842__ = ys__n18277 & new_new_n11130__;
  assign new_new_n11843__ = ys__n3214 & ~new_new_n11130__;
  assign new_new_n11844__ = ~new_new_n11842__ & ~new_new_n11843__;
  assign new_new_n11845__ = ~ys__n18271 & ~new_new_n11844__;
  assign new_new_n11846__ = ys__n18271 & ys__n18277;
  assign ys__n18278 = new_new_n11845__ | new_new_n11846__;
  assign new_new_n11848__ = ~new_new_n11841__ & ~ys__n18278;
  assign new_new_n11849__ = ys__n18885 & ys__n18278;
  assign ys__n796 = new_new_n11848__ | new_new_n11849__;
  assign new_new_n11851__ = ys__n18983 & ys__n18287;
  assign new_new_n11852__ = ~ys__n18284 & new_new_n11851__;
  assign new_new_n11853__ = ys__n56 & ~ys__n4764;
  assign new_new_n11854__ = ys__n24666 & ys__n4764;
  assign ys__n18818 = new_new_n11853__ | new_new_n11854__;
  assign new_new_n11856__ = ~ys__n18071 & ys__n18818;
  assign new_new_n11857__ = ys__n18071 & ys__n18819;
  assign new_new_n11858__ = ~new_new_n11856__ & ~new_new_n11857__;
  assign new_new_n11859__ = ~new_new_n11122__ & ~new_new_n11858__;
  assign new_new_n11860__ = ys__n24666 & ~ys__n24675;
  assign new_new_n11861__ = ys__n24675 & ys__n24706;
  assign ys__n18735 = new_new_n11860__ | new_new_n11861__;
  assign new_new_n11863__ = new_new_n11122__ & ys__n18735;
  assign ys__n18736 = new_new_n11859__ | new_new_n11863__;
  assign new_new_n11865__ = ys__n18284 & ys__n18736;
  assign new_new_n11866__ = ~new_new_n11852__ & ~new_new_n11865__;
  assign new_new_n11867__ = ~ys__n18281 & ~new_new_n11866__;
  assign new_new_n11868__ = ys__n18634 & ~new_new_n11125__;
  assign new_new_n11869__ = ys__n76 & new_new_n11125__;
  assign ys__n18635 = new_new_n11868__ | new_new_n11869__;
  assign new_new_n11871__ = ys__n18281 & ys__n18635;
  assign new_new_n11872__ = ~new_new_n11867__ & ~new_new_n11871__;
  assign new_new_n11873__ = ~ys__n18278 & ~new_new_n11872__;
  assign new_new_n11874__ = ys__n18883 & ys__n18278;
  assign ys__n798 = new_new_n11873__ | new_new_n11874__;
  assign new_new_n11876__ = ys__n18982 & ys__n18287;
  assign new_new_n11877__ = ~ys__n18284 & new_new_n11876__;
  assign new_new_n11878__ = ys__n58 & ~ys__n4764;
  assign new_new_n11879__ = ys__n24665 & ys__n4764;
  assign ys__n18816 = new_new_n11878__ | new_new_n11879__;
  assign new_new_n11881__ = ~ys__n18071 & ys__n18816;
  assign new_new_n11882__ = ys__n18071 & ys__n18817;
  assign new_new_n11883__ = ~new_new_n11881__ & ~new_new_n11882__;
  assign new_new_n11884__ = ~new_new_n11122__ & ~new_new_n11883__;
  assign new_new_n11885__ = ys__n24665 & ~ys__n24675;
  assign new_new_n11886__ = ys__n24675 & ys__n24705;
  assign ys__n18732 = new_new_n11885__ | new_new_n11886__;
  assign new_new_n11888__ = new_new_n11122__ & ys__n18732;
  assign ys__n18733 = new_new_n11884__ | new_new_n11888__;
  assign new_new_n11890__ = ys__n18284 & ys__n18733;
  assign new_new_n11891__ = ~new_new_n11877__ & ~new_new_n11890__;
  assign new_new_n11892__ = ~ys__n18281 & ~new_new_n11891__;
  assign new_new_n11893__ = ys__n18632 & ~new_new_n11125__;
  assign new_new_n11894__ = ys__n78 & new_new_n11125__;
  assign ys__n18633 = new_new_n11893__ | new_new_n11894__;
  assign new_new_n11896__ = ys__n18281 & ys__n18633;
  assign new_new_n11897__ = ~new_new_n11892__ & ~new_new_n11896__;
  assign new_new_n11898__ = ~ys__n18278 & ~new_new_n11897__;
  assign new_new_n11899__ = ys__n18881 & ys__n18278;
  assign ys__n800 = new_new_n11898__ | new_new_n11899__;
  assign new_new_n11901__ = ys__n18981 & ys__n18287;
  assign new_new_n11902__ = ~ys__n18284 & new_new_n11901__;
  assign new_new_n11903__ = ys__n60 & ~ys__n4764;
  assign new_new_n11904__ = ys__n24664 & ys__n4764;
  assign ys__n18814 = new_new_n11903__ | new_new_n11904__;
  assign new_new_n11906__ = ~ys__n18071 & ys__n18814;
  assign new_new_n11907__ = ys__n18071 & ys__n18815;
  assign new_new_n11908__ = ~new_new_n11906__ & ~new_new_n11907__;
  assign new_new_n11909__ = ~new_new_n11122__ & ~new_new_n11908__;
  assign new_new_n11910__ = ys__n24664 & ~ys__n24675;
  assign new_new_n11911__ = ys__n24675 & ys__n24704;
  assign ys__n18729 = new_new_n11910__ | new_new_n11911__;
  assign new_new_n11913__ = new_new_n11122__ & ys__n18729;
  assign ys__n18730 = new_new_n11909__ | new_new_n11913__;
  assign new_new_n11915__ = ys__n18284 & ys__n18730;
  assign new_new_n11916__ = ~new_new_n11902__ & ~new_new_n11915__;
  assign new_new_n11917__ = ~ys__n18281 & ~new_new_n11916__;
  assign new_new_n11918__ = ys__n18630 & ~new_new_n11125__;
  assign new_new_n11919__ = ys__n70 & new_new_n11125__;
  assign ys__n18631 = new_new_n11918__ | new_new_n11919__;
  assign new_new_n11921__ = ys__n18281 & ys__n18631;
  assign new_new_n11922__ = ~new_new_n11917__ & ~new_new_n11921__;
  assign new_new_n11923__ = ~ys__n18278 & ~new_new_n11922__;
  assign new_new_n11924__ = ys__n18879 & ys__n18278;
  assign ys__n802 = new_new_n11923__ | new_new_n11924__;
  assign new_new_n11926__ = ys__n18980 & ys__n18287;
  assign new_new_n11927__ = ~ys__n18284 & new_new_n11926__;
  assign new_new_n11928__ = ys__n62 & ~ys__n4764;
  assign new_new_n11929__ = ys__n24663 & ys__n4764;
  assign ys__n18812 = new_new_n11928__ | new_new_n11929__;
  assign new_new_n11931__ = ~ys__n18071 & ys__n18812;
  assign new_new_n11932__ = ys__n18071 & ys__n18813;
  assign new_new_n11933__ = ~new_new_n11931__ & ~new_new_n11932__;
  assign new_new_n11934__ = ~new_new_n11122__ & ~new_new_n11933__;
  assign new_new_n11935__ = ys__n24663 & ~ys__n24675;
  assign new_new_n11936__ = ys__n24675 & ys__n24703;
  assign ys__n18726 = new_new_n11935__ | new_new_n11936__;
  assign new_new_n11938__ = new_new_n11122__ & ys__n18726;
  assign ys__n18727 = new_new_n11934__ | new_new_n11938__;
  assign new_new_n11940__ = ys__n18284 & ys__n18727;
  assign new_new_n11941__ = ~new_new_n11927__ & ~new_new_n11940__;
  assign new_new_n11942__ = ~ys__n18281 & ~new_new_n11941__;
  assign new_new_n11943__ = ys__n18628 & ~new_new_n11125__;
  assign new_new_n11944__ = ys__n72 & new_new_n11125__;
  assign ys__n18629 = new_new_n11943__ | new_new_n11944__;
  assign new_new_n11946__ = ys__n18281 & ys__n18629;
  assign new_new_n11947__ = ~new_new_n11942__ & ~new_new_n11946__;
  assign new_new_n11948__ = ~ys__n18278 & ~new_new_n11947__;
  assign new_new_n11949__ = ys__n18877 & ys__n18278;
  assign ys__n804 = new_new_n11948__ | new_new_n11949__;
  assign new_new_n11951__ = ys__n18977 & ys__n18287;
  assign new_new_n11952__ = ~ys__n18284 & new_new_n11951__;
  assign new_new_n11953__ = ys__n24657 & ~ys__n4764;
  assign new_new_n11954__ = ys__n24658 & ys__n4764;
  assign ys__n18806 = new_new_n11953__ | new_new_n11954__;
  assign new_new_n11956__ = ~ys__n18071 & ys__n18806;
  assign new_new_n11957__ = ys__n18071 & ys__n18807;
  assign new_new_n11958__ = ~new_new_n11956__ & ~new_new_n11957__;
  assign new_new_n11959__ = ~new_new_n11122__ & ~new_new_n11958__;
  assign new_new_n11960__ = ys__n24658 & ~ys__n24675;
  assign new_new_n11961__ = ys__n24675 & ys__n24700;
  assign ys__n18717 = new_new_n11960__ | new_new_n11961__;
  assign new_new_n11963__ = new_new_n11122__ & ys__n18717;
  assign ys__n18718 = new_new_n11959__ | new_new_n11963__;
  assign new_new_n11965__ = ys__n18284 & ys__n18718;
  assign new_new_n11966__ = ~new_new_n11952__ & ~new_new_n11965__;
  assign new_new_n11967__ = ~ys__n18281 & ~new_new_n11966__;
  assign new_new_n11968__ = ys__n18619 & ~new_new_n11125__;
  assign new_new_n11969__ = ys__n18620 & new_new_n11125__;
  assign ys__n18621 = new_new_n11968__ | new_new_n11969__;
  assign new_new_n11971__ = ys__n18281 & ys__n18621;
  assign new_new_n11972__ = ~new_new_n11967__ & ~new_new_n11971__;
  assign new_new_n11973__ = ~ys__n18278 & ~new_new_n11972__;
  assign new_new_n11974__ = ys__n18871 & ys__n18278;
  assign ys__n806 = new_new_n11973__ | new_new_n11974__;
  assign new_new_n11976__ = ys__n18986 & ys__n18287;
  assign new_new_n11977__ = ~ys__n18284 & new_new_n11976__;
  assign new_new_n11978__ = ys__n24670 & ~ys__n4764;
  assign new_new_n11979__ = ys__n24671 & ys__n4764;
  assign ys__n18824 = new_new_n11978__ | new_new_n11979__;
  assign new_new_n11981__ = ~ys__n18071 & ys__n18824;
  assign new_new_n11982__ = ys__n18071 & ys__n18825;
  assign new_new_n11983__ = ~new_new_n11981__ & ~new_new_n11982__;
  assign new_new_n11984__ = ~new_new_n11122__ & ~new_new_n11983__;
  assign new_new_n11985__ = ys__n24671 & ~ys__n24675;
  assign new_new_n11986__ = ys__n24675 & ys__n24709;
  assign ys__n18744 = new_new_n11985__ | new_new_n11986__;
  assign new_new_n11988__ = new_new_n11122__ & ys__n18744;
  assign ys__n18745 = new_new_n11984__ | new_new_n11988__;
  assign new_new_n11990__ = ys__n18284 & ys__n18745;
  assign new_new_n11991__ = ~new_new_n11977__ & ~new_new_n11990__;
  assign new_new_n11992__ = ~ys__n18281 & ~new_new_n11991__;
  assign new_new_n11993__ = ys__n18641 & ~new_new_n11125__;
  assign new_new_n11994__ = ys__n18642 & new_new_n11125__;
  assign ys__n18643 = new_new_n11993__ | new_new_n11994__;
  assign new_new_n11996__ = ys__n18281 & ys__n18643;
  assign new_new_n11997__ = ~new_new_n11992__ & ~new_new_n11996__;
  assign new_new_n11998__ = ~ys__n18278 & ~new_new_n11997__;
  assign new_new_n11999__ = ys__n18889 & ys__n18278;
  assign ys__n808 = new_new_n11998__ | new_new_n11999__;
  assign new_new_n12001__ = ys__n18985 & ys__n18287;
  assign new_new_n12002__ = ~ys__n18284 & new_new_n12001__;
  assign new_new_n12003__ = ys__n24668 & ~ys__n4764;
  assign new_new_n12004__ = ys__n24669 & ys__n4764;
  assign ys__n18822 = new_new_n12003__ | new_new_n12004__;
  assign new_new_n12006__ = ~ys__n18071 & ys__n18822;
  assign new_new_n12007__ = ys__n18071 & ys__n18823;
  assign new_new_n12008__ = ~new_new_n12006__ & ~new_new_n12007__;
  assign new_new_n12009__ = ~new_new_n11122__ & ~new_new_n12008__;
  assign new_new_n12010__ = ys__n24669 & ~ys__n24675;
  assign new_new_n12011__ = ys__n24675 & ys__n24708;
  assign ys__n18741 = new_new_n12010__ | new_new_n12011__;
  assign new_new_n12013__ = new_new_n11122__ & ys__n18741;
  assign ys__n18742 = new_new_n12009__ | new_new_n12013__;
  assign new_new_n12015__ = ys__n18284 & ys__n18742;
  assign new_new_n12016__ = ~new_new_n12002__ & ~new_new_n12015__;
  assign new_new_n12017__ = ~ys__n18281 & ~new_new_n12016__;
  assign new_new_n12018__ = ys__n18638 & ~new_new_n11125__;
  assign new_new_n12019__ = ys__n18639 & new_new_n11125__;
  assign ys__n18640 = new_new_n12018__ | new_new_n12019__;
  assign new_new_n12021__ = ys__n18281 & ys__n18640;
  assign new_new_n12022__ = ~new_new_n12017__ & ~new_new_n12021__;
  assign new_new_n12023__ = ~ys__n18278 & ~new_new_n12022__;
  assign new_new_n12024__ = ys__n18887 & ys__n18278;
  assign ys__n810 = new_new_n12023__ | new_new_n12024__;
  assign new_new_n12026__ = ys__n18987 & ys__n18287;
  assign new_new_n12027__ = ~ys__n18284 & new_new_n12026__;
  assign new_new_n12028__ = ys__n24672 & ~ys__n4764;
  assign new_new_n12029__ = ys__n24673 & ys__n4764;
  assign ys__n18826 = new_new_n12028__ | new_new_n12029__;
  assign new_new_n12031__ = ~ys__n18071 & ys__n18826;
  assign new_new_n12032__ = ys__n18071 & ys__n18827;
  assign new_new_n12033__ = ~new_new_n12031__ & ~new_new_n12032__;
  assign new_new_n12034__ = ~new_new_n11122__ & ~new_new_n12033__;
  assign new_new_n12035__ = ys__n24673 & ~ys__n24675;
  assign new_new_n12036__ = ys__n24675 & ys__n24710;
  assign ys__n18747 = new_new_n12035__ | new_new_n12036__;
  assign new_new_n12038__ = new_new_n11122__ & ys__n18747;
  assign ys__n18748 = new_new_n12034__ | new_new_n12038__;
  assign new_new_n12040__ = ys__n18284 & ys__n18748;
  assign new_new_n12041__ = ~new_new_n12027__ & ~new_new_n12040__;
  assign new_new_n12042__ = ~ys__n18281 & ~new_new_n12041__;
  assign new_new_n12043__ = ys__n18644 & ~new_new_n11125__;
  assign new_new_n12044__ = ys__n18645 & new_new_n11125__;
  assign ys__n18646 = new_new_n12043__ | new_new_n12044__;
  assign new_new_n12046__ = ys__n18281 & ys__n18646;
  assign new_new_n12047__ = ~new_new_n12042__ & ~new_new_n12046__;
  assign new_new_n12048__ = ~ys__n18278 & ~new_new_n12047__;
  assign new_new_n12049__ = ys__n18891 & ys__n18278;
  assign ys__n812 = new_new_n12048__ | new_new_n12049__;
  assign new_new_n12051__ = ys__n20273 & ys__n738;
  assign ys__n814 = ~new_new_n10886__ & new_new_n12051__;
  assign new_new_n12053__ = ys__n29896 & ~new_new_n10603__;
  assign new_new_n12054__ = ~new_new_n10601__ & new_new_n12053__;
  assign new_new_n12055__ = ~ys__n23764 & new_new_n12054__;
  assign new_new_n12056__ = ys__n29912 & ~new_new_n10603__;
  assign new_new_n12057__ = ~new_new_n10601__ & new_new_n12056__;
  assign new_new_n12058__ = ~ys__n22466 & new_new_n12057__;
  assign new_new_n12059__ = ys__n22466 & new_new_n12054__;
  assign new_new_n12060__ = ~new_new_n12058__ & ~new_new_n12059__;
  assign new_new_n12061__ = ys__n23764 & ~new_new_n12060__;
  assign new_new_n12062__ = ~new_new_n12055__ & ~new_new_n12061__;
  assign new_new_n12063__ = ~new_new_n10859__ & ~new_new_n12062__;
  assign new_new_n12064__ = ys__n23764 & ~new_new_n10864__;
  assign new_new_n12065__ = ~new_new_n12063__ & ~new_new_n12064__;
  assign ys__n25435 = ~new_new_n10865__ & ~new_new_n12065__;
  assign new_new_n12067__ = ~ys__n19256 & ys__n25435;
  assign new_new_n12068__ = ys__n634 & ys__n19256;
  assign new_new_n12069__ = ~new_new_n12067__ & ~new_new_n12068__;
  assign new_new_n12070__ = ys__n874 & ~new_new_n12069__;
  assign ys__n862 = ys__n2 | ~new_new_n12070__;
  assign new_new_n12072__ = ys__n37703 & ~new_new_n11121__;
  assign new_new_n12073__ = ~ys__n37674 & ys__n37675;
  assign new_new_n12074__ = ys__n37674 & ~ys__n37675;
  assign new_new_n12075__ = ~new_new_n12073__ & ~new_new_n12074__;
  assign new_new_n12076__ = ~ys__n18393 & ~new_new_n12075__;
  assign new_new_n12077__ = ys__n18393 & new_new_n11149__;
  assign new_new_n12078__ = ~new_new_n11147__ & new_new_n12077__;
  assign new_new_n12079__ = ~new_new_n11147__ & ~new_new_n12078__;
  assign new_new_n12080__ = new_new_n11076__ & ~new_new_n11141__;
  assign new_new_n12081__ = ~new_new_n12079__ & new_new_n12080__;
  assign new_new_n12082__ = ys__n18393 & ys__n19203;
  assign new_new_n12083__ = ~ys__n19215 & new_new_n12082__;
  assign new_new_n12084__ = new_new_n11081__ & new_new_n12083__;
  assign new_new_n12085__ = new_new_n11143__ & new_new_n12084__;
  assign new_new_n12086__ = ~ys__n18393 & ~new_new_n11072__;
  assign new_new_n12087__ = ~new_new_n12085__ & ~new_new_n12086__;
  assign new_new_n12088__ = ~new_new_n12081__ & new_new_n12087__;
  assign new_new_n12089__ = ~new_new_n11076__ & ~new_new_n11081__;
  assign new_new_n12090__ = new_new_n11072__ & new_new_n12089__;
  assign ys__n27605 = ~new_new_n12088__ & ~new_new_n12090__;
  assign new_new_n12092__ = ys__n18393 & ys__n27605;
  assign new_new_n12093__ = ~new_new_n12076__ & ~new_new_n12092__;
  assign new_new_n12094__ = ys__n33300 & ys__n37692;
  assign new_new_n12095__ = new_new_n12093__ & ~new_new_n12094__;
  assign new_new_n12096__ = ~ys__n18317 & ~new_new_n12095__;
  assign new_new_n12097__ = ~ys__n33300 & ~ys__n37694;
  assign new_new_n12098__ = ~ys__n37696 & new_new_n12093__;
  assign new_new_n12099__ = ~new_new_n12097__ & ~new_new_n12098__;
  assign new_new_n12100__ = ys__n18271 & ys__n37692;
  assign new_new_n12101__ = ~new_new_n12099__ & ~new_new_n12100__;
  assign new_new_n12102__ = ys__n18317 & ~new_new_n12101__;
  assign new_new_n12103__ = ~new_new_n12096__ & ~new_new_n12102__;
  assign new_new_n12104__ = ~ys__n33309 & ~ys__n33311;
  assign new_new_n12105__ = ~ys__n33313 & new_new_n12104__;
  assign new_new_n12106__ = ~new_new_n12103__ & new_new_n12105__;
  assign ys__n863 = new_new_n12072__ & ~new_new_n12106__;
  assign new_new_n12108__ = ~new_new_n12072__ & new_new_n12106__;
  assign ys__n865 = ys__n863 | new_new_n12108__;
  assign ys__n866 = ~ys__n2 | new_new_n12070__;
  assign new_new_n12111__ = ys__n29895 & ~new_new_n10603__;
  assign new_new_n12112__ = ~new_new_n10601__ & new_new_n12111__;
  assign new_new_n12113__ = ~ys__n23764 & new_new_n12112__;
  assign new_new_n12114__ = ys__n29911 & ~new_new_n10603__;
  assign new_new_n12115__ = ~new_new_n10601__ & new_new_n12114__;
  assign new_new_n12116__ = ~ys__n22466 & new_new_n12115__;
  assign new_new_n12117__ = ys__n22466 & new_new_n12112__;
  assign new_new_n12118__ = ~new_new_n12116__ & ~new_new_n12117__;
  assign new_new_n12119__ = ys__n23764 & ~new_new_n12118__;
  assign new_new_n12120__ = ~new_new_n12113__ & ~new_new_n12119__;
  assign new_new_n12121__ = ~new_new_n10859__ & ~new_new_n12120__;
  assign new_new_n12122__ = ~new_new_n12064__ & ~new_new_n12121__;
  assign ys__n25434 = ~new_new_n10865__ & ~new_new_n12122__;
  assign new_new_n12124__ = ~ys__n19256 & ys__n25434;
  assign new_new_n12125__ = ys__n636 & ys__n19256;
  assign new_new_n12126__ = ~new_new_n12124__ & ~new_new_n12125__;
  assign new_new_n12127__ = ys__n874 & ~new_new_n12126__;
  assign ys__n868 = ys__n866 | new_new_n12127__;
  assign new_new_n12129__ = ys__n29894 & ~new_new_n10603__;
  assign new_new_n12130__ = ~new_new_n10601__ & new_new_n12129__;
  assign new_new_n12131__ = ~ys__n23764 & new_new_n12130__;
  assign new_new_n12132__ = ys__n29910 & ~new_new_n10603__;
  assign new_new_n12133__ = ~new_new_n10601__ & new_new_n12132__;
  assign new_new_n12134__ = ~ys__n22466 & new_new_n12133__;
  assign new_new_n12135__ = ys__n22466 & new_new_n12130__;
  assign new_new_n12136__ = ~new_new_n12134__ & ~new_new_n12135__;
  assign new_new_n12137__ = ys__n23764 & ~new_new_n12136__;
  assign new_new_n12138__ = ~new_new_n12131__ & ~new_new_n12137__;
  assign ys__n25433 = new_new_n10866__ & ~new_new_n12138__;
  assign new_new_n12140__ = ~ys__n19256 & ys__n25433;
  assign new_new_n12141__ = ys__n638 & ys__n19256;
  assign new_new_n12142__ = ~new_new_n12140__ & ~new_new_n12141__;
  assign new_new_n12143__ = ys__n874 & ~new_new_n12142__;
  assign new_new_n12144__ = new_new_n12127__ & new_new_n12143__;
  assign ys__n870 = ys__n862 | ~new_new_n12144__;
  assign new_new_n12146__ = ys__n18120 & ~ys__n740;
  assign ys__n871 = ~ys__n874 | new_new_n12146__;
  assign new_new_n12148__ = ~ys__n140 & ~ys__n214;
  assign new_new_n12149__ = ys__n216 & ~ys__n218;
  assign new_new_n12150__ = new_new_n12148__ & new_new_n12149__;
  assign new_new_n12151__ = ~ys__n216 & ys__n218;
  assign new_new_n12152__ = new_new_n12148__ & new_new_n12151__;
  assign new_new_n12153__ = ~new_new_n12150__ & ~new_new_n12152__;
  assign new_new_n12154__ = ~ys__n216 & ~ys__n218;
  assign new_new_n12155__ = ~ys__n140 & ys__n214;
  assign new_new_n12156__ = new_new_n12154__ & new_new_n12155__;
  assign new_new_n12157__ = new_new_n12153__ & ~new_new_n12156__;
  assign ys__n872 = ys__n871 | new_new_n12157__;
  assign new_new_n12159__ = ~ys__n140 & ~ys__n210;
  assign new_new_n12160__ = ys__n66 & ~ys__n212;
  assign new_new_n12161__ = new_new_n12159__ & new_new_n12160__;
  assign new_new_n12162__ = ~ys__n66 & ys__n212;
  assign new_new_n12163__ = new_new_n12159__ & new_new_n12162__;
  assign new_new_n12164__ = ~new_new_n12161__ & ~new_new_n12163__;
  assign new_new_n12165__ = ~ys__n66 & ~ys__n212;
  assign new_new_n12166__ = ~ys__n140 & ys__n210;
  assign new_new_n12167__ = new_new_n12165__ & new_new_n12166__;
  assign new_new_n12168__ = new_new_n12164__ & ~new_new_n12167__;
  assign ys__n873 = ys__n871 | new_new_n12168__;
  assign new_new_n12170__ = ~ys__n140 & ~ys__n298;
  assign new_new_n12171__ = ~ys__n300 & ys__n302;
  assign new_new_n12172__ = new_new_n12170__ & new_new_n12171__;
  assign new_new_n12173__ = ~ys__n140 & ~ys__n302;
  assign new_new_n12174__ = ~ys__n298 & ys__n300;
  assign new_new_n12175__ = new_new_n12173__ & new_new_n12174__;
  assign new_new_n12176__ = ys__n298 & ~ys__n300;
  assign new_new_n12177__ = new_new_n12173__ & new_new_n12176__;
  assign new_new_n12178__ = ~new_new_n12175__ & ~new_new_n12177__;
  assign new_new_n12179__ = ~new_new_n12172__ & new_new_n12178__;
  assign ys__n876 = ys__n874 & ~new_new_n12179__;
  assign new_new_n12181__ = ~ys__n140 & ~ys__n580;
  assign new_new_n12182__ = ~ys__n582 & ys__n584;
  assign new_new_n12183__ = new_new_n12181__ & new_new_n12182__;
  assign new_new_n12184__ = ~ys__n140 & ~ys__n584;
  assign new_new_n12185__ = ~ys__n580 & ys__n582;
  assign new_new_n12186__ = new_new_n12184__ & new_new_n12185__;
  assign new_new_n12187__ = ys__n580 & ~ys__n582;
  assign new_new_n12188__ = new_new_n12184__ & new_new_n12187__;
  assign new_new_n12189__ = ~new_new_n12186__ & ~new_new_n12188__;
  assign new_new_n12190__ = ~new_new_n12183__ & new_new_n12189__;
  assign ys__n878 = ys__n874 & ~new_new_n12190__;
  assign new_new_n12192__ = ~ys__n138 & ~ys__n140;
  assign new_new_n12193__ = ~ys__n120 & ys__n142;
  assign new_new_n12194__ = new_new_n12192__ & new_new_n12193__;
  assign new_new_n12195__ = ys__n120 & ~ys__n142;
  assign new_new_n12196__ = new_new_n12192__ & new_new_n12195__;
  assign new_new_n12197__ = ~new_new_n12194__ & ~new_new_n12196__;
  assign new_new_n12198__ = ~ys__n120 & ~ys__n142;
  assign new_new_n12199__ = ys__n138 & ~ys__n140;
  assign new_new_n12200__ = new_new_n12198__ & new_new_n12199__;
  assign new_new_n12201__ = new_new_n12197__ & ~new_new_n12200__;
  assign ys__n879 = ys__n871 | new_new_n12201__;
  assign new_new_n12203__ = ~ys__n140 & ~ys__n392;
  assign new_new_n12204__ = ~ys__n394 & ys__n396;
  assign new_new_n12205__ = new_new_n12203__ & new_new_n12204__;
  assign new_new_n12206__ = ~ys__n140 & ~ys__n396;
  assign new_new_n12207__ = ~ys__n392 & ys__n394;
  assign new_new_n12208__ = new_new_n12206__ & new_new_n12207__;
  assign new_new_n12209__ = ys__n392 & ~ys__n394;
  assign new_new_n12210__ = new_new_n12206__ & new_new_n12209__;
  assign new_new_n12211__ = ~new_new_n12208__ & ~new_new_n12210__;
  assign new_new_n12212__ = ~new_new_n12205__ & new_new_n12211__;
  assign ys__n881 = ys__n874 & ~new_new_n12212__;
  assign new_new_n12214__ = ~ys__n2779 & ~ys__n30816;
  assign new_new_n12215__ = ys__n30819 & new_new_n12214__;
  assign new_new_n12216__ = ys__n30815 & ys__n30816;
  assign new_new_n12217__ = ~new_new_n12215__ & ~new_new_n12216__;
  assign new_new_n12218__ = ~ys__n562 & ~new_new_n12217__;
  assign new_new_n12219__ = ys__n562 & new_new_n12217__;
  assign ys__n888 = new_new_n12218__ | new_new_n12219__;
  assign new_new_n12221__ = ~ys__n846 & ys__n874;
  assign new_new_n12222__ = ~ys__n889 & new_new_n12221__;
  assign new_new_n12223__ = ~ys__n4184 & ~ys__n4185;
  assign new_new_n12224__ = new_new_n11047__ & new_new_n12223__;
  assign new_new_n12225__ = ~ys__n4176 & ~ys__n4627;
  assign new_new_n12226__ = ~ys__n4177 & ~ys__n4698;
  assign new_new_n12227__ = new_new_n12225__ & new_new_n12226__;
  assign new_new_n12228__ = new_new_n12224__ & new_new_n12227__;
  assign ys__n900 = ~new_new_n12222__ | ~new_new_n12228__;
  assign ys__n902 = ~ys__n874 | ~new_new_n12103__;
  assign ys__n904 = ys__n30223 | ~ys__n740;
  assign new_new_n12232__ = ys__n38305 & ~ys__n738;
  assign ys__n911 = ~ys__n4566 & new_new_n12232__;
  assign new_new_n12234__ = ys__n30820 & new_new_n12214__;
  assign new_new_n12235__ = ys__n30816 & ys__n30818;
  assign new_new_n12236__ = ~new_new_n12234__ & ~new_new_n12235__;
  assign new_new_n12237__ = ~ys__n398 & ~new_new_n12236__;
  assign new_new_n12238__ = ys__n398 & new_new_n12236__;
  assign ys__n920 = new_new_n12237__ | new_new_n12238__;
  assign new_new_n12240__ = ys__n172 & ys__n338;
  assign new_new_n12241__ = ~ys__n172 & ~ys__n338;
  assign new_new_n12242__ = ~ys__n172 & ys__n338;
  assign new_new_n12243__ = ~new_new_n12241__ & ~new_new_n12242__;
  assign new_new_n12244__ = ~new_new_n12240__ & new_new_n12243__;
  assign new_new_n12245__ = ys__n22 & ~ys__n316;
  assign new_new_n12246__ = ~ys__n22 & ~ys__n316;
  assign new_new_n12247__ = ~new_new_n12245__ & ~new_new_n12246__;
  assign new_new_n12248__ = ~ys__n22 & ys__n316;
  assign new_new_n12249__ = new_new_n12247__ & ~new_new_n12248__;
  assign new_new_n12250__ = ys__n172 & ~ys__n338;
  assign new_new_n12251__ = ~new_new_n12249__ & new_new_n12250__;
  assign new_new_n12252__ = new_new_n12244__ & ~new_new_n12251__;
  assign new_new_n12253__ = ~ys__n35047 & ys__n46240;
  assign new_new_n12254__ = ~ys__n46230 & ys__n46239;
  assign new_new_n12255__ = ys__n46230 & ~ys__n46239;
  assign new_new_n12256__ = ~new_new_n12254__ & ~new_new_n12255__;
  assign new_new_n12257__ = ys__n46238 & ~new_new_n12256__;
  assign ys__n18210 = new_new_n12253__ | new_new_n12257__;
  assign new_new_n12259__ = ~ys__n44 & ys__n6115;
  assign new_new_n12260__ = ~ys__n44 & ~new_new_n12259__;
  assign new_new_n12261__ = ~ys__n18208 & new_new_n12260__;
  assign new_new_n12262__ = ys__n18210 & new_new_n12261__;
  assign new_new_n12263__ = ~ys__n6120 & ~ys__n6121;
  assign new_new_n12264__ = ~ys__n6123 & ~ys__n6124;
  assign new_new_n12265__ = new_new_n12263__ & new_new_n12264__;
  assign new_new_n12266__ = ~ys__n6118 & ~ys__n6119;
  assign new_new_n12267__ = ys__n46 & ~ys__n340;
  assign new_new_n12268__ = ys__n18317 & new_new_n12267__;
  assign new_new_n12269__ = new_new_n12266__ & new_new_n12268__;
  assign new_new_n12270__ = new_new_n12265__ & new_new_n12269__;
  assign new_new_n12271__ = ys__n40 & ys__n42;
  assign new_new_n12272__ = ~ys__n6133 & ~ys__n6134;
  assign new_new_n12273__ = new_new_n12271__ & new_new_n12272__;
  assign new_new_n12274__ = ~ys__n6126 & ~ys__n6127;
  assign new_new_n12275__ = ~ys__n6129 & ~ys__n6130;
  assign new_new_n12276__ = new_new_n12274__ & new_new_n12275__;
  assign new_new_n12277__ = new_new_n12273__ & new_new_n12276__;
  assign new_new_n12278__ = ys__n32 & ys__n34;
  assign new_new_n12279__ = ys__n36 & ys__n38;
  assign new_new_n12280__ = new_new_n12278__ & new_new_n12279__;
  assign new_new_n12281__ = ys__n24 & ys__n26;
  assign new_new_n12282__ = ys__n28 & ys__n30;
  assign new_new_n12283__ = new_new_n12281__ & new_new_n12282__;
  assign new_new_n12284__ = new_new_n12280__ & new_new_n12283__;
  assign new_new_n12285__ = new_new_n12277__ & new_new_n12284__;
  assign new_new_n12286__ = new_new_n12270__ & new_new_n12285__;
  assign new_new_n12287__ = new_new_n12262__ & new_new_n12286__;
  assign ys__n923 = new_new_n12252__ & new_new_n12287__;
  assign new_new_n12289__ = ys__n38307 & ~ys__n738;
  assign ys__n927 = ~ys__n4566 & new_new_n12289__;
  assign new_new_n12291__ = ys__n754 & ys__n756;
  assign new_new_n12292__ = ~ys__n738 & new_new_n12291__;
  assign new_new_n12293__ = ys__n478 & new_new_n12292__;
  assign new_new_n12294__ = ys__n482 & new_new_n12293__;
  assign ys__n929 = ~ys__n480 & new_new_n12294__;
  assign ys__n930 = ~ys__n738 & ys__n478;
  assign new_new_n12297__ = ys__n38220 & ~ys__n4566;
  assign new_new_n12298__ = ~ys__n935 & ~new_new_n12297__;
  assign ys__n932 = ~ys__n738 & ~new_new_n12298__;
  assign new_new_n12300__ = ys__n38221 & ~ys__n738;
  assign ys__n934 = ~ys__n4566 & new_new_n12300__;
  assign ys__n936 = ys__n935 & ~ys__n738;
  assign new_new_n12303__ = ~ys__n38407 & ~ys__n38408;
  assign new_new_n12304__ = ~ys__n226 & new_new_n12303__;
  assign new_new_n12305__ = ys__n478 & new_new_n12304__;
  assign new_new_n12306__ = ys__n226 & ys__n478;
  assign new_new_n12307__ = ~ys__n226 & ~new_new_n12303__;
  assign new_new_n12308__ = ys__n478 & new_new_n12307__;
  assign new_new_n12309__ = ~new_new_n12306__ & ~new_new_n12308__;
  assign new_new_n12310__ = ~new_new_n12305__ & new_new_n12309__;
  assign ys__n942 = ~ys__n738 & ~new_new_n12310__;
  assign new_new_n12312__ = ys__n326 & ~ys__n332;
  assign new_new_n12313__ = ~ys__n328 & ~ys__n330;
  assign new_new_n12314__ = ~ys__n336 & new_new_n12313__;
  assign new_new_n12315__ = new_new_n12312__ & new_new_n12314__;
  assign new_new_n12316__ = ys__n328 & ~ys__n330;
  assign new_new_n12317__ = ~ys__n336 & new_new_n12312__;
  assign new_new_n12318__ = new_new_n12316__ & new_new_n12317__;
  assign new_new_n12319__ = ~new_new_n12315__ & ~new_new_n12318__;
  assign new_new_n12320__ = ~ys__n328 & ys__n330;
  assign new_new_n12321__ = new_new_n12317__ & new_new_n12320__;
  assign new_new_n12322__ = ys__n328 & ys__n330;
  assign new_new_n12323__ = new_new_n12317__ & new_new_n12322__;
  assign new_new_n12324__ = ~new_new_n12321__ & ~new_new_n12323__;
  assign new_new_n12325__ = new_new_n12319__ & new_new_n12324__;
  assign new_new_n12326__ = ys__n326 & ys__n332;
  assign new_new_n12327__ = ys__n336 & new_new_n12326__;
  assign new_new_n12328__ = new_new_n12322__ & new_new_n12327__;
  assign new_new_n12329__ = new_new_n12325__ & ~new_new_n12328__;
  assign ys__n944 = ys__n602 & ~new_new_n12329__;
  assign new_new_n12331__ = ~ys__n4176 & new_new_n10613__;
  assign new_new_n12332__ = new_new_n10609__ & new_new_n12331__;
  assign new_new_n12333__ = new_new_n10608__ & new_new_n12332__;
  assign ys__n30832 = ys__n4698 | ~new_new_n12333__;
  assign ys__n948 = ~ys__n4566 & ~ys__n30832;
  assign new_new_n12336__ = ~ys__n160 & ys__n344;
  assign new_new_n12337__ = ys__n342 & ys__n350;
  assign new_new_n12338__ = new_new_n12336__ & new_new_n12337__;
  assign new_new_n12339__ = ys__n348 & ~ys__n2924;
  assign new_new_n12340__ = ~ys__n162 & ~ys__n346;
  assign new_new_n12341__ = new_new_n12339__ & new_new_n12340__;
  assign new_new_n12342__ = ys__n352 & new_new_n12341__;
  assign new_new_n12343__ = new_new_n12338__ & new_new_n12342__;
  assign new_new_n12344__ = ~ys__n342 & ys__n350;
  assign new_new_n12345__ = new_new_n12336__ & new_new_n12344__;
  assign new_new_n12346__ = ys__n352 & new_new_n12345__;
  assign new_new_n12347__ = new_new_n12341__ & new_new_n12346__;
  assign new_new_n12348__ = ys__n162 & ys__n346;
  assign new_new_n12349__ = new_new_n12339__ & new_new_n12348__;
  assign new_new_n12350__ = new_new_n12346__ & new_new_n12349__;
  assign new_new_n12351__ = ~new_new_n12347__ & ~new_new_n12350__;
  assign new_new_n12352__ = ~new_new_n12343__ & new_new_n12351__;
  assign ys__n949 = ys__n948 & ~new_new_n12352__;
  assign new_new_n12354__ = ~new_new_n12241__ & ~new_new_n12250__;
  assign new_new_n12355__ = ~new_new_n12242__ & new_new_n12354__;
  assign new_new_n12356__ = ys__n22 & ys__n316;
  assign new_new_n12357__ = ~new_new_n12246__ & ~new_new_n12248__;
  assign new_new_n12358__ = ~new_new_n12356__ & new_new_n12357__;
  assign new_new_n12359__ = new_new_n12240__ & ~new_new_n12358__;
  assign new_new_n12360__ = new_new_n12355__ & ~new_new_n12359__;
  assign new_new_n12361__ = ys__n46 & ys__n340;
  assign new_new_n12362__ = ys__n18317 & new_new_n12361__;
  assign new_new_n12363__ = new_new_n12266__ & new_new_n12362__;
  assign new_new_n12364__ = new_new_n12265__ & new_new_n12363__;
  assign new_new_n12365__ = new_new_n12285__ & new_new_n12364__;
  assign new_new_n12366__ = new_new_n12262__ & new_new_n12365__;
  assign ys__n970 = new_new_n12360__ & new_new_n12366__;
  assign new_new_n12368__ = ~new_new_n12245__ & ~new_new_n12248__;
  assign new_new_n12369__ = ~new_new_n12356__ & new_new_n12368__;
  assign new_new_n12370__ = new_new_n12240__ & ~new_new_n12369__;
  assign new_new_n12371__ = new_new_n12355__ & ~new_new_n12370__;
  assign ys__n972 = new_new_n12366__ & new_new_n12371__;
  assign new_new_n12373__ = new_new_n12247__ & ~new_new_n12356__;
  assign new_new_n12374__ = new_new_n12240__ & ~new_new_n12373__;
  assign new_new_n12375__ = new_new_n12355__ & ~new_new_n12374__;
  assign ys__n974 = new_new_n12366__ & new_new_n12375__;
  assign new_new_n12377__ = ~new_new_n12242__ & ~new_new_n12250__;
  assign new_new_n12378__ = ~new_new_n12240__ & new_new_n12377__;
  assign new_new_n12379__ = new_new_n12241__ & ~new_new_n12369__;
  assign new_new_n12380__ = new_new_n12378__ & ~new_new_n12379__;
  assign ys__n976 = new_new_n12366__ & new_new_n12380__;
  assign new_new_n12382__ = new_new_n12241__ & ~new_new_n12358__;
  assign new_new_n12383__ = new_new_n12378__ & ~new_new_n12382__;
  assign ys__n978 = new_new_n12366__ & new_new_n12383__;
  assign new_new_n12385__ = new_new_n12240__ & ~new_new_n12249__;
  assign new_new_n12386__ = new_new_n12355__ & ~new_new_n12385__;
  assign ys__n980 = new_new_n12366__ & new_new_n12386__;
  assign new_new_n12388__ = new_new_n12250__ & ~new_new_n12369__;
  assign new_new_n12389__ = new_new_n12244__ & ~new_new_n12388__;
  assign ys__n982 = new_new_n12366__ & new_new_n12389__;
  assign new_new_n12391__ = ~ys__n46 & ys__n340;
  assign new_new_n12392__ = ys__n18317 & new_new_n12391__;
  assign new_new_n12393__ = new_new_n12266__ & new_new_n12392__;
  assign new_new_n12394__ = new_new_n12265__ & new_new_n12393__;
  assign new_new_n12395__ = new_new_n12285__ & new_new_n12394__;
  assign new_new_n12396__ = new_new_n12262__ & new_new_n12395__;
  assign new_new_n12397__ = new_new_n12241__ & new_new_n12249__;
  assign ys__n989 = new_new_n12396__ & new_new_n12397__;
  assign ys__n991 = new_new_n12252__ & new_new_n12366__;
  assign new_new_n12400__ = new_new_n12250__ & ~new_new_n12373__;
  assign new_new_n12401__ = new_new_n12244__ & ~new_new_n12400__;
  assign ys__n993 = new_new_n12366__ & new_new_n12401__;
  assign new_new_n12403__ = new_new_n12241__ & ~new_new_n12249__;
  assign new_new_n12404__ = new_new_n12378__ & ~new_new_n12403__;
  assign ys__n995 = new_new_n12366__ & new_new_n12404__;
  assign new_new_n12406__ = new_new_n12242__ & ~new_new_n12358__;
  assign new_new_n12407__ = ~new_new_n12240__ & new_new_n12354__;
  assign new_new_n12408__ = ~new_new_n12406__ & new_new_n12407__;
  assign ys__n999 = new_new_n12366__ & new_new_n12408__;
  assign new_new_n12410__ = new_new_n12242__ & ~new_new_n12369__;
  assign new_new_n12411__ = new_new_n12407__ & ~new_new_n12410__;
  assign ys__n1001 = new_new_n12366__ & new_new_n12411__;
  assign new_new_n12413__ = new_new_n12242__ & ~new_new_n12249__;
  assign new_new_n12414__ = new_new_n12407__ & ~new_new_n12413__;
  assign ys__n1004 = new_new_n12366__ & new_new_n12414__;
  assign new_new_n12416__ = new_new_n12242__ & ~new_new_n12373__;
  assign new_new_n12417__ = new_new_n12407__ & ~new_new_n12416__;
  assign ys__n1007 = new_new_n12366__ & new_new_n12417__;
  assign new_new_n12419__ = new_new_n12241__ & ~new_new_n12373__;
  assign new_new_n12420__ = new_new_n12378__ & ~new_new_n12419__;
  assign ys__n1009 = new_new_n12366__ & new_new_n12420__;
  assign new_new_n12422__ = new_new_n12250__ & ~new_new_n12358__;
  assign new_new_n12423__ = new_new_n12244__ & ~new_new_n12422__;
  assign ys__n1013 = new_new_n12366__ & new_new_n12423__;
  assign new_new_n12425__ = ys__n1020 & new_new_n12156__;
  assign new_new_n12426__ = ~ys__n30223 & new_new_n12152__;
  assign ys__n16191 = new_new_n12425__ | new_new_n12426__;
  assign new_new_n12428__ = ys__n740 & new_new_n12150__;
  assign new_new_n12429__ = ~ys__n1020 & ~ys__n740;
  assign new_new_n12430__ = ~ys__n1020 & new_new_n12156__;
  assign new_new_n12431__ = ~new_new_n12429__ & new_new_n12430__;
  assign new_new_n12432__ = ~new_new_n12428__ & ~new_new_n12431__;
  assign ys__n1028 = ~ys__n16191 & new_new_n12432__;
  assign new_new_n12434__ = ~ys__n18121 & ~ys__n18122;
  assign ys__n1030 = ys__n18124 & ~new_new_n12434__;
  assign ys__n1031 = ys__n1029 | ys__n1030;
  assign ys__n1032 = ~ys__n874 | ys__n1029;
  assign ys__n1037 = ~ys__n874 | ys__n1036;
  assign new_new_n12439__ = ~ys__n1029 & ~ys__n1038;
  assign ys__n1040 = ys__n1037 | ~new_new_n12439__;
  assign ys__n3021 = ys__n874 & ys__n1048;
  assign ys__n1043 = ys__n140 | ~ys__n3021;
  assign new_new_n12443__ = new_new_n12242__ & new_new_n12369__;
  assign ys__n1046 = new_new_n12396__ & new_new_n12443__;
  assign ys__n1047 = ys__n140 | ~ys__n874;
  assign ys__n1049 = ys__n1048 | ys__n1047;
  assign new_new_n12447__ = ys__n1020 & new_new_n12167__;
  assign new_new_n12448__ = ~ys__n30223 & new_new_n12163__;
  assign ys__n16427 = new_new_n12447__ | new_new_n12448__;
  assign new_new_n12450__ = ys__n740 & new_new_n12161__;
  assign new_new_n12451__ = ~ys__n1020 & new_new_n12167__;
  assign new_new_n12452__ = ~new_new_n12429__ & new_new_n12451__;
  assign new_new_n12453__ = ~new_new_n12450__ & ~new_new_n12452__;
  assign ys__n1060 = ~ys__n16427 & new_new_n12453__;
  assign new_new_n12455__ = ys__n1020 & new_new_n12200__;
  assign new_new_n12456__ = ~ys__n30223 & new_new_n12196__;
  assign ys__n16721 = new_new_n12455__ | new_new_n12456__;
  assign new_new_n12458__ = ys__n740 & new_new_n12194__;
  assign new_new_n12459__ = ~ys__n1020 & new_new_n12200__;
  assign new_new_n12460__ = ~new_new_n12429__ & new_new_n12459__;
  assign new_new_n12461__ = ~new_new_n12458__ & ~new_new_n12460__;
  assign ys__n1071 = ~ys__n16721 & new_new_n12461__;
  assign ys__n1074 = ys__n1072 | ys__n1073;
  assign ys__n1075 = ~ys__n874 | ys__n1072;
  assign ys__n1077 = ~ys__n874 | ys__n1076;
  assign ys__n1079 = ys__n1072 | ys__n1078;
  assign ys__n1080 = ys__n1077 | ys__n1079;
  assign ys__n1448 = ys__n874 & ys__n1084;
  assign ys__n1083 = ys__n140 | ~ys__n1448;
  assign ys__n1085 = ys__n1084 | ys__n1047;
  assign ys__n1088 = ys__n1106 & ~ys__n33479;
  assign new_new_n12472__ = ~ys__n33481 & ys__n33495;
  assign new_new_n12473__ = ys__n1088 & new_new_n12472__;
  assign ys__n1087 = ys__n874 & new_new_n12473__;
  assign new_new_n12475__ = ~ys__n1098 & ~ys__n1107;
  assign new_new_n12476__ = ~ys__n1129 & new_new_n12475__;
  assign new_new_n12477__ = ~ys__n24463 & new_new_n12476__;
  assign ys__n1089 = ys__n24519 & ~new_new_n12477__;
  assign ys__n1090 = ys__n1088 | ys__n1089;
  assign ys__n1091 = ~ys__n874 | ys__n1088;
  assign ys__n1141 = ~ys__n874 | ys__n1094;
  assign ys__n1095 = ~ys__n1106 | ys__n1141;
  assign new_new_n12483__ = ~ys__n1094 & ~ys__n1106;
  assign new_new_n12484__ = ys__n874 & ~ys__n1098;
  assign new_new_n12485__ = ~ys__n1099 & ys__n1107;
  assign new_new_n12486__ = new_new_n12484__ & new_new_n12485__;
  assign ys__n1103 = ~new_new_n12483__ | ~new_new_n12486__;
  assign new_new_n12488__ = ~ys__n1109 & ~ys__n1110;
  assign new_new_n12489__ = ys__n1129 & new_new_n12488__;
  assign new_new_n12490__ = ~ys__n1099 & ~ys__n1107;
  assign new_new_n12491__ = new_new_n12484__ & new_new_n12490__;
  assign new_new_n12492__ = new_new_n12483__ & new_new_n12491__;
  assign ys__n1115 = ~new_new_n12489__ | ~new_new_n12492__;
  assign new_new_n12494__ = ~ys__n1098 & ~ys__n1106;
  assign new_new_n12495__ = ~ys__n1141 & new_new_n12494__;
  assign new_new_n12496__ = ~ys__n1107 & ~ys__n1109;
  assign new_new_n12497__ = ~ys__n1110 & ~ys__n1129;
  assign new_new_n12498__ = new_new_n12496__ & new_new_n12497__;
  assign new_new_n12499__ = new_new_n12495__ & new_new_n12498__;
  assign new_new_n12500__ = ~ys__n1119 & ~ys__n1120;
  assign new_new_n12501__ = ~ys__n1099 & ~ys__n1116;
  assign new_new_n12502__ = ~ys__n1117 & new_new_n12501__;
  assign new_new_n12503__ = new_new_n12500__ & new_new_n12502__;
  assign ys__n1125 = ~new_new_n12499__ | ~new_new_n12503__;
  assign new_new_n12505__ = ~ys__n1119 & new_new_n12501__;
  assign ys__n1128 = ~new_new_n12499__ | ~new_new_n12505__;
  assign new_new_n12507__ = ~ys__n1099 & ~ys__n1119;
  assign ys__n1135 = ~new_new_n12499__ | ~new_new_n12507__;
  assign new_new_n12509__ = ~ys__n1099 & ~ys__n1110;
  assign new_new_n12510__ = new_new_n12496__ & new_new_n12509__;
  assign ys__n1138 = ~new_new_n12495__ | ~new_new_n12510__;
  assign ys__n1142 = ~new_new_n12490__ | ~new_new_n12495__;
  assign ys__n1143 = ys__n1106 | ys__n1141;
  assign ys__n3118 = ys__n874 & ys__n1147;
  assign ys__n1146 = ys__n140 | ~ys__n3118;
  assign ys__n1148 = ys__n1147 | ys__n1047;
  assign new_new_n12517__ = ~ys__n1154 & ~ys__n1156;
  assign new_new_n12518__ = ~ys__n1157 & ys__n24591;
  assign new_new_n12519__ = new_new_n12517__ & new_new_n12518__;
  assign ys__n18137 = ys__n1151 | ys__n1153;
  assign new_new_n12521__ = ~ys__n1047 & ~ys__n18137;
  assign ys__n1161 = ~new_new_n12519__ | ~new_new_n12521__;
  assign ys__n1163 = new_new_n12287__ & new_new_n12414__;
  assign ys__n1164 = new_new_n12287__ & new_new_n12417__;
  assign ys__n1165 = new_new_n12287__ & new_new_n12408__;
  assign new_new_n12526__ = new_new_n12241__ & new_new_n12373__;
  assign ys__n1167 = new_new_n12396__ & new_new_n12526__;
  assign new_new_n12528__ = ~ys__n738 & new_new_n10820__;
  assign ys__n1170 = new_new_n11343__ & new_new_n12528__;
  assign ys__n1171 = ~ys__n874 | new_new_n12108__;
  assign ys__n1183 = ~ys__n858 | new_new_n12106__;
  assign ys__n1189 = ~ys__n856 | new_new_n12106__;
  assign ys__n1195 = ~ys__n854 | new_new_n12106__;
  assign ys__n1201 = ~ys__n852 | new_new_n12106__;
  assign ys__n1207 = ~ys__n850 | new_new_n12106__;
  assign ys__n1213 = ~ys__n848 | new_new_n12106__;
  assign ys__n1219 = ~ys__n846 | new_new_n12106__;
  assign ys__n1222 = ~ys__n844 | new_new_n12106__;
  assign ys__n1228 = ~ys__n842 | new_new_n12106__;
  assign ys__n1234 = ~ys__n840 | new_new_n12106__;
  assign ys__n1240 = ~ys__n838 | new_new_n12106__;
  assign ys__n1246 = ~ys__n836 | new_new_n12106__;
  assign ys__n1252 = ~ys__n834 | new_new_n12106__;
  assign ys__n1258 = ~ys__n832 | new_new_n12106__;
  assign ys__n1261 = ~ys__n830 | new_new_n12106__;
  assign ys__n1266 = ~ys__n828 | ~new_new_n11726__;
  assign ys__n1272 = ~ys__n826 | ~new_new_n11726__;
  assign ys__n1278 = ~ys__n824 | ~new_new_n11726__;
  assign ys__n1284 = ~ys__n822 | ~new_new_n11726__;
  assign ys__n1290 = ~ys__n820 | ~new_new_n11726__;
  assign ys__n1296 = ~ys__n818 | ~new_new_n11726__;
  assign ys__n1303 = ~ys__n816 | ~new_new_n11726__;
  assign new_new_n12553__ = new_new_n12250__ & new_new_n12373__;
  assign ys__n1377 = new_new_n12396__ & new_new_n12553__;
  assign new_new_n12555__ = ~ys__n536 & ~ys__n538;
  assign new_new_n12556__ = ys__n33403 & ~new_new_n12555__;
  assign new_new_n12557__ = ~ys__n935 & ys__n30863;
  assign new_new_n12558__ = ~ys__n33384 & new_new_n12557__;
  assign new_new_n12559__ = ~new_new_n12556__ & new_new_n12558__;
  assign new_new_n12560__ = ~ys__n738 & new_new_n12559__;
  assign ys__n1386 = ys__n4566 & new_new_n12560__;
  assign new_new_n12562__ = new_new_n12249__ & new_new_n12250__;
  assign ys__n1445 = new_new_n12396__ & new_new_n12562__;
  assign new_new_n12564__ = ~ys__n252 & ~ys__n254;
  assign new_new_n12565__ = ~ys__n250 & new_new_n12564__;
  assign new_new_n12566__ = ~ys__n246 & ~ys__n270;
  assign new_new_n12567__ = ys__n20273 & ys__n814;
  assign new_new_n12568__ = ~ys__n278 & new_new_n12567__;
  assign new_new_n12569__ = new_new_n12566__ & new_new_n12568__;
  assign ys__n1470 = ~new_new_n12565__ | ~new_new_n12569__;
  assign ys__n1591 = new_new_n12287__ & new_new_n12404__;
  assign ys__n1598 = ys__n44892 & ~ys__n4566;
  assign new_new_n12573__ = ~ys__n44840 & ~ys__n44842;
  assign new_new_n12574__ = ~ys__n4566 & ~new_new_n12573__;
  assign new_new_n12575__ = ys__n874 & ~ys__n1598;
  assign ys__n1601 = new_new_n12574__ | ~new_new_n12575__;
  assign ys__n1616 = new_new_n12287__ & new_new_n12389__;
  assign ys__n38453 = ~ys__n564 | ~new_new_n12555__;
  assign new_new_n12579__ = ~new_new_n10990__ & ~ys__n38453;
  assign new_new_n12580__ = ~new_new_n11005__ & ~new_new_n12579__;
  assign new_new_n12581__ = new_new_n11006__ & new_new_n12580__;
  assign new_new_n12582__ = ~new_new_n12559__ & new_new_n12579__;
  assign new_new_n12583__ = ~ys__n738 & ys__n4566;
  assign new_new_n12584__ = ~new_new_n12582__ & new_new_n12583__;
  assign new_new_n12585__ = ys__n738 & ~new_new_n12579__;
  assign new_new_n12586__ = ~new_new_n12584__ & ~new_new_n12585__;
  assign ys__n1790 = ~new_new_n12581__ & new_new_n12586__;
  assign new_new_n12588__ = ys__n33384 & ys__n38451;
  assign new_new_n12589__ = ~ys__n4177 & ~ys__n33394;
  assign ys__n26555 = ys__n34959 & new_new_n12589__;
  assign ys__n1802 = new_new_n12588__ | ys__n26555;
  assign new_new_n12592__ = ~ys__n348 & ~ys__n2924;
  assign new_new_n12593__ = ~ys__n162 & ys__n346;
  assign new_new_n12594__ = new_new_n12592__ & new_new_n12593__;
  assign new_new_n12595__ = ~ys__n342 & ~ys__n350;
  assign new_new_n12596__ = ys__n160 & ~ys__n344;
  assign new_new_n12597__ = new_new_n12595__ & new_new_n12596__;
  assign new_new_n12598__ = ys__n352 & new_new_n12597__;
  assign new_new_n12599__ = new_new_n12594__ & new_new_n12598__;
  assign new_new_n12600__ = ys__n342 & ~ys__n350;
  assign new_new_n12601__ = ys__n352 & new_new_n12596__;
  assign new_new_n12602__ = new_new_n12600__ & new_new_n12601__;
  assign new_new_n12603__ = new_new_n12594__ & new_new_n12602__;
  assign new_new_n12604__ = ~new_new_n12599__ & ~new_new_n12603__;
  assign new_new_n12605__ = ~ys__n160 & ~ys__n344;
  assign new_new_n12606__ = new_new_n12337__ & new_new_n12605__;
  assign new_new_n12607__ = ys__n352 & new_new_n12349__;
  assign new_new_n12608__ = new_new_n12606__ & new_new_n12607__;
  assign ys__n1817 = ~new_new_n12604__ | new_new_n12608__;
  assign new_new_n12610__ = new_new_n12242__ & new_new_n12249__;
  assign ys__n1835 = new_new_n12396__ & new_new_n12610__;
  assign new_new_n12612__ = ys__n480 & ~ys__n754;
  assign new_new_n12613__ = ~ys__n482 & ~ys__n756;
  assign new_new_n12614__ = new_new_n12612__ & new_new_n12613__;
  assign new_new_n12615__ = ys__n23652 & new_new_n12614__;
  assign new_new_n12616__ = new_new_n10973__ & new_new_n12614__;
  assign new_new_n12617__ = ys__n478 & new_new_n12616__;
  assign new_new_n12618__ = ~new_new_n12615__ & new_new_n12617__;
  assign new_new_n12619__ = ys__n478 & ~ys__n756;
  assign new_new_n12620__ = new_new_n10974__ & new_new_n12619__;
  assign new_new_n12621__ = ys__n482 & new_new_n12620__;
  assign new_new_n12622__ = new_new_n12612__ & new_new_n12621__;
  assign new_new_n12623__ = ~new_new_n12616__ & new_new_n12622__;
  assign new_new_n12624__ = ~new_new_n12615__ & new_new_n12623__;
  assign new_new_n12625__ = ~new_new_n12618__ & ~new_new_n12624__;
  assign new_new_n12626__ = ys__n478 & new_new_n12615__;
  assign new_new_n12627__ = new_new_n12625__ & ~new_new_n12626__;
  assign ys__n1837 = ~ys__n738 & ~new_new_n12627__;
  assign new_new_n12629__ = ys__n564 & ~new_new_n12555__;
  assign ys__n2152 = ys__n1386 | new_new_n12629__;
  assign new_new_n12631__ = new_new_n12250__ & new_new_n12358__;
  assign ys__n2365 = new_new_n12396__ & new_new_n12631__;
  assign new_new_n12633__ = new_new_n12250__ & new_new_n12369__;
  assign ys__n2400 = new_new_n12396__ & new_new_n12633__;
  assign new_new_n12635__ = ys__n38304 & ~ys__n4566;
  assign ys__n2423 = ~ys__n738 & new_new_n12635__;
  assign new_new_n12637__ = ys__n45046 & ys__n45580;
  assign new_new_n12638__ = ~ys__n45046 & ~ys__n45580;
  assign new_new_n12639__ = ~ys__n45622 & ~new_new_n12638__;
  assign new_new_n12640__ = ~new_new_n12637__ & new_new_n12639__;
  assign new_new_n12641__ = ys__n45049 & ys__n45582;
  assign new_new_n12642__ = ~ys__n45049 & ~ys__n45582;
  assign new_new_n12643__ = ~ys__n45623 & ~new_new_n12642__;
  assign new_new_n12644__ = ~new_new_n12641__ & new_new_n12643__;
  assign new_new_n12645__ = ~new_new_n12640__ & ~new_new_n12644__;
  assign new_new_n12646__ = ys__n45052 & ys__n45584;
  assign new_new_n12647__ = ~ys__n45052 & ~ys__n45584;
  assign new_new_n12648__ = ~ys__n45624 & ~new_new_n12647__;
  assign new_new_n12649__ = ~new_new_n12646__ & new_new_n12648__;
  assign new_new_n12650__ = ys__n45055 & ys__n45586;
  assign new_new_n12651__ = ~ys__n45055 & ~ys__n45586;
  assign new_new_n12652__ = ~ys__n45625 & ~new_new_n12651__;
  assign new_new_n12653__ = ~new_new_n12650__ & new_new_n12652__;
  assign new_new_n12654__ = ~new_new_n12649__ & ~new_new_n12653__;
  assign new_new_n12655__ = new_new_n12645__ & new_new_n12654__;
  assign new_new_n12656__ = ys__n45034 & ys__n45572;
  assign new_new_n12657__ = ~ys__n45034 & ~ys__n45572;
  assign new_new_n12658__ = ~ys__n45618 & ~new_new_n12657__;
  assign new_new_n12659__ = ~new_new_n12656__ & new_new_n12658__;
  assign new_new_n12660__ = ys__n45037 & ys__n45574;
  assign new_new_n12661__ = ~ys__n45037 & ~ys__n45574;
  assign new_new_n12662__ = ~ys__n45619 & ~new_new_n12661__;
  assign new_new_n12663__ = ~new_new_n12660__ & new_new_n12662__;
  assign new_new_n12664__ = ~new_new_n12659__ & ~new_new_n12663__;
  assign new_new_n12665__ = ys__n45040 & ys__n45576;
  assign new_new_n12666__ = ~ys__n45040 & ~ys__n45576;
  assign new_new_n12667__ = ~ys__n45620 & ~new_new_n12666__;
  assign new_new_n12668__ = ~new_new_n12665__ & new_new_n12667__;
  assign new_new_n12669__ = ys__n45043 & ys__n45578;
  assign new_new_n12670__ = ~ys__n45043 & ~ys__n45578;
  assign new_new_n12671__ = ~ys__n45621 & ~new_new_n12670__;
  assign new_new_n12672__ = ~new_new_n12669__ & new_new_n12671__;
  assign new_new_n12673__ = ~new_new_n12668__ & ~new_new_n12672__;
  assign new_new_n12674__ = new_new_n12664__ & new_new_n12673__;
  assign new_new_n12675__ = new_new_n12655__ & new_new_n12674__;
  assign new_new_n12676__ = ys__n45070 & ys__n45596;
  assign new_new_n12677__ = ~ys__n45070 & ~ys__n45596;
  assign new_new_n12678__ = ~ys__n45630 & ~new_new_n12677__;
  assign new_new_n12679__ = ~new_new_n12676__ & new_new_n12678__;
  assign new_new_n12680__ = ys__n45073 & ys__n45598;
  assign new_new_n12681__ = ~ys__n45073 & ~ys__n45598;
  assign new_new_n12682__ = ~ys__n45631 & ~new_new_n12681__;
  assign new_new_n12683__ = ~new_new_n12680__ & new_new_n12682__;
  assign new_new_n12684__ = ~new_new_n12679__ & ~new_new_n12683__;
  assign new_new_n12685__ = ys__n45076 & ys__n45600;
  assign new_new_n12686__ = ~ys__n45076 & ~ys__n45600;
  assign new_new_n12687__ = ~ys__n45632 & ~new_new_n12686__;
  assign new_new_n12688__ = ~new_new_n12685__ & new_new_n12687__;
  assign new_new_n12689__ = ys__n45079 & ys__n45602;
  assign new_new_n12690__ = ~ys__n45079 & ~ys__n45602;
  assign new_new_n12691__ = ~ys__n45633 & ~new_new_n12690__;
  assign new_new_n12692__ = ~new_new_n12689__ & new_new_n12691__;
  assign new_new_n12693__ = ~new_new_n12688__ & ~new_new_n12692__;
  assign new_new_n12694__ = new_new_n12684__ & new_new_n12693__;
  assign new_new_n12695__ = ys__n45058 & ys__n45588;
  assign new_new_n12696__ = ~ys__n45058 & ~ys__n45588;
  assign new_new_n12697__ = ~ys__n45626 & ~new_new_n12696__;
  assign new_new_n12698__ = ~new_new_n12695__ & new_new_n12697__;
  assign new_new_n12699__ = ys__n45061 & ys__n45590;
  assign new_new_n12700__ = ~ys__n45061 & ~ys__n45590;
  assign new_new_n12701__ = ~ys__n45627 & ~new_new_n12700__;
  assign new_new_n12702__ = ~new_new_n12699__ & new_new_n12701__;
  assign new_new_n12703__ = ~new_new_n12698__ & ~new_new_n12702__;
  assign new_new_n12704__ = ys__n45064 & ys__n45592;
  assign new_new_n12705__ = ~ys__n45064 & ~ys__n45592;
  assign new_new_n12706__ = ~ys__n45628 & ~new_new_n12705__;
  assign new_new_n12707__ = ~new_new_n12704__ & new_new_n12706__;
  assign new_new_n12708__ = ys__n45067 & ys__n45594;
  assign new_new_n12709__ = ~ys__n45067 & ~ys__n45594;
  assign new_new_n12710__ = ~ys__n45629 & ~new_new_n12709__;
  assign new_new_n12711__ = ~new_new_n12708__ & new_new_n12710__;
  assign new_new_n12712__ = ~new_new_n12707__ & ~new_new_n12711__;
  assign new_new_n12713__ = new_new_n12703__ & new_new_n12712__;
  assign new_new_n12714__ = new_new_n12694__ & new_new_n12713__;
  assign new_new_n12715__ = new_new_n12675__ & new_new_n12714__;
  assign new_new_n12716__ = ys__n44992 & ys__n45544;
  assign new_new_n12717__ = ~ys__n44992 & ~ys__n45544;
  assign new_new_n12718__ = ~ys__n45604 & ~new_new_n12717__;
  assign new_new_n12719__ = ~new_new_n12716__ & new_new_n12718__;
  assign new_new_n12720__ = ys__n44995 & ys__n45546;
  assign new_new_n12721__ = ~ys__n44995 & ~ys__n45546;
  assign new_new_n12722__ = ~ys__n45605 & ~new_new_n12721__;
  assign new_new_n12723__ = ~new_new_n12720__ & new_new_n12722__;
  assign new_new_n12724__ = ~new_new_n12719__ & ~new_new_n12723__;
  assign new_new_n12725__ = ys__n44998 & ys__n45548;
  assign new_new_n12726__ = ~ys__n44998 & ~ys__n45548;
  assign new_new_n12727__ = ~ys__n45606 & ~new_new_n12726__;
  assign new_new_n12728__ = ~new_new_n12725__ & new_new_n12727__;
  assign new_new_n12729__ = ys__n45001 & ys__n45550;
  assign new_new_n12730__ = ~ys__n45001 & ~ys__n45550;
  assign new_new_n12731__ = ~ys__n45607 & ~new_new_n12730__;
  assign new_new_n12732__ = ~new_new_n12729__ & new_new_n12731__;
  assign new_new_n12733__ = ~new_new_n12728__ & ~new_new_n12732__;
  assign new_new_n12734__ = ys__n45004 & ys__n45552;
  assign new_new_n12735__ = ~ys__n45004 & ~ys__n45552;
  assign new_new_n12736__ = ~ys__n45608 & ~new_new_n12735__;
  assign new_new_n12737__ = ~new_new_n12734__ & new_new_n12736__;
  assign new_new_n12738__ = ys__n45007 & ys__n45554;
  assign new_new_n12739__ = ~ys__n45007 & ~ys__n45554;
  assign new_new_n12740__ = ~ys__n45609 & ~new_new_n12739__;
  assign new_new_n12741__ = ~new_new_n12738__ & new_new_n12740__;
  assign new_new_n12742__ = ~new_new_n12737__ & ~new_new_n12741__;
  assign new_new_n12743__ = new_new_n12733__ & new_new_n12742__;
  assign new_new_n12744__ = new_new_n12724__ & new_new_n12743__;
  assign new_new_n12745__ = ys__n45022 & ys__n45564;
  assign new_new_n12746__ = ~ys__n45022 & ~ys__n45564;
  assign new_new_n12747__ = ~ys__n45614 & ~new_new_n12746__;
  assign new_new_n12748__ = ~new_new_n12745__ & new_new_n12747__;
  assign new_new_n12749__ = ys__n45025 & ys__n45566;
  assign new_new_n12750__ = ~ys__n45025 & ~ys__n45566;
  assign new_new_n12751__ = ~ys__n45615 & ~new_new_n12750__;
  assign new_new_n12752__ = ~new_new_n12749__ & new_new_n12751__;
  assign new_new_n12753__ = ~new_new_n12748__ & ~new_new_n12752__;
  assign new_new_n12754__ = ys__n45028 & ys__n45568;
  assign new_new_n12755__ = ~ys__n45028 & ~ys__n45568;
  assign new_new_n12756__ = ~ys__n45616 & ~new_new_n12755__;
  assign new_new_n12757__ = ~new_new_n12754__ & new_new_n12756__;
  assign new_new_n12758__ = ys__n45031 & ys__n45570;
  assign new_new_n12759__ = ~ys__n45031 & ~ys__n45570;
  assign new_new_n12760__ = ~ys__n45617 & ~new_new_n12759__;
  assign new_new_n12761__ = ~new_new_n12758__ & new_new_n12760__;
  assign new_new_n12762__ = ~new_new_n12757__ & ~new_new_n12761__;
  assign new_new_n12763__ = new_new_n12753__ & new_new_n12762__;
  assign new_new_n12764__ = ys__n45010 & ys__n45556;
  assign new_new_n12765__ = ~ys__n45010 & ~ys__n45556;
  assign new_new_n12766__ = ~ys__n45610 & ~new_new_n12765__;
  assign new_new_n12767__ = ~new_new_n12764__ & new_new_n12766__;
  assign new_new_n12768__ = ys__n45013 & ys__n45558;
  assign new_new_n12769__ = ~ys__n45013 & ~ys__n45558;
  assign new_new_n12770__ = ~ys__n45611 & ~new_new_n12769__;
  assign new_new_n12771__ = ~new_new_n12768__ & new_new_n12770__;
  assign new_new_n12772__ = ~new_new_n12767__ & ~new_new_n12771__;
  assign new_new_n12773__ = ys__n45016 & ys__n45560;
  assign new_new_n12774__ = ~ys__n45016 & ~ys__n45560;
  assign new_new_n12775__ = ~ys__n45612 & ~new_new_n12774__;
  assign new_new_n12776__ = ~new_new_n12773__ & new_new_n12775__;
  assign new_new_n12777__ = ys__n45019 & ys__n45562;
  assign new_new_n12778__ = ~ys__n45019 & ~ys__n45562;
  assign new_new_n12779__ = ~ys__n45613 & ~new_new_n12778__;
  assign new_new_n12780__ = ~new_new_n12777__ & new_new_n12779__;
  assign new_new_n12781__ = ~new_new_n12776__ & ~new_new_n12780__;
  assign new_new_n12782__ = new_new_n12772__ & new_new_n12781__;
  assign new_new_n12783__ = new_new_n12763__ & new_new_n12782__;
  assign new_new_n12784__ = new_new_n12744__ & new_new_n12783__;
  assign new_new_n12785__ = new_new_n12715__ & new_new_n12784__;
  assign new_new_n12786__ = ys__n45172 & ys__n45674;
  assign new_new_n12787__ = ~ys__n45172 & ~ys__n45674;
  assign new_new_n12788__ = ~ys__n45700 & ~new_new_n12787__;
  assign new_new_n12789__ = ~new_new_n12786__ & new_new_n12788__;
  assign new_new_n12790__ = ys__n45175 & ys__n45676;
  assign new_new_n12791__ = ~ys__n45175 & ~ys__n45676;
  assign new_new_n12792__ = ~ys__n45700 & ~new_new_n12791__;
  assign new_new_n12793__ = ~new_new_n12790__ & new_new_n12792__;
  assign new_new_n12794__ = ~new_new_n12789__ & ~new_new_n12793__;
  assign new_new_n12795__ = ys__n45178 & ys__n45678;
  assign new_new_n12796__ = ~ys__n45178 & ~ys__n45678;
  assign new_new_n12797__ = ~ys__n45700 & ~new_new_n12796__;
  assign new_new_n12798__ = ~new_new_n12795__ & new_new_n12797__;
  assign new_new_n12799__ = ys__n45181 & ys__n45680;
  assign new_new_n12800__ = ~ys__n45181 & ~ys__n45680;
  assign new_new_n12801__ = ~ys__n45700 & ~new_new_n12800__;
  assign new_new_n12802__ = ~new_new_n12799__ & new_new_n12801__;
  assign new_new_n12803__ = ~new_new_n12798__ & ~new_new_n12802__;
  assign new_new_n12804__ = new_new_n12794__ & new_new_n12803__;
  assign new_new_n12805__ = ys__n45160 & ys__n45666;
  assign new_new_n12806__ = ~ys__n45160 & ~ys__n45666;
  assign new_new_n12807__ = ~ys__n45700 & ~new_new_n12806__;
  assign new_new_n12808__ = ~new_new_n12805__ & new_new_n12807__;
  assign new_new_n12809__ = ys__n45163 & ys__n45668;
  assign new_new_n12810__ = ~ys__n45163 & ~ys__n45668;
  assign new_new_n12811__ = ~ys__n45700 & ~new_new_n12810__;
  assign new_new_n12812__ = ~new_new_n12809__ & new_new_n12811__;
  assign new_new_n12813__ = ~new_new_n12808__ & ~new_new_n12812__;
  assign new_new_n12814__ = ys__n45166 & ys__n45670;
  assign new_new_n12815__ = ~ys__n45166 & ~ys__n45670;
  assign new_new_n12816__ = ~ys__n45700 & ~new_new_n12815__;
  assign new_new_n12817__ = ~new_new_n12814__ & new_new_n12816__;
  assign new_new_n12818__ = ys__n45169 & ys__n45672;
  assign new_new_n12819__ = ~ys__n45169 & ~ys__n45672;
  assign new_new_n12820__ = ~ys__n45700 & ~new_new_n12819__;
  assign new_new_n12821__ = ~new_new_n12818__ & new_new_n12820__;
  assign new_new_n12822__ = ~new_new_n12817__ & ~new_new_n12821__;
  assign new_new_n12823__ = new_new_n12813__ & new_new_n12822__;
  assign new_new_n12824__ = new_new_n12804__ & new_new_n12823__;
  assign new_new_n12825__ = ys__n45196 & ys__n45690;
  assign new_new_n12826__ = ~ys__n45196 & ~ys__n45690;
  assign new_new_n12827__ = ~ys__n45701 & ~new_new_n12826__;
  assign new_new_n12828__ = ~new_new_n12825__ & new_new_n12827__;
  assign new_new_n12829__ = ys__n45199 & ys__n45692;
  assign new_new_n12830__ = ~ys__n45199 & ~ys__n45692;
  assign new_new_n12831__ = ~ys__n45701 & ~new_new_n12830__;
  assign new_new_n12832__ = ~new_new_n12829__ & new_new_n12831__;
  assign new_new_n12833__ = ~new_new_n12828__ & ~new_new_n12832__;
  assign new_new_n12834__ = ys__n45202 & ys__n45694;
  assign new_new_n12835__ = ~ys__n45202 & ~ys__n45694;
  assign new_new_n12836__ = ~ys__n45701 & ~new_new_n12835__;
  assign new_new_n12837__ = ~new_new_n12834__ & new_new_n12836__;
  assign new_new_n12838__ = ys__n45205 & ys__n45696;
  assign new_new_n12839__ = ~ys__n45205 & ~ys__n45696;
  assign new_new_n12840__ = ~ys__n45701 & ~new_new_n12839__;
  assign new_new_n12841__ = ~new_new_n12838__ & new_new_n12840__;
  assign new_new_n12842__ = ~new_new_n12837__ & ~new_new_n12841__;
  assign new_new_n12843__ = new_new_n12833__ & new_new_n12842__;
  assign new_new_n12844__ = ys__n45184 & ys__n45682;
  assign new_new_n12845__ = ~ys__n45184 & ~ys__n45682;
  assign new_new_n12846__ = ~ys__n45701 & ~new_new_n12845__;
  assign new_new_n12847__ = ~new_new_n12844__ & new_new_n12846__;
  assign new_new_n12848__ = ys__n45187 & ys__n45684;
  assign new_new_n12849__ = ~ys__n45187 & ~ys__n45684;
  assign new_new_n12850__ = ~ys__n45701 & ~new_new_n12849__;
  assign new_new_n12851__ = ~new_new_n12848__ & new_new_n12850__;
  assign new_new_n12852__ = ~new_new_n12847__ & ~new_new_n12851__;
  assign new_new_n12853__ = ys__n45190 & ys__n45686;
  assign new_new_n12854__ = ~ys__n45190 & ~ys__n45686;
  assign new_new_n12855__ = ~ys__n45701 & ~new_new_n12854__;
  assign new_new_n12856__ = ~new_new_n12853__ & new_new_n12855__;
  assign new_new_n12857__ = ys__n45193 & ys__n45688;
  assign new_new_n12858__ = ~ys__n45193 & ~ys__n45688;
  assign new_new_n12859__ = ~ys__n45701 & ~new_new_n12858__;
  assign new_new_n12860__ = ~new_new_n12857__ & new_new_n12859__;
  assign new_new_n12861__ = ~new_new_n12856__ & ~new_new_n12860__;
  assign new_new_n12862__ = new_new_n12852__ & new_new_n12861__;
  assign new_new_n12863__ = new_new_n12843__ & new_new_n12862__;
  assign new_new_n12864__ = new_new_n12824__ & new_new_n12863__;
  assign new_new_n12865__ = ys__n45124 & ys__n45642;
  assign new_new_n12866__ = ~ys__n45124 & ~ys__n45642;
  assign new_new_n12867__ = ~ys__n45698 & ~new_new_n12866__;
  assign new_new_n12868__ = ~new_new_n12865__ & new_new_n12867__;
  assign new_new_n12869__ = ys__n45127 & ys__n45644;
  assign new_new_n12870__ = ~ys__n45127 & ~ys__n45644;
  assign new_new_n12871__ = ~ys__n45698 & ~new_new_n12870__;
  assign new_new_n12872__ = ~new_new_n12869__ & new_new_n12871__;
  assign new_new_n12873__ = ~new_new_n12868__ & ~new_new_n12872__;
  assign new_new_n12874__ = ys__n45130 & ys__n45646;
  assign new_new_n12875__ = ~ys__n45130 & ~ys__n45646;
  assign new_new_n12876__ = ~ys__n45698 & ~new_new_n12875__;
  assign new_new_n12877__ = ~new_new_n12874__ & new_new_n12876__;
  assign new_new_n12878__ = ys__n45133 & ys__n45648;
  assign new_new_n12879__ = ~ys__n45133 & ~ys__n45648;
  assign new_new_n12880__ = ~ys__n45698 & ~new_new_n12879__;
  assign new_new_n12881__ = ~new_new_n12878__ & new_new_n12880__;
  assign new_new_n12882__ = ~new_new_n12877__ & ~new_new_n12881__;
  assign new_new_n12883__ = new_new_n12873__ & new_new_n12882__;
  assign new_new_n12884__ = ys__n45112 & ys__n45634;
  assign new_new_n12885__ = ~ys__n45112 & ~ys__n45634;
  assign new_new_n12886__ = ~ys__n45698 & ~new_new_n12885__;
  assign new_new_n12887__ = ~new_new_n12884__ & new_new_n12886__;
  assign new_new_n12888__ = ys__n45115 & ys__n45636;
  assign new_new_n12889__ = ~ys__n45115 & ~ys__n45636;
  assign new_new_n12890__ = ~ys__n45698 & ~new_new_n12889__;
  assign new_new_n12891__ = ~new_new_n12888__ & new_new_n12890__;
  assign new_new_n12892__ = ~new_new_n12887__ & ~new_new_n12891__;
  assign new_new_n12893__ = ys__n45118 & ys__n45638;
  assign new_new_n12894__ = ~ys__n45118 & ~ys__n45638;
  assign new_new_n12895__ = ~ys__n45698 & ~new_new_n12894__;
  assign new_new_n12896__ = ~new_new_n12893__ & new_new_n12895__;
  assign new_new_n12897__ = ys__n45121 & ys__n45640;
  assign new_new_n12898__ = ~ys__n45121 & ~ys__n45640;
  assign new_new_n12899__ = ~ys__n45698 & ~new_new_n12898__;
  assign new_new_n12900__ = ~new_new_n12897__ & new_new_n12899__;
  assign new_new_n12901__ = ~new_new_n12896__ & ~new_new_n12900__;
  assign new_new_n12902__ = new_new_n12892__ & new_new_n12901__;
  assign new_new_n12903__ = new_new_n12883__ & new_new_n12902__;
  assign new_new_n12904__ = ys__n45148 & ys__n45658;
  assign new_new_n12905__ = ~ys__n45148 & ~ys__n45658;
  assign new_new_n12906__ = ~ys__n45699 & ~new_new_n12905__;
  assign new_new_n12907__ = ~new_new_n12904__ & new_new_n12906__;
  assign new_new_n12908__ = ys__n45151 & ys__n45660;
  assign new_new_n12909__ = ~ys__n45151 & ~ys__n45660;
  assign new_new_n12910__ = ~ys__n45699 & ~new_new_n12909__;
  assign new_new_n12911__ = ~new_new_n12908__ & new_new_n12910__;
  assign new_new_n12912__ = ~new_new_n12907__ & ~new_new_n12911__;
  assign new_new_n12913__ = ys__n45154 & ys__n45662;
  assign new_new_n12914__ = ~ys__n45154 & ~ys__n45662;
  assign new_new_n12915__ = ~ys__n45699 & ~new_new_n12914__;
  assign new_new_n12916__ = ~new_new_n12913__ & new_new_n12915__;
  assign new_new_n12917__ = ys__n45157 & ys__n45664;
  assign new_new_n12918__ = ~ys__n45157 & ~ys__n45664;
  assign new_new_n12919__ = ~ys__n45699 & ~new_new_n12918__;
  assign new_new_n12920__ = ~new_new_n12917__ & new_new_n12919__;
  assign new_new_n12921__ = ~new_new_n12916__ & ~new_new_n12920__;
  assign new_new_n12922__ = new_new_n12912__ & new_new_n12921__;
  assign new_new_n12923__ = ys__n45136 & ys__n45650;
  assign new_new_n12924__ = ~ys__n45136 & ~ys__n45650;
  assign new_new_n12925__ = ~ys__n45699 & ~new_new_n12924__;
  assign new_new_n12926__ = ~new_new_n12923__ & new_new_n12925__;
  assign new_new_n12927__ = ys__n45139 & ys__n45652;
  assign new_new_n12928__ = ~ys__n45139 & ~ys__n45652;
  assign new_new_n12929__ = ~ys__n45699 & ~new_new_n12928__;
  assign new_new_n12930__ = ~new_new_n12927__ & new_new_n12929__;
  assign new_new_n12931__ = ~new_new_n12926__ & ~new_new_n12930__;
  assign new_new_n12932__ = ys__n45142 & ys__n45654;
  assign new_new_n12933__ = ~ys__n45142 & ~ys__n45654;
  assign new_new_n12934__ = ~ys__n45699 & ~new_new_n12933__;
  assign new_new_n12935__ = ~new_new_n12932__ & new_new_n12934__;
  assign new_new_n12936__ = ys__n45145 & ys__n45656;
  assign new_new_n12937__ = ~ys__n45145 & ~ys__n45656;
  assign new_new_n12938__ = ~ys__n45699 & ~new_new_n12937__;
  assign new_new_n12939__ = ~new_new_n12936__ & new_new_n12938__;
  assign new_new_n12940__ = ~new_new_n12935__ & ~new_new_n12939__;
  assign new_new_n12941__ = new_new_n12931__ & new_new_n12940__;
  assign new_new_n12942__ = new_new_n12922__ & new_new_n12941__;
  assign new_new_n12943__ = new_new_n12903__ & new_new_n12942__;
  assign new_new_n12944__ = new_new_n12864__ & new_new_n12943__;
  assign new_new_n12945__ = new_new_n12785__ & new_new_n12944__;
  assign new_new_n12946__ = ys__n45702 & new_new_n12945__;
  assign new_new_n12947__ = ys__n45046 & ys__n45416;
  assign new_new_n12948__ = ~ys__n45046 & ~ys__n45416;
  assign new_new_n12949__ = ~ys__n45458 & ~new_new_n12948__;
  assign new_new_n12950__ = ~new_new_n12947__ & new_new_n12949__;
  assign new_new_n12951__ = ys__n45049 & ys__n45418;
  assign new_new_n12952__ = ~ys__n45049 & ~ys__n45418;
  assign new_new_n12953__ = ~ys__n45459 & ~new_new_n12952__;
  assign new_new_n12954__ = ~new_new_n12951__ & new_new_n12953__;
  assign new_new_n12955__ = ~new_new_n12950__ & ~new_new_n12954__;
  assign new_new_n12956__ = ys__n45052 & ys__n45420;
  assign new_new_n12957__ = ~ys__n45052 & ~ys__n45420;
  assign new_new_n12958__ = ~ys__n45460 & ~new_new_n12957__;
  assign new_new_n12959__ = ~new_new_n12956__ & new_new_n12958__;
  assign new_new_n12960__ = ys__n45055 & ys__n45422;
  assign new_new_n12961__ = ~ys__n45055 & ~ys__n45422;
  assign new_new_n12962__ = ~ys__n45461 & ~new_new_n12961__;
  assign new_new_n12963__ = ~new_new_n12960__ & new_new_n12962__;
  assign new_new_n12964__ = ~new_new_n12959__ & ~new_new_n12963__;
  assign new_new_n12965__ = new_new_n12955__ & new_new_n12964__;
  assign new_new_n12966__ = ys__n45034 & ys__n45408;
  assign new_new_n12967__ = ~ys__n45034 & ~ys__n45408;
  assign new_new_n12968__ = ~ys__n45454 & ~new_new_n12967__;
  assign new_new_n12969__ = ~new_new_n12966__ & new_new_n12968__;
  assign new_new_n12970__ = ys__n45037 & ys__n45410;
  assign new_new_n12971__ = ~ys__n45037 & ~ys__n45410;
  assign new_new_n12972__ = ~ys__n45455 & ~new_new_n12971__;
  assign new_new_n12973__ = ~new_new_n12970__ & new_new_n12972__;
  assign new_new_n12974__ = ~new_new_n12969__ & ~new_new_n12973__;
  assign new_new_n12975__ = ys__n45040 & ys__n45412;
  assign new_new_n12976__ = ~ys__n45040 & ~ys__n45412;
  assign new_new_n12977__ = ~ys__n45456 & ~new_new_n12976__;
  assign new_new_n12978__ = ~new_new_n12975__ & new_new_n12977__;
  assign new_new_n12979__ = ys__n45043 & ys__n45414;
  assign new_new_n12980__ = ~ys__n45043 & ~ys__n45414;
  assign new_new_n12981__ = ~ys__n45457 & ~new_new_n12980__;
  assign new_new_n12982__ = ~new_new_n12979__ & new_new_n12981__;
  assign new_new_n12983__ = ~new_new_n12978__ & ~new_new_n12982__;
  assign new_new_n12984__ = new_new_n12974__ & new_new_n12983__;
  assign new_new_n12985__ = new_new_n12965__ & new_new_n12984__;
  assign new_new_n12986__ = ys__n45070 & ys__n45432;
  assign new_new_n12987__ = ~ys__n45070 & ~ys__n45432;
  assign new_new_n12988__ = ~ys__n45466 & ~new_new_n12987__;
  assign new_new_n12989__ = ~new_new_n12986__ & new_new_n12988__;
  assign new_new_n12990__ = ys__n45073 & ys__n45434;
  assign new_new_n12991__ = ~ys__n45073 & ~ys__n45434;
  assign new_new_n12992__ = ~ys__n45467 & ~new_new_n12991__;
  assign new_new_n12993__ = ~new_new_n12990__ & new_new_n12992__;
  assign new_new_n12994__ = ~new_new_n12989__ & ~new_new_n12993__;
  assign new_new_n12995__ = ys__n45076 & ys__n45436;
  assign new_new_n12996__ = ~ys__n45076 & ~ys__n45436;
  assign new_new_n12997__ = ~ys__n45468 & ~new_new_n12996__;
  assign new_new_n12998__ = ~new_new_n12995__ & new_new_n12997__;
  assign new_new_n12999__ = ys__n45079 & ys__n45438;
  assign new_new_n13000__ = ~ys__n45079 & ~ys__n45438;
  assign new_new_n13001__ = ~ys__n45469 & ~new_new_n13000__;
  assign new_new_n13002__ = ~new_new_n12999__ & new_new_n13001__;
  assign new_new_n13003__ = ~new_new_n12998__ & ~new_new_n13002__;
  assign new_new_n13004__ = new_new_n12994__ & new_new_n13003__;
  assign new_new_n13005__ = ys__n45058 & ys__n45424;
  assign new_new_n13006__ = ~ys__n45058 & ~ys__n45424;
  assign new_new_n13007__ = ~ys__n45462 & ~new_new_n13006__;
  assign new_new_n13008__ = ~new_new_n13005__ & new_new_n13007__;
  assign new_new_n13009__ = ys__n45061 & ys__n45426;
  assign new_new_n13010__ = ~ys__n45061 & ~ys__n45426;
  assign new_new_n13011__ = ~ys__n45463 & ~new_new_n13010__;
  assign new_new_n13012__ = ~new_new_n13009__ & new_new_n13011__;
  assign new_new_n13013__ = ~new_new_n13008__ & ~new_new_n13012__;
  assign new_new_n13014__ = ys__n45064 & ys__n45428;
  assign new_new_n13015__ = ~ys__n45064 & ~ys__n45428;
  assign new_new_n13016__ = ~ys__n45464 & ~new_new_n13015__;
  assign new_new_n13017__ = ~new_new_n13014__ & new_new_n13016__;
  assign new_new_n13018__ = ys__n45067 & ys__n45430;
  assign new_new_n13019__ = ~ys__n45067 & ~ys__n45430;
  assign new_new_n13020__ = ~ys__n45465 & ~new_new_n13019__;
  assign new_new_n13021__ = ~new_new_n13018__ & new_new_n13020__;
  assign new_new_n13022__ = ~new_new_n13017__ & ~new_new_n13021__;
  assign new_new_n13023__ = new_new_n13013__ & new_new_n13022__;
  assign new_new_n13024__ = new_new_n13004__ & new_new_n13023__;
  assign new_new_n13025__ = new_new_n12985__ & new_new_n13024__;
  assign new_new_n13026__ = ys__n44992 & ys__n45380;
  assign new_new_n13027__ = ~ys__n44992 & ~ys__n45380;
  assign new_new_n13028__ = ~ys__n45440 & ~new_new_n13027__;
  assign new_new_n13029__ = ~new_new_n13026__ & new_new_n13028__;
  assign new_new_n13030__ = ys__n44995 & ys__n45382;
  assign new_new_n13031__ = ~ys__n44995 & ~ys__n45382;
  assign new_new_n13032__ = ~ys__n45441 & ~new_new_n13031__;
  assign new_new_n13033__ = ~new_new_n13030__ & new_new_n13032__;
  assign new_new_n13034__ = ~new_new_n13029__ & ~new_new_n13033__;
  assign new_new_n13035__ = ys__n44998 & ys__n45384;
  assign new_new_n13036__ = ~ys__n44998 & ~ys__n45384;
  assign new_new_n13037__ = ~ys__n45442 & ~new_new_n13036__;
  assign new_new_n13038__ = ~new_new_n13035__ & new_new_n13037__;
  assign new_new_n13039__ = ys__n45001 & ys__n45386;
  assign new_new_n13040__ = ~ys__n45001 & ~ys__n45386;
  assign new_new_n13041__ = ~ys__n45443 & ~new_new_n13040__;
  assign new_new_n13042__ = ~new_new_n13039__ & new_new_n13041__;
  assign new_new_n13043__ = ~new_new_n13038__ & ~new_new_n13042__;
  assign new_new_n13044__ = ys__n45004 & ys__n45388;
  assign new_new_n13045__ = ~ys__n45004 & ~ys__n45388;
  assign new_new_n13046__ = ~ys__n45444 & ~new_new_n13045__;
  assign new_new_n13047__ = ~new_new_n13044__ & new_new_n13046__;
  assign new_new_n13048__ = ys__n45007 & ys__n45390;
  assign new_new_n13049__ = ~ys__n45007 & ~ys__n45390;
  assign new_new_n13050__ = ~ys__n45445 & ~new_new_n13049__;
  assign new_new_n13051__ = ~new_new_n13048__ & new_new_n13050__;
  assign new_new_n13052__ = ~new_new_n13047__ & ~new_new_n13051__;
  assign new_new_n13053__ = new_new_n13043__ & new_new_n13052__;
  assign new_new_n13054__ = new_new_n13034__ & new_new_n13053__;
  assign new_new_n13055__ = ys__n45022 & ys__n45400;
  assign new_new_n13056__ = ~ys__n45022 & ~ys__n45400;
  assign new_new_n13057__ = ~ys__n45450 & ~new_new_n13056__;
  assign new_new_n13058__ = ~new_new_n13055__ & new_new_n13057__;
  assign new_new_n13059__ = ys__n45025 & ys__n45402;
  assign new_new_n13060__ = ~ys__n45025 & ~ys__n45402;
  assign new_new_n13061__ = ~ys__n45451 & ~new_new_n13060__;
  assign new_new_n13062__ = ~new_new_n13059__ & new_new_n13061__;
  assign new_new_n13063__ = ~new_new_n13058__ & ~new_new_n13062__;
  assign new_new_n13064__ = ys__n45028 & ys__n45404;
  assign new_new_n13065__ = ~ys__n45028 & ~ys__n45404;
  assign new_new_n13066__ = ~ys__n45452 & ~new_new_n13065__;
  assign new_new_n13067__ = ~new_new_n13064__ & new_new_n13066__;
  assign new_new_n13068__ = ys__n45031 & ys__n45406;
  assign new_new_n13069__ = ~ys__n45031 & ~ys__n45406;
  assign new_new_n13070__ = ~ys__n45453 & ~new_new_n13069__;
  assign new_new_n13071__ = ~new_new_n13068__ & new_new_n13070__;
  assign new_new_n13072__ = ~new_new_n13067__ & ~new_new_n13071__;
  assign new_new_n13073__ = new_new_n13063__ & new_new_n13072__;
  assign new_new_n13074__ = ys__n45010 & ys__n45392;
  assign new_new_n13075__ = ~ys__n45010 & ~ys__n45392;
  assign new_new_n13076__ = ~ys__n45446 & ~new_new_n13075__;
  assign new_new_n13077__ = ~new_new_n13074__ & new_new_n13076__;
  assign new_new_n13078__ = ys__n45013 & ys__n45394;
  assign new_new_n13079__ = ~ys__n45013 & ~ys__n45394;
  assign new_new_n13080__ = ~ys__n45447 & ~new_new_n13079__;
  assign new_new_n13081__ = ~new_new_n13078__ & new_new_n13080__;
  assign new_new_n13082__ = ~new_new_n13077__ & ~new_new_n13081__;
  assign new_new_n13083__ = ys__n45016 & ys__n45396;
  assign new_new_n13084__ = ~ys__n45016 & ~ys__n45396;
  assign new_new_n13085__ = ~ys__n45448 & ~new_new_n13084__;
  assign new_new_n13086__ = ~new_new_n13083__ & new_new_n13085__;
  assign new_new_n13087__ = ys__n45019 & ys__n45398;
  assign new_new_n13088__ = ~ys__n45019 & ~ys__n45398;
  assign new_new_n13089__ = ~ys__n45449 & ~new_new_n13088__;
  assign new_new_n13090__ = ~new_new_n13087__ & new_new_n13089__;
  assign new_new_n13091__ = ~new_new_n13086__ & ~new_new_n13090__;
  assign new_new_n13092__ = new_new_n13082__ & new_new_n13091__;
  assign new_new_n13093__ = new_new_n13073__ & new_new_n13092__;
  assign new_new_n13094__ = new_new_n13054__ & new_new_n13093__;
  assign new_new_n13095__ = new_new_n13025__ & new_new_n13094__;
  assign new_new_n13096__ = ys__n45172 & ys__n45510;
  assign new_new_n13097__ = ~ys__n45172 & ~ys__n45510;
  assign new_new_n13098__ = ~ys__n45536 & ~new_new_n13097__;
  assign new_new_n13099__ = ~new_new_n13096__ & new_new_n13098__;
  assign new_new_n13100__ = ys__n45175 & ys__n45512;
  assign new_new_n13101__ = ~ys__n45175 & ~ys__n45512;
  assign new_new_n13102__ = ~ys__n45536 & ~new_new_n13101__;
  assign new_new_n13103__ = ~new_new_n13100__ & new_new_n13102__;
  assign new_new_n13104__ = ~new_new_n13099__ & ~new_new_n13103__;
  assign new_new_n13105__ = ys__n45178 & ys__n45514;
  assign new_new_n13106__ = ~ys__n45178 & ~ys__n45514;
  assign new_new_n13107__ = ~ys__n45536 & ~new_new_n13106__;
  assign new_new_n13108__ = ~new_new_n13105__ & new_new_n13107__;
  assign new_new_n13109__ = ys__n45181 & ys__n45516;
  assign new_new_n13110__ = ~ys__n45181 & ~ys__n45516;
  assign new_new_n13111__ = ~ys__n45536 & ~new_new_n13110__;
  assign new_new_n13112__ = ~new_new_n13109__ & new_new_n13111__;
  assign new_new_n13113__ = ~new_new_n13108__ & ~new_new_n13112__;
  assign new_new_n13114__ = new_new_n13104__ & new_new_n13113__;
  assign new_new_n13115__ = ys__n45160 & ys__n45502;
  assign new_new_n13116__ = ~ys__n45160 & ~ys__n45502;
  assign new_new_n13117__ = ~ys__n45536 & ~new_new_n13116__;
  assign new_new_n13118__ = ~new_new_n13115__ & new_new_n13117__;
  assign new_new_n13119__ = ys__n45163 & ys__n45504;
  assign new_new_n13120__ = ~ys__n45163 & ~ys__n45504;
  assign new_new_n13121__ = ~ys__n45536 & ~new_new_n13120__;
  assign new_new_n13122__ = ~new_new_n13119__ & new_new_n13121__;
  assign new_new_n13123__ = ~new_new_n13118__ & ~new_new_n13122__;
  assign new_new_n13124__ = ys__n45166 & ys__n45506;
  assign new_new_n13125__ = ~ys__n45166 & ~ys__n45506;
  assign new_new_n13126__ = ~ys__n45536 & ~new_new_n13125__;
  assign new_new_n13127__ = ~new_new_n13124__ & new_new_n13126__;
  assign new_new_n13128__ = ys__n45169 & ys__n45508;
  assign new_new_n13129__ = ~ys__n45169 & ~ys__n45508;
  assign new_new_n13130__ = ~ys__n45536 & ~new_new_n13129__;
  assign new_new_n13131__ = ~new_new_n13128__ & new_new_n13130__;
  assign new_new_n13132__ = ~new_new_n13127__ & ~new_new_n13131__;
  assign new_new_n13133__ = new_new_n13123__ & new_new_n13132__;
  assign new_new_n13134__ = new_new_n13114__ & new_new_n13133__;
  assign new_new_n13135__ = ys__n45196 & ys__n45526;
  assign new_new_n13136__ = ~ys__n45196 & ~ys__n45526;
  assign new_new_n13137__ = ~ys__n45537 & ~new_new_n13136__;
  assign new_new_n13138__ = ~new_new_n13135__ & new_new_n13137__;
  assign new_new_n13139__ = ys__n45199 & ys__n45528;
  assign new_new_n13140__ = ~ys__n45199 & ~ys__n45528;
  assign new_new_n13141__ = ~ys__n45537 & ~new_new_n13140__;
  assign new_new_n13142__ = ~new_new_n13139__ & new_new_n13141__;
  assign new_new_n13143__ = ~new_new_n13138__ & ~new_new_n13142__;
  assign new_new_n13144__ = ys__n45202 & ys__n45530;
  assign new_new_n13145__ = ~ys__n45202 & ~ys__n45530;
  assign new_new_n13146__ = ~ys__n45537 & ~new_new_n13145__;
  assign new_new_n13147__ = ~new_new_n13144__ & new_new_n13146__;
  assign new_new_n13148__ = ys__n45205 & ys__n45532;
  assign new_new_n13149__ = ~ys__n45205 & ~ys__n45532;
  assign new_new_n13150__ = ~ys__n45537 & ~new_new_n13149__;
  assign new_new_n13151__ = ~new_new_n13148__ & new_new_n13150__;
  assign new_new_n13152__ = ~new_new_n13147__ & ~new_new_n13151__;
  assign new_new_n13153__ = new_new_n13143__ & new_new_n13152__;
  assign new_new_n13154__ = ys__n45184 & ys__n45518;
  assign new_new_n13155__ = ~ys__n45184 & ~ys__n45518;
  assign new_new_n13156__ = ~ys__n45537 & ~new_new_n13155__;
  assign new_new_n13157__ = ~new_new_n13154__ & new_new_n13156__;
  assign new_new_n13158__ = ys__n45187 & ys__n45520;
  assign new_new_n13159__ = ~ys__n45187 & ~ys__n45520;
  assign new_new_n13160__ = ~ys__n45537 & ~new_new_n13159__;
  assign new_new_n13161__ = ~new_new_n13158__ & new_new_n13160__;
  assign new_new_n13162__ = ~new_new_n13157__ & ~new_new_n13161__;
  assign new_new_n13163__ = ys__n45190 & ys__n45522;
  assign new_new_n13164__ = ~ys__n45190 & ~ys__n45522;
  assign new_new_n13165__ = ~ys__n45537 & ~new_new_n13164__;
  assign new_new_n13166__ = ~new_new_n13163__ & new_new_n13165__;
  assign new_new_n13167__ = ys__n45193 & ys__n45524;
  assign new_new_n13168__ = ~ys__n45193 & ~ys__n45524;
  assign new_new_n13169__ = ~ys__n45537 & ~new_new_n13168__;
  assign new_new_n13170__ = ~new_new_n13167__ & new_new_n13169__;
  assign new_new_n13171__ = ~new_new_n13166__ & ~new_new_n13170__;
  assign new_new_n13172__ = new_new_n13162__ & new_new_n13171__;
  assign new_new_n13173__ = new_new_n13153__ & new_new_n13172__;
  assign new_new_n13174__ = new_new_n13134__ & new_new_n13173__;
  assign new_new_n13175__ = ys__n45124 & ys__n45478;
  assign new_new_n13176__ = ~ys__n45124 & ~ys__n45478;
  assign new_new_n13177__ = ~ys__n45534 & ~new_new_n13176__;
  assign new_new_n13178__ = ~new_new_n13175__ & new_new_n13177__;
  assign new_new_n13179__ = ys__n45127 & ys__n45480;
  assign new_new_n13180__ = ~ys__n45127 & ~ys__n45480;
  assign new_new_n13181__ = ~ys__n45534 & ~new_new_n13180__;
  assign new_new_n13182__ = ~new_new_n13179__ & new_new_n13181__;
  assign new_new_n13183__ = ~new_new_n13178__ & ~new_new_n13182__;
  assign new_new_n13184__ = ys__n45130 & ys__n45482;
  assign new_new_n13185__ = ~ys__n45130 & ~ys__n45482;
  assign new_new_n13186__ = ~ys__n45534 & ~new_new_n13185__;
  assign new_new_n13187__ = ~new_new_n13184__ & new_new_n13186__;
  assign new_new_n13188__ = ys__n45133 & ys__n45484;
  assign new_new_n13189__ = ~ys__n45133 & ~ys__n45484;
  assign new_new_n13190__ = ~ys__n45534 & ~new_new_n13189__;
  assign new_new_n13191__ = ~new_new_n13188__ & new_new_n13190__;
  assign new_new_n13192__ = ~new_new_n13187__ & ~new_new_n13191__;
  assign new_new_n13193__ = new_new_n13183__ & new_new_n13192__;
  assign new_new_n13194__ = ys__n45112 & ys__n45470;
  assign new_new_n13195__ = ~ys__n45112 & ~ys__n45470;
  assign new_new_n13196__ = ~ys__n45534 & ~new_new_n13195__;
  assign new_new_n13197__ = ~new_new_n13194__ & new_new_n13196__;
  assign new_new_n13198__ = ys__n45115 & ys__n45472;
  assign new_new_n13199__ = ~ys__n45115 & ~ys__n45472;
  assign new_new_n13200__ = ~ys__n45534 & ~new_new_n13199__;
  assign new_new_n13201__ = ~new_new_n13198__ & new_new_n13200__;
  assign new_new_n13202__ = ~new_new_n13197__ & ~new_new_n13201__;
  assign new_new_n13203__ = ys__n45118 & ys__n45474;
  assign new_new_n13204__ = ~ys__n45118 & ~ys__n45474;
  assign new_new_n13205__ = ~ys__n45534 & ~new_new_n13204__;
  assign new_new_n13206__ = ~new_new_n13203__ & new_new_n13205__;
  assign new_new_n13207__ = ys__n45121 & ys__n45476;
  assign new_new_n13208__ = ~ys__n45121 & ~ys__n45476;
  assign new_new_n13209__ = ~ys__n45534 & ~new_new_n13208__;
  assign new_new_n13210__ = ~new_new_n13207__ & new_new_n13209__;
  assign new_new_n13211__ = ~new_new_n13206__ & ~new_new_n13210__;
  assign new_new_n13212__ = new_new_n13202__ & new_new_n13211__;
  assign new_new_n13213__ = new_new_n13193__ & new_new_n13212__;
  assign new_new_n13214__ = ys__n45148 & ys__n45494;
  assign new_new_n13215__ = ~ys__n45148 & ~ys__n45494;
  assign new_new_n13216__ = ~ys__n45535 & ~new_new_n13215__;
  assign new_new_n13217__ = ~new_new_n13214__ & new_new_n13216__;
  assign new_new_n13218__ = ys__n45151 & ys__n45496;
  assign new_new_n13219__ = ~ys__n45151 & ~ys__n45496;
  assign new_new_n13220__ = ~ys__n45535 & ~new_new_n13219__;
  assign new_new_n13221__ = ~new_new_n13218__ & new_new_n13220__;
  assign new_new_n13222__ = ~new_new_n13217__ & ~new_new_n13221__;
  assign new_new_n13223__ = ys__n45154 & ys__n45498;
  assign new_new_n13224__ = ~ys__n45154 & ~ys__n45498;
  assign new_new_n13225__ = ~ys__n45535 & ~new_new_n13224__;
  assign new_new_n13226__ = ~new_new_n13223__ & new_new_n13225__;
  assign new_new_n13227__ = ys__n45157 & ys__n45500;
  assign new_new_n13228__ = ~ys__n45157 & ~ys__n45500;
  assign new_new_n13229__ = ~ys__n45535 & ~new_new_n13228__;
  assign new_new_n13230__ = ~new_new_n13227__ & new_new_n13229__;
  assign new_new_n13231__ = ~new_new_n13226__ & ~new_new_n13230__;
  assign new_new_n13232__ = new_new_n13222__ & new_new_n13231__;
  assign new_new_n13233__ = ys__n45136 & ys__n45486;
  assign new_new_n13234__ = ~ys__n45136 & ~ys__n45486;
  assign new_new_n13235__ = ~ys__n45535 & ~new_new_n13234__;
  assign new_new_n13236__ = ~new_new_n13233__ & new_new_n13235__;
  assign new_new_n13237__ = ys__n45139 & ys__n45488;
  assign new_new_n13238__ = ~ys__n45139 & ~ys__n45488;
  assign new_new_n13239__ = ~ys__n45535 & ~new_new_n13238__;
  assign new_new_n13240__ = ~new_new_n13237__ & new_new_n13239__;
  assign new_new_n13241__ = ~new_new_n13236__ & ~new_new_n13240__;
  assign new_new_n13242__ = ys__n45142 & ys__n45490;
  assign new_new_n13243__ = ~ys__n45142 & ~ys__n45490;
  assign new_new_n13244__ = ~ys__n45535 & ~new_new_n13243__;
  assign new_new_n13245__ = ~new_new_n13242__ & new_new_n13244__;
  assign new_new_n13246__ = ys__n45145 & ys__n45492;
  assign new_new_n13247__ = ~ys__n45145 & ~ys__n45492;
  assign new_new_n13248__ = ~ys__n45535 & ~new_new_n13247__;
  assign new_new_n13249__ = ~new_new_n13246__ & new_new_n13248__;
  assign new_new_n13250__ = ~new_new_n13245__ & ~new_new_n13249__;
  assign new_new_n13251__ = new_new_n13241__ & new_new_n13250__;
  assign new_new_n13252__ = new_new_n13232__ & new_new_n13251__;
  assign new_new_n13253__ = new_new_n13213__ & new_new_n13252__;
  assign new_new_n13254__ = new_new_n13174__ & new_new_n13253__;
  assign new_new_n13255__ = new_new_n13095__ & new_new_n13254__;
  assign new_new_n13256__ = ys__n45538 & new_new_n13255__;
  assign new_new_n13257__ = ~new_new_n12946__ & ~new_new_n13256__;
  assign new_new_n13258__ = ys__n45046 & ys__n45252;
  assign new_new_n13259__ = ~ys__n45046 & ~ys__n45252;
  assign new_new_n13260__ = ~ys__n45294 & ~new_new_n13259__;
  assign new_new_n13261__ = ~new_new_n13258__ & new_new_n13260__;
  assign new_new_n13262__ = ys__n45049 & ys__n45254;
  assign new_new_n13263__ = ~ys__n45049 & ~ys__n45254;
  assign new_new_n13264__ = ~ys__n45295 & ~new_new_n13263__;
  assign new_new_n13265__ = ~new_new_n13262__ & new_new_n13264__;
  assign new_new_n13266__ = ~new_new_n13261__ & ~new_new_n13265__;
  assign new_new_n13267__ = ys__n45052 & ys__n45256;
  assign new_new_n13268__ = ~ys__n45052 & ~ys__n45256;
  assign new_new_n13269__ = ~ys__n45296 & ~new_new_n13268__;
  assign new_new_n13270__ = ~new_new_n13267__ & new_new_n13269__;
  assign new_new_n13271__ = ys__n45055 & ys__n45258;
  assign new_new_n13272__ = ~ys__n45055 & ~ys__n45258;
  assign new_new_n13273__ = ~ys__n45297 & ~new_new_n13272__;
  assign new_new_n13274__ = ~new_new_n13271__ & new_new_n13273__;
  assign new_new_n13275__ = ~new_new_n13270__ & ~new_new_n13274__;
  assign new_new_n13276__ = new_new_n13266__ & new_new_n13275__;
  assign new_new_n13277__ = ys__n45034 & ys__n45244;
  assign new_new_n13278__ = ~ys__n45034 & ~ys__n45244;
  assign new_new_n13279__ = ~ys__n45290 & ~new_new_n13278__;
  assign new_new_n13280__ = ~new_new_n13277__ & new_new_n13279__;
  assign new_new_n13281__ = ys__n45037 & ys__n45246;
  assign new_new_n13282__ = ~ys__n45037 & ~ys__n45246;
  assign new_new_n13283__ = ~ys__n45291 & ~new_new_n13282__;
  assign new_new_n13284__ = ~new_new_n13281__ & new_new_n13283__;
  assign new_new_n13285__ = ~new_new_n13280__ & ~new_new_n13284__;
  assign new_new_n13286__ = ys__n45040 & ys__n45248;
  assign new_new_n13287__ = ~ys__n45040 & ~ys__n45248;
  assign new_new_n13288__ = ~ys__n45292 & ~new_new_n13287__;
  assign new_new_n13289__ = ~new_new_n13286__ & new_new_n13288__;
  assign new_new_n13290__ = ys__n45043 & ys__n45250;
  assign new_new_n13291__ = ~ys__n45043 & ~ys__n45250;
  assign new_new_n13292__ = ~ys__n45293 & ~new_new_n13291__;
  assign new_new_n13293__ = ~new_new_n13290__ & new_new_n13292__;
  assign new_new_n13294__ = ~new_new_n13289__ & ~new_new_n13293__;
  assign new_new_n13295__ = new_new_n13285__ & new_new_n13294__;
  assign new_new_n13296__ = new_new_n13276__ & new_new_n13295__;
  assign new_new_n13297__ = ys__n45070 & ys__n45268;
  assign new_new_n13298__ = ~ys__n45070 & ~ys__n45268;
  assign new_new_n13299__ = ~ys__n45302 & ~new_new_n13298__;
  assign new_new_n13300__ = ~new_new_n13297__ & new_new_n13299__;
  assign new_new_n13301__ = ys__n45073 & ys__n45270;
  assign new_new_n13302__ = ~ys__n45073 & ~ys__n45270;
  assign new_new_n13303__ = ~ys__n45303 & ~new_new_n13302__;
  assign new_new_n13304__ = ~new_new_n13301__ & new_new_n13303__;
  assign new_new_n13305__ = ~new_new_n13300__ & ~new_new_n13304__;
  assign new_new_n13306__ = ys__n45076 & ys__n45272;
  assign new_new_n13307__ = ~ys__n45076 & ~ys__n45272;
  assign new_new_n13308__ = ~ys__n45304 & ~new_new_n13307__;
  assign new_new_n13309__ = ~new_new_n13306__ & new_new_n13308__;
  assign new_new_n13310__ = ys__n45079 & ys__n45274;
  assign new_new_n13311__ = ~ys__n45079 & ~ys__n45274;
  assign new_new_n13312__ = ~ys__n45305 & ~new_new_n13311__;
  assign new_new_n13313__ = ~new_new_n13310__ & new_new_n13312__;
  assign new_new_n13314__ = ~new_new_n13309__ & ~new_new_n13313__;
  assign new_new_n13315__ = new_new_n13305__ & new_new_n13314__;
  assign new_new_n13316__ = ys__n45058 & ys__n45260;
  assign new_new_n13317__ = ~ys__n45058 & ~ys__n45260;
  assign new_new_n13318__ = ~ys__n45298 & ~new_new_n13317__;
  assign new_new_n13319__ = ~new_new_n13316__ & new_new_n13318__;
  assign new_new_n13320__ = ys__n45061 & ys__n45262;
  assign new_new_n13321__ = ~ys__n45061 & ~ys__n45262;
  assign new_new_n13322__ = ~ys__n45299 & ~new_new_n13321__;
  assign new_new_n13323__ = ~new_new_n13320__ & new_new_n13322__;
  assign new_new_n13324__ = ~new_new_n13319__ & ~new_new_n13323__;
  assign new_new_n13325__ = ys__n45064 & ys__n45264;
  assign new_new_n13326__ = ~ys__n45064 & ~ys__n45264;
  assign new_new_n13327__ = ~ys__n45300 & ~new_new_n13326__;
  assign new_new_n13328__ = ~new_new_n13325__ & new_new_n13327__;
  assign new_new_n13329__ = ys__n45067 & ys__n45266;
  assign new_new_n13330__ = ~ys__n45067 & ~ys__n45266;
  assign new_new_n13331__ = ~ys__n45301 & ~new_new_n13330__;
  assign new_new_n13332__ = ~new_new_n13329__ & new_new_n13331__;
  assign new_new_n13333__ = ~new_new_n13328__ & ~new_new_n13332__;
  assign new_new_n13334__ = new_new_n13324__ & new_new_n13333__;
  assign new_new_n13335__ = new_new_n13315__ & new_new_n13334__;
  assign new_new_n13336__ = new_new_n13296__ & new_new_n13335__;
  assign new_new_n13337__ = ys__n44992 & ys__n45216;
  assign new_new_n13338__ = ~ys__n44992 & ~ys__n45216;
  assign new_new_n13339__ = ~ys__n45276 & ~new_new_n13338__;
  assign new_new_n13340__ = ~new_new_n13337__ & new_new_n13339__;
  assign new_new_n13341__ = ys__n44995 & ys__n45218;
  assign new_new_n13342__ = ~ys__n44995 & ~ys__n45218;
  assign new_new_n13343__ = ~ys__n45277 & ~new_new_n13342__;
  assign new_new_n13344__ = ~new_new_n13341__ & new_new_n13343__;
  assign new_new_n13345__ = ~new_new_n13340__ & ~new_new_n13344__;
  assign new_new_n13346__ = ys__n44998 & ys__n45220;
  assign new_new_n13347__ = ~ys__n44998 & ~ys__n45220;
  assign new_new_n13348__ = ~ys__n45278 & ~new_new_n13347__;
  assign new_new_n13349__ = ~new_new_n13346__ & new_new_n13348__;
  assign new_new_n13350__ = ys__n45001 & ys__n45222;
  assign new_new_n13351__ = ~ys__n45001 & ~ys__n45222;
  assign new_new_n13352__ = ~ys__n45279 & ~new_new_n13351__;
  assign new_new_n13353__ = ~new_new_n13350__ & new_new_n13352__;
  assign new_new_n13354__ = ~new_new_n13349__ & ~new_new_n13353__;
  assign new_new_n13355__ = ys__n45004 & ys__n45224;
  assign new_new_n13356__ = ~ys__n45004 & ~ys__n45224;
  assign new_new_n13357__ = ~ys__n45280 & ~new_new_n13356__;
  assign new_new_n13358__ = ~new_new_n13355__ & new_new_n13357__;
  assign new_new_n13359__ = ys__n45007 & ys__n45226;
  assign new_new_n13360__ = ~ys__n45007 & ~ys__n45226;
  assign new_new_n13361__ = ~ys__n45281 & ~new_new_n13360__;
  assign new_new_n13362__ = ~new_new_n13359__ & new_new_n13361__;
  assign new_new_n13363__ = ~new_new_n13358__ & ~new_new_n13362__;
  assign new_new_n13364__ = new_new_n13354__ & new_new_n13363__;
  assign new_new_n13365__ = new_new_n13345__ & new_new_n13364__;
  assign new_new_n13366__ = ys__n45022 & ys__n45236;
  assign new_new_n13367__ = ~ys__n45022 & ~ys__n45236;
  assign new_new_n13368__ = ~ys__n45286 & ~new_new_n13367__;
  assign new_new_n13369__ = ~new_new_n13366__ & new_new_n13368__;
  assign new_new_n13370__ = ys__n45025 & ys__n45238;
  assign new_new_n13371__ = ~ys__n45025 & ~ys__n45238;
  assign new_new_n13372__ = ~ys__n45287 & ~new_new_n13371__;
  assign new_new_n13373__ = ~new_new_n13370__ & new_new_n13372__;
  assign new_new_n13374__ = ~new_new_n13369__ & ~new_new_n13373__;
  assign new_new_n13375__ = ys__n45028 & ys__n45240;
  assign new_new_n13376__ = ~ys__n45028 & ~ys__n45240;
  assign new_new_n13377__ = ~ys__n45288 & ~new_new_n13376__;
  assign new_new_n13378__ = ~new_new_n13375__ & new_new_n13377__;
  assign new_new_n13379__ = ys__n45031 & ys__n45242;
  assign new_new_n13380__ = ~ys__n45031 & ~ys__n45242;
  assign new_new_n13381__ = ~ys__n45289 & ~new_new_n13380__;
  assign new_new_n13382__ = ~new_new_n13379__ & new_new_n13381__;
  assign new_new_n13383__ = ~new_new_n13378__ & ~new_new_n13382__;
  assign new_new_n13384__ = new_new_n13374__ & new_new_n13383__;
  assign new_new_n13385__ = ys__n45010 & ys__n45228;
  assign new_new_n13386__ = ~ys__n45010 & ~ys__n45228;
  assign new_new_n13387__ = ~ys__n45282 & ~new_new_n13386__;
  assign new_new_n13388__ = ~new_new_n13385__ & new_new_n13387__;
  assign new_new_n13389__ = ys__n45013 & ys__n45230;
  assign new_new_n13390__ = ~ys__n45013 & ~ys__n45230;
  assign new_new_n13391__ = ~ys__n45283 & ~new_new_n13390__;
  assign new_new_n13392__ = ~new_new_n13389__ & new_new_n13391__;
  assign new_new_n13393__ = ~new_new_n13388__ & ~new_new_n13392__;
  assign new_new_n13394__ = ys__n45016 & ys__n45232;
  assign new_new_n13395__ = ~ys__n45016 & ~ys__n45232;
  assign new_new_n13396__ = ~ys__n45284 & ~new_new_n13395__;
  assign new_new_n13397__ = ~new_new_n13394__ & new_new_n13396__;
  assign new_new_n13398__ = ys__n45019 & ys__n45234;
  assign new_new_n13399__ = ~ys__n45019 & ~ys__n45234;
  assign new_new_n13400__ = ~ys__n45285 & ~new_new_n13399__;
  assign new_new_n13401__ = ~new_new_n13398__ & new_new_n13400__;
  assign new_new_n13402__ = ~new_new_n13397__ & ~new_new_n13401__;
  assign new_new_n13403__ = new_new_n13393__ & new_new_n13402__;
  assign new_new_n13404__ = new_new_n13384__ & new_new_n13403__;
  assign new_new_n13405__ = new_new_n13365__ & new_new_n13404__;
  assign new_new_n13406__ = new_new_n13336__ & new_new_n13405__;
  assign new_new_n13407__ = ys__n45172 & ys__n45346;
  assign new_new_n13408__ = ~ys__n45172 & ~ys__n45346;
  assign new_new_n13409__ = ~ys__n45372 & ~new_new_n13408__;
  assign new_new_n13410__ = ~new_new_n13407__ & new_new_n13409__;
  assign new_new_n13411__ = ys__n45175 & ys__n45348;
  assign new_new_n13412__ = ~ys__n45175 & ~ys__n45348;
  assign new_new_n13413__ = ~ys__n45372 & ~new_new_n13412__;
  assign new_new_n13414__ = ~new_new_n13411__ & new_new_n13413__;
  assign new_new_n13415__ = ~new_new_n13410__ & ~new_new_n13414__;
  assign new_new_n13416__ = ys__n45178 & ys__n45350;
  assign new_new_n13417__ = ~ys__n45178 & ~ys__n45350;
  assign new_new_n13418__ = ~ys__n45372 & ~new_new_n13417__;
  assign new_new_n13419__ = ~new_new_n13416__ & new_new_n13418__;
  assign new_new_n13420__ = ys__n45181 & ys__n45352;
  assign new_new_n13421__ = ~ys__n45181 & ~ys__n45352;
  assign new_new_n13422__ = ~ys__n45372 & ~new_new_n13421__;
  assign new_new_n13423__ = ~new_new_n13420__ & new_new_n13422__;
  assign new_new_n13424__ = ~new_new_n13419__ & ~new_new_n13423__;
  assign new_new_n13425__ = new_new_n13415__ & new_new_n13424__;
  assign new_new_n13426__ = ys__n45160 & ys__n45338;
  assign new_new_n13427__ = ~ys__n45160 & ~ys__n45338;
  assign new_new_n13428__ = ~ys__n45372 & ~new_new_n13427__;
  assign new_new_n13429__ = ~new_new_n13426__ & new_new_n13428__;
  assign new_new_n13430__ = ys__n45163 & ys__n45340;
  assign new_new_n13431__ = ~ys__n45163 & ~ys__n45340;
  assign new_new_n13432__ = ~ys__n45372 & ~new_new_n13431__;
  assign new_new_n13433__ = ~new_new_n13430__ & new_new_n13432__;
  assign new_new_n13434__ = ~new_new_n13429__ & ~new_new_n13433__;
  assign new_new_n13435__ = ys__n45166 & ys__n45342;
  assign new_new_n13436__ = ~ys__n45166 & ~ys__n45342;
  assign new_new_n13437__ = ~ys__n45372 & ~new_new_n13436__;
  assign new_new_n13438__ = ~new_new_n13435__ & new_new_n13437__;
  assign new_new_n13439__ = ys__n45169 & ys__n45344;
  assign new_new_n13440__ = ~ys__n45169 & ~ys__n45344;
  assign new_new_n13441__ = ~ys__n45372 & ~new_new_n13440__;
  assign new_new_n13442__ = ~new_new_n13439__ & new_new_n13441__;
  assign new_new_n13443__ = ~new_new_n13438__ & ~new_new_n13442__;
  assign new_new_n13444__ = new_new_n13434__ & new_new_n13443__;
  assign new_new_n13445__ = new_new_n13425__ & new_new_n13444__;
  assign new_new_n13446__ = ys__n45196 & ys__n45362;
  assign new_new_n13447__ = ~ys__n45196 & ~ys__n45362;
  assign new_new_n13448__ = ~ys__n45373 & ~new_new_n13447__;
  assign new_new_n13449__ = ~new_new_n13446__ & new_new_n13448__;
  assign new_new_n13450__ = ys__n45199 & ys__n45364;
  assign new_new_n13451__ = ~ys__n45199 & ~ys__n45364;
  assign new_new_n13452__ = ~ys__n45373 & ~new_new_n13451__;
  assign new_new_n13453__ = ~new_new_n13450__ & new_new_n13452__;
  assign new_new_n13454__ = ~new_new_n13449__ & ~new_new_n13453__;
  assign new_new_n13455__ = ys__n45202 & ys__n45366;
  assign new_new_n13456__ = ~ys__n45202 & ~ys__n45366;
  assign new_new_n13457__ = ~ys__n45373 & ~new_new_n13456__;
  assign new_new_n13458__ = ~new_new_n13455__ & new_new_n13457__;
  assign new_new_n13459__ = ys__n45205 & ys__n45368;
  assign new_new_n13460__ = ~ys__n45205 & ~ys__n45368;
  assign new_new_n13461__ = ~ys__n45373 & ~new_new_n13460__;
  assign new_new_n13462__ = ~new_new_n13459__ & new_new_n13461__;
  assign new_new_n13463__ = ~new_new_n13458__ & ~new_new_n13462__;
  assign new_new_n13464__ = new_new_n13454__ & new_new_n13463__;
  assign new_new_n13465__ = ys__n45184 & ys__n45354;
  assign new_new_n13466__ = ~ys__n45184 & ~ys__n45354;
  assign new_new_n13467__ = ~ys__n45373 & ~new_new_n13466__;
  assign new_new_n13468__ = ~new_new_n13465__ & new_new_n13467__;
  assign new_new_n13469__ = ys__n45187 & ys__n45356;
  assign new_new_n13470__ = ~ys__n45187 & ~ys__n45356;
  assign new_new_n13471__ = ~ys__n45373 & ~new_new_n13470__;
  assign new_new_n13472__ = ~new_new_n13469__ & new_new_n13471__;
  assign new_new_n13473__ = ~new_new_n13468__ & ~new_new_n13472__;
  assign new_new_n13474__ = ys__n45190 & ys__n45358;
  assign new_new_n13475__ = ~ys__n45190 & ~ys__n45358;
  assign new_new_n13476__ = ~ys__n45373 & ~new_new_n13475__;
  assign new_new_n13477__ = ~new_new_n13474__ & new_new_n13476__;
  assign new_new_n13478__ = ys__n45193 & ys__n45360;
  assign new_new_n13479__ = ~ys__n45193 & ~ys__n45360;
  assign new_new_n13480__ = ~ys__n45373 & ~new_new_n13479__;
  assign new_new_n13481__ = ~new_new_n13478__ & new_new_n13480__;
  assign new_new_n13482__ = ~new_new_n13477__ & ~new_new_n13481__;
  assign new_new_n13483__ = new_new_n13473__ & new_new_n13482__;
  assign new_new_n13484__ = new_new_n13464__ & new_new_n13483__;
  assign new_new_n13485__ = new_new_n13445__ & new_new_n13484__;
  assign new_new_n13486__ = ys__n45124 & ys__n45314;
  assign new_new_n13487__ = ~ys__n45124 & ~ys__n45314;
  assign new_new_n13488__ = ~ys__n45370 & ~new_new_n13487__;
  assign new_new_n13489__ = ~new_new_n13486__ & new_new_n13488__;
  assign new_new_n13490__ = ys__n45127 & ys__n45316;
  assign new_new_n13491__ = ~ys__n45127 & ~ys__n45316;
  assign new_new_n13492__ = ~ys__n45370 & ~new_new_n13491__;
  assign new_new_n13493__ = ~new_new_n13490__ & new_new_n13492__;
  assign new_new_n13494__ = ~new_new_n13489__ & ~new_new_n13493__;
  assign new_new_n13495__ = ys__n45130 & ys__n45318;
  assign new_new_n13496__ = ~ys__n45130 & ~ys__n45318;
  assign new_new_n13497__ = ~ys__n45370 & ~new_new_n13496__;
  assign new_new_n13498__ = ~new_new_n13495__ & new_new_n13497__;
  assign new_new_n13499__ = ys__n45133 & ys__n45320;
  assign new_new_n13500__ = ~ys__n45133 & ~ys__n45320;
  assign new_new_n13501__ = ~ys__n45370 & ~new_new_n13500__;
  assign new_new_n13502__ = ~new_new_n13499__ & new_new_n13501__;
  assign new_new_n13503__ = ~new_new_n13498__ & ~new_new_n13502__;
  assign new_new_n13504__ = new_new_n13494__ & new_new_n13503__;
  assign new_new_n13505__ = ys__n45112 & ys__n45306;
  assign new_new_n13506__ = ~ys__n45112 & ~ys__n45306;
  assign new_new_n13507__ = ~ys__n45370 & ~new_new_n13506__;
  assign new_new_n13508__ = ~new_new_n13505__ & new_new_n13507__;
  assign new_new_n13509__ = ys__n45115 & ys__n45308;
  assign new_new_n13510__ = ~ys__n45115 & ~ys__n45308;
  assign new_new_n13511__ = ~ys__n45370 & ~new_new_n13510__;
  assign new_new_n13512__ = ~new_new_n13509__ & new_new_n13511__;
  assign new_new_n13513__ = ~new_new_n13508__ & ~new_new_n13512__;
  assign new_new_n13514__ = ys__n45118 & ys__n45310;
  assign new_new_n13515__ = ~ys__n45118 & ~ys__n45310;
  assign new_new_n13516__ = ~ys__n45370 & ~new_new_n13515__;
  assign new_new_n13517__ = ~new_new_n13514__ & new_new_n13516__;
  assign new_new_n13518__ = ys__n45121 & ys__n45312;
  assign new_new_n13519__ = ~ys__n45121 & ~ys__n45312;
  assign new_new_n13520__ = ~ys__n45370 & ~new_new_n13519__;
  assign new_new_n13521__ = ~new_new_n13518__ & new_new_n13520__;
  assign new_new_n13522__ = ~new_new_n13517__ & ~new_new_n13521__;
  assign new_new_n13523__ = new_new_n13513__ & new_new_n13522__;
  assign new_new_n13524__ = new_new_n13504__ & new_new_n13523__;
  assign new_new_n13525__ = ys__n45148 & ys__n45330;
  assign new_new_n13526__ = ~ys__n45148 & ~ys__n45330;
  assign new_new_n13527__ = ~ys__n45371 & ~new_new_n13526__;
  assign new_new_n13528__ = ~new_new_n13525__ & new_new_n13527__;
  assign new_new_n13529__ = ys__n45151 & ys__n45332;
  assign new_new_n13530__ = ~ys__n45151 & ~ys__n45332;
  assign new_new_n13531__ = ~ys__n45371 & ~new_new_n13530__;
  assign new_new_n13532__ = ~new_new_n13529__ & new_new_n13531__;
  assign new_new_n13533__ = ~new_new_n13528__ & ~new_new_n13532__;
  assign new_new_n13534__ = ys__n45154 & ys__n45334;
  assign new_new_n13535__ = ~ys__n45154 & ~ys__n45334;
  assign new_new_n13536__ = ~ys__n45371 & ~new_new_n13535__;
  assign new_new_n13537__ = ~new_new_n13534__ & new_new_n13536__;
  assign new_new_n13538__ = ys__n45157 & ys__n45336;
  assign new_new_n13539__ = ~ys__n45157 & ~ys__n45336;
  assign new_new_n13540__ = ~ys__n45371 & ~new_new_n13539__;
  assign new_new_n13541__ = ~new_new_n13538__ & new_new_n13540__;
  assign new_new_n13542__ = ~new_new_n13537__ & ~new_new_n13541__;
  assign new_new_n13543__ = new_new_n13533__ & new_new_n13542__;
  assign new_new_n13544__ = ys__n45136 & ys__n45322;
  assign new_new_n13545__ = ~ys__n45136 & ~ys__n45322;
  assign new_new_n13546__ = ~ys__n45371 & ~new_new_n13545__;
  assign new_new_n13547__ = ~new_new_n13544__ & new_new_n13546__;
  assign new_new_n13548__ = ys__n45139 & ys__n45324;
  assign new_new_n13549__ = ~ys__n45139 & ~ys__n45324;
  assign new_new_n13550__ = ~ys__n45371 & ~new_new_n13549__;
  assign new_new_n13551__ = ~new_new_n13548__ & new_new_n13550__;
  assign new_new_n13552__ = ~new_new_n13547__ & ~new_new_n13551__;
  assign new_new_n13553__ = ys__n45142 & ys__n45326;
  assign new_new_n13554__ = ~ys__n45142 & ~ys__n45326;
  assign new_new_n13555__ = ~ys__n45371 & ~new_new_n13554__;
  assign new_new_n13556__ = ~new_new_n13553__ & new_new_n13555__;
  assign new_new_n13557__ = ys__n45145 & ys__n45328;
  assign new_new_n13558__ = ~ys__n45145 & ~ys__n45328;
  assign new_new_n13559__ = ~ys__n45371 & ~new_new_n13558__;
  assign new_new_n13560__ = ~new_new_n13557__ & new_new_n13559__;
  assign new_new_n13561__ = ~new_new_n13556__ & ~new_new_n13560__;
  assign new_new_n13562__ = new_new_n13552__ & new_new_n13561__;
  assign new_new_n13563__ = new_new_n13543__ & new_new_n13562__;
  assign new_new_n13564__ = new_new_n13524__ & new_new_n13563__;
  assign new_new_n13565__ = new_new_n13485__ & new_new_n13564__;
  assign new_new_n13566__ = new_new_n13406__ & new_new_n13565__;
  assign new_new_n13567__ = ys__n45374 & new_new_n13566__;
  assign new_new_n13568__ = ys__n45046 & ys__n45047;
  assign new_new_n13569__ = ~ys__n45046 & ~ys__n45047;
  assign new_new_n13570__ = ~ys__n45100 & ~new_new_n13569__;
  assign new_new_n13571__ = ~new_new_n13568__ & new_new_n13570__;
  assign new_new_n13572__ = ys__n45049 & ys__n45050;
  assign new_new_n13573__ = ~ys__n45049 & ~ys__n45050;
  assign new_new_n13574__ = ~ys__n45101 & ~new_new_n13573__;
  assign new_new_n13575__ = ~new_new_n13572__ & new_new_n13574__;
  assign new_new_n13576__ = ~new_new_n13571__ & ~new_new_n13575__;
  assign new_new_n13577__ = ys__n45052 & ys__n45053;
  assign new_new_n13578__ = ~ys__n45052 & ~ys__n45053;
  assign new_new_n13579__ = ~ys__n45102 & ~new_new_n13578__;
  assign new_new_n13580__ = ~new_new_n13577__ & new_new_n13579__;
  assign new_new_n13581__ = ys__n45055 & ys__n45056;
  assign new_new_n13582__ = ~ys__n45055 & ~ys__n45056;
  assign new_new_n13583__ = ~ys__n45103 & ~new_new_n13582__;
  assign new_new_n13584__ = ~new_new_n13581__ & new_new_n13583__;
  assign new_new_n13585__ = ~new_new_n13580__ & ~new_new_n13584__;
  assign new_new_n13586__ = new_new_n13576__ & new_new_n13585__;
  assign new_new_n13587__ = ys__n45034 & ys__n45035;
  assign new_new_n13588__ = ~ys__n45034 & ~ys__n45035;
  assign new_new_n13589__ = ~ys__n45096 & ~new_new_n13588__;
  assign new_new_n13590__ = ~new_new_n13587__ & new_new_n13589__;
  assign new_new_n13591__ = ys__n45037 & ys__n45038;
  assign new_new_n13592__ = ~ys__n45037 & ~ys__n45038;
  assign new_new_n13593__ = ~ys__n45097 & ~new_new_n13592__;
  assign new_new_n13594__ = ~new_new_n13591__ & new_new_n13593__;
  assign new_new_n13595__ = ~new_new_n13590__ & ~new_new_n13594__;
  assign new_new_n13596__ = ys__n45040 & ys__n45041;
  assign new_new_n13597__ = ~ys__n45040 & ~ys__n45041;
  assign new_new_n13598__ = ~ys__n45098 & ~new_new_n13597__;
  assign new_new_n13599__ = ~new_new_n13596__ & new_new_n13598__;
  assign new_new_n13600__ = ys__n45043 & ys__n45044;
  assign new_new_n13601__ = ~ys__n45043 & ~ys__n45044;
  assign new_new_n13602__ = ~ys__n45099 & ~new_new_n13601__;
  assign new_new_n13603__ = ~new_new_n13600__ & new_new_n13602__;
  assign new_new_n13604__ = ~new_new_n13599__ & ~new_new_n13603__;
  assign new_new_n13605__ = new_new_n13595__ & new_new_n13604__;
  assign new_new_n13606__ = new_new_n13586__ & new_new_n13605__;
  assign new_new_n13607__ = ys__n45070 & ys__n45071;
  assign new_new_n13608__ = ~ys__n45070 & ~ys__n45071;
  assign new_new_n13609__ = ~ys__n45108 & ~new_new_n13608__;
  assign new_new_n13610__ = ~new_new_n13607__ & new_new_n13609__;
  assign new_new_n13611__ = ys__n45073 & ys__n45074;
  assign new_new_n13612__ = ~ys__n45073 & ~ys__n45074;
  assign new_new_n13613__ = ~ys__n45109 & ~new_new_n13612__;
  assign new_new_n13614__ = ~new_new_n13611__ & new_new_n13613__;
  assign new_new_n13615__ = ~new_new_n13610__ & ~new_new_n13614__;
  assign new_new_n13616__ = ys__n45076 & ys__n45077;
  assign new_new_n13617__ = ~ys__n45076 & ~ys__n45077;
  assign new_new_n13618__ = ~ys__n45110 & ~new_new_n13617__;
  assign new_new_n13619__ = ~new_new_n13616__ & new_new_n13618__;
  assign new_new_n13620__ = ys__n45079 & ys__n45080;
  assign new_new_n13621__ = ~ys__n45079 & ~ys__n45080;
  assign new_new_n13622__ = ~ys__n45111 & ~new_new_n13621__;
  assign new_new_n13623__ = ~new_new_n13620__ & new_new_n13622__;
  assign new_new_n13624__ = ~new_new_n13619__ & ~new_new_n13623__;
  assign new_new_n13625__ = new_new_n13615__ & new_new_n13624__;
  assign new_new_n13626__ = ys__n45058 & ys__n45059;
  assign new_new_n13627__ = ~ys__n45058 & ~ys__n45059;
  assign new_new_n13628__ = ~ys__n45104 & ~new_new_n13627__;
  assign new_new_n13629__ = ~new_new_n13626__ & new_new_n13628__;
  assign new_new_n13630__ = ys__n45061 & ys__n45062;
  assign new_new_n13631__ = ~ys__n45061 & ~ys__n45062;
  assign new_new_n13632__ = ~ys__n45105 & ~new_new_n13631__;
  assign new_new_n13633__ = ~new_new_n13630__ & new_new_n13632__;
  assign new_new_n13634__ = ~new_new_n13629__ & ~new_new_n13633__;
  assign new_new_n13635__ = ys__n45064 & ys__n45065;
  assign new_new_n13636__ = ~ys__n45064 & ~ys__n45065;
  assign new_new_n13637__ = ~ys__n45106 & ~new_new_n13636__;
  assign new_new_n13638__ = ~new_new_n13635__ & new_new_n13637__;
  assign new_new_n13639__ = ys__n45067 & ys__n45068;
  assign new_new_n13640__ = ~ys__n45067 & ~ys__n45068;
  assign new_new_n13641__ = ~ys__n45107 & ~new_new_n13640__;
  assign new_new_n13642__ = ~new_new_n13639__ & new_new_n13641__;
  assign new_new_n13643__ = ~new_new_n13638__ & ~new_new_n13642__;
  assign new_new_n13644__ = new_new_n13634__ & new_new_n13643__;
  assign new_new_n13645__ = new_new_n13625__ & new_new_n13644__;
  assign new_new_n13646__ = new_new_n13606__ & new_new_n13645__;
  assign new_new_n13647__ = ys__n44992 & ys__n44993;
  assign new_new_n13648__ = ~ys__n44992 & ~ys__n44993;
  assign new_new_n13649__ = ~ys__n45082 & ~new_new_n13648__;
  assign new_new_n13650__ = ~new_new_n13647__ & new_new_n13649__;
  assign new_new_n13651__ = ys__n44995 & ys__n44996;
  assign new_new_n13652__ = ~ys__n44995 & ~ys__n44996;
  assign new_new_n13653__ = ~ys__n45083 & ~new_new_n13652__;
  assign new_new_n13654__ = ~new_new_n13651__ & new_new_n13653__;
  assign new_new_n13655__ = ~new_new_n13650__ & ~new_new_n13654__;
  assign new_new_n13656__ = ys__n44998 & ys__n44999;
  assign new_new_n13657__ = ~ys__n44998 & ~ys__n44999;
  assign new_new_n13658__ = ~ys__n45084 & ~new_new_n13657__;
  assign new_new_n13659__ = ~new_new_n13656__ & new_new_n13658__;
  assign new_new_n13660__ = ys__n45001 & ys__n45002;
  assign new_new_n13661__ = ~ys__n45001 & ~ys__n45002;
  assign new_new_n13662__ = ~ys__n45085 & ~new_new_n13661__;
  assign new_new_n13663__ = ~new_new_n13660__ & new_new_n13662__;
  assign new_new_n13664__ = ~new_new_n13659__ & ~new_new_n13663__;
  assign new_new_n13665__ = ys__n45004 & ys__n45005;
  assign new_new_n13666__ = ~ys__n45004 & ~ys__n45005;
  assign new_new_n13667__ = ~ys__n45086 & ~new_new_n13666__;
  assign new_new_n13668__ = ~new_new_n13665__ & new_new_n13667__;
  assign new_new_n13669__ = ys__n45007 & ys__n45008;
  assign new_new_n13670__ = ~ys__n45007 & ~ys__n45008;
  assign new_new_n13671__ = ~ys__n45087 & ~new_new_n13670__;
  assign new_new_n13672__ = ~new_new_n13669__ & new_new_n13671__;
  assign new_new_n13673__ = ~new_new_n13668__ & ~new_new_n13672__;
  assign new_new_n13674__ = new_new_n13664__ & new_new_n13673__;
  assign new_new_n13675__ = new_new_n13655__ & new_new_n13674__;
  assign new_new_n13676__ = ys__n45022 & ys__n45023;
  assign new_new_n13677__ = ~ys__n45022 & ~ys__n45023;
  assign new_new_n13678__ = ~ys__n45092 & ~new_new_n13677__;
  assign new_new_n13679__ = ~new_new_n13676__ & new_new_n13678__;
  assign new_new_n13680__ = ys__n45025 & ys__n45026;
  assign new_new_n13681__ = ~ys__n45025 & ~ys__n45026;
  assign new_new_n13682__ = ~ys__n45093 & ~new_new_n13681__;
  assign new_new_n13683__ = ~new_new_n13680__ & new_new_n13682__;
  assign new_new_n13684__ = ~new_new_n13679__ & ~new_new_n13683__;
  assign new_new_n13685__ = ys__n45028 & ys__n45029;
  assign new_new_n13686__ = ~ys__n45028 & ~ys__n45029;
  assign new_new_n13687__ = ~ys__n45094 & ~new_new_n13686__;
  assign new_new_n13688__ = ~new_new_n13685__ & new_new_n13687__;
  assign new_new_n13689__ = ys__n45031 & ys__n45032;
  assign new_new_n13690__ = ~ys__n45031 & ~ys__n45032;
  assign new_new_n13691__ = ~ys__n45095 & ~new_new_n13690__;
  assign new_new_n13692__ = ~new_new_n13689__ & new_new_n13691__;
  assign new_new_n13693__ = ~new_new_n13688__ & ~new_new_n13692__;
  assign new_new_n13694__ = new_new_n13684__ & new_new_n13693__;
  assign new_new_n13695__ = ys__n45010 & ys__n45011;
  assign new_new_n13696__ = ~ys__n45010 & ~ys__n45011;
  assign new_new_n13697__ = ~ys__n45088 & ~new_new_n13696__;
  assign new_new_n13698__ = ~new_new_n13695__ & new_new_n13697__;
  assign new_new_n13699__ = ys__n45013 & ys__n45014;
  assign new_new_n13700__ = ~ys__n45013 & ~ys__n45014;
  assign new_new_n13701__ = ~ys__n45089 & ~new_new_n13700__;
  assign new_new_n13702__ = ~new_new_n13699__ & new_new_n13701__;
  assign new_new_n13703__ = ~new_new_n13698__ & ~new_new_n13702__;
  assign new_new_n13704__ = ys__n45016 & ys__n45017;
  assign new_new_n13705__ = ~ys__n45016 & ~ys__n45017;
  assign new_new_n13706__ = ~ys__n45090 & ~new_new_n13705__;
  assign new_new_n13707__ = ~new_new_n13704__ & new_new_n13706__;
  assign new_new_n13708__ = ys__n45019 & ys__n45020;
  assign new_new_n13709__ = ~ys__n45019 & ~ys__n45020;
  assign new_new_n13710__ = ~ys__n45091 & ~new_new_n13709__;
  assign new_new_n13711__ = ~new_new_n13708__ & new_new_n13710__;
  assign new_new_n13712__ = ~new_new_n13707__ & ~new_new_n13711__;
  assign new_new_n13713__ = new_new_n13703__ & new_new_n13712__;
  assign new_new_n13714__ = new_new_n13694__ & new_new_n13713__;
  assign new_new_n13715__ = new_new_n13675__ & new_new_n13714__;
  assign new_new_n13716__ = new_new_n13646__ & new_new_n13715__;
  assign new_new_n13717__ = ys__n45172 & ys__n45173;
  assign new_new_n13718__ = ~ys__n45172 & ~ys__n45173;
  assign new_new_n13719__ = ~ys__n45210 & ~new_new_n13718__;
  assign new_new_n13720__ = ~new_new_n13717__ & new_new_n13719__;
  assign new_new_n13721__ = ys__n45175 & ys__n45176;
  assign new_new_n13722__ = ~ys__n45175 & ~ys__n45176;
  assign new_new_n13723__ = ~ys__n45210 & ~new_new_n13722__;
  assign new_new_n13724__ = ~new_new_n13721__ & new_new_n13723__;
  assign new_new_n13725__ = ~new_new_n13720__ & ~new_new_n13724__;
  assign new_new_n13726__ = ys__n45178 & ys__n45179;
  assign new_new_n13727__ = ~ys__n45178 & ~ys__n45179;
  assign new_new_n13728__ = ~ys__n45210 & ~new_new_n13727__;
  assign new_new_n13729__ = ~new_new_n13726__ & new_new_n13728__;
  assign new_new_n13730__ = ys__n45181 & ys__n45182;
  assign new_new_n13731__ = ~ys__n45181 & ~ys__n45182;
  assign new_new_n13732__ = ~ys__n45210 & ~new_new_n13731__;
  assign new_new_n13733__ = ~new_new_n13730__ & new_new_n13732__;
  assign new_new_n13734__ = ~new_new_n13729__ & ~new_new_n13733__;
  assign new_new_n13735__ = new_new_n13725__ & new_new_n13734__;
  assign new_new_n13736__ = ys__n45160 & ys__n45161;
  assign new_new_n13737__ = ~ys__n45160 & ~ys__n45161;
  assign new_new_n13738__ = ~ys__n45210 & ~new_new_n13737__;
  assign new_new_n13739__ = ~new_new_n13736__ & new_new_n13738__;
  assign new_new_n13740__ = ys__n45163 & ys__n45164;
  assign new_new_n13741__ = ~ys__n45163 & ~ys__n45164;
  assign new_new_n13742__ = ~ys__n45210 & ~new_new_n13741__;
  assign new_new_n13743__ = ~new_new_n13740__ & new_new_n13742__;
  assign new_new_n13744__ = ~new_new_n13739__ & ~new_new_n13743__;
  assign new_new_n13745__ = ys__n45166 & ys__n45167;
  assign new_new_n13746__ = ~ys__n45166 & ~ys__n45167;
  assign new_new_n13747__ = ~ys__n45210 & ~new_new_n13746__;
  assign new_new_n13748__ = ~new_new_n13745__ & new_new_n13747__;
  assign new_new_n13749__ = ys__n45169 & ys__n45170;
  assign new_new_n13750__ = ~ys__n45169 & ~ys__n45170;
  assign new_new_n13751__ = ~ys__n45210 & ~new_new_n13750__;
  assign new_new_n13752__ = ~new_new_n13749__ & new_new_n13751__;
  assign new_new_n13753__ = ~new_new_n13748__ & ~new_new_n13752__;
  assign new_new_n13754__ = new_new_n13744__ & new_new_n13753__;
  assign new_new_n13755__ = new_new_n13735__ & new_new_n13754__;
  assign new_new_n13756__ = ys__n45196 & ys__n45197;
  assign new_new_n13757__ = ~ys__n45196 & ~ys__n45197;
  assign new_new_n13758__ = ~ys__n45211 & ~new_new_n13757__;
  assign new_new_n13759__ = ~new_new_n13756__ & new_new_n13758__;
  assign new_new_n13760__ = ys__n45199 & ys__n45200;
  assign new_new_n13761__ = ~ys__n45199 & ~ys__n45200;
  assign new_new_n13762__ = ~ys__n45211 & ~new_new_n13761__;
  assign new_new_n13763__ = ~new_new_n13760__ & new_new_n13762__;
  assign new_new_n13764__ = ~new_new_n13759__ & ~new_new_n13763__;
  assign new_new_n13765__ = ys__n45202 & ys__n45203;
  assign new_new_n13766__ = ~ys__n45202 & ~ys__n45203;
  assign new_new_n13767__ = ~ys__n45211 & ~new_new_n13766__;
  assign new_new_n13768__ = ~new_new_n13765__ & new_new_n13767__;
  assign new_new_n13769__ = ys__n45205 & ys__n45206;
  assign new_new_n13770__ = ~ys__n45205 & ~ys__n45206;
  assign new_new_n13771__ = ~ys__n45211 & ~new_new_n13770__;
  assign new_new_n13772__ = ~new_new_n13769__ & new_new_n13771__;
  assign new_new_n13773__ = ~new_new_n13768__ & ~new_new_n13772__;
  assign new_new_n13774__ = new_new_n13764__ & new_new_n13773__;
  assign new_new_n13775__ = ys__n45184 & ys__n45185;
  assign new_new_n13776__ = ~ys__n45184 & ~ys__n45185;
  assign new_new_n13777__ = ~ys__n45211 & ~new_new_n13776__;
  assign new_new_n13778__ = ~new_new_n13775__ & new_new_n13777__;
  assign new_new_n13779__ = ys__n45187 & ys__n45188;
  assign new_new_n13780__ = ~ys__n45187 & ~ys__n45188;
  assign new_new_n13781__ = ~ys__n45211 & ~new_new_n13780__;
  assign new_new_n13782__ = ~new_new_n13779__ & new_new_n13781__;
  assign new_new_n13783__ = ~new_new_n13778__ & ~new_new_n13782__;
  assign new_new_n13784__ = ys__n45190 & ys__n45191;
  assign new_new_n13785__ = ~ys__n45190 & ~ys__n45191;
  assign new_new_n13786__ = ~ys__n45211 & ~new_new_n13785__;
  assign new_new_n13787__ = ~new_new_n13784__ & new_new_n13786__;
  assign new_new_n13788__ = ys__n45193 & ys__n45194;
  assign new_new_n13789__ = ~ys__n45193 & ~ys__n45194;
  assign new_new_n13790__ = ~ys__n45211 & ~new_new_n13789__;
  assign new_new_n13791__ = ~new_new_n13788__ & new_new_n13790__;
  assign new_new_n13792__ = ~new_new_n13787__ & ~new_new_n13791__;
  assign new_new_n13793__ = new_new_n13783__ & new_new_n13792__;
  assign new_new_n13794__ = new_new_n13774__ & new_new_n13793__;
  assign new_new_n13795__ = new_new_n13755__ & new_new_n13794__;
  assign new_new_n13796__ = ys__n45124 & ys__n45125;
  assign new_new_n13797__ = ~ys__n45124 & ~ys__n45125;
  assign new_new_n13798__ = ~ys__n45208 & ~new_new_n13797__;
  assign new_new_n13799__ = ~new_new_n13796__ & new_new_n13798__;
  assign new_new_n13800__ = ys__n45127 & ys__n45128;
  assign new_new_n13801__ = ~ys__n45127 & ~ys__n45128;
  assign new_new_n13802__ = ~ys__n45208 & ~new_new_n13801__;
  assign new_new_n13803__ = ~new_new_n13800__ & new_new_n13802__;
  assign new_new_n13804__ = ~new_new_n13799__ & ~new_new_n13803__;
  assign new_new_n13805__ = ys__n45130 & ys__n45131;
  assign new_new_n13806__ = ~ys__n45130 & ~ys__n45131;
  assign new_new_n13807__ = ~ys__n45208 & ~new_new_n13806__;
  assign new_new_n13808__ = ~new_new_n13805__ & new_new_n13807__;
  assign new_new_n13809__ = ys__n45133 & ys__n45134;
  assign new_new_n13810__ = ~ys__n45133 & ~ys__n45134;
  assign new_new_n13811__ = ~ys__n45208 & ~new_new_n13810__;
  assign new_new_n13812__ = ~new_new_n13809__ & new_new_n13811__;
  assign new_new_n13813__ = ~new_new_n13808__ & ~new_new_n13812__;
  assign new_new_n13814__ = new_new_n13804__ & new_new_n13813__;
  assign new_new_n13815__ = ys__n45112 & ys__n45113;
  assign new_new_n13816__ = ~ys__n45112 & ~ys__n45113;
  assign new_new_n13817__ = ~ys__n45208 & ~new_new_n13816__;
  assign new_new_n13818__ = ~new_new_n13815__ & new_new_n13817__;
  assign new_new_n13819__ = ys__n45115 & ys__n45116;
  assign new_new_n13820__ = ~ys__n45115 & ~ys__n45116;
  assign new_new_n13821__ = ~ys__n45208 & ~new_new_n13820__;
  assign new_new_n13822__ = ~new_new_n13819__ & new_new_n13821__;
  assign new_new_n13823__ = ~new_new_n13818__ & ~new_new_n13822__;
  assign new_new_n13824__ = ys__n45118 & ys__n45119;
  assign new_new_n13825__ = ~ys__n45118 & ~ys__n45119;
  assign new_new_n13826__ = ~ys__n45208 & ~new_new_n13825__;
  assign new_new_n13827__ = ~new_new_n13824__ & new_new_n13826__;
  assign new_new_n13828__ = ys__n45121 & ys__n45122;
  assign new_new_n13829__ = ~ys__n45121 & ~ys__n45122;
  assign new_new_n13830__ = ~ys__n45208 & ~new_new_n13829__;
  assign new_new_n13831__ = ~new_new_n13828__ & new_new_n13830__;
  assign new_new_n13832__ = ~new_new_n13827__ & ~new_new_n13831__;
  assign new_new_n13833__ = new_new_n13823__ & new_new_n13832__;
  assign new_new_n13834__ = new_new_n13814__ & new_new_n13833__;
  assign new_new_n13835__ = ys__n45148 & ys__n45149;
  assign new_new_n13836__ = ~ys__n45148 & ~ys__n45149;
  assign new_new_n13837__ = ~ys__n45209 & ~new_new_n13836__;
  assign new_new_n13838__ = ~new_new_n13835__ & new_new_n13837__;
  assign new_new_n13839__ = ys__n45151 & ys__n45152;
  assign new_new_n13840__ = ~ys__n45151 & ~ys__n45152;
  assign new_new_n13841__ = ~ys__n45209 & ~new_new_n13840__;
  assign new_new_n13842__ = ~new_new_n13839__ & new_new_n13841__;
  assign new_new_n13843__ = ~new_new_n13838__ & ~new_new_n13842__;
  assign new_new_n13844__ = ys__n45154 & ys__n45155;
  assign new_new_n13845__ = ~ys__n45154 & ~ys__n45155;
  assign new_new_n13846__ = ~ys__n45209 & ~new_new_n13845__;
  assign new_new_n13847__ = ~new_new_n13844__ & new_new_n13846__;
  assign new_new_n13848__ = ys__n45157 & ys__n45158;
  assign new_new_n13849__ = ~ys__n45157 & ~ys__n45158;
  assign new_new_n13850__ = ~ys__n45209 & ~new_new_n13849__;
  assign new_new_n13851__ = ~new_new_n13848__ & new_new_n13850__;
  assign new_new_n13852__ = ~new_new_n13847__ & ~new_new_n13851__;
  assign new_new_n13853__ = new_new_n13843__ & new_new_n13852__;
  assign new_new_n13854__ = ys__n45136 & ys__n45137;
  assign new_new_n13855__ = ~ys__n45136 & ~ys__n45137;
  assign new_new_n13856__ = ~ys__n45209 & ~new_new_n13855__;
  assign new_new_n13857__ = ~new_new_n13854__ & new_new_n13856__;
  assign new_new_n13858__ = ys__n45139 & ys__n45140;
  assign new_new_n13859__ = ~ys__n45139 & ~ys__n45140;
  assign new_new_n13860__ = ~ys__n45209 & ~new_new_n13859__;
  assign new_new_n13861__ = ~new_new_n13858__ & new_new_n13860__;
  assign new_new_n13862__ = ~new_new_n13857__ & ~new_new_n13861__;
  assign new_new_n13863__ = ys__n45142 & ys__n45143;
  assign new_new_n13864__ = ~ys__n45142 & ~ys__n45143;
  assign new_new_n13865__ = ~ys__n45209 & ~new_new_n13864__;
  assign new_new_n13866__ = ~new_new_n13863__ & new_new_n13865__;
  assign new_new_n13867__ = ys__n45145 & ys__n45146;
  assign new_new_n13868__ = ~ys__n45145 & ~ys__n45146;
  assign new_new_n13869__ = ~ys__n45209 & ~new_new_n13868__;
  assign new_new_n13870__ = ~new_new_n13867__ & new_new_n13869__;
  assign new_new_n13871__ = ~new_new_n13866__ & ~new_new_n13870__;
  assign new_new_n13872__ = new_new_n13862__ & new_new_n13871__;
  assign new_new_n13873__ = new_new_n13853__ & new_new_n13872__;
  assign new_new_n13874__ = new_new_n13834__ & new_new_n13873__;
  assign new_new_n13875__ = new_new_n13795__ & new_new_n13874__;
  assign new_new_n13876__ = new_new_n13716__ & new_new_n13875__;
  assign new_new_n13877__ = ys__n45212 & new_new_n13876__;
  assign new_new_n13878__ = ~new_new_n13567__ & ~new_new_n13877__;
  assign new_new_n13879__ = new_new_n13257__ & new_new_n13878__;
  assign new_new_n13880__ = ~ys__n23850 & ~ys__n30214;
  assign new_new_n13881__ = ys__n38906 & new_new_n13880__;
  assign new_new_n13882__ = ~ys__n38902 & ~ys__n38904;
  assign new_new_n13883__ = ~new_new_n13881__ & new_new_n13882__;
  assign new_new_n13884__ = ~new_new_n13879__ & ~new_new_n13883__;
  assign new_new_n13885__ = ~ys__n262 & ~ys__n18101;
  assign new_new_n13886__ = ~ys__n18106 & new_new_n13885__;
  assign new_new_n13887__ = ~ys__n4566 & new_new_n13886__;
  assign new_new_n13888__ = ~ys__n22799 & ys__n38272;
  assign new_new_n13889__ = ys__n22794 & ~ys__n33359;
  assign new_new_n13890__ = ~ys__n33375 & ~ys__n33389;
  assign new_new_n13891__ = new_new_n13889__ & new_new_n13890__;
  assign ys__n33357 = ~new_new_n13888__ & new_new_n13891__;
  assign new_new_n13893__ = ~ys__n33375 & ~ys__n33357;
  assign new_new_n13894__ = ~ys__n33350 & ~ys__n33352;
  assign new_new_n13895__ = new_new_n13893__ & new_new_n13894__;
  assign new_new_n13896__ = ys__n38259 & new_new_n13895__;
  assign new_new_n13897__ = new_new_n13895__ & ~new_new_n13896__;
  assign new_new_n13898__ = ys__n38257 & new_new_n13897__;
  assign new_new_n13899__ = ~ys__n38278 & ~ys__n38279;
  assign new_new_n13900__ = ~ys__n38277 & new_new_n13899__;
  assign new_new_n13901__ = new_new_n13897__ & ~new_new_n13900__;
  assign new_new_n13902__ = ~new_new_n13898__ & new_new_n13901__;
  assign new_new_n13903__ = ys__n33350 & new_new_n13893__;
  assign new_new_n13904__ = ys__n33352 & new_new_n13893__;
  assign new_new_n13905__ = ~ys__n33357 & ~new_new_n13904__;
  assign new_new_n13906__ = ~new_new_n13903__ & new_new_n13905__;
  assign new_new_n13907__ = ~new_new_n13896__ & new_new_n13906__;
  assign new_new_n13908__ = ~new_new_n13898__ & new_new_n13907__;
  assign new_new_n13909__ = ~new_new_n13902__ & new_new_n13908__;
  assign new_new_n13910__ = new_new_n13887__ & ~new_new_n13909__;
  assign new_new_n13911__ = ~ys__n738 & new_new_n13910__;
  assign new_new_n13912__ = ~new_new_n13884__ & new_new_n13911__;
  assign new_new_n13913__ = ys__n38236 & new_new_n13893__;
  assign new_new_n13914__ = ys__n38237 & new_new_n13893__;
  assign new_new_n13915__ = ~new_new_n13913__ & ~new_new_n13914__;
  assign new_new_n13916__ = new_new_n13906__ & new_new_n13915__;
  assign new_new_n13917__ = new_new_n13887__ & ~new_new_n13916__;
  assign new_new_n13918__ = ~ys__n738 & new_new_n13917__;
  assign new_new_n13919__ = new_new_n13884__ & new_new_n13918__;
  assign new_new_n13920__ = ~new_new_n13912__ & ~new_new_n13919__;
  assign new_new_n13921__ = ys__n874 & ~ys__n738;
  assign new_new_n13922__ = new_new_n13896__ & new_new_n13921__;
  assign new_new_n13923__ = ~new_new_n13884__ & new_new_n13922__;
  assign ys__n2491 = ~new_new_n13920__ & new_new_n13923__;
  assign ys__n2535 = ys__n196 & ~ys__n4566;
  assign ys__n2536 = ys__n874 & ys__n2535;
  assign new_new_n13927__ = ~ys__n768 & ~ys__n776;
  assign new_new_n13928__ = ~ys__n778 & ~ys__n4168;
  assign new_new_n13929__ = new_new_n13927__ & new_new_n13928__;
  assign new_new_n13930__ = ~ys__n600 & ~ys__n602;
  assign new_new_n13931__ = ~ys__n604 & ~ys__n698;
  assign new_new_n13932__ = new_new_n13930__ & new_new_n13931__;
  assign new_new_n13933__ = ~ys__n598 & ~ys__n774;
  assign new_new_n13934__ = ~ys__n770 & ~ys__n784;
  assign new_new_n13935__ = new_new_n13933__ & ~new_new_n13934__;
  assign new_new_n13936__ = new_new_n13932__ & new_new_n13935__;
  assign ys__n2582 = new_new_n13929__ & new_new_n13936__;
  assign new_new_n13938__ = new_new_n12242__ & new_new_n12358__;
  assign ys__n2635 = new_new_n12396__ & new_new_n13938__;
  assign new_new_n13940__ = ~ys__n4832 & ~ys__n4833;
  assign new_new_n13941__ = ys__n164 & ~ys__n4826;
  assign new_new_n13942__ = ys__n354 & new_new_n13941__;
  assign ys__n2651 = new_new_n13940__ & new_new_n13942__;
  assign ys__n2653 = ys__n2652 | ys__n2651;
  assign new_new_n13945__ = new_new_n12241__ & new_new_n12358__;
  assign ys__n2655 = new_new_n12396__ & new_new_n13945__;
  assign new_new_n13947__ = new_new_n12241__ & new_new_n12369__;
  assign ys__n2674 = new_new_n12396__ & new_new_n13947__;
  assign ys__n2684 = new_new_n12287__ & new_new_n12411__;
  assign new_new_n13950__ = ~ys__n738 & new_new_n13893__;
  assign new_new_n13951__ = new_new_n13887__ & new_new_n13950__;
  assign ys__n2733 = ~ys__n874 | new_new_n13951__;
  assign ys__n2776 = new_new_n12287__ & new_new_n12375__;
  assign new_new_n13954__ = ys__n38219 & ~ys__n738;
  assign ys__n2778 = ~ys__n4566 & new_new_n13954__;
  assign ys__n2780 = ys__n874 & ys__n2779;
  assign ys__n2782 = ~ys__n740 | new_new_n12210__;
  assign new_new_n13958__ = ~ys__n738 & ~new_new_n13915__;
  assign new_new_n13959__ = ~new_new_n13920__ & new_new_n13958__;
  assign new_new_n13960__ = ~new_new_n13903__ & ~new_new_n13904__;
  assign new_new_n13961__ = ~ys__n738 & ~new_new_n13960__;
  assign new_new_n13962__ = ~new_new_n13920__ & new_new_n13961__;
  assign ys__n2804 = new_new_n13959__ | new_new_n13962__;
  assign new_new_n13964__ = ys__n874 & ~ys__n34959;
  assign ys__n2806 = ys__n740 & new_new_n13964__;
  assign new_new_n13966__ = ~new_new_n11071__ & ~new_new_n11078__;
  assign new_new_n13967__ = new_new_n11078__ & ~new_new_n11708__;
  assign ys__n2845 = ~new_new_n13966__ & ~new_new_n13967__;
  assign new_new_n13969__ = ys__n828 & ~new_new_n11727__;
  assign new_new_n13970__ = ~new_new_n11727__ & ~new_new_n13969__;
  assign new_new_n13971__ = ~new_new_n11731__ & ~new_new_n13970__;
  assign new_new_n13972__ = ys__n826 & new_new_n11731__;
  assign ys__n4603 = new_new_n13971__ | new_new_n13972__;
  assign new_new_n13974__ = ~new_new_n11726__ & ~ys__n4603;
  assign new_new_n13975__ = new_new_n11727__ & ys__n730;
  assign new_new_n13976__ = ~ys__n732 & new_new_n11726__;
  assign new_new_n13977__ = ~new_new_n13975__ & ~new_new_n13976__;
  assign ys__n2855 = ~new_new_n13974__ & new_new_n13977__;
  assign ys__n3024 = new_new_n12287__ & new_new_n12383__;
  assign ys__n3035 = ~ys__n740 | new_new_n12177__;
  assign new_new_n13981__ = ~ys__n452 & ys__n24427;
  assign new_new_n13982__ = ys__n452 & ~ys__n24427;
  assign new_new_n13983__ = ~new_new_n13981__ & ~new_new_n13982__;
  assign new_new_n13984__ = ~ys__n35426 & ys__n38695;
  assign new_new_n13985__ = ys__n35426 & ~ys__n38695;
  assign new_new_n13986__ = ~new_new_n13984__ & ~new_new_n13985__;
  assign new_new_n13987__ = new_new_n13983__ & new_new_n13986__;
  assign new_new_n13988__ = ys__n1098 & ys__n24519;
  assign new_new_n13989__ = new_new_n13987__ & new_new_n13988__;
  assign new_new_n13990__ = ys__n24463 & ys__n24519;
  assign new_new_n13991__ = ~ys__n1110 & ~ys__n1120;
  assign new_new_n13992__ = ~new_new_n13990__ & new_new_n13991__;
  assign ys__n3039 = new_new_n13989__ | ~new_new_n13992__;
  assign ys__n3040 = ~ys__n740 | ys__n3039;
  assign ys__n3051 = new_new_n12287__ & new_new_n12380__;
  assign ys__n3061 = new_new_n12287__ & new_new_n12401__;
  assign ys__n3068 = new_new_n11727__ | new_new_n11731__;
  assign ys__n3083 = new_new_n12287__ & new_new_n12423__;
  assign new_new_n13999__ = ~ys__n164 & ~ys__n354;
  assign new_new_n14000__ = ~ys__n4826 & new_new_n13999__;
  assign new_new_n14001__ = new_new_n13940__ & new_new_n14000__;
  assign new_new_n14002__ = ~ys__n402 & new_new_n14001__;
  assign new_new_n14003__ = ys__n402 & ~ys__n408;
  assign new_new_n14004__ = ~ys__n404 & new_new_n14003__;
  assign ys__n3085 = new_new_n14002__ | ~new_new_n14004__;
  assign new_new_n14006__ = new_new_n12242__ & new_new_n12373__;
  assign ys__n3097 = new_new_n12396__ & new_new_n14006__;
  assign ys__n3106 = new_new_n12287__ & new_new_n12386__;
  assign ys__n3114 = new_new_n12287__ & new_new_n12360__;
  assign ys__n3115 = new_new_n12287__ & new_new_n12420__;
  assign ys__n3121 = new_new_n12287__ & new_new_n12371__;
  assign new_new_n14012__ = ~ys__n46 & ~ys__n340;
  assign new_new_n14013__ = new_new_n12266__ & new_new_n14012__;
  assign new_new_n14014__ = new_new_n12265__ & new_new_n14013__;
  assign new_new_n14015__ = ~ys__n44 & ~ys__n6115;
  assign new_new_n14016__ = new_new_n12246__ & new_new_n14015__;
  assign new_new_n14017__ = ~ys__n6112 & ~ys__n6113;
  assign new_new_n14018__ = ys__n18317 & new_new_n12241__;
  assign new_new_n14019__ = new_new_n14017__ & new_new_n14018__;
  assign new_new_n14020__ = new_new_n14016__ & new_new_n14019__;
  assign new_new_n14021__ = new_new_n14014__ & new_new_n14020__;
  assign new_new_n14022__ = new_new_n12285__ & new_new_n14021__;
  assign ys__n3195 = ~ys__n874 | new_new_n14022__;
  assign new_new_n14024__ = ~ys__n18821 & ~ys__n38090;
  assign new_new_n14025__ = ys__n18821 & ys__n38090;
  assign new_new_n14026__ = ~new_new_n14024__ & ~new_new_n14025__;
  assign new_new_n14027__ = ~ys__n18823 & ~ys__n38091;
  assign new_new_n14028__ = ys__n18823 & ys__n38091;
  assign new_new_n14029__ = ~new_new_n14027__ & ~new_new_n14028__;
  assign new_new_n14030__ = ~new_new_n14026__ & ~new_new_n14029__;
  assign new_new_n14031__ = ~ys__n18825 & ~ys__n38092;
  assign new_new_n14032__ = ys__n18825 & ys__n38092;
  assign new_new_n14033__ = ~new_new_n14031__ & ~new_new_n14032__;
  assign new_new_n14034__ = ~ys__n18827 & ~ys__n38093;
  assign new_new_n14035__ = ys__n18827 & ys__n38093;
  assign new_new_n14036__ = ~new_new_n14034__ & ~new_new_n14035__;
  assign new_new_n14037__ = ~new_new_n14033__ & ~new_new_n14036__;
  assign new_new_n14038__ = new_new_n14030__ & new_new_n14037__;
  assign new_new_n14039__ = ~ys__n18813 & ~ys__n38086;
  assign new_new_n14040__ = ys__n18813 & ys__n38086;
  assign new_new_n14041__ = ~new_new_n14039__ & ~new_new_n14040__;
  assign new_new_n14042__ = ~ys__n18815 & ~ys__n38087;
  assign new_new_n14043__ = ys__n18815 & ys__n38087;
  assign new_new_n14044__ = ~new_new_n14042__ & ~new_new_n14043__;
  assign new_new_n14045__ = ~new_new_n14041__ & ~new_new_n14044__;
  assign new_new_n14046__ = ~ys__n18817 & ~ys__n38088;
  assign new_new_n14047__ = ys__n18817 & ys__n38088;
  assign new_new_n14048__ = ~new_new_n14046__ & ~new_new_n14047__;
  assign new_new_n14049__ = ~ys__n18819 & ~ys__n38089;
  assign new_new_n14050__ = ys__n18819 & ys__n38089;
  assign new_new_n14051__ = ~new_new_n14049__ & ~new_new_n14050__;
  assign new_new_n14052__ = ~new_new_n14048__ & ~new_new_n14051__;
  assign new_new_n14053__ = new_new_n14045__ & new_new_n14052__;
  assign new_new_n14054__ = ~ys__n18805 & ~ys__n38082;
  assign new_new_n14055__ = ys__n18805 & ys__n38082;
  assign new_new_n14056__ = ~new_new_n14054__ & ~new_new_n14055__;
  assign new_new_n14057__ = ~ys__n18807 & ~ys__n38083;
  assign new_new_n14058__ = ys__n18807 & ys__n38083;
  assign new_new_n14059__ = ~new_new_n14057__ & ~new_new_n14058__;
  assign new_new_n14060__ = ~new_new_n14056__ & ~new_new_n14059__;
  assign new_new_n14061__ = ~ys__n18809 & ~ys__n38084;
  assign new_new_n14062__ = ys__n18809 & ys__n38084;
  assign new_new_n14063__ = ~new_new_n14061__ & ~new_new_n14062__;
  assign new_new_n14064__ = ~ys__n18811 & ~ys__n38085;
  assign new_new_n14065__ = ys__n18811 & ys__n38085;
  assign new_new_n14066__ = ~new_new_n14064__ & ~new_new_n14065__;
  assign new_new_n14067__ = ~new_new_n14063__ & ~new_new_n14066__;
  assign new_new_n14068__ = new_new_n14060__ & new_new_n14067__;
  assign new_new_n14069__ = new_new_n14053__ & new_new_n14068__;
  assign new_new_n14070__ = new_new_n14038__ & new_new_n14069__;
  assign new_new_n14071__ = ~ys__n18781 & ~ys__n38070;
  assign new_new_n14072__ = ys__n18781 & ys__n38070;
  assign new_new_n14073__ = ~new_new_n14071__ & ~new_new_n14072__;
  assign new_new_n14074__ = ~ys__n18783 & ~ys__n38071;
  assign new_new_n14075__ = ys__n18783 & ys__n38071;
  assign new_new_n14076__ = ~new_new_n14074__ & ~new_new_n14075__;
  assign new_new_n14077__ = ~new_new_n14073__ & ~new_new_n14076__;
  assign new_new_n14078__ = ~ys__n18785 & ~ys__n38072;
  assign new_new_n14079__ = ys__n18785 & ys__n38072;
  assign new_new_n14080__ = ~new_new_n14078__ & ~new_new_n14079__;
  assign new_new_n14081__ = ~ys__n18787 & ~ys__n38073;
  assign new_new_n14082__ = ys__n18787 & ys__n38073;
  assign new_new_n14083__ = ~new_new_n14081__ & ~new_new_n14082__;
  assign new_new_n14084__ = ~new_new_n14080__ & ~new_new_n14083__;
  assign new_new_n14085__ = new_new_n14077__ & new_new_n14084__;
  assign new_new_n14086__ = ~ys__n18773 & ~ys__n38066;
  assign new_new_n14087__ = ys__n18773 & ys__n38066;
  assign new_new_n14088__ = ~new_new_n14086__ & ~new_new_n14087__;
  assign new_new_n14089__ = ~ys__n18775 & ~ys__n38067;
  assign new_new_n14090__ = ys__n18775 & ys__n38067;
  assign new_new_n14091__ = ~new_new_n14089__ & ~new_new_n14090__;
  assign new_new_n14092__ = ~new_new_n14088__ & ~new_new_n14091__;
  assign new_new_n14093__ = ~ys__n18777 & ~ys__n38068;
  assign new_new_n14094__ = ys__n18777 & ys__n38068;
  assign new_new_n14095__ = ~new_new_n14093__ & ~new_new_n14094__;
  assign new_new_n14096__ = ~ys__n18779 & ~ys__n38069;
  assign new_new_n14097__ = ys__n18779 & ys__n38069;
  assign new_new_n14098__ = ~new_new_n14096__ & ~new_new_n14097__;
  assign new_new_n14099__ = ~new_new_n14095__ & ~new_new_n14098__;
  assign new_new_n14100__ = new_new_n14092__ & new_new_n14099__;
  assign new_new_n14101__ = new_new_n14085__ & new_new_n14100__;
  assign new_new_n14102__ = ~ys__n18797 & ~ys__n38078;
  assign new_new_n14103__ = ys__n18797 & ys__n38078;
  assign new_new_n14104__ = ~new_new_n14102__ & ~new_new_n14103__;
  assign new_new_n14105__ = ~ys__n18799 & ~ys__n38079;
  assign new_new_n14106__ = ys__n18799 & ys__n38079;
  assign new_new_n14107__ = ~new_new_n14105__ & ~new_new_n14106__;
  assign new_new_n14108__ = ~new_new_n14104__ & ~new_new_n14107__;
  assign new_new_n14109__ = ~ys__n18801 & ~ys__n38080;
  assign new_new_n14110__ = ys__n18801 & ys__n38080;
  assign new_new_n14111__ = ~new_new_n14109__ & ~new_new_n14110__;
  assign new_new_n14112__ = ~ys__n18803 & ~ys__n38081;
  assign new_new_n14113__ = ys__n18803 & ys__n38081;
  assign new_new_n14114__ = ~new_new_n14112__ & ~new_new_n14113__;
  assign new_new_n14115__ = ~new_new_n14111__ & ~new_new_n14114__;
  assign new_new_n14116__ = new_new_n14108__ & new_new_n14115__;
  assign new_new_n14117__ = ~ys__n18789 & ~ys__n38074;
  assign new_new_n14118__ = ys__n18789 & ys__n38074;
  assign new_new_n14119__ = ~new_new_n14117__ & ~new_new_n14118__;
  assign new_new_n14120__ = ~ys__n18791 & ~ys__n38075;
  assign new_new_n14121__ = ys__n18791 & ys__n38075;
  assign new_new_n14122__ = ~new_new_n14120__ & ~new_new_n14121__;
  assign new_new_n14123__ = ~new_new_n14119__ & ~new_new_n14122__;
  assign new_new_n14124__ = ~ys__n18793 & ~ys__n38076;
  assign new_new_n14125__ = ys__n18793 & ys__n38076;
  assign new_new_n14126__ = ~new_new_n14124__ & ~new_new_n14125__;
  assign new_new_n14127__ = ~ys__n18795 & ~ys__n38077;
  assign new_new_n14128__ = ys__n18795 & ys__n38077;
  assign new_new_n14129__ = ~new_new_n14127__ & ~new_new_n14128__;
  assign new_new_n14130__ = ~new_new_n14126__ & ~new_new_n14129__;
  assign new_new_n14131__ = new_new_n14123__ & new_new_n14130__;
  assign new_new_n14132__ = new_new_n14116__ & new_new_n14131__;
  assign new_new_n14133__ = new_new_n14101__ & new_new_n14132__;
  assign new_new_n14134__ = new_new_n14070__ & new_new_n14133__;
  assign new_new_n14135__ = ~ys__n37746 & ~new_new_n14134__;
  assign new_new_n14136__ = ys__n836 & ~new_new_n14135__;
  assign new_new_n14137__ = ~ys__n18821 & ~ys__n38062;
  assign new_new_n14138__ = ys__n18821 & ys__n38062;
  assign new_new_n14139__ = ~new_new_n14137__ & ~new_new_n14138__;
  assign new_new_n14140__ = ~ys__n18823 & ~ys__n38063;
  assign new_new_n14141__ = ys__n18823 & ys__n38063;
  assign new_new_n14142__ = ~new_new_n14140__ & ~new_new_n14141__;
  assign new_new_n14143__ = ~new_new_n14139__ & ~new_new_n14142__;
  assign new_new_n14144__ = ~ys__n18825 & ~ys__n38064;
  assign new_new_n14145__ = ys__n18825 & ys__n38064;
  assign new_new_n14146__ = ~new_new_n14144__ & ~new_new_n14145__;
  assign new_new_n14147__ = ~ys__n18827 & ~ys__n38065;
  assign new_new_n14148__ = ys__n18827 & ys__n38065;
  assign new_new_n14149__ = ~new_new_n14147__ & ~new_new_n14148__;
  assign new_new_n14150__ = ~new_new_n14146__ & ~new_new_n14149__;
  assign new_new_n14151__ = new_new_n14143__ & new_new_n14150__;
  assign new_new_n14152__ = ~ys__n18813 & ~ys__n38058;
  assign new_new_n14153__ = ys__n18813 & ys__n38058;
  assign new_new_n14154__ = ~new_new_n14152__ & ~new_new_n14153__;
  assign new_new_n14155__ = ~ys__n18815 & ~ys__n38059;
  assign new_new_n14156__ = ys__n18815 & ys__n38059;
  assign new_new_n14157__ = ~new_new_n14155__ & ~new_new_n14156__;
  assign new_new_n14158__ = ~new_new_n14154__ & ~new_new_n14157__;
  assign new_new_n14159__ = ~ys__n18817 & ~ys__n38060;
  assign new_new_n14160__ = ys__n18817 & ys__n38060;
  assign new_new_n14161__ = ~new_new_n14159__ & ~new_new_n14160__;
  assign new_new_n14162__ = ~ys__n18819 & ~ys__n38061;
  assign new_new_n14163__ = ys__n18819 & ys__n38061;
  assign new_new_n14164__ = ~new_new_n14162__ & ~new_new_n14163__;
  assign new_new_n14165__ = ~new_new_n14161__ & ~new_new_n14164__;
  assign new_new_n14166__ = new_new_n14158__ & new_new_n14165__;
  assign new_new_n14167__ = ~ys__n18805 & ~ys__n38054;
  assign new_new_n14168__ = ys__n18805 & ys__n38054;
  assign new_new_n14169__ = ~new_new_n14167__ & ~new_new_n14168__;
  assign new_new_n14170__ = ~ys__n18807 & ~ys__n38055;
  assign new_new_n14171__ = ys__n18807 & ys__n38055;
  assign new_new_n14172__ = ~new_new_n14170__ & ~new_new_n14171__;
  assign new_new_n14173__ = ~new_new_n14169__ & ~new_new_n14172__;
  assign new_new_n14174__ = ~ys__n18809 & ~ys__n38056;
  assign new_new_n14175__ = ys__n18809 & ys__n38056;
  assign new_new_n14176__ = ~new_new_n14174__ & ~new_new_n14175__;
  assign new_new_n14177__ = ~ys__n18811 & ~ys__n38057;
  assign new_new_n14178__ = ys__n18811 & ys__n38057;
  assign new_new_n14179__ = ~new_new_n14177__ & ~new_new_n14178__;
  assign new_new_n14180__ = ~new_new_n14176__ & ~new_new_n14179__;
  assign new_new_n14181__ = new_new_n14173__ & new_new_n14180__;
  assign new_new_n14182__ = new_new_n14166__ & new_new_n14181__;
  assign new_new_n14183__ = new_new_n14151__ & new_new_n14182__;
  assign new_new_n14184__ = ~ys__n18781 & ~ys__n38042;
  assign new_new_n14185__ = ys__n18781 & ys__n38042;
  assign new_new_n14186__ = ~new_new_n14184__ & ~new_new_n14185__;
  assign new_new_n14187__ = ~ys__n18783 & ~ys__n38043;
  assign new_new_n14188__ = ys__n18783 & ys__n38043;
  assign new_new_n14189__ = ~new_new_n14187__ & ~new_new_n14188__;
  assign new_new_n14190__ = ~new_new_n14186__ & ~new_new_n14189__;
  assign new_new_n14191__ = ~ys__n18785 & ~ys__n38044;
  assign new_new_n14192__ = ys__n18785 & ys__n38044;
  assign new_new_n14193__ = ~new_new_n14191__ & ~new_new_n14192__;
  assign new_new_n14194__ = ~ys__n18787 & ~ys__n38045;
  assign new_new_n14195__ = ys__n18787 & ys__n38045;
  assign new_new_n14196__ = ~new_new_n14194__ & ~new_new_n14195__;
  assign new_new_n14197__ = ~new_new_n14193__ & ~new_new_n14196__;
  assign new_new_n14198__ = new_new_n14190__ & new_new_n14197__;
  assign new_new_n14199__ = ~ys__n18773 & ~ys__n38038;
  assign new_new_n14200__ = ys__n18773 & ys__n38038;
  assign new_new_n14201__ = ~new_new_n14199__ & ~new_new_n14200__;
  assign new_new_n14202__ = ~ys__n18775 & ~ys__n38039;
  assign new_new_n14203__ = ys__n18775 & ys__n38039;
  assign new_new_n14204__ = ~new_new_n14202__ & ~new_new_n14203__;
  assign new_new_n14205__ = ~new_new_n14201__ & ~new_new_n14204__;
  assign new_new_n14206__ = ~ys__n18777 & ~ys__n38040;
  assign new_new_n14207__ = ys__n18777 & ys__n38040;
  assign new_new_n14208__ = ~new_new_n14206__ & ~new_new_n14207__;
  assign new_new_n14209__ = ~ys__n18779 & ~ys__n38041;
  assign new_new_n14210__ = ys__n18779 & ys__n38041;
  assign new_new_n14211__ = ~new_new_n14209__ & ~new_new_n14210__;
  assign new_new_n14212__ = ~new_new_n14208__ & ~new_new_n14211__;
  assign new_new_n14213__ = new_new_n14205__ & new_new_n14212__;
  assign new_new_n14214__ = new_new_n14198__ & new_new_n14213__;
  assign new_new_n14215__ = ~ys__n18797 & ~ys__n38050;
  assign new_new_n14216__ = ys__n18797 & ys__n38050;
  assign new_new_n14217__ = ~new_new_n14215__ & ~new_new_n14216__;
  assign new_new_n14218__ = ~ys__n18799 & ~ys__n38051;
  assign new_new_n14219__ = ys__n18799 & ys__n38051;
  assign new_new_n14220__ = ~new_new_n14218__ & ~new_new_n14219__;
  assign new_new_n14221__ = ~new_new_n14217__ & ~new_new_n14220__;
  assign new_new_n14222__ = ~ys__n18801 & ~ys__n38052;
  assign new_new_n14223__ = ys__n18801 & ys__n38052;
  assign new_new_n14224__ = ~new_new_n14222__ & ~new_new_n14223__;
  assign new_new_n14225__ = ~ys__n18803 & ~ys__n38053;
  assign new_new_n14226__ = ys__n18803 & ys__n38053;
  assign new_new_n14227__ = ~new_new_n14225__ & ~new_new_n14226__;
  assign new_new_n14228__ = ~new_new_n14224__ & ~new_new_n14227__;
  assign new_new_n14229__ = new_new_n14221__ & new_new_n14228__;
  assign new_new_n14230__ = ~ys__n18789 & ~ys__n38046;
  assign new_new_n14231__ = ys__n18789 & ys__n38046;
  assign new_new_n14232__ = ~new_new_n14230__ & ~new_new_n14231__;
  assign new_new_n14233__ = ~ys__n18791 & ~ys__n38047;
  assign new_new_n14234__ = ys__n18791 & ys__n38047;
  assign new_new_n14235__ = ~new_new_n14233__ & ~new_new_n14234__;
  assign new_new_n14236__ = ~new_new_n14232__ & ~new_new_n14235__;
  assign new_new_n14237__ = ~ys__n18793 & ~ys__n38048;
  assign new_new_n14238__ = ys__n18793 & ys__n38048;
  assign new_new_n14239__ = ~new_new_n14237__ & ~new_new_n14238__;
  assign new_new_n14240__ = ~ys__n18795 & ~ys__n38049;
  assign new_new_n14241__ = ys__n18795 & ys__n38049;
  assign new_new_n14242__ = ~new_new_n14240__ & ~new_new_n14241__;
  assign new_new_n14243__ = ~new_new_n14239__ & ~new_new_n14242__;
  assign new_new_n14244__ = new_new_n14236__ & new_new_n14243__;
  assign new_new_n14245__ = new_new_n14229__ & new_new_n14244__;
  assign new_new_n14246__ = new_new_n14214__ & new_new_n14245__;
  assign new_new_n14247__ = new_new_n14183__ & new_new_n14246__;
  assign new_new_n14248__ = ~ys__n37747 & ~new_new_n14247__;
  assign new_new_n14249__ = ys__n834 & ~new_new_n14248__;
  assign new_new_n14250__ = ~new_new_n14136__ & ~new_new_n14249__;
  assign new_new_n14251__ = ~ys__n18821 & ~ys__n38034;
  assign new_new_n14252__ = ys__n18821 & ys__n38034;
  assign new_new_n14253__ = ~new_new_n14251__ & ~new_new_n14252__;
  assign new_new_n14254__ = ~ys__n18823 & ~ys__n38035;
  assign new_new_n14255__ = ys__n18823 & ys__n38035;
  assign new_new_n14256__ = ~new_new_n14254__ & ~new_new_n14255__;
  assign new_new_n14257__ = ~new_new_n14253__ & ~new_new_n14256__;
  assign new_new_n14258__ = ~ys__n18825 & ~ys__n38036;
  assign new_new_n14259__ = ys__n18825 & ys__n38036;
  assign new_new_n14260__ = ~new_new_n14258__ & ~new_new_n14259__;
  assign new_new_n14261__ = ~ys__n18827 & ~ys__n38037;
  assign new_new_n14262__ = ys__n18827 & ys__n38037;
  assign new_new_n14263__ = ~new_new_n14261__ & ~new_new_n14262__;
  assign new_new_n14264__ = ~new_new_n14260__ & ~new_new_n14263__;
  assign new_new_n14265__ = new_new_n14257__ & new_new_n14264__;
  assign new_new_n14266__ = ~ys__n18813 & ~ys__n38030;
  assign new_new_n14267__ = ys__n18813 & ys__n38030;
  assign new_new_n14268__ = ~new_new_n14266__ & ~new_new_n14267__;
  assign new_new_n14269__ = ~ys__n18815 & ~ys__n38031;
  assign new_new_n14270__ = ys__n18815 & ys__n38031;
  assign new_new_n14271__ = ~new_new_n14269__ & ~new_new_n14270__;
  assign new_new_n14272__ = ~new_new_n14268__ & ~new_new_n14271__;
  assign new_new_n14273__ = ~ys__n18817 & ~ys__n38032;
  assign new_new_n14274__ = ys__n18817 & ys__n38032;
  assign new_new_n14275__ = ~new_new_n14273__ & ~new_new_n14274__;
  assign new_new_n14276__ = ~ys__n18819 & ~ys__n38033;
  assign new_new_n14277__ = ys__n18819 & ys__n38033;
  assign new_new_n14278__ = ~new_new_n14276__ & ~new_new_n14277__;
  assign new_new_n14279__ = ~new_new_n14275__ & ~new_new_n14278__;
  assign new_new_n14280__ = new_new_n14272__ & new_new_n14279__;
  assign new_new_n14281__ = ~ys__n18805 & ~ys__n38026;
  assign new_new_n14282__ = ys__n18805 & ys__n38026;
  assign new_new_n14283__ = ~new_new_n14281__ & ~new_new_n14282__;
  assign new_new_n14284__ = ~ys__n18807 & ~ys__n38027;
  assign new_new_n14285__ = ys__n18807 & ys__n38027;
  assign new_new_n14286__ = ~new_new_n14284__ & ~new_new_n14285__;
  assign new_new_n14287__ = ~new_new_n14283__ & ~new_new_n14286__;
  assign new_new_n14288__ = ~ys__n18809 & ~ys__n38028;
  assign new_new_n14289__ = ys__n18809 & ys__n38028;
  assign new_new_n14290__ = ~new_new_n14288__ & ~new_new_n14289__;
  assign new_new_n14291__ = ~ys__n18811 & ~ys__n38029;
  assign new_new_n14292__ = ys__n18811 & ys__n38029;
  assign new_new_n14293__ = ~new_new_n14291__ & ~new_new_n14292__;
  assign new_new_n14294__ = ~new_new_n14290__ & ~new_new_n14293__;
  assign new_new_n14295__ = new_new_n14287__ & new_new_n14294__;
  assign new_new_n14296__ = new_new_n14280__ & new_new_n14295__;
  assign new_new_n14297__ = new_new_n14265__ & new_new_n14296__;
  assign new_new_n14298__ = ~ys__n18781 & ~ys__n38014;
  assign new_new_n14299__ = ys__n18781 & ys__n38014;
  assign new_new_n14300__ = ~new_new_n14298__ & ~new_new_n14299__;
  assign new_new_n14301__ = ~ys__n18783 & ~ys__n38015;
  assign new_new_n14302__ = ys__n18783 & ys__n38015;
  assign new_new_n14303__ = ~new_new_n14301__ & ~new_new_n14302__;
  assign new_new_n14304__ = ~new_new_n14300__ & ~new_new_n14303__;
  assign new_new_n14305__ = ~ys__n18785 & ~ys__n38016;
  assign new_new_n14306__ = ys__n18785 & ys__n38016;
  assign new_new_n14307__ = ~new_new_n14305__ & ~new_new_n14306__;
  assign new_new_n14308__ = ~ys__n18787 & ~ys__n38017;
  assign new_new_n14309__ = ys__n18787 & ys__n38017;
  assign new_new_n14310__ = ~new_new_n14308__ & ~new_new_n14309__;
  assign new_new_n14311__ = ~new_new_n14307__ & ~new_new_n14310__;
  assign new_new_n14312__ = new_new_n14304__ & new_new_n14311__;
  assign new_new_n14313__ = ~ys__n18773 & ~ys__n38010;
  assign new_new_n14314__ = ys__n18773 & ys__n38010;
  assign new_new_n14315__ = ~new_new_n14313__ & ~new_new_n14314__;
  assign new_new_n14316__ = ~ys__n18775 & ~ys__n38011;
  assign new_new_n14317__ = ys__n18775 & ys__n38011;
  assign new_new_n14318__ = ~new_new_n14316__ & ~new_new_n14317__;
  assign new_new_n14319__ = ~new_new_n14315__ & ~new_new_n14318__;
  assign new_new_n14320__ = ~ys__n18777 & ~ys__n38012;
  assign new_new_n14321__ = ys__n18777 & ys__n38012;
  assign new_new_n14322__ = ~new_new_n14320__ & ~new_new_n14321__;
  assign new_new_n14323__ = ~ys__n18779 & ~ys__n38013;
  assign new_new_n14324__ = ys__n18779 & ys__n38013;
  assign new_new_n14325__ = ~new_new_n14323__ & ~new_new_n14324__;
  assign new_new_n14326__ = ~new_new_n14322__ & ~new_new_n14325__;
  assign new_new_n14327__ = new_new_n14319__ & new_new_n14326__;
  assign new_new_n14328__ = new_new_n14312__ & new_new_n14327__;
  assign new_new_n14329__ = ~ys__n18797 & ~ys__n38022;
  assign new_new_n14330__ = ys__n18797 & ys__n38022;
  assign new_new_n14331__ = ~new_new_n14329__ & ~new_new_n14330__;
  assign new_new_n14332__ = ~ys__n18799 & ~ys__n38023;
  assign new_new_n14333__ = ys__n18799 & ys__n38023;
  assign new_new_n14334__ = ~new_new_n14332__ & ~new_new_n14333__;
  assign new_new_n14335__ = ~new_new_n14331__ & ~new_new_n14334__;
  assign new_new_n14336__ = ~ys__n18801 & ~ys__n38024;
  assign new_new_n14337__ = ys__n18801 & ys__n38024;
  assign new_new_n14338__ = ~new_new_n14336__ & ~new_new_n14337__;
  assign new_new_n14339__ = ~ys__n18803 & ~ys__n38025;
  assign new_new_n14340__ = ys__n18803 & ys__n38025;
  assign new_new_n14341__ = ~new_new_n14339__ & ~new_new_n14340__;
  assign new_new_n14342__ = ~new_new_n14338__ & ~new_new_n14341__;
  assign new_new_n14343__ = new_new_n14335__ & new_new_n14342__;
  assign new_new_n14344__ = ~ys__n18789 & ~ys__n38018;
  assign new_new_n14345__ = ys__n18789 & ys__n38018;
  assign new_new_n14346__ = ~new_new_n14344__ & ~new_new_n14345__;
  assign new_new_n14347__ = ~ys__n18791 & ~ys__n38019;
  assign new_new_n14348__ = ys__n18791 & ys__n38019;
  assign new_new_n14349__ = ~new_new_n14347__ & ~new_new_n14348__;
  assign new_new_n14350__ = ~new_new_n14346__ & ~new_new_n14349__;
  assign new_new_n14351__ = ~ys__n18793 & ~ys__n38020;
  assign new_new_n14352__ = ys__n18793 & ys__n38020;
  assign new_new_n14353__ = ~new_new_n14351__ & ~new_new_n14352__;
  assign new_new_n14354__ = ~ys__n18795 & ~ys__n38021;
  assign new_new_n14355__ = ys__n18795 & ys__n38021;
  assign new_new_n14356__ = ~new_new_n14354__ & ~new_new_n14355__;
  assign new_new_n14357__ = ~new_new_n14353__ & ~new_new_n14356__;
  assign new_new_n14358__ = new_new_n14350__ & new_new_n14357__;
  assign new_new_n14359__ = new_new_n14343__ & new_new_n14358__;
  assign new_new_n14360__ = new_new_n14328__ & new_new_n14359__;
  assign new_new_n14361__ = new_new_n14297__ & new_new_n14360__;
  assign new_new_n14362__ = ~ys__n37748 & ~new_new_n14361__;
  assign new_new_n14363__ = ys__n832 & ~new_new_n14362__;
  assign new_new_n14364__ = ~ys__n18821 & ~ys__n38006;
  assign new_new_n14365__ = ys__n18821 & ys__n38006;
  assign new_new_n14366__ = ~new_new_n14364__ & ~new_new_n14365__;
  assign new_new_n14367__ = ~ys__n18823 & ~ys__n38007;
  assign new_new_n14368__ = ys__n18823 & ys__n38007;
  assign new_new_n14369__ = ~new_new_n14367__ & ~new_new_n14368__;
  assign new_new_n14370__ = ~new_new_n14366__ & ~new_new_n14369__;
  assign new_new_n14371__ = ~ys__n18825 & ~ys__n38008;
  assign new_new_n14372__ = ys__n18825 & ys__n38008;
  assign new_new_n14373__ = ~new_new_n14371__ & ~new_new_n14372__;
  assign new_new_n14374__ = ~ys__n18827 & ~ys__n38009;
  assign new_new_n14375__ = ys__n18827 & ys__n38009;
  assign new_new_n14376__ = ~new_new_n14374__ & ~new_new_n14375__;
  assign new_new_n14377__ = ~new_new_n14373__ & ~new_new_n14376__;
  assign new_new_n14378__ = new_new_n14370__ & new_new_n14377__;
  assign new_new_n14379__ = ~ys__n18813 & ~ys__n38002;
  assign new_new_n14380__ = ys__n18813 & ys__n38002;
  assign new_new_n14381__ = ~new_new_n14379__ & ~new_new_n14380__;
  assign new_new_n14382__ = ~ys__n18815 & ~ys__n38003;
  assign new_new_n14383__ = ys__n18815 & ys__n38003;
  assign new_new_n14384__ = ~new_new_n14382__ & ~new_new_n14383__;
  assign new_new_n14385__ = ~new_new_n14381__ & ~new_new_n14384__;
  assign new_new_n14386__ = ~ys__n18817 & ~ys__n38004;
  assign new_new_n14387__ = ys__n18817 & ys__n38004;
  assign new_new_n14388__ = ~new_new_n14386__ & ~new_new_n14387__;
  assign new_new_n14389__ = ~ys__n18819 & ~ys__n38005;
  assign new_new_n14390__ = ys__n18819 & ys__n38005;
  assign new_new_n14391__ = ~new_new_n14389__ & ~new_new_n14390__;
  assign new_new_n14392__ = ~new_new_n14388__ & ~new_new_n14391__;
  assign new_new_n14393__ = new_new_n14385__ & new_new_n14392__;
  assign new_new_n14394__ = ~ys__n18805 & ~ys__n37998;
  assign new_new_n14395__ = ys__n18805 & ys__n37998;
  assign new_new_n14396__ = ~new_new_n14394__ & ~new_new_n14395__;
  assign new_new_n14397__ = ~ys__n18807 & ~ys__n37999;
  assign new_new_n14398__ = ys__n18807 & ys__n37999;
  assign new_new_n14399__ = ~new_new_n14397__ & ~new_new_n14398__;
  assign new_new_n14400__ = ~new_new_n14396__ & ~new_new_n14399__;
  assign new_new_n14401__ = ~ys__n18809 & ~ys__n38000;
  assign new_new_n14402__ = ys__n18809 & ys__n38000;
  assign new_new_n14403__ = ~new_new_n14401__ & ~new_new_n14402__;
  assign new_new_n14404__ = ~ys__n18811 & ~ys__n38001;
  assign new_new_n14405__ = ys__n18811 & ys__n38001;
  assign new_new_n14406__ = ~new_new_n14404__ & ~new_new_n14405__;
  assign new_new_n14407__ = ~new_new_n14403__ & ~new_new_n14406__;
  assign new_new_n14408__ = new_new_n14400__ & new_new_n14407__;
  assign new_new_n14409__ = new_new_n14393__ & new_new_n14408__;
  assign new_new_n14410__ = new_new_n14378__ & new_new_n14409__;
  assign new_new_n14411__ = ~ys__n18781 & ~ys__n37986;
  assign new_new_n14412__ = ys__n18781 & ys__n37986;
  assign new_new_n14413__ = ~new_new_n14411__ & ~new_new_n14412__;
  assign new_new_n14414__ = ~ys__n18783 & ~ys__n37987;
  assign new_new_n14415__ = ys__n18783 & ys__n37987;
  assign new_new_n14416__ = ~new_new_n14414__ & ~new_new_n14415__;
  assign new_new_n14417__ = ~new_new_n14413__ & ~new_new_n14416__;
  assign new_new_n14418__ = ~ys__n18785 & ~ys__n37988;
  assign new_new_n14419__ = ys__n18785 & ys__n37988;
  assign new_new_n14420__ = ~new_new_n14418__ & ~new_new_n14419__;
  assign new_new_n14421__ = ~ys__n18787 & ~ys__n37989;
  assign new_new_n14422__ = ys__n18787 & ys__n37989;
  assign new_new_n14423__ = ~new_new_n14421__ & ~new_new_n14422__;
  assign new_new_n14424__ = ~new_new_n14420__ & ~new_new_n14423__;
  assign new_new_n14425__ = new_new_n14417__ & new_new_n14424__;
  assign new_new_n14426__ = ~ys__n18773 & ~ys__n37982;
  assign new_new_n14427__ = ys__n18773 & ys__n37982;
  assign new_new_n14428__ = ~new_new_n14426__ & ~new_new_n14427__;
  assign new_new_n14429__ = ~ys__n18775 & ~ys__n37983;
  assign new_new_n14430__ = ys__n18775 & ys__n37983;
  assign new_new_n14431__ = ~new_new_n14429__ & ~new_new_n14430__;
  assign new_new_n14432__ = ~new_new_n14428__ & ~new_new_n14431__;
  assign new_new_n14433__ = ~ys__n18777 & ~ys__n37984;
  assign new_new_n14434__ = ys__n18777 & ys__n37984;
  assign new_new_n14435__ = ~new_new_n14433__ & ~new_new_n14434__;
  assign new_new_n14436__ = ~ys__n18779 & ~ys__n37985;
  assign new_new_n14437__ = ys__n18779 & ys__n37985;
  assign new_new_n14438__ = ~new_new_n14436__ & ~new_new_n14437__;
  assign new_new_n14439__ = ~new_new_n14435__ & ~new_new_n14438__;
  assign new_new_n14440__ = new_new_n14432__ & new_new_n14439__;
  assign new_new_n14441__ = new_new_n14425__ & new_new_n14440__;
  assign new_new_n14442__ = ~ys__n18797 & ~ys__n37994;
  assign new_new_n14443__ = ys__n18797 & ys__n37994;
  assign new_new_n14444__ = ~new_new_n14442__ & ~new_new_n14443__;
  assign new_new_n14445__ = ~ys__n18799 & ~ys__n37995;
  assign new_new_n14446__ = ys__n18799 & ys__n37995;
  assign new_new_n14447__ = ~new_new_n14445__ & ~new_new_n14446__;
  assign new_new_n14448__ = ~new_new_n14444__ & ~new_new_n14447__;
  assign new_new_n14449__ = ~ys__n18801 & ~ys__n37996;
  assign new_new_n14450__ = ys__n18801 & ys__n37996;
  assign new_new_n14451__ = ~new_new_n14449__ & ~new_new_n14450__;
  assign new_new_n14452__ = ~ys__n18803 & ~ys__n37997;
  assign new_new_n14453__ = ys__n18803 & ys__n37997;
  assign new_new_n14454__ = ~new_new_n14452__ & ~new_new_n14453__;
  assign new_new_n14455__ = ~new_new_n14451__ & ~new_new_n14454__;
  assign new_new_n14456__ = new_new_n14448__ & new_new_n14455__;
  assign new_new_n14457__ = ~ys__n18789 & ~ys__n37990;
  assign new_new_n14458__ = ys__n18789 & ys__n37990;
  assign new_new_n14459__ = ~new_new_n14457__ & ~new_new_n14458__;
  assign new_new_n14460__ = ~ys__n18791 & ~ys__n37991;
  assign new_new_n14461__ = ys__n18791 & ys__n37991;
  assign new_new_n14462__ = ~new_new_n14460__ & ~new_new_n14461__;
  assign new_new_n14463__ = ~new_new_n14459__ & ~new_new_n14462__;
  assign new_new_n14464__ = ~ys__n18793 & ~ys__n37992;
  assign new_new_n14465__ = ys__n18793 & ys__n37992;
  assign new_new_n14466__ = ~new_new_n14464__ & ~new_new_n14465__;
  assign new_new_n14467__ = ~ys__n18795 & ~ys__n37993;
  assign new_new_n14468__ = ys__n18795 & ys__n37993;
  assign new_new_n14469__ = ~new_new_n14467__ & ~new_new_n14468__;
  assign new_new_n14470__ = ~new_new_n14466__ & ~new_new_n14469__;
  assign new_new_n14471__ = new_new_n14463__ & new_new_n14470__;
  assign new_new_n14472__ = new_new_n14456__ & new_new_n14471__;
  assign new_new_n14473__ = new_new_n14441__ & new_new_n14472__;
  assign new_new_n14474__ = new_new_n14410__ & new_new_n14473__;
  assign new_new_n14475__ = ~ys__n37749 & ~new_new_n14474__;
  assign new_new_n14476__ = ys__n830 & ~new_new_n14475__;
  assign new_new_n14477__ = ~new_new_n14363__ & ~new_new_n14476__;
  assign new_new_n14478__ = new_new_n14250__ & new_new_n14477__;
  assign new_new_n14479__ = ~ys__n18821 & ~ys__n18984;
  assign new_new_n14480__ = ys__n18821 & ys__n18984;
  assign new_new_n14481__ = ~new_new_n14479__ & ~new_new_n14480__;
  assign new_new_n14482__ = ~ys__n18823 & ~ys__n18985;
  assign new_new_n14483__ = ys__n18823 & ys__n18985;
  assign new_new_n14484__ = ~new_new_n14482__ & ~new_new_n14483__;
  assign new_new_n14485__ = ~new_new_n14481__ & ~new_new_n14484__;
  assign new_new_n14486__ = ~ys__n18825 & ~ys__n18986;
  assign new_new_n14487__ = ys__n18825 & ys__n18986;
  assign new_new_n14488__ = ~new_new_n14486__ & ~new_new_n14487__;
  assign new_new_n14489__ = ~ys__n18827 & ~ys__n18987;
  assign new_new_n14490__ = ys__n18827 & ys__n18987;
  assign new_new_n14491__ = ~new_new_n14489__ & ~new_new_n14490__;
  assign new_new_n14492__ = ~new_new_n14488__ & ~new_new_n14491__;
  assign new_new_n14493__ = new_new_n14485__ & new_new_n14492__;
  assign new_new_n14494__ = ~ys__n18813 & ~ys__n18980;
  assign new_new_n14495__ = ys__n18813 & ys__n18980;
  assign new_new_n14496__ = ~new_new_n14494__ & ~new_new_n14495__;
  assign new_new_n14497__ = ~ys__n18815 & ~ys__n18981;
  assign new_new_n14498__ = ys__n18815 & ys__n18981;
  assign new_new_n14499__ = ~new_new_n14497__ & ~new_new_n14498__;
  assign new_new_n14500__ = ~new_new_n14496__ & ~new_new_n14499__;
  assign new_new_n14501__ = ~ys__n18817 & ~ys__n18982;
  assign new_new_n14502__ = ys__n18817 & ys__n18982;
  assign new_new_n14503__ = ~new_new_n14501__ & ~new_new_n14502__;
  assign new_new_n14504__ = ~ys__n18819 & ~ys__n18983;
  assign new_new_n14505__ = ys__n18819 & ys__n18983;
  assign new_new_n14506__ = ~new_new_n14504__ & ~new_new_n14505__;
  assign new_new_n14507__ = ~new_new_n14503__ & ~new_new_n14506__;
  assign new_new_n14508__ = new_new_n14500__ & new_new_n14507__;
  assign new_new_n14509__ = ~ys__n18805 & ~ys__n18976;
  assign new_new_n14510__ = ys__n18805 & ys__n18976;
  assign new_new_n14511__ = ~new_new_n14509__ & ~new_new_n14510__;
  assign new_new_n14512__ = ~ys__n18807 & ~ys__n18977;
  assign new_new_n14513__ = ys__n18807 & ys__n18977;
  assign new_new_n14514__ = ~new_new_n14512__ & ~new_new_n14513__;
  assign new_new_n14515__ = ~new_new_n14511__ & ~new_new_n14514__;
  assign new_new_n14516__ = ~ys__n18809 & ~ys__n18978;
  assign new_new_n14517__ = ys__n18809 & ys__n18978;
  assign new_new_n14518__ = ~new_new_n14516__ & ~new_new_n14517__;
  assign new_new_n14519__ = ~ys__n18811 & ~ys__n18979;
  assign new_new_n14520__ = ys__n18811 & ys__n18979;
  assign new_new_n14521__ = ~new_new_n14519__ & ~new_new_n14520__;
  assign new_new_n14522__ = ~new_new_n14518__ & ~new_new_n14521__;
  assign new_new_n14523__ = new_new_n14515__ & new_new_n14522__;
  assign new_new_n14524__ = new_new_n14508__ & new_new_n14523__;
  assign new_new_n14525__ = new_new_n14493__ & new_new_n14524__;
  assign new_new_n14526__ = ~ys__n18781 & ~ys__n18964;
  assign new_new_n14527__ = ys__n18781 & ys__n18964;
  assign new_new_n14528__ = ~new_new_n14526__ & ~new_new_n14527__;
  assign new_new_n14529__ = ~ys__n18783 & ~ys__n18965;
  assign new_new_n14530__ = ys__n18783 & ys__n18965;
  assign new_new_n14531__ = ~new_new_n14529__ & ~new_new_n14530__;
  assign new_new_n14532__ = ~new_new_n14528__ & ~new_new_n14531__;
  assign new_new_n14533__ = ~ys__n18785 & ~ys__n18966;
  assign new_new_n14534__ = ys__n18785 & ys__n18966;
  assign new_new_n14535__ = ~new_new_n14533__ & ~new_new_n14534__;
  assign new_new_n14536__ = ~ys__n18787 & ~ys__n18967;
  assign new_new_n14537__ = ys__n18787 & ys__n18967;
  assign new_new_n14538__ = ~new_new_n14536__ & ~new_new_n14537__;
  assign new_new_n14539__ = ~new_new_n14535__ & ~new_new_n14538__;
  assign new_new_n14540__ = new_new_n14532__ & new_new_n14539__;
  assign new_new_n14541__ = ~ys__n18773 & ~ys__n18960;
  assign new_new_n14542__ = ys__n18773 & ys__n18960;
  assign new_new_n14543__ = ~new_new_n14541__ & ~new_new_n14542__;
  assign new_new_n14544__ = ~ys__n18775 & ~ys__n18961;
  assign new_new_n14545__ = ys__n18775 & ys__n18961;
  assign new_new_n14546__ = ~new_new_n14544__ & ~new_new_n14545__;
  assign new_new_n14547__ = ~new_new_n14543__ & ~new_new_n14546__;
  assign new_new_n14548__ = ~ys__n18777 & ~ys__n18962;
  assign new_new_n14549__ = ys__n18777 & ys__n18962;
  assign new_new_n14550__ = ~new_new_n14548__ & ~new_new_n14549__;
  assign new_new_n14551__ = ~ys__n18779 & ~ys__n18963;
  assign new_new_n14552__ = ys__n18779 & ys__n18963;
  assign new_new_n14553__ = ~new_new_n14551__ & ~new_new_n14552__;
  assign new_new_n14554__ = ~new_new_n14550__ & ~new_new_n14553__;
  assign new_new_n14555__ = new_new_n14547__ & new_new_n14554__;
  assign new_new_n14556__ = new_new_n14540__ & new_new_n14555__;
  assign new_new_n14557__ = ~ys__n18797 & ~ys__n18972;
  assign new_new_n14558__ = ys__n18797 & ys__n18972;
  assign new_new_n14559__ = ~new_new_n14557__ & ~new_new_n14558__;
  assign new_new_n14560__ = ~ys__n18799 & ~ys__n18973;
  assign new_new_n14561__ = ys__n18799 & ys__n18973;
  assign new_new_n14562__ = ~new_new_n14560__ & ~new_new_n14561__;
  assign new_new_n14563__ = ~new_new_n14559__ & ~new_new_n14562__;
  assign new_new_n14564__ = ~ys__n18801 & ~ys__n18974;
  assign new_new_n14565__ = ys__n18801 & ys__n18974;
  assign new_new_n14566__ = ~new_new_n14564__ & ~new_new_n14565__;
  assign new_new_n14567__ = ~ys__n18803 & ~ys__n18975;
  assign new_new_n14568__ = ys__n18803 & ys__n18975;
  assign new_new_n14569__ = ~new_new_n14567__ & ~new_new_n14568__;
  assign new_new_n14570__ = ~new_new_n14566__ & ~new_new_n14569__;
  assign new_new_n14571__ = new_new_n14563__ & new_new_n14570__;
  assign new_new_n14572__ = ~ys__n18789 & ~ys__n18968;
  assign new_new_n14573__ = ys__n18789 & ys__n18968;
  assign new_new_n14574__ = ~new_new_n14572__ & ~new_new_n14573__;
  assign new_new_n14575__ = ~ys__n18791 & ~ys__n18969;
  assign new_new_n14576__ = ys__n18791 & ys__n18969;
  assign new_new_n14577__ = ~new_new_n14575__ & ~new_new_n14576__;
  assign new_new_n14578__ = ~new_new_n14574__ & ~new_new_n14577__;
  assign new_new_n14579__ = ~ys__n18793 & ~ys__n18970;
  assign new_new_n14580__ = ys__n18793 & ys__n18970;
  assign new_new_n14581__ = ~new_new_n14579__ & ~new_new_n14580__;
  assign new_new_n14582__ = ~ys__n18795 & ~ys__n18971;
  assign new_new_n14583__ = ys__n18795 & ys__n18971;
  assign new_new_n14584__ = ~new_new_n14582__ & ~new_new_n14583__;
  assign new_new_n14585__ = ~new_new_n14581__ & ~new_new_n14584__;
  assign new_new_n14586__ = new_new_n14578__ & new_new_n14585__;
  assign new_new_n14587__ = new_new_n14571__ & new_new_n14586__;
  assign new_new_n14588__ = new_new_n14556__ & new_new_n14587__;
  assign new_new_n14589__ = new_new_n14525__ & new_new_n14588__;
  assign new_new_n14590__ = ~ys__n19166 & ~new_new_n14589__;
  assign new_new_n14591__ = ys__n844 & ~new_new_n14590__;
  assign new_new_n14592__ = ~ys__n18821 & ~ys__n38174;
  assign new_new_n14593__ = ys__n18821 & ys__n38174;
  assign new_new_n14594__ = ~new_new_n14592__ & ~new_new_n14593__;
  assign new_new_n14595__ = ~ys__n18823 & ~ys__n38175;
  assign new_new_n14596__ = ys__n18823 & ys__n38175;
  assign new_new_n14597__ = ~new_new_n14595__ & ~new_new_n14596__;
  assign new_new_n14598__ = ~new_new_n14594__ & ~new_new_n14597__;
  assign new_new_n14599__ = ~ys__n18825 & ~ys__n38176;
  assign new_new_n14600__ = ys__n18825 & ys__n38176;
  assign new_new_n14601__ = ~new_new_n14599__ & ~new_new_n14600__;
  assign new_new_n14602__ = ~ys__n18827 & ~ys__n38177;
  assign new_new_n14603__ = ys__n18827 & ys__n38177;
  assign new_new_n14604__ = ~new_new_n14602__ & ~new_new_n14603__;
  assign new_new_n14605__ = ~new_new_n14601__ & ~new_new_n14604__;
  assign new_new_n14606__ = new_new_n14598__ & new_new_n14605__;
  assign new_new_n14607__ = ~ys__n18813 & ~ys__n38170;
  assign new_new_n14608__ = ys__n18813 & ys__n38170;
  assign new_new_n14609__ = ~new_new_n14607__ & ~new_new_n14608__;
  assign new_new_n14610__ = ~ys__n18815 & ~ys__n38171;
  assign new_new_n14611__ = ys__n18815 & ys__n38171;
  assign new_new_n14612__ = ~new_new_n14610__ & ~new_new_n14611__;
  assign new_new_n14613__ = ~new_new_n14609__ & ~new_new_n14612__;
  assign new_new_n14614__ = ~ys__n18817 & ~ys__n38172;
  assign new_new_n14615__ = ys__n18817 & ys__n38172;
  assign new_new_n14616__ = ~new_new_n14614__ & ~new_new_n14615__;
  assign new_new_n14617__ = ~ys__n18819 & ~ys__n38173;
  assign new_new_n14618__ = ys__n18819 & ys__n38173;
  assign new_new_n14619__ = ~new_new_n14617__ & ~new_new_n14618__;
  assign new_new_n14620__ = ~new_new_n14616__ & ~new_new_n14619__;
  assign new_new_n14621__ = new_new_n14613__ & new_new_n14620__;
  assign new_new_n14622__ = ~ys__n18805 & ~ys__n38166;
  assign new_new_n14623__ = ys__n18805 & ys__n38166;
  assign new_new_n14624__ = ~new_new_n14622__ & ~new_new_n14623__;
  assign new_new_n14625__ = ~ys__n18807 & ~ys__n38167;
  assign new_new_n14626__ = ys__n18807 & ys__n38167;
  assign new_new_n14627__ = ~new_new_n14625__ & ~new_new_n14626__;
  assign new_new_n14628__ = ~new_new_n14624__ & ~new_new_n14627__;
  assign new_new_n14629__ = ~ys__n18809 & ~ys__n38168;
  assign new_new_n14630__ = ys__n18809 & ys__n38168;
  assign new_new_n14631__ = ~new_new_n14629__ & ~new_new_n14630__;
  assign new_new_n14632__ = ~ys__n18811 & ~ys__n38169;
  assign new_new_n14633__ = ys__n18811 & ys__n38169;
  assign new_new_n14634__ = ~new_new_n14632__ & ~new_new_n14633__;
  assign new_new_n14635__ = ~new_new_n14631__ & ~new_new_n14634__;
  assign new_new_n14636__ = new_new_n14628__ & new_new_n14635__;
  assign new_new_n14637__ = new_new_n14621__ & new_new_n14636__;
  assign new_new_n14638__ = new_new_n14606__ & new_new_n14637__;
  assign new_new_n14639__ = ~ys__n18781 & ~ys__n38154;
  assign new_new_n14640__ = ys__n18781 & ys__n38154;
  assign new_new_n14641__ = ~new_new_n14639__ & ~new_new_n14640__;
  assign new_new_n14642__ = ~ys__n18783 & ~ys__n38155;
  assign new_new_n14643__ = ys__n18783 & ys__n38155;
  assign new_new_n14644__ = ~new_new_n14642__ & ~new_new_n14643__;
  assign new_new_n14645__ = ~new_new_n14641__ & ~new_new_n14644__;
  assign new_new_n14646__ = ~ys__n18785 & ~ys__n38156;
  assign new_new_n14647__ = ys__n18785 & ys__n38156;
  assign new_new_n14648__ = ~new_new_n14646__ & ~new_new_n14647__;
  assign new_new_n14649__ = ~ys__n18787 & ~ys__n38157;
  assign new_new_n14650__ = ys__n18787 & ys__n38157;
  assign new_new_n14651__ = ~new_new_n14649__ & ~new_new_n14650__;
  assign new_new_n14652__ = ~new_new_n14648__ & ~new_new_n14651__;
  assign new_new_n14653__ = new_new_n14645__ & new_new_n14652__;
  assign new_new_n14654__ = ~ys__n18773 & ~ys__n38150;
  assign new_new_n14655__ = ys__n18773 & ys__n38150;
  assign new_new_n14656__ = ~new_new_n14654__ & ~new_new_n14655__;
  assign new_new_n14657__ = ~ys__n18775 & ~ys__n38151;
  assign new_new_n14658__ = ys__n18775 & ys__n38151;
  assign new_new_n14659__ = ~new_new_n14657__ & ~new_new_n14658__;
  assign new_new_n14660__ = ~new_new_n14656__ & ~new_new_n14659__;
  assign new_new_n14661__ = ~ys__n18777 & ~ys__n38152;
  assign new_new_n14662__ = ys__n18777 & ys__n38152;
  assign new_new_n14663__ = ~new_new_n14661__ & ~new_new_n14662__;
  assign new_new_n14664__ = ~ys__n18779 & ~ys__n38153;
  assign new_new_n14665__ = ys__n18779 & ys__n38153;
  assign new_new_n14666__ = ~new_new_n14664__ & ~new_new_n14665__;
  assign new_new_n14667__ = ~new_new_n14663__ & ~new_new_n14666__;
  assign new_new_n14668__ = new_new_n14660__ & new_new_n14667__;
  assign new_new_n14669__ = new_new_n14653__ & new_new_n14668__;
  assign new_new_n14670__ = ~ys__n18797 & ~ys__n38162;
  assign new_new_n14671__ = ys__n18797 & ys__n38162;
  assign new_new_n14672__ = ~new_new_n14670__ & ~new_new_n14671__;
  assign new_new_n14673__ = ~ys__n18799 & ~ys__n38163;
  assign new_new_n14674__ = ys__n18799 & ys__n38163;
  assign new_new_n14675__ = ~new_new_n14673__ & ~new_new_n14674__;
  assign new_new_n14676__ = ~new_new_n14672__ & ~new_new_n14675__;
  assign new_new_n14677__ = ~ys__n18801 & ~ys__n38164;
  assign new_new_n14678__ = ys__n18801 & ys__n38164;
  assign new_new_n14679__ = ~new_new_n14677__ & ~new_new_n14678__;
  assign new_new_n14680__ = ~ys__n18803 & ~ys__n38165;
  assign new_new_n14681__ = ys__n18803 & ys__n38165;
  assign new_new_n14682__ = ~new_new_n14680__ & ~new_new_n14681__;
  assign new_new_n14683__ = ~new_new_n14679__ & ~new_new_n14682__;
  assign new_new_n14684__ = new_new_n14676__ & new_new_n14683__;
  assign new_new_n14685__ = ~ys__n18789 & ~ys__n38158;
  assign new_new_n14686__ = ys__n18789 & ys__n38158;
  assign new_new_n14687__ = ~new_new_n14685__ & ~new_new_n14686__;
  assign new_new_n14688__ = ~ys__n18791 & ~ys__n38159;
  assign new_new_n14689__ = ys__n18791 & ys__n38159;
  assign new_new_n14690__ = ~new_new_n14688__ & ~new_new_n14689__;
  assign new_new_n14691__ = ~new_new_n14687__ & ~new_new_n14690__;
  assign new_new_n14692__ = ~ys__n18793 & ~ys__n38160;
  assign new_new_n14693__ = ys__n18793 & ys__n38160;
  assign new_new_n14694__ = ~new_new_n14692__ & ~new_new_n14693__;
  assign new_new_n14695__ = ~ys__n18795 & ~ys__n38161;
  assign new_new_n14696__ = ys__n18795 & ys__n38161;
  assign new_new_n14697__ = ~new_new_n14695__ & ~new_new_n14696__;
  assign new_new_n14698__ = ~new_new_n14694__ & ~new_new_n14697__;
  assign new_new_n14699__ = new_new_n14691__ & new_new_n14698__;
  assign new_new_n14700__ = new_new_n14684__ & new_new_n14699__;
  assign new_new_n14701__ = new_new_n14669__ & new_new_n14700__;
  assign new_new_n14702__ = new_new_n14638__ & new_new_n14701__;
  assign new_new_n14703__ = ~ys__n37743 & ~new_new_n14702__;
  assign new_new_n14704__ = ys__n842 & ~new_new_n14703__;
  assign new_new_n14705__ = ~new_new_n14591__ & ~new_new_n14704__;
  assign new_new_n14706__ = ~ys__n18821 & ~ys__n38146;
  assign new_new_n14707__ = ys__n18821 & ys__n38146;
  assign new_new_n14708__ = ~new_new_n14706__ & ~new_new_n14707__;
  assign new_new_n14709__ = ~ys__n18823 & ~ys__n38147;
  assign new_new_n14710__ = ys__n18823 & ys__n38147;
  assign new_new_n14711__ = ~new_new_n14709__ & ~new_new_n14710__;
  assign new_new_n14712__ = ~new_new_n14708__ & ~new_new_n14711__;
  assign new_new_n14713__ = ~ys__n18825 & ~ys__n38148;
  assign new_new_n14714__ = ys__n18825 & ys__n38148;
  assign new_new_n14715__ = ~new_new_n14713__ & ~new_new_n14714__;
  assign new_new_n14716__ = ~ys__n18827 & ~ys__n38149;
  assign new_new_n14717__ = ys__n18827 & ys__n38149;
  assign new_new_n14718__ = ~new_new_n14716__ & ~new_new_n14717__;
  assign new_new_n14719__ = ~new_new_n14715__ & ~new_new_n14718__;
  assign new_new_n14720__ = new_new_n14712__ & new_new_n14719__;
  assign new_new_n14721__ = ~ys__n18813 & ~ys__n38142;
  assign new_new_n14722__ = ys__n18813 & ys__n38142;
  assign new_new_n14723__ = ~new_new_n14721__ & ~new_new_n14722__;
  assign new_new_n14724__ = ~ys__n18815 & ~ys__n38143;
  assign new_new_n14725__ = ys__n18815 & ys__n38143;
  assign new_new_n14726__ = ~new_new_n14724__ & ~new_new_n14725__;
  assign new_new_n14727__ = ~new_new_n14723__ & ~new_new_n14726__;
  assign new_new_n14728__ = ~ys__n18817 & ~ys__n38144;
  assign new_new_n14729__ = ys__n18817 & ys__n38144;
  assign new_new_n14730__ = ~new_new_n14728__ & ~new_new_n14729__;
  assign new_new_n14731__ = ~ys__n18819 & ~ys__n38145;
  assign new_new_n14732__ = ys__n18819 & ys__n38145;
  assign new_new_n14733__ = ~new_new_n14731__ & ~new_new_n14732__;
  assign new_new_n14734__ = ~new_new_n14730__ & ~new_new_n14733__;
  assign new_new_n14735__ = new_new_n14727__ & new_new_n14734__;
  assign new_new_n14736__ = ~ys__n18805 & ~ys__n38138;
  assign new_new_n14737__ = ys__n18805 & ys__n38138;
  assign new_new_n14738__ = ~new_new_n14736__ & ~new_new_n14737__;
  assign new_new_n14739__ = ~ys__n18807 & ~ys__n38139;
  assign new_new_n14740__ = ys__n18807 & ys__n38139;
  assign new_new_n14741__ = ~new_new_n14739__ & ~new_new_n14740__;
  assign new_new_n14742__ = ~new_new_n14738__ & ~new_new_n14741__;
  assign new_new_n14743__ = ~ys__n18809 & ~ys__n38140;
  assign new_new_n14744__ = ys__n18809 & ys__n38140;
  assign new_new_n14745__ = ~new_new_n14743__ & ~new_new_n14744__;
  assign new_new_n14746__ = ~ys__n18811 & ~ys__n38141;
  assign new_new_n14747__ = ys__n18811 & ys__n38141;
  assign new_new_n14748__ = ~new_new_n14746__ & ~new_new_n14747__;
  assign new_new_n14749__ = ~new_new_n14745__ & ~new_new_n14748__;
  assign new_new_n14750__ = new_new_n14742__ & new_new_n14749__;
  assign new_new_n14751__ = new_new_n14735__ & new_new_n14750__;
  assign new_new_n14752__ = new_new_n14720__ & new_new_n14751__;
  assign new_new_n14753__ = ~ys__n18781 & ~ys__n38126;
  assign new_new_n14754__ = ys__n18781 & ys__n38126;
  assign new_new_n14755__ = ~new_new_n14753__ & ~new_new_n14754__;
  assign new_new_n14756__ = ~ys__n18783 & ~ys__n38127;
  assign new_new_n14757__ = ys__n18783 & ys__n38127;
  assign new_new_n14758__ = ~new_new_n14756__ & ~new_new_n14757__;
  assign new_new_n14759__ = ~new_new_n14755__ & ~new_new_n14758__;
  assign new_new_n14760__ = ~ys__n18785 & ~ys__n38128;
  assign new_new_n14761__ = ys__n18785 & ys__n38128;
  assign new_new_n14762__ = ~new_new_n14760__ & ~new_new_n14761__;
  assign new_new_n14763__ = ~ys__n18787 & ~ys__n38129;
  assign new_new_n14764__ = ys__n18787 & ys__n38129;
  assign new_new_n14765__ = ~new_new_n14763__ & ~new_new_n14764__;
  assign new_new_n14766__ = ~new_new_n14762__ & ~new_new_n14765__;
  assign new_new_n14767__ = new_new_n14759__ & new_new_n14766__;
  assign new_new_n14768__ = ~ys__n18773 & ~ys__n38122;
  assign new_new_n14769__ = ys__n18773 & ys__n38122;
  assign new_new_n14770__ = ~new_new_n14768__ & ~new_new_n14769__;
  assign new_new_n14771__ = ~ys__n18775 & ~ys__n38123;
  assign new_new_n14772__ = ys__n18775 & ys__n38123;
  assign new_new_n14773__ = ~new_new_n14771__ & ~new_new_n14772__;
  assign new_new_n14774__ = ~new_new_n14770__ & ~new_new_n14773__;
  assign new_new_n14775__ = ~ys__n18777 & ~ys__n38124;
  assign new_new_n14776__ = ys__n18777 & ys__n38124;
  assign new_new_n14777__ = ~new_new_n14775__ & ~new_new_n14776__;
  assign new_new_n14778__ = ~ys__n18779 & ~ys__n38125;
  assign new_new_n14779__ = ys__n18779 & ys__n38125;
  assign new_new_n14780__ = ~new_new_n14778__ & ~new_new_n14779__;
  assign new_new_n14781__ = ~new_new_n14777__ & ~new_new_n14780__;
  assign new_new_n14782__ = new_new_n14774__ & new_new_n14781__;
  assign new_new_n14783__ = new_new_n14767__ & new_new_n14782__;
  assign new_new_n14784__ = ~ys__n18797 & ~ys__n38134;
  assign new_new_n14785__ = ys__n18797 & ys__n38134;
  assign new_new_n14786__ = ~new_new_n14784__ & ~new_new_n14785__;
  assign new_new_n14787__ = ~ys__n18799 & ~ys__n38135;
  assign new_new_n14788__ = ys__n18799 & ys__n38135;
  assign new_new_n14789__ = ~new_new_n14787__ & ~new_new_n14788__;
  assign new_new_n14790__ = ~new_new_n14786__ & ~new_new_n14789__;
  assign new_new_n14791__ = ~ys__n18801 & ~ys__n38136;
  assign new_new_n14792__ = ys__n18801 & ys__n38136;
  assign new_new_n14793__ = ~new_new_n14791__ & ~new_new_n14792__;
  assign new_new_n14794__ = ~ys__n18803 & ~ys__n38137;
  assign new_new_n14795__ = ys__n18803 & ys__n38137;
  assign new_new_n14796__ = ~new_new_n14794__ & ~new_new_n14795__;
  assign new_new_n14797__ = ~new_new_n14793__ & ~new_new_n14796__;
  assign new_new_n14798__ = new_new_n14790__ & new_new_n14797__;
  assign new_new_n14799__ = ~ys__n18789 & ~ys__n38130;
  assign new_new_n14800__ = ys__n18789 & ys__n38130;
  assign new_new_n14801__ = ~new_new_n14799__ & ~new_new_n14800__;
  assign new_new_n14802__ = ~ys__n18791 & ~ys__n38131;
  assign new_new_n14803__ = ys__n18791 & ys__n38131;
  assign new_new_n14804__ = ~new_new_n14802__ & ~new_new_n14803__;
  assign new_new_n14805__ = ~new_new_n14801__ & ~new_new_n14804__;
  assign new_new_n14806__ = ~ys__n18793 & ~ys__n38132;
  assign new_new_n14807__ = ys__n18793 & ys__n38132;
  assign new_new_n14808__ = ~new_new_n14806__ & ~new_new_n14807__;
  assign new_new_n14809__ = ~ys__n18795 & ~ys__n38133;
  assign new_new_n14810__ = ys__n18795 & ys__n38133;
  assign new_new_n14811__ = ~new_new_n14809__ & ~new_new_n14810__;
  assign new_new_n14812__ = ~new_new_n14808__ & ~new_new_n14811__;
  assign new_new_n14813__ = new_new_n14805__ & new_new_n14812__;
  assign new_new_n14814__ = new_new_n14798__ & new_new_n14813__;
  assign new_new_n14815__ = new_new_n14783__ & new_new_n14814__;
  assign new_new_n14816__ = new_new_n14752__ & new_new_n14815__;
  assign new_new_n14817__ = ~ys__n37744 & ~new_new_n14816__;
  assign new_new_n14818__ = ys__n840 & ~new_new_n14817__;
  assign new_new_n14819__ = ~ys__n18821 & ~ys__n38118;
  assign new_new_n14820__ = ys__n18821 & ys__n38118;
  assign new_new_n14821__ = ~new_new_n14819__ & ~new_new_n14820__;
  assign new_new_n14822__ = ~ys__n18823 & ~ys__n38119;
  assign new_new_n14823__ = ys__n18823 & ys__n38119;
  assign new_new_n14824__ = ~new_new_n14822__ & ~new_new_n14823__;
  assign new_new_n14825__ = ~new_new_n14821__ & ~new_new_n14824__;
  assign new_new_n14826__ = ~ys__n18825 & ~ys__n38120;
  assign new_new_n14827__ = ys__n18825 & ys__n38120;
  assign new_new_n14828__ = ~new_new_n14826__ & ~new_new_n14827__;
  assign new_new_n14829__ = ~ys__n18827 & ~ys__n38121;
  assign new_new_n14830__ = ys__n18827 & ys__n38121;
  assign new_new_n14831__ = ~new_new_n14829__ & ~new_new_n14830__;
  assign new_new_n14832__ = ~new_new_n14828__ & ~new_new_n14831__;
  assign new_new_n14833__ = new_new_n14825__ & new_new_n14832__;
  assign new_new_n14834__ = ~ys__n18813 & ~ys__n38114;
  assign new_new_n14835__ = ys__n18813 & ys__n38114;
  assign new_new_n14836__ = ~new_new_n14834__ & ~new_new_n14835__;
  assign new_new_n14837__ = ~ys__n18815 & ~ys__n38115;
  assign new_new_n14838__ = ys__n18815 & ys__n38115;
  assign new_new_n14839__ = ~new_new_n14837__ & ~new_new_n14838__;
  assign new_new_n14840__ = ~new_new_n14836__ & ~new_new_n14839__;
  assign new_new_n14841__ = ~ys__n18817 & ~ys__n38116;
  assign new_new_n14842__ = ys__n18817 & ys__n38116;
  assign new_new_n14843__ = ~new_new_n14841__ & ~new_new_n14842__;
  assign new_new_n14844__ = ~ys__n18819 & ~ys__n38117;
  assign new_new_n14845__ = ys__n18819 & ys__n38117;
  assign new_new_n14846__ = ~new_new_n14844__ & ~new_new_n14845__;
  assign new_new_n14847__ = ~new_new_n14843__ & ~new_new_n14846__;
  assign new_new_n14848__ = new_new_n14840__ & new_new_n14847__;
  assign new_new_n14849__ = ~ys__n18805 & ~ys__n38110;
  assign new_new_n14850__ = ys__n18805 & ys__n38110;
  assign new_new_n14851__ = ~new_new_n14849__ & ~new_new_n14850__;
  assign new_new_n14852__ = ~ys__n18807 & ~ys__n38111;
  assign new_new_n14853__ = ys__n18807 & ys__n38111;
  assign new_new_n14854__ = ~new_new_n14852__ & ~new_new_n14853__;
  assign new_new_n14855__ = ~new_new_n14851__ & ~new_new_n14854__;
  assign new_new_n14856__ = ~ys__n18809 & ~ys__n38112;
  assign new_new_n14857__ = ys__n18809 & ys__n38112;
  assign new_new_n14858__ = ~new_new_n14856__ & ~new_new_n14857__;
  assign new_new_n14859__ = ~ys__n18811 & ~ys__n38113;
  assign new_new_n14860__ = ys__n18811 & ys__n38113;
  assign new_new_n14861__ = ~new_new_n14859__ & ~new_new_n14860__;
  assign new_new_n14862__ = ~new_new_n14858__ & ~new_new_n14861__;
  assign new_new_n14863__ = new_new_n14855__ & new_new_n14862__;
  assign new_new_n14864__ = new_new_n14848__ & new_new_n14863__;
  assign new_new_n14865__ = new_new_n14833__ & new_new_n14864__;
  assign new_new_n14866__ = ~ys__n18781 & ~ys__n38098;
  assign new_new_n14867__ = ys__n18781 & ys__n38098;
  assign new_new_n14868__ = ~new_new_n14866__ & ~new_new_n14867__;
  assign new_new_n14869__ = ~ys__n18783 & ~ys__n38099;
  assign new_new_n14870__ = ys__n18783 & ys__n38099;
  assign new_new_n14871__ = ~new_new_n14869__ & ~new_new_n14870__;
  assign new_new_n14872__ = ~new_new_n14868__ & ~new_new_n14871__;
  assign new_new_n14873__ = ~ys__n18785 & ~ys__n38100;
  assign new_new_n14874__ = ys__n18785 & ys__n38100;
  assign new_new_n14875__ = ~new_new_n14873__ & ~new_new_n14874__;
  assign new_new_n14876__ = ~ys__n18787 & ~ys__n38101;
  assign new_new_n14877__ = ys__n18787 & ys__n38101;
  assign new_new_n14878__ = ~new_new_n14876__ & ~new_new_n14877__;
  assign new_new_n14879__ = ~new_new_n14875__ & ~new_new_n14878__;
  assign new_new_n14880__ = new_new_n14872__ & new_new_n14879__;
  assign new_new_n14881__ = ~ys__n18773 & ~ys__n38094;
  assign new_new_n14882__ = ys__n18773 & ys__n38094;
  assign new_new_n14883__ = ~new_new_n14881__ & ~new_new_n14882__;
  assign new_new_n14884__ = ~ys__n18775 & ~ys__n38095;
  assign new_new_n14885__ = ys__n18775 & ys__n38095;
  assign new_new_n14886__ = ~new_new_n14884__ & ~new_new_n14885__;
  assign new_new_n14887__ = ~new_new_n14883__ & ~new_new_n14886__;
  assign new_new_n14888__ = ~ys__n18777 & ~ys__n38096;
  assign new_new_n14889__ = ys__n18777 & ys__n38096;
  assign new_new_n14890__ = ~new_new_n14888__ & ~new_new_n14889__;
  assign new_new_n14891__ = ~ys__n18779 & ~ys__n38097;
  assign new_new_n14892__ = ys__n18779 & ys__n38097;
  assign new_new_n14893__ = ~new_new_n14891__ & ~new_new_n14892__;
  assign new_new_n14894__ = ~new_new_n14890__ & ~new_new_n14893__;
  assign new_new_n14895__ = new_new_n14887__ & new_new_n14894__;
  assign new_new_n14896__ = new_new_n14880__ & new_new_n14895__;
  assign new_new_n14897__ = ~ys__n18797 & ~ys__n38106;
  assign new_new_n14898__ = ys__n18797 & ys__n38106;
  assign new_new_n14899__ = ~new_new_n14897__ & ~new_new_n14898__;
  assign new_new_n14900__ = ~ys__n18799 & ~ys__n38107;
  assign new_new_n14901__ = ys__n18799 & ys__n38107;
  assign new_new_n14902__ = ~new_new_n14900__ & ~new_new_n14901__;
  assign new_new_n14903__ = ~new_new_n14899__ & ~new_new_n14902__;
  assign new_new_n14904__ = ~ys__n18801 & ~ys__n38108;
  assign new_new_n14905__ = ys__n18801 & ys__n38108;
  assign new_new_n14906__ = ~new_new_n14904__ & ~new_new_n14905__;
  assign new_new_n14907__ = ~ys__n18803 & ~ys__n38109;
  assign new_new_n14908__ = ys__n18803 & ys__n38109;
  assign new_new_n14909__ = ~new_new_n14907__ & ~new_new_n14908__;
  assign new_new_n14910__ = ~new_new_n14906__ & ~new_new_n14909__;
  assign new_new_n14911__ = new_new_n14903__ & new_new_n14910__;
  assign new_new_n14912__ = ~ys__n18789 & ~ys__n38102;
  assign new_new_n14913__ = ys__n18789 & ys__n38102;
  assign new_new_n14914__ = ~new_new_n14912__ & ~new_new_n14913__;
  assign new_new_n14915__ = ~ys__n18791 & ~ys__n38103;
  assign new_new_n14916__ = ys__n18791 & ys__n38103;
  assign new_new_n14917__ = ~new_new_n14915__ & ~new_new_n14916__;
  assign new_new_n14918__ = ~new_new_n14914__ & ~new_new_n14917__;
  assign new_new_n14919__ = ~ys__n18793 & ~ys__n38104;
  assign new_new_n14920__ = ys__n18793 & ys__n38104;
  assign new_new_n14921__ = ~new_new_n14919__ & ~new_new_n14920__;
  assign new_new_n14922__ = ~ys__n18795 & ~ys__n38105;
  assign new_new_n14923__ = ys__n18795 & ys__n38105;
  assign new_new_n14924__ = ~new_new_n14922__ & ~new_new_n14923__;
  assign new_new_n14925__ = ~new_new_n14921__ & ~new_new_n14924__;
  assign new_new_n14926__ = new_new_n14918__ & new_new_n14925__;
  assign new_new_n14927__ = new_new_n14911__ & new_new_n14926__;
  assign new_new_n14928__ = new_new_n14896__ & new_new_n14927__;
  assign new_new_n14929__ = new_new_n14865__ & new_new_n14928__;
  assign new_new_n14930__ = ~ys__n37745 & ~new_new_n14929__;
  assign new_new_n14931__ = ys__n838 & ~new_new_n14930__;
  assign new_new_n14932__ = ~new_new_n14818__ & ~new_new_n14931__;
  assign new_new_n14933__ = new_new_n14705__ & new_new_n14932__;
  assign new_new_n14934__ = new_new_n14478__ & new_new_n14933__;
  assign new_new_n14935__ = ~ys__n18821 & ~ys__n37866;
  assign new_new_n14936__ = ys__n18821 & ys__n37866;
  assign new_new_n14937__ = ~new_new_n14935__ & ~new_new_n14936__;
  assign new_new_n14938__ = ~ys__n18823 & ~ys__n37867;
  assign new_new_n14939__ = ys__n18823 & ys__n37867;
  assign new_new_n14940__ = ~new_new_n14938__ & ~new_new_n14939__;
  assign new_new_n14941__ = ~new_new_n14937__ & ~new_new_n14940__;
  assign new_new_n14942__ = ~ys__n18825 & ~ys__n37868;
  assign new_new_n14943__ = ys__n18825 & ys__n37868;
  assign new_new_n14944__ = ~new_new_n14942__ & ~new_new_n14943__;
  assign new_new_n14945__ = ~ys__n18827 & ~ys__n37869;
  assign new_new_n14946__ = ys__n18827 & ys__n37869;
  assign new_new_n14947__ = ~new_new_n14945__ & ~new_new_n14946__;
  assign new_new_n14948__ = ~new_new_n14944__ & ~new_new_n14947__;
  assign new_new_n14949__ = new_new_n14941__ & new_new_n14948__;
  assign new_new_n14950__ = ~ys__n18813 & ~ys__n37862;
  assign new_new_n14951__ = ys__n18813 & ys__n37862;
  assign new_new_n14952__ = ~new_new_n14950__ & ~new_new_n14951__;
  assign new_new_n14953__ = ~ys__n18815 & ~ys__n37863;
  assign new_new_n14954__ = ys__n18815 & ys__n37863;
  assign new_new_n14955__ = ~new_new_n14953__ & ~new_new_n14954__;
  assign new_new_n14956__ = ~new_new_n14952__ & ~new_new_n14955__;
  assign new_new_n14957__ = ~ys__n18817 & ~ys__n37864;
  assign new_new_n14958__ = ys__n18817 & ys__n37864;
  assign new_new_n14959__ = ~new_new_n14957__ & ~new_new_n14958__;
  assign new_new_n14960__ = ~ys__n18819 & ~ys__n37865;
  assign new_new_n14961__ = ys__n18819 & ys__n37865;
  assign new_new_n14962__ = ~new_new_n14960__ & ~new_new_n14961__;
  assign new_new_n14963__ = ~new_new_n14959__ & ~new_new_n14962__;
  assign new_new_n14964__ = new_new_n14956__ & new_new_n14963__;
  assign new_new_n14965__ = ~ys__n18805 & ~ys__n37858;
  assign new_new_n14966__ = ys__n18805 & ys__n37858;
  assign new_new_n14967__ = ~new_new_n14965__ & ~new_new_n14966__;
  assign new_new_n14968__ = ~ys__n18807 & ~ys__n37859;
  assign new_new_n14969__ = ys__n18807 & ys__n37859;
  assign new_new_n14970__ = ~new_new_n14968__ & ~new_new_n14969__;
  assign new_new_n14971__ = ~new_new_n14967__ & ~new_new_n14970__;
  assign new_new_n14972__ = ~ys__n18809 & ~ys__n37860;
  assign new_new_n14973__ = ys__n18809 & ys__n37860;
  assign new_new_n14974__ = ~new_new_n14972__ & ~new_new_n14973__;
  assign new_new_n14975__ = ~ys__n18811 & ~ys__n37861;
  assign new_new_n14976__ = ys__n18811 & ys__n37861;
  assign new_new_n14977__ = ~new_new_n14975__ & ~new_new_n14976__;
  assign new_new_n14978__ = ~new_new_n14974__ & ~new_new_n14977__;
  assign new_new_n14979__ = new_new_n14971__ & new_new_n14978__;
  assign new_new_n14980__ = new_new_n14964__ & new_new_n14979__;
  assign new_new_n14981__ = new_new_n14949__ & new_new_n14980__;
  assign new_new_n14982__ = ~ys__n18781 & ~ys__n37846;
  assign new_new_n14983__ = ys__n18781 & ys__n37846;
  assign new_new_n14984__ = ~new_new_n14982__ & ~new_new_n14983__;
  assign new_new_n14985__ = ~ys__n18783 & ~ys__n37847;
  assign new_new_n14986__ = ys__n18783 & ys__n37847;
  assign new_new_n14987__ = ~new_new_n14985__ & ~new_new_n14986__;
  assign new_new_n14988__ = ~new_new_n14984__ & ~new_new_n14987__;
  assign new_new_n14989__ = ~ys__n18785 & ~ys__n37848;
  assign new_new_n14990__ = ys__n18785 & ys__n37848;
  assign new_new_n14991__ = ~new_new_n14989__ & ~new_new_n14990__;
  assign new_new_n14992__ = ~ys__n18787 & ~ys__n37849;
  assign new_new_n14993__ = ys__n18787 & ys__n37849;
  assign new_new_n14994__ = ~new_new_n14992__ & ~new_new_n14993__;
  assign new_new_n14995__ = ~new_new_n14991__ & ~new_new_n14994__;
  assign new_new_n14996__ = new_new_n14988__ & new_new_n14995__;
  assign new_new_n14997__ = ~ys__n18773 & ~ys__n37842;
  assign new_new_n14998__ = ys__n18773 & ys__n37842;
  assign new_new_n14999__ = ~new_new_n14997__ & ~new_new_n14998__;
  assign new_new_n15000__ = ~ys__n18775 & ~ys__n37843;
  assign new_new_n15001__ = ys__n18775 & ys__n37843;
  assign new_new_n15002__ = ~new_new_n15000__ & ~new_new_n15001__;
  assign new_new_n15003__ = ~new_new_n14999__ & ~new_new_n15002__;
  assign new_new_n15004__ = ~ys__n18777 & ~ys__n37844;
  assign new_new_n15005__ = ys__n18777 & ys__n37844;
  assign new_new_n15006__ = ~new_new_n15004__ & ~new_new_n15005__;
  assign new_new_n15007__ = ~ys__n18779 & ~ys__n37845;
  assign new_new_n15008__ = ys__n18779 & ys__n37845;
  assign new_new_n15009__ = ~new_new_n15007__ & ~new_new_n15008__;
  assign new_new_n15010__ = ~new_new_n15006__ & ~new_new_n15009__;
  assign new_new_n15011__ = new_new_n15003__ & new_new_n15010__;
  assign new_new_n15012__ = new_new_n14996__ & new_new_n15011__;
  assign new_new_n15013__ = ~ys__n18797 & ~ys__n37854;
  assign new_new_n15014__ = ys__n18797 & ys__n37854;
  assign new_new_n15015__ = ~new_new_n15013__ & ~new_new_n15014__;
  assign new_new_n15016__ = ~ys__n18799 & ~ys__n37855;
  assign new_new_n15017__ = ys__n18799 & ys__n37855;
  assign new_new_n15018__ = ~new_new_n15016__ & ~new_new_n15017__;
  assign new_new_n15019__ = ~new_new_n15015__ & ~new_new_n15018__;
  assign new_new_n15020__ = ~ys__n18801 & ~ys__n37856;
  assign new_new_n15021__ = ys__n18801 & ys__n37856;
  assign new_new_n15022__ = ~new_new_n15020__ & ~new_new_n15021__;
  assign new_new_n15023__ = ~ys__n18803 & ~ys__n37857;
  assign new_new_n15024__ = ys__n18803 & ys__n37857;
  assign new_new_n15025__ = ~new_new_n15023__ & ~new_new_n15024__;
  assign new_new_n15026__ = ~new_new_n15022__ & ~new_new_n15025__;
  assign new_new_n15027__ = new_new_n15019__ & new_new_n15026__;
  assign new_new_n15028__ = ~ys__n18789 & ~ys__n37850;
  assign new_new_n15029__ = ys__n18789 & ys__n37850;
  assign new_new_n15030__ = ~new_new_n15028__ & ~new_new_n15029__;
  assign new_new_n15031__ = ~ys__n18791 & ~ys__n37851;
  assign new_new_n15032__ = ys__n18791 & ys__n37851;
  assign new_new_n15033__ = ~new_new_n15031__ & ~new_new_n15032__;
  assign new_new_n15034__ = ~new_new_n15030__ & ~new_new_n15033__;
  assign new_new_n15035__ = ~ys__n18793 & ~ys__n37852;
  assign new_new_n15036__ = ys__n18793 & ys__n37852;
  assign new_new_n15037__ = ~new_new_n15035__ & ~new_new_n15036__;
  assign new_new_n15038__ = ~ys__n18795 & ~ys__n37853;
  assign new_new_n15039__ = ys__n18795 & ys__n37853;
  assign new_new_n15040__ = ~new_new_n15038__ & ~new_new_n15039__;
  assign new_new_n15041__ = ~new_new_n15037__ & ~new_new_n15040__;
  assign new_new_n15042__ = new_new_n15034__ & new_new_n15041__;
  assign new_new_n15043__ = new_new_n15027__ & new_new_n15042__;
  assign new_new_n15044__ = new_new_n15012__ & new_new_n15043__;
  assign new_new_n15045__ = new_new_n14981__ & new_new_n15044__;
  assign new_new_n15046__ = ~ys__n37754 & ~new_new_n15045__;
  assign new_new_n15047__ = ys__n850 & ~new_new_n15046__;
  assign new_new_n15048__ = ~ys__n18821 & ~ys__n37838;
  assign new_new_n15049__ = ys__n18821 & ys__n37838;
  assign new_new_n15050__ = ~new_new_n15048__ & ~new_new_n15049__;
  assign new_new_n15051__ = ~ys__n18823 & ~ys__n37839;
  assign new_new_n15052__ = ys__n18823 & ys__n37839;
  assign new_new_n15053__ = ~new_new_n15051__ & ~new_new_n15052__;
  assign new_new_n15054__ = ~new_new_n15050__ & ~new_new_n15053__;
  assign new_new_n15055__ = ~ys__n18825 & ~ys__n37840;
  assign new_new_n15056__ = ys__n18825 & ys__n37840;
  assign new_new_n15057__ = ~new_new_n15055__ & ~new_new_n15056__;
  assign new_new_n15058__ = ~ys__n18827 & ~ys__n37841;
  assign new_new_n15059__ = ys__n18827 & ys__n37841;
  assign new_new_n15060__ = ~new_new_n15058__ & ~new_new_n15059__;
  assign new_new_n15061__ = ~new_new_n15057__ & ~new_new_n15060__;
  assign new_new_n15062__ = new_new_n15054__ & new_new_n15061__;
  assign new_new_n15063__ = ~ys__n18813 & ~ys__n37834;
  assign new_new_n15064__ = ys__n18813 & ys__n37834;
  assign new_new_n15065__ = ~new_new_n15063__ & ~new_new_n15064__;
  assign new_new_n15066__ = ~ys__n18815 & ~ys__n37835;
  assign new_new_n15067__ = ys__n18815 & ys__n37835;
  assign new_new_n15068__ = ~new_new_n15066__ & ~new_new_n15067__;
  assign new_new_n15069__ = ~new_new_n15065__ & ~new_new_n15068__;
  assign new_new_n15070__ = ~ys__n18817 & ~ys__n37836;
  assign new_new_n15071__ = ys__n18817 & ys__n37836;
  assign new_new_n15072__ = ~new_new_n15070__ & ~new_new_n15071__;
  assign new_new_n15073__ = ~ys__n18819 & ~ys__n37837;
  assign new_new_n15074__ = ys__n18819 & ys__n37837;
  assign new_new_n15075__ = ~new_new_n15073__ & ~new_new_n15074__;
  assign new_new_n15076__ = ~new_new_n15072__ & ~new_new_n15075__;
  assign new_new_n15077__ = new_new_n15069__ & new_new_n15076__;
  assign new_new_n15078__ = ~ys__n18805 & ~ys__n37830;
  assign new_new_n15079__ = ys__n18805 & ys__n37830;
  assign new_new_n15080__ = ~new_new_n15078__ & ~new_new_n15079__;
  assign new_new_n15081__ = ~ys__n18807 & ~ys__n37831;
  assign new_new_n15082__ = ys__n18807 & ys__n37831;
  assign new_new_n15083__ = ~new_new_n15081__ & ~new_new_n15082__;
  assign new_new_n15084__ = ~new_new_n15080__ & ~new_new_n15083__;
  assign new_new_n15085__ = ~ys__n18809 & ~ys__n37832;
  assign new_new_n15086__ = ys__n18809 & ys__n37832;
  assign new_new_n15087__ = ~new_new_n15085__ & ~new_new_n15086__;
  assign new_new_n15088__ = ~ys__n18811 & ~ys__n37833;
  assign new_new_n15089__ = ys__n18811 & ys__n37833;
  assign new_new_n15090__ = ~new_new_n15088__ & ~new_new_n15089__;
  assign new_new_n15091__ = ~new_new_n15087__ & ~new_new_n15090__;
  assign new_new_n15092__ = new_new_n15084__ & new_new_n15091__;
  assign new_new_n15093__ = new_new_n15077__ & new_new_n15092__;
  assign new_new_n15094__ = new_new_n15062__ & new_new_n15093__;
  assign new_new_n15095__ = ~ys__n18781 & ~ys__n37818;
  assign new_new_n15096__ = ys__n18781 & ys__n37818;
  assign new_new_n15097__ = ~new_new_n15095__ & ~new_new_n15096__;
  assign new_new_n15098__ = ~ys__n18783 & ~ys__n37819;
  assign new_new_n15099__ = ys__n18783 & ys__n37819;
  assign new_new_n15100__ = ~new_new_n15098__ & ~new_new_n15099__;
  assign new_new_n15101__ = ~new_new_n15097__ & ~new_new_n15100__;
  assign new_new_n15102__ = ~ys__n18785 & ~ys__n37820;
  assign new_new_n15103__ = ys__n18785 & ys__n37820;
  assign new_new_n15104__ = ~new_new_n15102__ & ~new_new_n15103__;
  assign new_new_n15105__ = ~ys__n18787 & ~ys__n37821;
  assign new_new_n15106__ = ys__n18787 & ys__n37821;
  assign new_new_n15107__ = ~new_new_n15105__ & ~new_new_n15106__;
  assign new_new_n15108__ = ~new_new_n15104__ & ~new_new_n15107__;
  assign new_new_n15109__ = new_new_n15101__ & new_new_n15108__;
  assign new_new_n15110__ = ~ys__n18773 & ~ys__n37814;
  assign new_new_n15111__ = ys__n18773 & ys__n37814;
  assign new_new_n15112__ = ~new_new_n15110__ & ~new_new_n15111__;
  assign new_new_n15113__ = ~ys__n18775 & ~ys__n37815;
  assign new_new_n15114__ = ys__n18775 & ys__n37815;
  assign new_new_n15115__ = ~new_new_n15113__ & ~new_new_n15114__;
  assign new_new_n15116__ = ~new_new_n15112__ & ~new_new_n15115__;
  assign new_new_n15117__ = ~ys__n18777 & ~ys__n37816;
  assign new_new_n15118__ = ys__n18777 & ys__n37816;
  assign new_new_n15119__ = ~new_new_n15117__ & ~new_new_n15118__;
  assign new_new_n15120__ = ~ys__n18779 & ~ys__n37817;
  assign new_new_n15121__ = ys__n18779 & ys__n37817;
  assign new_new_n15122__ = ~new_new_n15120__ & ~new_new_n15121__;
  assign new_new_n15123__ = ~new_new_n15119__ & ~new_new_n15122__;
  assign new_new_n15124__ = new_new_n15116__ & new_new_n15123__;
  assign new_new_n15125__ = new_new_n15109__ & new_new_n15124__;
  assign new_new_n15126__ = ~ys__n18797 & ~ys__n37826;
  assign new_new_n15127__ = ys__n18797 & ys__n37826;
  assign new_new_n15128__ = ~new_new_n15126__ & ~new_new_n15127__;
  assign new_new_n15129__ = ~ys__n18799 & ~ys__n37827;
  assign new_new_n15130__ = ys__n18799 & ys__n37827;
  assign new_new_n15131__ = ~new_new_n15129__ & ~new_new_n15130__;
  assign new_new_n15132__ = ~new_new_n15128__ & ~new_new_n15131__;
  assign new_new_n15133__ = ~ys__n18801 & ~ys__n37828;
  assign new_new_n15134__ = ys__n18801 & ys__n37828;
  assign new_new_n15135__ = ~new_new_n15133__ & ~new_new_n15134__;
  assign new_new_n15136__ = ~ys__n18803 & ~ys__n37829;
  assign new_new_n15137__ = ys__n18803 & ys__n37829;
  assign new_new_n15138__ = ~new_new_n15136__ & ~new_new_n15137__;
  assign new_new_n15139__ = ~new_new_n15135__ & ~new_new_n15138__;
  assign new_new_n15140__ = new_new_n15132__ & new_new_n15139__;
  assign new_new_n15141__ = ~ys__n18789 & ~ys__n37822;
  assign new_new_n15142__ = ys__n18789 & ys__n37822;
  assign new_new_n15143__ = ~new_new_n15141__ & ~new_new_n15142__;
  assign new_new_n15144__ = ~ys__n18791 & ~ys__n37823;
  assign new_new_n15145__ = ys__n18791 & ys__n37823;
  assign new_new_n15146__ = ~new_new_n15144__ & ~new_new_n15145__;
  assign new_new_n15147__ = ~new_new_n15143__ & ~new_new_n15146__;
  assign new_new_n15148__ = ~ys__n18793 & ~ys__n37824;
  assign new_new_n15149__ = ys__n18793 & ys__n37824;
  assign new_new_n15150__ = ~new_new_n15148__ & ~new_new_n15149__;
  assign new_new_n15151__ = ~ys__n18795 & ~ys__n37825;
  assign new_new_n15152__ = ys__n18795 & ys__n37825;
  assign new_new_n15153__ = ~new_new_n15151__ & ~new_new_n15152__;
  assign new_new_n15154__ = ~new_new_n15150__ & ~new_new_n15153__;
  assign new_new_n15155__ = new_new_n15147__ & new_new_n15154__;
  assign new_new_n15156__ = new_new_n15140__ & new_new_n15155__;
  assign new_new_n15157__ = new_new_n15125__ & new_new_n15156__;
  assign new_new_n15158__ = new_new_n15094__ & new_new_n15157__;
  assign new_new_n15159__ = ~ys__n37755 & ~new_new_n15158__;
  assign new_new_n15160__ = ys__n848 & ~new_new_n15159__;
  assign new_new_n15161__ = ~new_new_n15047__ & ~new_new_n15160__;
  assign new_new_n15162__ = ~ys__n18821 & ~ys__n37810;
  assign new_new_n15163__ = ys__n18821 & ys__n37810;
  assign new_new_n15164__ = ~new_new_n15162__ & ~new_new_n15163__;
  assign new_new_n15165__ = ~ys__n18823 & ~ys__n37811;
  assign new_new_n15166__ = ys__n18823 & ys__n37811;
  assign new_new_n15167__ = ~new_new_n15165__ & ~new_new_n15166__;
  assign new_new_n15168__ = ~new_new_n15164__ & ~new_new_n15167__;
  assign new_new_n15169__ = ~ys__n18825 & ~ys__n37812;
  assign new_new_n15170__ = ys__n18825 & ys__n37812;
  assign new_new_n15171__ = ~new_new_n15169__ & ~new_new_n15170__;
  assign new_new_n15172__ = ~ys__n18827 & ~ys__n37813;
  assign new_new_n15173__ = ys__n18827 & ys__n37813;
  assign new_new_n15174__ = ~new_new_n15172__ & ~new_new_n15173__;
  assign new_new_n15175__ = ~new_new_n15171__ & ~new_new_n15174__;
  assign new_new_n15176__ = new_new_n15168__ & new_new_n15175__;
  assign new_new_n15177__ = ~ys__n18813 & ~ys__n37806;
  assign new_new_n15178__ = ys__n18813 & ys__n37806;
  assign new_new_n15179__ = ~new_new_n15177__ & ~new_new_n15178__;
  assign new_new_n15180__ = ~ys__n18815 & ~ys__n37807;
  assign new_new_n15181__ = ys__n18815 & ys__n37807;
  assign new_new_n15182__ = ~new_new_n15180__ & ~new_new_n15181__;
  assign new_new_n15183__ = ~new_new_n15179__ & ~new_new_n15182__;
  assign new_new_n15184__ = ~ys__n18817 & ~ys__n37808;
  assign new_new_n15185__ = ys__n18817 & ys__n37808;
  assign new_new_n15186__ = ~new_new_n15184__ & ~new_new_n15185__;
  assign new_new_n15187__ = ~ys__n18819 & ~ys__n37809;
  assign new_new_n15188__ = ys__n18819 & ys__n37809;
  assign new_new_n15189__ = ~new_new_n15187__ & ~new_new_n15188__;
  assign new_new_n15190__ = ~new_new_n15186__ & ~new_new_n15189__;
  assign new_new_n15191__ = new_new_n15183__ & new_new_n15190__;
  assign new_new_n15192__ = ~ys__n18805 & ~ys__n37802;
  assign new_new_n15193__ = ys__n18805 & ys__n37802;
  assign new_new_n15194__ = ~new_new_n15192__ & ~new_new_n15193__;
  assign new_new_n15195__ = ~ys__n18807 & ~ys__n37803;
  assign new_new_n15196__ = ys__n18807 & ys__n37803;
  assign new_new_n15197__ = ~new_new_n15195__ & ~new_new_n15196__;
  assign new_new_n15198__ = ~new_new_n15194__ & ~new_new_n15197__;
  assign new_new_n15199__ = ~ys__n18809 & ~ys__n37804;
  assign new_new_n15200__ = ys__n18809 & ys__n37804;
  assign new_new_n15201__ = ~new_new_n15199__ & ~new_new_n15200__;
  assign new_new_n15202__ = ~ys__n18811 & ~ys__n37805;
  assign new_new_n15203__ = ys__n18811 & ys__n37805;
  assign new_new_n15204__ = ~new_new_n15202__ & ~new_new_n15203__;
  assign new_new_n15205__ = ~new_new_n15201__ & ~new_new_n15204__;
  assign new_new_n15206__ = new_new_n15198__ & new_new_n15205__;
  assign new_new_n15207__ = new_new_n15191__ & new_new_n15206__;
  assign new_new_n15208__ = new_new_n15176__ & new_new_n15207__;
  assign new_new_n15209__ = ~ys__n18781 & ~ys__n37790;
  assign new_new_n15210__ = ys__n18781 & ys__n37790;
  assign new_new_n15211__ = ~new_new_n15209__ & ~new_new_n15210__;
  assign new_new_n15212__ = ~ys__n18783 & ~ys__n37791;
  assign new_new_n15213__ = ys__n18783 & ys__n37791;
  assign new_new_n15214__ = ~new_new_n15212__ & ~new_new_n15213__;
  assign new_new_n15215__ = ~new_new_n15211__ & ~new_new_n15214__;
  assign new_new_n15216__ = ~ys__n18785 & ~ys__n37792;
  assign new_new_n15217__ = ys__n18785 & ys__n37792;
  assign new_new_n15218__ = ~new_new_n15216__ & ~new_new_n15217__;
  assign new_new_n15219__ = ~ys__n18787 & ~ys__n37793;
  assign new_new_n15220__ = ys__n18787 & ys__n37793;
  assign new_new_n15221__ = ~new_new_n15219__ & ~new_new_n15220__;
  assign new_new_n15222__ = ~new_new_n15218__ & ~new_new_n15221__;
  assign new_new_n15223__ = new_new_n15215__ & new_new_n15222__;
  assign new_new_n15224__ = ~ys__n18773 & ~ys__n37786;
  assign new_new_n15225__ = ys__n18773 & ys__n37786;
  assign new_new_n15226__ = ~new_new_n15224__ & ~new_new_n15225__;
  assign new_new_n15227__ = ~ys__n18775 & ~ys__n37787;
  assign new_new_n15228__ = ys__n18775 & ys__n37787;
  assign new_new_n15229__ = ~new_new_n15227__ & ~new_new_n15228__;
  assign new_new_n15230__ = ~new_new_n15226__ & ~new_new_n15229__;
  assign new_new_n15231__ = ~ys__n18777 & ~ys__n37788;
  assign new_new_n15232__ = ys__n18777 & ys__n37788;
  assign new_new_n15233__ = ~new_new_n15231__ & ~new_new_n15232__;
  assign new_new_n15234__ = ~ys__n18779 & ~ys__n37789;
  assign new_new_n15235__ = ys__n18779 & ys__n37789;
  assign new_new_n15236__ = ~new_new_n15234__ & ~new_new_n15235__;
  assign new_new_n15237__ = ~new_new_n15233__ & ~new_new_n15236__;
  assign new_new_n15238__ = new_new_n15230__ & new_new_n15237__;
  assign new_new_n15239__ = new_new_n15223__ & new_new_n15238__;
  assign new_new_n15240__ = ~ys__n18797 & ~ys__n37798;
  assign new_new_n15241__ = ys__n18797 & ys__n37798;
  assign new_new_n15242__ = ~new_new_n15240__ & ~new_new_n15241__;
  assign new_new_n15243__ = ~ys__n18799 & ~ys__n37799;
  assign new_new_n15244__ = ys__n18799 & ys__n37799;
  assign new_new_n15245__ = ~new_new_n15243__ & ~new_new_n15244__;
  assign new_new_n15246__ = ~new_new_n15242__ & ~new_new_n15245__;
  assign new_new_n15247__ = ~ys__n18801 & ~ys__n37800;
  assign new_new_n15248__ = ys__n18801 & ys__n37800;
  assign new_new_n15249__ = ~new_new_n15247__ & ~new_new_n15248__;
  assign new_new_n15250__ = ~ys__n18803 & ~ys__n37801;
  assign new_new_n15251__ = ys__n18803 & ys__n37801;
  assign new_new_n15252__ = ~new_new_n15250__ & ~new_new_n15251__;
  assign new_new_n15253__ = ~new_new_n15249__ & ~new_new_n15252__;
  assign new_new_n15254__ = new_new_n15246__ & new_new_n15253__;
  assign new_new_n15255__ = ~ys__n18789 & ~ys__n37794;
  assign new_new_n15256__ = ys__n18789 & ys__n37794;
  assign new_new_n15257__ = ~new_new_n15255__ & ~new_new_n15256__;
  assign new_new_n15258__ = ~ys__n18791 & ~ys__n37795;
  assign new_new_n15259__ = ys__n18791 & ys__n37795;
  assign new_new_n15260__ = ~new_new_n15258__ & ~new_new_n15259__;
  assign new_new_n15261__ = ~new_new_n15257__ & ~new_new_n15260__;
  assign new_new_n15262__ = ~ys__n18793 & ~ys__n37796;
  assign new_new_n15263__ = ys__n18793 & ys__n37796;
  assign new_new_n15264__ = ~new_new_n15262__ & ~new_new_n15263__;
  assign new_new_n15265__ = ~ys__n18795 & ~ys__n37797;
  assign new_new_n15266__ = ys__n18795 & ys__n37797;
  assign new_new_n15267__ = ~new_new_n15265__ & ~new_new_n15266__;
  assign new_new_n15268__ = ~new_new_n15264__ & ~new_new_n15267__;
  assign new_new_n15269__ = new_new_n15261__ & new_new_n15268__;
  assign new_new_n15270__ = new_new_n15254__ & new_new_n15269__;
  assign new_new_n15271__ = new_new_n15239__ & new_new_n15270__;
  assign new_new_n15272__ = new_new_n15208__ & new_new_n15271__;
  assign new_new_n15273__ = ~ys__n37756 & ~new_new_n15272__;
  assign new_new_n15274__ = ys__n846 & ~new_new_n15273__;
  assign new_new_n15275__ = ~ys__n18821 & ~ys__n37782;
  assign new_new_n15276__ = ys__n18821 & ys__n37782;
  assign new_new_n15277__ = ~new_new_n15275__ & ~new_new_n15276__;
  assign new_new_n15278__ = ~ys__n18823 & ~ys__n37783;
  assign new_new_n15279__ = ys__n18823 & ys__n37783;
  assign new_new_n15280__ = ~new_new_n15278__ & ~new_new_n15279__;
  assign new_new_n15281__ = ~new_new_n15277__ & ~new_new_n15280__;
  assign new_new_n15282__ = ~ys__n18825 & ~ys__n37784;
  assign new_new_n15283__ = ys__n18825 & ys__n37784;
  assign new_new_n15284__ = ~new_new_n15282__ & ~new_new_n15283__;
  assign new_new_n15285__ = ~ys__n18827 & ~ys__n37785;
  assign new_new_n15286__ = ys__n18827 & ys__n37785;
  assign new_new_n15287__ = ~new_new_n15285__ & ~new_new_n15286__;
  assign new_new_n15288__ = ~new_new_n15284__ & ~new_new_n15287__;
  assign new_new_n15289__ = new_new_n15281__ & new_new_n15288__;
  assign new_new_n15290__ = ~ys__n18813 & ~ys__n37778;
  assign new_new_n15291__ = ys__n18813 & ys__n37778;
  assign new_new_n15292__ = ~new_new_n15290__ & ~new_new_n15291__;
  assign new_new_n15293__ = ~ys__n18815 & ~ys__n37779;
  assign new_new_n15294__ = ys__n18815 & ys__n37779;
  assign new_new_n15295__ = ~new_new_n15293__ & ~new_new_n15294__;
  assign new_new_n15296__ = ~new_new_n15292__ & ~new_new_n15295__;
  assign new_new_n15297__ = ~ys__n18817 & ~ys__n37780;
  assign new_new_n15298__ = ys__n18817 & ys__n37780;
  assign new_new_n15299__ = ~new_new_n15297__ & ~new_new_n15298__;
  assign new_new_n15300__ = ~ys__n18819 & ~ys__n37781;
  assign new_new_n15301__ = ys__n18819 & ys__n37781;
  assign new_new_n15302__ = ~new_new_n15300__ & ~new_new_n15301__;
  assign new_new_n15303__ = ~new_new_n15299__ & ~new_new_n15302__;
  assign new_new_n15304__ = new_new_n15296__ & new_new_n15303__;
  assign new_new_n15305__ = ~ys__n18805 & ~ys__n37774;
  assign new_new_n15306__ = ys__n18805 & ys__n37774;
  assign new_new_n15307__ = ~new_new_n15305__ & ~new_new_n15306__;
  assign new_new_n15308__ = ~ys__n18807 & ~ys__n37775;
  assign new_new_n15309__ = ys__n18807 & ys__n37775;
  assign new_new_n15310__ = ~new_new_n15308__ & ~new_new_n15309__;
  assign new_new_n15311__ = ~new_new_n15307__ & ~new_new_n15310__;
  assign new_new_n15312__ = ~ys__n18809 & ~ys__n37776;
  assign new_new_n15313__ = ys__n18809 & ys__n37776;
  assign new_new_n15314__ = ~new_new_n15312__ & ~new_new_n15313__;
  assign new_new_n15315__ = ~ys__n18811 & ~ys__n37777;
  assign new_new_n15316__ = ys__n18811 & ys__n37777;
  assign new_new_n15317__ = ~new_new_n15315__ & ~new_new_n15316__;
  assign new_new_n15318__ = ~new_new_n15314__ & ~new_new_n15317__;
  assign new_new_n15319__ = new_new_n15311__ & new_new_n15318__;
  assign new_new_n15320__ = new_new_n15304__ & new_new_n15319__;
  assign new_new_n15321__ = new_new_n15289__ & new_new_n15320__;
  assign new_new_n15322__ = ~ys__n18781 & ~ys__n37762;
  assign new_new_n15323__ = ys__n18781 & ys__n37762;
  assign new_new_n15324__ = ~new_new_n15322__ & ~new_new_n15323__;
  assign new_new_n15325__ = ~ys__n18783 & ~ys__n37763;
  assign new_new_n15326__ = ys__n18783 & ys__n37763;
  assign new_new_n15327__ = ~new_new_n15325__ & ~new_new_n15326__;
  assign new_new_n15328__ = ~new_new_n15324__ & ~new_new_n15327__;
  assign new_new_n15329__ = ~ys__n18785 & ~ys__n37764;
  assign new_new_n15330__ = ys__n18785 & ys__n37764;
  assign new_new_n15331__ = ~new_new_n15329__ & ~new_new_n15330__;
  assign new_new_n15332__ = ~ys__n18787 & ~ys__n37765;
  assign new_new_n15333__ = ys__n18787 & ys__n37765;
  assign new_new_n15334__ = ~new_new_n15332__ & ~new_new_n15333__;
  assign new_new_n15335__ = ~new_new_n15331__ & ~new_new_n15334__;
  assign new_new_n15336__ = new_new_n15328__ & new_new_n15335__;
  assign new_new_n15337__ = ~ys__n18773 & ~ys__n37758;
  assign new_new_n15338__ = ys__n18773 & ys__n37758;
  assign new_new_n15339__ = ~new_new_n15337__ & ~new_new_n15338__;
  assign new_new_n15340__ = ~ys__n18775 & ~ys__n37759;
  assign new_new_n15341__ = ys__n18775 & ys__n37759;
  assign new_new_n15342__ = ~new_new_n15340__ & ~new_new_n15341__;
  assign new_new_n15343__ = ~new_new_n15339__ & ~new_new_n15342__;
  assign new_new_n15344__ = ~ys__n18777 & ~ys__n37760;
  assign new_new_n15345__ = ys__n18777 & ys__n37760;
  assign new_new_n15346__ = ~new_new_n15344__ & ~new_new_n15345__;
  assign new_new_n15347__ = ~ys__n18779 & ~ys__n37761;
  assign new_new_n15348__ = ys__n18779 & ys__n37761;
  assign new_new_n15349__ = ~new_new_n15347__ & ~new_new_n15348__;
  assign new_new_n15350__ = ~new_new_n15346__ & ~new_new_n15349__;
  assign new_new_n15351__ = new_new_n15343__ & new_new_n15350__;
  assign new_new_n15352__ = new_new_n15336__ & new_new_n15351__;
  assign new_new_n15353__ = ~ys__n18797 & ~ys__n37770;
  assign new_new_n15354__ = ys__n18797 & ys__n37770;
  assign new_new_n15355__ = ~new_new_n15353__ & ~new_new_n15354__;
  assign new_new_n15356__ = ~ys__n18799 & ~ys__n37771;
  assign new_new_n15357__ = ys__n18799 & ys__n37771;
  assign new_new_n15358__ = ~new_new_n15356__ & ~new_new_n15357__;
  assign new_new_n15359__ = ~new_new_n15355__ & ~new_new_n15358__;
  assign new_new_n15360__ = ~ys__n18801 & ~ys__n37772;
  assign new_new_n15361__ = ys__n18801 & ys__n37772;
  assign new_new_n15362__ = ~new_new_n15360__ & ~new_new_n15361__;
  assign new_new_n15363__ = ~ys__n18803 & ~ys__n37773;
  assign new_new_n15364__ = ys__n18803 & ys__n37773;
  assign new_new_n15365__ = ~new_new_n15363__ & ~new_new_n15364__;
  assign new_new_n15366__ = ~new_new_n15362__ & ~new_new_n15365__;
  assign new_new_n15367__ = new_new_n15359__ & new_new_n15366__;
  assign new_new_n15368__ = ~ys__n18789 & ~ys__n37766;
  assign new_new_n15369__ = ys__n18789 & ys__n37766;
  assign new_new_n15370__ = ~new_new_n15368__ & ~new_new_n15369__;
  assign new_new_n15371__ = ~ys__n18791 & ~ys__n37767;
  assign new_new_n15372__ = ys__n18791 & ys__n37767;
  assign new_new_n15373__ = ~new_new_n15371__ & ~new_new_n15372__;
  assign new_new_n15374__ = ~new_new_n15370__ & ~new_new_n15373__;
  assign new_new_n15375__ = ~ys__n18793 & ~ys__n37768;
  assign new_new_n15376__ = ys__n18793 & ys__n37768;
  assign new_new_n15377__ = ~new_new_n15375__ & ~new_new_n15376__;
  assign new_new_n15378__ = ~ys__n18795 & ~ys__n37769;
  assign new_new_n15379__ = ys__n18795 & ys__n37769;
  assign new_new_n15380__ = ~new_new_n15378__ & ~new_new_n15379__;
  assign new_new_n15381__ = ~new_new_n15377__ & ~new_new_n15380__;
  assign new_new_n15382__ = new_new_n15374__ & new_new_n15381__;
  assign new_new_n15383__ = new_new_n15367__ & new_new_n15382__;
  assign new_new_n15384__ = new_new_n15352__ & new_new_n15383__;
  assign new_new_n15385__ = new_new_n15321__ & new_new_n15384__;
  assign new_new_n15386__ = ~ys__n37757 & ~new_new_n15385__;
  assign new_new_n15387__ = ys__n116 & ~new_new_n15386__;
  assign new_new_n15388__ = ~new_new_n15274__ & ~new_new_n15387__;
  assign new_new_n15389__ = new_new_n15161__ & new_new_n15388__;
  assign new_new_n15390__ = ~ys__n18821 & ~ys__n37978;
  assign new_new_n15391__ = ys__n18821 & ys__n37978;
  assign new_new_n15392__ = ~new_new_n15390__ & ~new_new_n15391__;
  assign new_new_n15393__ = ~ys__n18823 & ~ys__n37979;
  assign new_new_n15394__ = ys__n18823 & ys__n37979;
  assign new_new_n15395__ = ~new_new_n15393__ & ~new_new_n15394__;
  assign new_new_n15396__ = ~new_new_n15392__ & ~new_new_n15395__;
  assign new_new_n15397__ = ~ys__n18825 & ~ys__n37980;
  assign new_new_n15398__ = ys__n18825 & ys__n37980;
  assign new_new_n15399__ = ~new_new_n15397__ & ~new_new_n15398__;
  assign new_new_n15400__ = ~ys__n18827 & ~ys__n37981;
  assign new_new_n15401__ = ys__n18827 & ys__n37981;
  assign new_new_n15402__ = ~new_new_n15400__ & ~new_new_n15401__;
  assign new_new_n15403__ = ~new_new_n15399__ & ~new_new_n15402__;
  assign new_new_n15404__ = new_new_n15396__ & new_new_n15403__;
  assign new_new_n15405__ = ~ys__n18813 & ~ys__n37974;
  assign new_new_n15406__ = ys__n18813 & ys__n37974;
  assign new_new_n15407__ = ~new_new_n15405__ & ~new_new_n15406__;
  assign new_new_n15408__ = ~ys__n18815 & ~ys__n37975;
  assign new_new_n15409__ = ys__n18815 & ys__n37975;
  assign new_new_n15410__ = ~new_new_n15408__ & ~new_new_n15409__;
  assign new_new_n15411__ = ~new_new_n15407__ & ~new_new_n15410__;
  assign new_new_n15412__ = ~ys__n18817 & ~ys__n37976;
  assign new_new_n15413__ = ys__n18817 & ys__n37976;
  assign new_new_n15414__ = ~new_new_n15412__ & ~new_new_n15413__;
  assign new_new_n15415__ = ~ys__n18819 & ~ys__n37977;
  assign new_new_n15416__ = ys__n18819 & ys__n37977;
  assign new_new_n15417__ = ~new_new_n15415__ & ~new_new_n15416__;
  assign new_new_n15418__ = ~new_new_n15414__ & ~new_new_n15417__;
  assign new_new_n15419__ = new_new_n15411__ & new_new_n15418__;
  assign new_new_n15420__ = ~ys__n18805 & ~ys__n37970;
  assign new_new_n15421__ = ys__n18805 & ys__n37970;
  assign new_new_n15422__ = ~new_new_n15420__ & ~new_new_n15421__;
  assign new_new_n15423__ = ~ys__n18807 & ~ys__n37971;
  assign new_new_n15424__ = ys__n18807 & ys__n37971;
  assign new_new_n15425__ = ~new_new_n15423__ & ~new_new_n15424__;
  assign new_new_n15426__ = ~new_new_n15422__ & ~new_new_n15425__;
  assign new_new_n15427__ = ~ys__n18809 & ~ys__n37972;
  assign new_new_n15428__ = ys__n18809 & ys__n37972;
  assign new_new_n15429__ = ~new_new_n15427__ & ~new_new_n15428__;
  assign new_new_n15430__ = ~ys__n18811 & ~ys__n37973;
  assign new_new_n15431__ = ys__n18811 & ys__n37973;
  assign new_new_n15432__ = ~new_new_n15430__ & ~new_new_n15431__;
  assign new_new_n15433__ = ~new_new_n15429__ & ~new_new_n15432__;
  assign new_new_n15434__ = new_new_n15426__ & new_new_n15433__;
  assign new_new_n15435__ = new_new_n15419__ & new_new_n15434__;
  assign new_new_n15436__ = new_new_n15404__ & new_new_n15435__;
  assign new_new_n15437__ = ~ys__n18781 & ~ys__n37958;
  assign new_new_n15438__ = ys__n18781 & ys__n37958;
  assign new_new_n15439__ = ~new_new_n15437__ & ~new_new_n15438__;
  assign new_new_n15440__ = ~ys__n18783 & ~ys__n37959;
  assign new_new_n15441__ = ys__n18783 & ys__n37959;
  assign new_new_n15442__ = ~new_new_n15440__ & ~new_new_n15441__;
  assign new_new_n15443__ = ~new_new_n15439__ & ~new_new_n15442__;
  assign new_new_n15444__ = ~ys__n18785 & ~ys__n37960;
  assign new_new_n15445__ = ys__n18785 & ys__n37960;
  assign new_new_n15446__ = ~new_new_n15444__ & ~new_new_n15445__;
  assign new_new_n15447__ = ~ys__n18787 & ~ys__n37961;
  assign new_new_n15448__ = ys__n18787 & ys__n37961;
  assign new_new_n15449__ = ~new_new_n15447__ & ~new_new_n15448__;
  assign new_new_n15450__ = ~new_new_n15446__ & ~new_new_n15449__;
  assign new_new_n15451__ = new_new_n15443__ & new_new_n15450__;
  assign new_new_n15452__ = ~ys__n18773 & ~ys__n37954;
  assign new_new_n15453__ = ys__n18773 & ys__n37954;
  assign new_new_n15454__ = ~new_new_n15452__ & ~new_new_n15453__;
  assign new_new_n15455__ = ~ys__n18775 & ~ys__n37955;
  assign new_new_n15456__ = ys__n18775 & ys__n37955;
  assign new_new_n15457__ = ~new_new_n15455__ & ~new_new_n15456__;
  assign new_new_n15458__ = ~new_new_n15454__ & ~new_new_n15457__;
  assign new_new_n15459__ = ~ys__n18777 & ~ys__n37956;
  assign new_new_n15460__ = ys__n18777 & ys__n37956;
  assign new_new_n15461__ = ~new_new_n15459__ & ~new_new_n15460__;
  assign new_new_n15462__ = ~ys__n18779 & ~ys__n37957;
  assign new_new_n15463__ = ys__n18779 & ys__n37957;
  assign new_new_n15464__ = ~new_new_n15462__ & ~new_new_n15463__;
  assign new_new_n15465__ = ~new_new_n15461__ & ~new_new_n15464__;
  assign new_new_n15466__ = new_new_n15458__ & new_new_n15465__;
  assign new_new_n15467__ = new_new_n15451__ & new_new_n15466__;
  assign new_new_n15468__ = ~ys__n18797 & ~ys__n37966;
  assign new_new_n15469__ = ys__n18797 & ys__n37966;
  assign new_new_n15470__ = ~new_new_n15468__ & ~new_new_n15469__;
  assign new_new_n15471__ = ~ys__n18799 & ~ys__n37967;
  assign new_new_n15472__ = ys__n18799 & ys__n37967;
  assign new_new_n15473__ = ~new_new_n15471__ & ~new_new_n15472__;
  assign new_new_n15474__ = ~new_new_n15470__ & ~new_new_n15473__;
  assign new_new_n15475__ = ~ys__n18801 & ~ys__n37968;
  assign new_new_n15476__ = ys__n18801 & ys__n37968;
  assign new_new_n15477__ = ~new_new_n15475__ & ~new_new_n15476__;
  assign new_new_n15478__ = ~ys__n18803 & ~ys__n37969;
  assign new_new_n15479__ = ys__n18803 & ys__n37969;
  assign new_new_n15480__ = ~new_new_n15478__ & ~new_new_n15479__;
  assign new_new_n15481__ = ~new_new_n15477__ & ~new_new_n15480__;
  assign new_new_n15482__ = new_new_n15474__ & new_new_n15481__;
  assign new_new_n15483__ = ~ys__n18789 & ~ys__n37962;
  assign new_new_n15484__ = ys__n18789 & ys__n37962;
  assign new_new_n15485__ = ~new_new_n15483__ & ~new_new_n15484__;
  assign new_new_n15486__ = ~ys__n18791 & ~ys__n37963;
  assign new_new_n15487__ = ys__n18791 & ys__n37963;
  assign new_new_n15488__ = ~new_new_n15486__ & ~new_new_n15487__;
  assign new_new_n15489__ = ~new_new_n15485__ & ~new_new_n15488__;
  assign new_new_n15490__ = ~ys__n18793 & ~ys__n37964;
  assign new_new_n15491__ = ys__n18793 & ys__n37964;
  assign new_new_n15492__ = ~new_new_n15490__ & ~new_new_n15491__;
  assign new_new_n15493__ = ~ys__n18795 & ~ys__n37965;
  assign new_new_n15494__ = ys__n18795 & ys__n37965;
  assign new_new_n15495__ = ~new_new_n15493__ & ~new_new_n15494__;
  assign new_new_n15496__ = ~new_new_n15492__ & ~new_new_n15495__;
  assign new_new_n15497__ = new_new_n15489__ & new_new_n15496__;
  assign new_new_n15498__ = new_new_n15482__ & new_new_n15497__;
  assign new_new_n15499__ = new_new_n15467__ & new_new_n15498__;
  assign new_new_n15500__ = new_new_n15436__ & new_new_n15499__;
  assign new_new_n15501__ = ~ys__n37750 & ~new_new_n15500__;
  assign new_new_n15502__ = ys__n858 & ~new_new_n15501__;
  assign new_new_n15503__ = ~ys__n18821 & ~ys__n37950;
  assign new_new_n15504__ = ys__n18821 & ys__n37950;
  assign new_new_n15505__ = ~new_new_n15503__ & ~new_new_n15504__;
  assign new_new_n15506__ = ~ys__n18823 & ~ys__n37951;
  assign new_new_n15507__ = ys__n18823 & ys__n37951;
  assign new_new_n15508__ = ~new_new_n15506__ & ~new_new_n15507__;
  assign new_new_n15509__ = ~new_new_n15505__ & ~new_new_n15508__;
  assign new_new_n15510__ = ~ys__n18825 & ~ys__n37952;
  assign new_new_n15511__ = ys__n18825 & ys__n37952;
  assign new_new_n15512__ = ~new_new_n15510__ & ~new_new_n15511__;
  assign new_new_n15513__ = ~ys__n18827 & ~ys__n37953;
  assign new_new_n15514__ = ys__n18827 & ys__n37953;
  assign new_new_n15515__ = ~new_new_n15513__ & ~new_new_n15514__;
  assign new_new_n15516__ = ~new_new_n15512__ & ~new_new_n15515__;
  assign new_new_n15517__ = new_new_n15509__ & new_new_n15516__;
  assign new_new_n15518__ = ~ys__n18813 & ~ys__n37946;
  assign new_new_n15519__ = ys__n18813 & ys__n37946;
  assign new_new_n15520__ = ~new_new_n15518__ & ~new_new_n15519__;
  assign new_new_n15521__ = ~ys__n18815 & ~ys__n37947;
  assign new_new_n15522__ = ys__n18815 & ys__n37947;
  assign new_new_n15523__ = ~new_new_n15521__ & ~new_new_n15522__;
  assign new_new_n15524__ = ~new_new_n15520__ & ~new_new_n15523__;
  assign new_new_n15525__ = ~ys__n18817 & ~ys__n37948;
  assign new_new_n15526__ = ys__n18817 & ys__n37948;
  assign new_new_n15527__ = ~new_new_n15525__ & ~new_new_n15526__;
  assign new_new_n15528__ = ~ys__n18819 & ~ys__n37949;
  assign new_new_n15529__ = ys__n18819 & ys__n37949;
  assign new_new_n15530__ = ~new_new_n15528__ & ~new_new_n15529__;
  assign new_new_n15531__ = ~new_new_n15527__ & ~new_new_n15530__;
  assign new_new_n15532__ = new_new_n15524__ & new_new_n15531__;
  assign new_new_n15533__ = ~ys__n18805 & ~ys__n37942;
  assign new_new_n15534__ = ys__n18805 & ys__n37942;
  assign new_new_n15535__ = ~new_new_n15533__ & ~new_new_n15534__;
  assign new_new_n15536__ = ~ys__n18807 & ~ys__n37943;
  assign new_new_n15537__ = ys__n18807 & ys__n37943;
  assign new_new_n15538__ = ~new_new_n15536__ & ~new_new_n15537__;
  assign new_new_n15539__ = ~new_new_n15535__ & ~new_new_n15538__;
  assign new_new_n15540__ = ~ys__n18809 & ~ys__n37944;
  assign new_new_n15541__ = ys__n18809 & ys__n37944;
  assign new_new_n15542__ = ~new_new_n15540__ & ~new_new_n15541__;
  assign new_new_n15543__ = ~ys__n18811 & ~ys__n37945;
  assign new_new_n15544__ = ys__n18811 & ys__n37945;
  assign new_new_n15545__ = ~new_new_n15543__ & ~new_new_n15544__;
  assign new_new_n15546__ = ~new_new_n15542__ & ~new_new_n15545__;
  assign new_new_n15547__ = new_new_n15539__ & new_new_n15546__;
  assign new_new_n15548__ = new_new_n15532__ & new_new_n15547__;
  assign new_new_n15549__ = new_new_n15517__ & new_new_n15548__;
  assign new_new_n15550__ = ~ys__n18781 & ~ys__n37930;
  assign new_new_n15551__ = ys__n18781 & ys__n37930;
  assign new_new_n15552__ = ~new_new_n15550__ & ~new_new_n15551__;
  assign new_new_n15553__ = ~ys__n18783 & ~ys__n37931;
  assign new_new_n15554__ = ys__n18783 & ys__n37931;
  assign new_new_n15555__ = ~new_new_n15553__ & ~new_new_n15554__;
  assign new_new_n15556__ = ~new_new_n15552__ & ~new_new_n15555__;
  assign new_new_n15557__ = ~ys__n18785 & ~ys__n37932;
  assign new_new_n15558__ = ys__n18785 & ys__n37932;
  assign new_new_n15559__ = ~new_new_n15557__ & ~new_new_n15558__;
  assign new_new_n15560__ = ~ys__n18787 & ~ys__n37933;
  assign new_new_n15561__ = ys__n18787 & ys__n37933;
  assign new_new_n15562__ = ~new_new_n15560__ & ~new_new_n15561__;
  assign new_new_n15563__ = ~new_new_n15559__ & ~new_new_n15562__;
  assign new_new_n15564__ = new_new_n15556__ & new_new_n15563__;
  assign new_new_n15565__ = ~ys__n18773 & ~ys__n37926;
  assign new_new_n15566__ = ys__n18773 & ys__n37926;
  assign new_new_n15567__ = ~new_new_n15565__ & ~new_new_n15566__;
  assign new_new_n15568__ = ~ys__n18775 & ~ys__n37927;
  assign new_new_n15569__ = ys__n18775 & ys__n37927;
  assign new_new_n15570__ = ~new_new_n15568__ & ~new_new_n15569__;
  assign new_new_n15571__ = ~new_new_n15567__ & ~new_new_n15570__;
  assign new_new_n15572__ = ~ys__n18777 & ~ys__n37928;
  assign new_new_n15573__ = ys__n18777 & ys__n37928;
  assign new_new_n15574__ = ~new_new_n15572__ & ~new_new_n15573__;
  assign new_new_n15575__ = ~ys__n18779 & ~ys__n37929;
  assign new_new_n15576__ = ys__n18779 & ys__n37929;
  assign new_new_n15577__ = ~new_new_n15575__ & ~new_new_n15576__;
  assign new_new_n15578__ = ~new_new_n15574__ & ~new_new_n15577__;
  assign new_new_n15579__ = new_new_n15571__ & new_new_n15578__;
  assign new_new_n15580__ = new_new_n15564__ & new_new_n15579__;
  assign new_new_n15581__ = ~ys__n18797 & ~ys__n37938;
  assign new_new_n15582__ = ys__n18797 & ys__n37938;
  assign new_new_n15583__ = ~new_new_n15581__ & ~new_new_n15582__;
  assign new_new_n15584__ = ~ys__n18799 & ~ys__n37939;
  assign new_new_n15585__ = ys__n18799 & ys__n37939;
  assign new_new_n15586__ = ~new_new_n15584__ & ~new_new_n15585__;
  assign new_new_n15587__ = ~new_new_n15583__ & ~new_new_n15586__;
  assign new_new_n15588__ = ~ys__n18801 & ~ys__n37940;
  assign new_new_n15589__ = ys__n18801 & ys__n37940;
  assign new_new_n15590__ = ~new_new_n15588__ & ~new_new_n15589__;
  assign new_new_n15591__ = ~ys__n18803 & ~ys__n37941;
  assign new_new_n15592__ = ys__n18803 & ys__n37941;
  assign new_new_n15593__ = ~new_new_n15591__ & ~new_new_n15592__;
  assign new_new_n15594__ = ~new_new_n15590__ & ~new_new_n15593__;
  assign new_new_n15595__ = new_new_n15587__ & new_new_n15594__;
  assign new_new_n15596__ = ~ys__n18789 & ~ys__n37934;
  assign new_new_n15597__ = ys__n18789 & ys__n37934;
  assign new_new_n15598__ = ~new_new_n15596__ & ~new_new_n15597__;
  assign new_new_n15599__ = ~ys__n18791 & ~ys__n37935;
  assign new_new_n15600__ = ys__n18791 & ys__n37935;
  assign new_new_n15601__ = ~new_new_n15599__ & ~new_new_n15600__;
  assign new_new_n15602__ = ~new_new_n15598__ & ~new_new_n15601__;
  assign new_new_n15603__ = ~ys__n18793 & ~ys__n37936;
  assign new_new_n15604__ = ys__n18793 & ys__n37936;
  assign new_new_n15605__ = ~new_new_n15603__ & ~new_new_n15604__;
  assign new_new_n15606__ = ~ys__n18795 & ~ys__n37937;
  assign new_new_n15607__ = ys__n18795 & ys__n37937;
  assign new_new_n15608__ = ~new_new_n15606__ & ~new_new_n15607__;
  assign new_new_n15609__ = ~new_new_n15605__ & ~new_new_n15608__;
  assign new_new_n15610__ = new_new_n15602__ & new_new_n15609__;
  assign new_new_n15611__ = new_new_n15595__ & new_new_n15610__;
  assign new_new_n15612__ = new_new_n15580__ & new_new_n15611__;
  assign new_new_n15613__ = new_new_n15549__ & new_new_n15612__;
  assign new_new_n15614__ = ~ys__n37751 & ~new_new_n15613__;
  assign new_new_n15615__ = ys__n856 & ~new_new_n15614__;
  assign new_new_n15616__ = ~new_new_n15502__ & ~new_new_n15615__;
  assign new_new_n15617__ = ~ys__n18821 & ~ys__n37922;
  assign new_new_n15618__ = ys__n18821 & ys__n37922;
  assign new_new_n15619__ = ~new_new_n15617__ & ~new_new_n15618__;
  assign new_new_n15620__ = ~ys__n18823 & ~ys__n37923;
  assign new_new_n15621__ = ys__n18823 & ys__n37923;
  assign new_new_n15622__ = ~new_new_n15620__ & ~new_new_n15621__;
  assign new_new_n15623__ = ~new_new_n15619__ & ~new_new_n15622__;
  assign new_new_n15624__ = ~ys__n18825 & ~ys__n37924;
  assign new_new_n15625__ = ys__n18825 & ys__n37924;
  assign new_new_n15626__ = ~new_new_n15624__ & ~new_new_n15625__;
  assign new_new_n15627__ = ~ys__n18827 & ~ys__n37925;
  assign new_new_n15628__ = ys__n18827 & ys__n37925;
  assign new_new_n15629__ = ~new_new_n15627__ & ~new_new_n15628__;
  assign new_new_n15630__ = ~new_new_n15626__ & ~new_new_n15629__;
  assign new_new_n15631__ = new_new_n15623__ & new_new_n15630__;
  assign new_new_n15632__ = ~ys__n18813 & ~ys__n37918;
  assign new_new_n15633__ = ys__n18813 & ys__n37918;
  assign new_new_n15634__ = ~new_new_n15632__ & ~new_new_n15633__;
  assign new_new_n15635__ = ~ys__n18815 & ~ys__n37919;
  assign new_new_n15636__ = ys__n18815 & ys__n37919;
  assign new_new_n15637__ = ~new_new_n15635__ & ~new_new_n15636__;
  assign new_new_n15638__ = ~new_new_n15634__ & ~new_new_n15637__;
  assign new_new_n15639__ = ~ys__n18817 & ~ys__n37920;
  assign new_new_n15640__ = ys__n18817 & ys__n37920;
  assign new_new_n15641__ = ~new_new_n15639__ & ~new_new_n15640__;
  assign new_new_n15642__ = ~ys__n18819 & ~ys__n37921;
  assign new_new_n15643__ = ys__n18819 & ys__n37921;
  assign new_new_n15644__ = ~new_new_n15642__ & ~new_new_n15643__;
  assign new_new_n15645__ = ~new_new_n15641__ & ~new_new_n15644__;
  assign new_new_n15646__ = new_new_n15638__ & new_new_n15645__;
  assign new_new_n15647__ = ~ys__n18805 & ~ys__n37914;
  assign new_new_n15648__ = ys__n18805 & ys__n37914;
  assign new_new_n15649__ = ~new_new_n15647__ & ~new_new_n15648__;
  assign new_new_n15650__ = ~ys__n18807 & ~ys__n37915;
  assign new_new_n15651__ = ys__n18807 & ys__n37915;
  assign new_new_n15652__ = ~new_new_n15650__ & ~new_new_n15651__;
  assign new_new_n15653__ = ~new_new_n15649__ & ~new_new_n15652__;
  assign new_new_n15654__ = ~ys__n18809 & ~ys__n37916;
  assign new_new_n15655__ = ys__n18809 & ys__n37916;
  assign new_new_n15656__ = ~new_new_n15654__ & ~new_new_n15655__;
  assign new_new_n15657__ = ~ys__n18811 & ~ys__n37917;
  assign new_new_n15658__ = ys__n18811 & ys__n37917;
  assign new_new_n15659__ = ~new_new_n15657__ & ~new_new_n15658__;
  assign new_new_n15660__ = ~new_new_n15656__ & ~new_new_n15659__;
  assign new_new_n15661__ = new_new_n15653__ & new_new_n15660__;
  assign new_new_n15662__ = new_new_n15646__ & new_new_n15661__;
  assign new_new_n15663__ = new_new_n15631__ & new_new_n15662__;
  assign new_new_n15664__ = ~ys__n18781 & ~ys__n37902;
  assign new_new_n15665__ = ys__n18781 & ys__n37902;
  assign new_new_n15666__ = ~new_new_n15664__ & ~new_new_n15665__;
  assign new_new_n15667__ = ~ys__n18783 & ~ys__n37903;
  assign new_new_n15668__ = ys__n18783 & ys__n37903;
  assign new_new_n15669__ = ~new_new_n15667__ & ~new_new_n15668__;
  assign new_new_n15670__ = ~new_new_n15666__ & ~new_new_n15669__;
  assign new_new_n15671__ = ~ys__n18785 & ~ys__n37904;
  assign new_new_n15672__ = ys__n18785 & ys__n37904;
  assign new_new_n15673__ = ~new_new_n15671__ & ~new_new_n15672__;
  assign new_new_n15674__ = ~ys__n18787 & ~ys__n37905;
  assign new_new_n15675__ = ys__n18787 & ys__n37905;
  assign new_new_n15676__ = ~new_new_n15674__ & ~new_new_n15675__;
  assign new_new_n15677__ = ~new_new_n15673__ & ~new_new_n15676__;
  assign new_new_n15678__ = new_new_n15670__ & new_new_n15677__;
  assign new_new_n15679__ = ~ys__n18773 & ~ys__n37898;
  assign new_new_n15680__ = ys__n18773 & ys__n37898;
  assign new_new_n15681__ = ~new_new_n15679__ & ~new_new_n15680__;
  assign new_new_n15682__ = ~ys__n18775 & ~ys__n37899;
  assign new_new_n15683__ = ys__n18775 & ys__n37899;
  assign new_new_n15684__ = ~new_new_n15682__ & ~new_new_n15683__;
  assign new_new_n15685__ = ~new_new_n15681__ & ~new_new_n15684__;
  assign new_new_n15686__ = ~ys__n18777 & ~ys__n37900;
  assign new_new_n15687__ = ys__n18777 & ys__n37900;
  assign new_new_n15688__ = ~new_new_n15686__ & ~new_new_n15687__;
  assign new_new_n15689__ = ~ys__n18779 & ~ys__n37901;
  assign new_new_n15690__ = ys__n18779 & ys__n37901;
  assign new_new_n15691__ = ~new_new_n15689__ & ~new_new_n15690__;
  assign new_new_n15692__ = ~new_new_n15688__ & ~new_new_n15691__;
  assign new_new_n15693__ = new_new_n15685__ & new_new_n15692__;
  assign new_new_n15694__ = new_new_n15678__ & new_new_n15693__;
  assign new_new_n15695__ = ~ys__n18797 & ~ys__n37910;
  assign new_new_n15696__ = ys__n18797 & ys__n37910;
  assign new_new_n15697__ = ~new_new_n15695__ & ~new_new_n15696__;
  assign new_new_n15698__ = ~ys__n18799 & ~ys__n37911;
  assign new_new_n15699__ = ys__n18799 & ys__n37911;
  assign new_new_n15700__ = ~new_new_n15698__ & ~new_new_n15699__;
  assign new_new_n15701__ = ~new_new_n15697__ & ~new_new_n15700__;
  assign new_new_n15702__ = ~ys__n18801 & ~ys__n37912;
  assign new_new_n15703__ = ys__n18801 & ys__n37912;
  assign new_new_n15704__ = ~new_new_n15702__ & ~new_new_n15703__;
  assign new_new_n15705__ = ~ys__n18803 & ~ys__n37913;
  assign new_new_n15706__ = ys__n18803 & ys__n37913;
  assign new_new_n15707__ = ~new_new_n15705__ & ~new_new_n15706__;
  assign new_new_n15708__ = ~new_new_n15704__ & ~new_new_n15707__;
  assign new_new_n15709__ = new_new_n15701__ & new_new_n15708__;
  assign new_new_n15710__ = ~ys__n18789 & ~ys__n37906;
  assign new_new_n15711__ = ys__n18789 & ys__n37906;
  assign new_new_n15712__ = ~new_new_n15710__ & ~new_new_n15711__;
  assign new_new_n15713__ = ~ys__n18791 & ~ys__n37907;
  assign new_new_n15714__ = ys__n18791 & ys__n37907;
  assign new_new_n15715__ = ~new_new_n15713__ & ~new_new_n15714__;
  assign new_new_n15716__ = ~new_new_n15712__ & ~new_new_n15715__;
  assign new_new_n15717__ = ~ys__n18793 & ~ys__n37908;
  assign new_new_n15718__ = ys__n18793 & ys__n37908;
  assign new_new_n15719__ = ~new_new_n15717__ & ~new_new_n15718__;
  assign new_new_n15720__ = ~ys__n18795 & ~ys__n37909;
  assign new_new_n15721__ = ys__n18795 & ys__n37909;
  assign new_new_n15722__ = ~new_new_n15720__ & ~new_new_n15721__;
  assign new_new_n15723__ = ~new_new_n15719__ & ~new_new_n15722__;
  assign new_new_n15724__ = new_new_n15716__ & new_new_n15723__;
  assign new_new_n15725__ = new_new_n15709__ & new_new_n15724__;
  assign new_new_n15726__ = new_new_n15694__ & new_new_n15725__;
  assign new_new_n15727__ = new_new_n15663__ & new_new_n15726__;
  assign new_new_n15728__ = ~ys__n37752 & ~new_new_n15727__;
  assign new_new_n15729__ = ys__n854 & ~new_new_n15728__;
  assign new_new_n15730__ = ~ys__n18821 & ~ys__n37894;
  assign new_new_n15731__ = ys__n18821 & ys__n37894;
  assign new_new_n15732__ = ~new_new_n15730__ & ~new_new_n15731__;
  assign new_new_n15733__ = ~ys__n18823 & ~ys__n37895;
  assign new_new_n15734__ = ys__n18823 & ys__n37895;
  assign new_new_n15735__ = ~new_new_n15733__ & ~new_new_n15734__;
  assign new_new_n15736__ = ~new_new_n15732__ & ~new_new_n15735__;
  assign new_new_n15737__ = ~ys__n18825 & ~ys__n37896;
  assign new_new_n15738__ = ys__n18825 & ys__n37896;
  assign new_new_n15739__ = ~new_new_n15737__ & ~new_new_n15738__;
  assign new_new_n15740__ = ~ys__n18827 & ~ys__n37897;
  assign new_new_n15741__ = ys__n18827 & ys__n37897;
  assign new_new_n15742__ = ~new_new_n15740__ & ~new_new_n15741__;
  assign new_new_n15743__ = ~new_new_n15739__ & ~new_new_n15742__;
  assign new_new_n15744__ = new_new_n15736__ & new_new_n15743__;
  assign new_new_n15745__ = ~ys__n18813 & ~ys__n37890;
  assign new_new_n15746__ = ys__n18813 & ys__n37890;
  assign new_new_n15747__ = ~new_new_n15745__ & ~new_new_n15746__;
  assign new_new_n15748__ = ~ys__n18815 & ~ys__n37891;
  assign new_new_n15749__ = ys__n18815 & ys__n37891;
  assign new_new_n15750__ = ~new_new_n15748__ & ~new_new_n15749__;
  assign new_new_n15751__ = ~new_new_n15747__ & ~new_new_n15750__;
  assign new_new_n15752__ = ~ys__n18817 & ~ys__n37892;
  assign new_new_n15753__ = ys__n18817 & ys__n37892;
  assign new_new_n15754__ = ~new_new_n15752__ & ~new_new_n15753__;
  assign new_new_n15755__ = ~ys__n18819 & ~ys__n37893;
  assign new_new_n15756__ = ys__n18819 & ys__n37893;
  assign new_new_n15757__ = ~new_new_n15755__ & ~new_new_n15756__;
  assign new_new_n15758__ = ~new_new_n15754__ & ~new_new_n15757__;
  assign new_new_n15759__ = new_new_n15751__ & new_new_n15758__;
  assign new_new_n15760__ = ~ys__n18805 & ~ys__n37886;
  assign new_new_n15761__ = ys__n18805 & ys__n37886;
  assign new_new_n15762__ = ~new_new_n15760__ & ~new_new_n15761__;
  assign new_new_n15763__ = ~ys__n18807 & ~ys__n37887;
  assign new_new_n15764__ = ys__n18807 & ys__n37887;
  assign new_new_n15765__ = ~new_new_n15763__ & ~new_new_n15764__;
  assign new_new_n15766__ = ~new_new_n15762__ & ~new_new_n15765__;
  assign new_new_n15767__ = ~ys__n18809 & ~ys__n37888;
  assign new_new_n15768__ = ys__n18809 & ys__n37888;
  assign new_new_n15769__ = ~new_new_n15767__ & ~new_new_n15768__;
  assign new_new_n15770__ = ~ys__n18811 & ~ys__n37889;
  assign new_new_n15771__ = ys__n18811 & ys__n37889;
  assign new_new_n15772__ = ~new_new_n15770__ & ~new_new_n15771__;
  assign new_new_n15773__ = ~new_new_n15769__ & ~new_new_n15772__;
  assign new_new_n15774__ = new_new_n15766__ & new_new_n15773__;
  assign new_new_n15775__ = new_new_n15759__ & new_new_n15774__;
  assign new_new_n15776__ = new_new_n15744__ & new_new_n15775__;
  assign new_new_n15777__ = ~ys__n18781 & ~ys__n37874;
  assign new_new_n15778__ = ys__n18781 & ys__n37874;
  assign new_new_n15779__ = ~new_new_n15777__ & ~new_new_n15778__;
  assign new_new_n15780__ = ~ys__n18783 & ~ys__n37875;
  assign new_new_n15781__ = ys__n18783 & ys__n37875;
  assign new_new_n15782__ = ~new_new_n15780__ & ~new_new_n15781__;
  assign new_new_n15783__ = ~new_new_n15779__ & ~new_new_n15782__;
  assign new_new_n15784__ = ~ys__n18785 & ~ys__n37876;
  assign new_new_n15785__ = ys__n18785 & ys__n37876;
  assign new_new_n15786__ = ~new_new_n15784__ & ~new_new_n15785__;
  assign new_new_n15787__ = ~ys__n18787 & ~ys__n37877;
  assign new_new_n15788__ = ys__n18787 & ys__n37877;
  assign new_new_n15789__ = ~new_new_n15787__ & ~new_new_n15788__;
  assign new_new_n15790__ = ~new_new_n15786__ & ~new_new_n15789__;
  assign new_new_n15791__ = new_new_n15783__ & new_new_n15790__;
  assign new_new_n15792__ = ~ys__n18773 & ~ys__n37870;
  assign new_new_n15793__ = ys__n18773 & ys__n37870;
  assign new_new_n15794__ = ~new_new_n15792__ & ~new_new_n15793__;
  assign new_new_n15795__ = ~ys__n18775 & ~ys__n37871;
  assign new_new_n15796__ = ys__n18775 & ys__n37871;
  assign new_new_n15797__ = ~new_new_n15795__ & ~new_new_n15796__;
  assign new_new_n15798__ = ~new_new_n15794__ & ~new_new_n15797__;
  assign new_new_n15799__ = ~ys__n18777 & ~ys__n37872;
  assign new_new_n15800__ = ys__n18777 & ys__n37872;
  assign new_new_n15801__ = ~new_new_n15799__ & ~new_new_n15800__;
  assign new_new_n15802__ = ~ys__n18779 & ~ys__n37873;
  assign new_new_n15803__ = ys__n18779 & ys__n37873;
  assign new_new_n15804__ = ~new_new_n15802__ & ~new_new_n15803__;
  assign new_new_n15805__ = ~new_new_n15801__ & ~new_new_n15804__;
  assign new_new_n15806__ = new_new_n15798__ & new_new_n15805__;
  assign new_new_n15807__ = new_new_n15791__ & new_new_n15806__;
  assign new_new_n15808__ = ~ys__n18797 & ~ys__n37882;
  assign new_new_n15809__ = ys__n18797 & ys__n37882;
  assign new_new_n15810__ = ~new_new_n15808__ & ~new_new_n15809__;
  assign new_new_n15811__ = ~ys__n18799 & ~ys__n37883;
  assign new_new_n15812__ = ys__n18799 & ys__n37883;
  assign new_new_n15813__ = ~new_new_n15811__ & ~new_new_n15812__;
  assign new_new_n15814__ = ~new_new_n15810__ & ~new_new_n15813__;
  assign new_new_n15815__ = ~ys__n18801 & ~ys__n37884;
  assign new_new_n15816__ = ys__n18801 & ys__n37884;
  assign new_new_n15817__ = ~new_new_n15815__ & ~new_new_n15816__;
  assign new_new_n15818__ = ~ys__n18803 & ~ys__n37885;
  assign new_new_n15819__ = ys__n18803 & ys__n37885;
  assign new_new_n15820__ = ~new_new_n15818__ & ~new_new_n15819__;
  assign new_new_n15821__ = ~new_new_n15817__ & ~new_new_n15820__;
  assign new_new_n15822__ = new_new_n15814__ & new_new_n15821__;
  assign new_new_n15823__ = ~ys__n18789 & ~ys__n37878;
  assign new_new_n15824__ = ys__n18789 & ys__n37878;
  assign new_new_n15825__ = ~new_new_n15823__ & ~new_new_n15824__;
  assign new_new_n15826__ = ~ys__n18791 & ~ys__n37879;
  assign new_new_n15827__ = ys__n18791 & ys__n37879;
  assign new_new_n15828__ = ~new_new_n15826__ & ~new_new_n15827__;
  assign new_new_n15829__ = ~new_new_n15825__ & ~new_new_n15828__;
  assign new_new_n15830__ = ~ys__n18793 & ~ys__n37880;
  assign new_new_n15831__ = ys__n18793 & ys__n37880;
  assign new_new_n15832__ = ~new_new_n15830__ & ~new_new_n15831__;
  assign new_new_n15833__ = ~ys__n18795 & ~ys__n37881;
  assign new_new_n15834__ = ys__n18795 & ys__n37881;
  assign new_new_n15835__ = ~new_new_n15833__ & ~new_new_n15834__;
  assign new_new_n15836__ = ~new_new_n15832__ & ~new_new_n15835__;
  assign new_new_n15837__ = new_new_n15829__ & new_new_n15836__;
  assign new_new_n15838__ = new_new_n15822__ & new_new_n15837__;
  assign new_new_n15839__ = new_new_n15807__ & new_new_n15838__;
  assign new_new_n15840__ = new_new_n15776__ & new_new_n15839__;
  assign new_new_n15841__ = ~ys__n37753 & ~new_new_n15840__;
  assign new_new_n15842__ = ys__n852 & ~new_new_n15841__;
  assign new_new_n15843__ = ~new_new_n15729__ & ~new_new_n15842__;
  assign new_new_n15844__ = new_new_n15616__ & new_new_n15843__;
  assign new_new_n15845__ = new_new_n15389__ & new_new_n15844__;
  assign ys__n3249 = ~new_new_n14934__ | ~new_new_n15845__;
  assign new_new_n15847__ = ys__n18978 & ys__n18287;
  assign new_new_n15848__ = ~ys__n18284 & new_new_n15847__;
  assign new_new_n15849__ = ys__n24659 & ~ys__n4764;
  assign new_new_n15850__ = ys__n24660 & ys__n4764;
  assign ys__n18808 = new_new_n15849__ | new_new_n15850__;
  assign new_new_n15852__ = ~ys__n18071 & ys__n18808;
  assign new_new_n15853__ = ys__n18071 & ys__n18809;
  assign new_new_n15854__ = ~new_new_n15852__ & ~new_new_n15853__;
  assign new_new_n15855__ = ~new_new_n11122__ & ~new_new_n15854__;
  assign new_new_n15856__ = ys__n24660 & ~ys__n24675;
  assign new_new_n15857__ = ys__n24675 & ys__n24701;
  assign ys__n18720 = new_new_n15856__ | new_new_n15857__;
  assign new_new_n15859__ = new_new_n11122__ & ys__n18720;
  assign ys__n18721 = new_new_n15855__ | new_new_n15859__;
  assign new_new_n15861__ = ys__n18284 & ys__n18721;
  assign new_new_n15862__ = ~new_new_n15848__ & ~new_new_n15861__;
  assign new_new_n15863__ = ~ys__n18281 & ~new_new_n15862__;
  assign new_new_n15864__ = ys__n18622 & ~new_new_n11125__;
  assign new_new_n15865__ = ys__n18623 & new_new_n11125__;
  assign ys__n18624 = new_new_n15864__ | new_new_n15865__;
  assign new_new_n15867__ = ys__n18281 & ys__n18624;
  assign new_new_n15868__ = ~new_new_n15863__ & ~new_new_n15867__;
  assign new_new_n15869__ = ~ys__n18278 & ~new_new_n15868__;
  assign new_new_n15870__ = ys__n18873 & ys__n18278;
  assign ys__n3250 = new_new_n15869__ | new_new_n15870__;
  assign new_new_n15872__ = ys__n18979 & ys__n18287;
  assign new_new_n15873__ = ~ys__n18284 & new_new_n15872__;
  assign new_new_n15874__ = ys__n24661 & ~ys__n4764;
  assign new_new_n15875__ = ys__n24662 & ys__n4764;
  assign ys__n18810 = new_new_n15874__ | new_new_n15875__;
  assign new_new_n15877__ = ~ys__n18071 & ys__n18810;
  assign new_new_n15878__ = ys__n18071 & ys__n18811;
  assign new_new_n15879__ = ~new_new_n15877__ & ~new_new_n15878__;
  assign new_new_n15880__ = ~new_new_n11122__ & ~new_new_n15879__;
  assign new_new_n15881__ = ys__n24662 & ~ys__n24675;
  assign new_new_n15882__ = ys__n24675 & ys__n24702;
  assign ys__n18723 = new_new_n15881__ | new_new_n15882__;
  assign new_new_n15884__ = new_new_n11122__ & ys__n18723;
  assign ys__n18724 = new_new_n15880__ | new_new_n15884__;
  assign new_new_n15886__ = ys__n18284 & ys__n18724;
  assign new_new_n15887__ = ~new_new_n15873__ & ~new_new_n15886__;
  assign new_new_n15888__ = ~ys__n18281 & ~new_new_n15887__;
  assign new_new_n15889__ = ys__n18625 & ~new_new_n11125__;
  assign new_new_n15890__ = ys__n18626 & new_new_n11125__;
  assign ys__n18627 = new_new_n15889__ | new_new_n15890__;
  assign new_new_n15892__ = ys__n18281 & ys__n18627;
  assign new_new_n15893__ = ~new_new_n15888__ & ~new_new_n15892__;
  assign new_new_n15894__ = ~ys__n18278 & ~new_new_n15893__;
  assign new_new_n15895__ = ys__n18875 & ys__n18278;
  assign ys__n3252 = new_new_n15894__ | new_new_n15895__;
  assign new_new_n15897__ = ~ys__n846 & new_new_n11047__;
  assign new_new_n15898__ = new_new_n12223__ & new_new_n15897__;
  assign ys__n4189 = ~new_new_n12227__ | ~new_new_n15898__;
  assign new_new_n15900__ = ~ys__n776 & ~ys__n4168;
  assign new_new_n15901__ = ~ys__n604 & ~ys__n778;
  assign new_new_n15902__ = new_new_n15900__ & new_new_n15901__;
  assign new_new_n15903__ = ~ys__n698 & ~ys__n768;
  assign new_new_n15904__ = new_new_n13930__ & new_new_n15903__;
  assign new_new_n15905__ = new_new_n15902__ & new_new_n15904__;
  assign new_new_n15906__ = new_new_n13933__ & new_new_n13934__;
  assign new_new_n15907__ = ys__n772 & new_new_n15906__;
  assign new_new_n15908__ = new_new_n15905__ & new_new_n15907__;
  assign new_new_n15909__ = ~ys__n598 & ys__n774;
  assign new_new_n15910__ = new_new_n15905__ & new_new_n15909__;
  assign new_new_n15911__ = ys__n770 & ~ys__n784;
  assign new_new_n15912__ = new_new_n13933__ & new_new_n15911__;
  assign new_new_n15913__ = new_new_n15905__ & new_new_n15912__;
  assign new_new_n15914__ = ~new_new_n15910__ & ~new_new_n15913__;
  assign new_new_n15915__ = ~new_new_n15908__ & new_new_n15914__;
  assign new_new_n15916__ = ~ys__n772 & ~ys__n780;
  assign new_new_n15917__ = ys__n782 & new_new_n15916__;
  assign new_new_n15918__ = new_new_n15906__ & new_new_n15917__;
  assign new_new_n15919__ = new_new_n15905__ & new_new_n15918__;
  assign new_new_n15920__ = ~ys__n772 & ys__n780;
  assign new_new_n15921__ = new_new_n15906__ & new_new_n15920__;
  assign new_new_n15922__ = new_new_n15905__ & new_new_n15921__;
  assign new_new_n15923__ = ~new_new_n15919__ & ~new_new_n15922__;
  assign new_new_n15924__ = ~ys__n782 & ~ys__n2644;
  assign new_new_n15925__ = new_new_n15916__ & new_new_n15924__;
  assign new_new_n15926__ = new_new_n15906__ & new_new_n15925__;
  assign new_new_n15927__ = new_new_n15905__ & new_new_n15926__;
  assign new_new_n15928__ = ys__n598 & new_new_n15905__;
  assign new_new_n15929__ = ~new_new_n15927__ & ~new_new_n15928__;
  assign new_new_n15930__ = new_new_n15923__ & new_new_n15929__;
  assign new_new_n15931__ = ys__n602 & new_new_n15902__;
  assign new_new_n15932__ = ys__n698 & new_new_n13930__;
  assign new_new_n15933__ = new_new_n15902__ & new_new_n15932__;
  assign new_new_n15934__ = ~new_new_n15931__ & ~new_new_n15933__;
  assign new_new_n15935__ = ys__n600 & ~ys__n602;
  assign new_new_n15936__ = new_new_n15902__ & new_new_n15935__;
  assign new_new_n15937__ = ~ys__n698 & ys__n768;
  assign new_new_n15938__ = new_new_n13930__ & new_new_n15937__;
  assign new_new_n15939__ = new_new_n15902__ & new_new_n15938__;
  assign new_new_n15940__ = ~new_new_n15936__ & ~new_new_n15939__;
  assign new_new_n15941__ = new_new_n15934__ & new_new_n15940__;
  assign new_new_n15942__ = ys__n784 & new_new_n13933__;
  assign new_new_n15943__ = new_new_n15905__ & new_new_n15942__;
  assign new_new_n15944__ = ys__n604 & new_new_n15900__;
  assign new_new_n15945__ = ~ys__n604 & ys__n778;
  assign new_new_n15946__ = new_new_n15900__ & new_new_n15945__;
  assign new_new_n15947__ = ys__n776 & ~ys__n4168;
  assign new_new_n15948__ = ~new_new_n15946__ & ~new_new_n15947__;
  assign new_new_n15949__ = ~new_new_n15944__ & new_new_n15948__;
  assign new_new_n15950__ = ~new_new_n15943__ & new_new_n15949__;
  assign new_new_n15951__ = new_new_n15941__ & new_new_n15950__;
  assign new_new_n15952__ = new_new_n15930__ & new_new_n15951__;
  assign ys__n4320 = new_new_n15915__ & new_new_n15952__;
  assign ys__n4414 = ~ys__n18271 & ~new_new_n11130__;
  assign ys__n4521 = ~ys__n740 | new_new_n12188__;
  assign new_new_n15956__ = new_new_n11193__ & ~new_new_n11230__;
  assign new_new_n15957__ = ~new_new_n11203__ & ~new_new_n11205__;
  assign new_new_n15958__ = ~ys__n530 & ~ys__n752;
  assign new_new_n15959__ = ~ys__n526 & ys__n528;
  assign new_new_n15960__ = ys__n522 & ~ys__n524;
  assign new_new_n15961__ = new_new_n15959__ & new_new_n15960__;
  assign new_new_n15962__ = new_new_n15958__ & new_new_n15961__;
  assign new_new_n15963__ = new_new_n10632__ & new_new_n10657__;
  assign new_new_n15964__ = new_new_n15962__ & new_new_n15963__;
  assign new_new_n15965__ = new_new_n15957__ & ~new_new_n15964__;
  assign new_new_n15966__ = ~new_new_n15956__ & new_new_n15965__;
  assign new_new_n15967__ = ~new_new_n11193__ & ~new_new_n15963__;
  assign new_new_n15968__ = new_new_n15957__ & new_new_n15967__;
  assign new_new_n15969__ = ~ys__n28243 & ~new_new_n15968__;
  assign new_new_n15970__ = ~new_new_n15966__ & new_new_n15969__;
  assign new_new_n15971__ = new_new_n11250__ & new_new_n11260__;
  assign new_new_n15972__ = ys__n736 & ~ys__n752;
  assign new_new_n15973__ = ~ys__n4488 & ~ys__n23730;
  assign new_new_n15974__ = new_new_n15972__ & new_new_n15973__;
  assign new_new_n15975__ = new_new_n15971__ & new_new_n15974__;
  assign new_new_n15976__ = ~ys__n23730 & ~new_new_n15975__;
  assign new_new_n15977__ = ys__n28243 & ~new_new_n15976__;
  assign new_new_n15978__ = ~new_new_n15970__ & ~new_new_n15977__;
  assign ys__n4588 = ~ys__n738 & ~new_new_n15978__;
  assign new_new_n15980__ = ~ys__n23627 & ys__n23629;
  assign new_new_n15981__ = ~new_new_n11175__ & new_new_n15980__;
  assign new_new_n15982__ = ys__n22882 & new_new_n11175__;
  assign new_new_n15983__ = ~new_new_n15981__ & ~new_new_n15982__;
  assign new_new_n15984__ = ~new_new_n11180__ & ~new_new_n15983__;
  assign new_new_n15985__ = ys__n23330 & new_new_n11180__;
  assign new_new_n15986__ = ~new_new_n15984__ & ~new_new_n15985__;
  assign new_new_n15987__ = ~new_new_n11186__ & ~new_new_n15986__;
  assign new_new_n15988__ = ys__n424 & new_new_n11186__;
  assign new_new_n15989__ = ~new_new_n15987__ & ~new_new_n15988__;
  assign new_new_n15990__ = ~new_new_n11270__ & ~new_new_n15989__;
  assign new_new_n15991__ = ys__n424 & ~new_new_n11292__;
  assign new_new_n15992__ = ~ys__n424 & new_new_n11664__;
  assign new_new_n15993__ = ys__n424 & ~new_new_n11664__;
  assign new_new_n15994__ = ~new_new_n15992__ & ~new_new_n15993__;
  assign new_new_n15995__ = new_new_n11292__ & ~new_new_n15994__;
  assign ys__n23541 = new_new_n15991__ | new_new_n15995__;
  assign new_new_n15997__ = new_new_n11270__ & ys__n23541;
  assign new_new_n15998__ = ~new_new_n15990__ & ~new_new_n15997__;
  assign new_new_n15999__ = new_new_n11324__ & ~new_new_n15998__;
  assign new_new_n16000__ = ys__n424 & ~new_new_n11324__;
  assign new_new_n16001__ = ~new_new_n15999__ & ~new_new_n16000__;
  assign new_new_n16002__ = ~new_new_n11343__ & ~new_new_n16001__;
  assign new_new_n16003__ = ys__n424 & ~new_new_n11569__;
  assign new_new_n16004__ = ~ys__n450 & ~new_new_n11599__;
  assign new_new_n16005__ = ~ys__n450 & ~new_new_n16004__;
  assign new_new_n16006__ = ys__n424 & ~new_new_n16005__;
  assign new_new_n16007__ = ~ys__n424 & new_new_n16005__;
  assign new_new_n16008__ = ~new_new_n16006__ & ~new_new_n16007__;
  assign new_new_n16009__ = new_new_n11603__ & ~new_new_n16008__;
  assign new_new_n16010__ = ys__n450 & new_new_n11615__;
  assign new_new_n16011__ = ~ys__n424 & new_new_n16010__;
  assign new_new_n16012__ = ys__n424 & ~new_new_n16010__;
  assign new_new_n16013__ = ~new_new_n16011__ & ~new_new_n16012__;
  assign new_new_n16014__ = new_new_n11619__ & ~new_new_n16013__;
  assign new_new_n16015__ = ~new_new_n16009__ & ~new_new_n16014__;
  assign new_new_n16016__ = ~new_new_n16003__ & new_new_n16015__;
  assign new_new_n16017__ = new_new_n11625__ & ~new_new_n16016__;
  assign new_new_n16018__ = ~new_new_n16002__ & ~new_new_n16017__;
  assign new_new_n16019__ = new_new_n11629__ & ~new_new_n16018__;
  assign new_new_n16020__ = ys__n935 & ys__n23629;
  assign new_new_n16021__ = new_new_n11628__ & new_new_n16020__;
  assign new_new_n16022__ = ys__n47691 & new_new_n11634__;
  assign new_new_n16023__ = ~new_new_n16021__ & ~new_new_n16022__;
  assign new_new_n16024__ = ~new_new_n16019__ & new_new_n16023__;
  assign new_new_n16025__ = new_new_n11640__ & ~new_new_n16024__;
  assign new_new_n16026__ = new_new_n11642__ & ~new_new_n16018__;
  assign new_new_n16027__ = ys__n47691 & new_new_n11644__;
  assign new_new_n16028__ = ~new_new_n16021__ & ~new_new_n16027__;
  assign new_new_n16029__ = ~new_new_n16026__ & new_new_n16028__;
  assign new_new_n16030__ = new_new_n11650__ & ~new_new_n16029__;
  assign ys__n4615 = new_new_n16025__ | new_new_n16030__;
  assign new_new_n16032__ = ~ys__n35098 & ~ys__n35423;
  assign new_new_n16033__ = ys__n35098 & ys__n35423;
  assign new_new_n16034__ = ~new_new_n16032__ & ~new_new_n16033__;
  assign new_new_n16035__ = ~ys__n35096 & ~ys__n35421;
  assign new_new_n16036__ = ys__n35096 & ys__n35421;
  assign new_new_n16037__ = ~new_new_n16035__ & ~new_new_n16036__;
  assign new_new_n16038__ = ~new_new_n16034__ & ~new_new_n16037__;
  assign new_new_n16039__ = ~ys__n35094 & ~ys__n35419;
  assign new_new_n16040__ = ys__n35094 & ys__n35419;
  assign new_new_n16041__ = ~new_new_n16039__ & ~new_new_n16040__;
  assign new_new_n16042__ = ~ys__n35092 & ~ys__n35417;
  assign new_new_n16043__ = ys__n35092 & ys__n35417;
  assign new_new_n16044__ = ~new_new_n16042__ & ~new_new_n16043__;
  assign new_new_n16045__ = ~new_new_n16041__ & ~new_new_n16044__;
  assign new_new_n16046__ = new_new_n16038__ & new_new_n16045__;
  assign new_new_n16047__ = ~ys__n35090 & ~ys__n35415;
  assign new_new_n16048__ = ys__n35090 & ys__n35415;
  assign new_new_n16049__ = ~new_new_n16047__ & ~new_new_n16048__;
  assign new_new_n16050__ = ~ys__n35088 & ~ys__n35413;
  assign new_new_n16051__ = ys__n35088 & ys__n35413;
  assign new_new_n16052__ = ~new_new_n16050__ & ~new_new_n16051__;
  assign new_new_n16053__ = ~new_new_n16049__ & ~new_new_n16052__;
  assign new_new_n16054__ = ~ys__n35086 & ~ys__n48335;
  assign new_new_n16055__ = ys__n35086 & ys__n48335;
  assign new_new_n16056__ = ~new_new_n16054__ & ~new_new_n16055__;
  assign new_new_n16057__ = ~ys__n35084 & ~ys__n48334;
  assign new_new_n16058__ = ys__n35084 & ys__n48334;
  assign new_new_n16059__ = ~new_new_n16057__ & ~new_new_n16058__;
  assign new_new_n16060__ = ~new_new_n16056__ & ~new_new_n16059__;
  assign new_new_n16061__ = new_new_n16053__ & new_new_n16060__;
  assign new_new_n16062__ = ~ys__n35082 & ~ys__n48333;
  assign new_new_n16063__ = ys__n35082 & ys__n48333;
  assign new_new_n16064__ = ~new_new_n16062__ & ~new_new_n16063__;
  assign new_new_n16065__ = ~ys__n35080 & ~ys__n48332;
  assign new_new_n16066__ = ys__n35080 & ys__n48332;
  assign new_new_n16067__ = ~new_new_n16065__ & ~new_new_n16066__;
  assign new_new_n16068__ = ~new_new_n16064__ & ~new_new_n16067__;
  assign new_new_n16069__ = ~ys__n35078 & ys__n48331;
  assign new_new_n16070__ = ~ys__n35078 & ~ys__n48331;
  assign new_new_n16071__ = ys__n35078 & ys__n48331;
  assign new_new_n16072__ = ~new_new_n16070__ & ~new_new_n16071__;
  assign new_new_n16073__ = ~ys__n35076 & ys__n48330;
  assign new_new_n16074__ = ~ys__n35076 & ~ys__n48330;
  assign new_new_n16075__ = ys__n35076 & ys__n48330;
  assign new_new_n16076__ = ~new_new_n16074__ & ~new_new_n16075__;
  assign new_new_n16077__ = ~new_new_n16073__ & new_new_n16076__;
  assign new_new_n16078__ = ~new_new_n16072__ & ~new_new_n16077__;
  assign new_new_n16079__ = ~new_new_n16069__ & ~new_new_n16078__;
  assign new_new_n16080__ = new_new_n16068__ & ~new_new_n16079__;
  assign new_new_n16081__ = ~ys__n35082 & ys__n48333;
  assign new_new_n16082__ = ~ys__n35080 & ys__n48332;
  assign new_new_n16083__ = ~new_new_n16064__ & new_new_n16082__;
  assign new_new_n16084__ = ~new_new_n16081__ & ~new_new_n16083__;
  assign new_new_n16085__ = ~new_new_n16080__ & new_new_n16084__;
  assign new_new_n16086__ = new_new_n16061__ & ~new_new_n16085__;
  assign new_new_n16087__ = ~ys__n35086 & ys__n48335;
  assign new_new_n16088__ = ~ys__n35084 & ys__n48334;
  assign new_new_n16089__ = ~new_new_n16056__ & new_new_n16088__;
  assign new_new_n16090__ = ~new_new_n16087__ & ~new_new_n16089__;
  assign new_new_n16091__ = new_new_n16053__ & ~new_new_n16090__;
  assign new_new_n16092__ = ~ys__n35090 & ys__n35415;
  assign new_new_n16093__ = ~ys__n35088 & ys__n35413;
  assign new_new_n16094__ = ~new_new_n16049__ & new_new_n16093__;
  assign new_new_n16095__ = ~new_new_n16092__ & ~new_new_n16094__;
  assign new_new_n16096__ = ~new_new_n16091__ & new_new_n16095__;
  assign new_new_n16097__ = ~new_new_n16086__ & new_new_n16096__;
  assign new_new_n16098__ = new_new_n16046__ & ~new_new_n16097__;
  assign new_new_n16099__ = ~ys__n35094 & ys__n35419;
  assign new_new_n16100__ = ~ys__n35092 & ys__n35417;
  assign new_new_n16101__ = ~new_new_n16041__ & new_new_n16100__;
  assign new_new_n16102__ = ~new_new_n16099__ & ~new_new_n16101__;
  assign new_new_n16103__ = new_new_n16038__ & ~new_new_n16102__;
  assign new_new_n16104__ = ~ys__n35098 & ys__n35423;
  assign new_new_n16105__ = ~ys__n35096 & ys__n35421;
  assign new_new_n16106__ = ~new_new_n16034__ & new_new_n16105__;
  assign new_new_n16107__ = ~new_new_n16104__ & ~new_new_n16106__;
  assign new_new_n16108__ = ~new_new_n16103__ & new_new_n16107__;
  assign new_new_n16109__ = ~new_new_n16098__ & new_new_n16108__;
  assign new_new_n16110__ = ~new_new_n16072__ & ~new_new_n16076__;
  assign new_new_n16111__ = new_new_n16068__ & new_new_n16110__;
  assign new_new_n16112__ = new_new_n16046__ & new_new_n16111__;
  assign new_new_n16113__ = new_new_n16061__ & new_new_n16112__;
  assign new_new_n16114__ = ~new_new_n16109__ & ~new_new_n16113__;
  assign new_new_n16115__ = ~ys__n33218 & ~ys__n35419;
  assign new_new_n16116__ = ys__n33218 & ys__n35419;
  assign new_new_n16117__ = ~new_new_n16115__ & ~new_new_n16116__;
  assign new_new_n16118__ = ~ys__n33216 & ~ys__n35417;
  assign new_new_n16119__ = ys__n33216 & ys__n35417;
  assign new_new_n16120__ = ~new_new_n16118__ & ~new_new_n16119__;
  assign new_new_n16121__ = ~new_new_n16117__ & ~new_new_n16120__;
  assign new_new_n16122__ = ~ys__n33222 & ~ys__n35423;
  assign new_new_n16123__ = ys__n33222 & ys__n35423;
  assign new_new_n16124__ = ~new_new_n16122__ & ~new_new_n16123__;
  assign new_new_n16125__ = ~ys__n33220 & ~ys__n35421;
  assign new_new_n16126__ = ys__n33220 & ys__n35421;
  assign new_new_n16127__ = ~new_new_n16125__ & ~new_new_n16126__;
  assign new_new_n16128__ = ~new_new_n16124__ & ~new_new_n16127__;
  assign new_new_n16129__ = ~ys__n33214 & ~ys__n35415;
  assign new_new_n16130__ = ys__n33214 & ys__n35415;
  assign new_new_n16131__ = ~new_new_n16129__ & ~new_new_n16130__;
  assign new_new_n16132__ = ~ys__n33212 & ~ys__n35413;
  assign new_new_n16133__ = ys__n33212 & ys__n35413;
  assign new_new_n16134__ = ~new_new_n16132__ & ~new_new_n16133__;
  assign new_new_n16135__ = ~new_new_n16131__ & ~new_new_n16134__;
  assign new_new_n16136__ = new_new_n16128__ & new_new_n16135__;
  assign new_new_n16137__ = new_new_n16121__ & new_new_n16136__;
  assign new_new_n16138__ = ~ys__n33214 & ys__n35415;
  assign new_new_n16139__ = ~ys__n33212 & ys__n35413;
  assign new_new_n16140__ = new_new_n16134__ & ~new_new_n16139__;
  assign new_new_n16141__ = ~new_new_n16131__ & ~new_new_n16140__;
  assign new_new_n16142__ = ~new_new_n16138__ & ~new_new_n16141__;
  assign new_new_n16143__ = new_new_n16121__ & ~new_new_n16142__;
  assign new_new_n16144__ = ~ys__n33218 & ys__n35419;
  assign new_new_n16145__ = ~ys__n33216 & ys__n35417;
  assign new_new_n16146__ = ~new_new_n16117__ & new_new_n16145__;
  assign new_new_n16147__ = ~new_new_n16144__ & ~new_new_n16146__;
  assign new_new_n16148__ = ~new_new_n16143__ & new_new_n16147__;
  assign new_new_n16149__ = new_new_n16128__ & ~new_new_n16148__;
  assign new_new_n16150__ = ~ys__n33222 & ys__n35423;
  assign new_new_n16151__ = ~ys__n33220 & ys__n35421;
  assign new_new_n16152__ = ~new_new_n16124__ & new_new_n16151__;
  assign new_new_n16153__ = ~new_new_n16150__ & ~new_new_n16152__;
  assign new_new_n16154__ = ~new_new_n16149__ & new_new_n16153__;
  assign new_new_n16155__ = ~new_new_n16137__ & ~new_new_n16154__;
  assign new_new_n16156__ = ~new_new_n16137__ & ~new_new_n16155__;
  assign new_new_n16157__ = ~ys__n38847 & ys__n38848;
  assign new_new_n16158__ = ys__n38847 & ~ys__n38848;
  assign new_new_n16159__ = ~new_new_n16157__ & ~new_new_n16158__;
  assign new_new_n16160__ = ~ys__n38849 & ys__n38850;
  assign new_new_n16161__ = ys__n38849 & ~ys__n38850;
  assign new_new_n16162__ = ~new_new_n16160__ & ~new_new_n16161__;
  assign new_new_n16163__ = new_new_n16159__ & new_new_n16162__;
  assign new_new_n16164__ = ~ys__n38843 & ys__n38844;
  assign new_new_n16165__ = ys__n38843 & ~ys__n38844;
  assign new_new_n16166__ = ~new_new_n16164__ & ~new_new_n16165__;
  assign new_new_n16167__ = ~ys__n38845 & ys__n38846;
  assign new_new_n16168__ = ys__n38845 & ~ys__n38846;
  assign new_new_n16169__ = ~new_new_n16167__ & ~new_new_n16168__;
  assign new_new_n16170__ = new_new_n16166__ & new_new_n16169__;
  assign new_new_n16171__ = new_new_n16163__ & new_new_n16170__;
  assign new_new_n16172__ = ~ys__n38855 & ys__n38856;
  assign new_new_n16173__ = ys__n38855 & ~ys__n38856;
  assign new_new_n16174__ = ~new_new_n16172__ & ~new_new_n16173__;
  assign new_new_n16175__ = ~ys__n38857 & ys__n38858;
  assign new_new_n16176__ = ys__n38857 & ~ys__n38858;
  assign new_new_n16177__ = ~new_new_n16175__ & ~new_new_n16176__;
  assign new_new_n16178__ = new_new_n16174__ & new_new_n16177__;
  assign new_new_n16179__ = ~ys__n38851 & ys__n38852;
  assign new_new_n16180__ = ys__n38851 & ~ys__n38852;
  assign new_new_n16181__ = ~new_new_n16179__ & ~new_new_n16180__;
  assign new_new_n16182__ = ~ys__n38853 & ys__n38854;
  assign new_new_n16183__ = ys__n38853 & ~ys__n38854;
  assign new_new_n16184__ = ~new_new_n16182__ & ~new_new_n16183__;
  assign new_new_n16185__ = new_new_n16181__ & new_new_n16184__;
  assign new_new_n16186__ = new_new_n16178__ & new_new_n16185__;
  assign new_new_n16187__ = new_new_n16171__ & new_new_n16186__;
  assign new_new_n16188__ = ~ys__n38831 & ys__n38832;
  assign new_new_n16189__ = ys__n38831 & ~ys__n38832;
  assign new_new_n16190__ = ~new_new_n16188__ & ~new_new_n16189__;
  assign new_new_n16191__ = ~ys__n38833 & ys__n38834;
  assign new_new_n16192__ = ys__n38833 & ~ys__n38834;
  assign new_new_n16193__ = ~new_new_n16191__ & ~new_new_n16192__;
  assign new_new_n16194__ = new_new_n16190__ & new_new_n16193__;
  assign new_new_n16195__ = ~ys__n38827 & ys__n38828;
  assign new_new_n16196__ = ys__n38827 & ~ys__n38828;
  assign new_new_n16197__ = ~new_new_n16195__ & ~new_new_n16196__;
  assign new_new_n16198__ = ~ys__n38829 & ys__n38830;
  assign new_new_n16199__ = ys__n38829 & ~ys__n38830;
  assign new_new_n16200__ = ~new_new_n16198__ & ~new_new_n16199__;
  assign new_new_n16201__ = new_new_n16197__ & new_new_n16200__;
  assign new_new_n16202__ = new_new_n16194__ & new_new_n16201__;
  assign new_new_n16203__ = ~ys__n38839 & ys__n38840;
  assign new_new_n16204__ = ys__n38839 & ~ys__n38840;
  assign new_new_n16205__ = ~new_new_n16203__ & ~new_new_n16204__;
  assign new_new_n16206__ = ~ys__n38841 & ys__n38842;
  assign new_new_n16207__ = ys__n38841 & ~ys__n38842;
  assign new_new_n16208__ = ~new_new_n16206__ & ~new_new_n16207__;
  assign new_new_n16209__ = new_new_n16205__ & new_new_n16208__;
  assign new_new_n16210__ = ~ys__n38835 & ys__n38836;
  assign new_new_n16211__ = ys__n38835 & ~ys__n38836;
  assign new_new_n16212__ = ~new_new_n16210__ & ~new_new_n16211__;
  assign new_new_n16213__ = ~ys__n38837 & ys__n38838;
  assign new_new_n16214__ = ys__n38837 & ~ys__n38838;
  assign new_new_n16215__ = ~new_new_n16213__ & ~new_new_n16214__;
  assign new_new_n16216__ = new_new_n16212__ & new_new_n16215__;
  assign new_new_n16217__ = new_new_n16209__ & new_new_n16216__;
  assign new_new_n16218__ = new_new_n16202__ & new_new_n16217__;
  assign new_new_n16219__ = new_new_n16187__ & new_new_n16218__;
  assign new_new_n16220__ = ~new_new_n16156__ & new_new_n16219__;
  assign new_new_n16221__ = ~new_new_n16114__ & new_new_n16220__;
  assign new_new_n16222__ = ~ys__n18149 & ~ys__n18150;
  assign new_new_n16223__ = ys__n18137 & ~new_new_n16222__;
  assign ys__n4696 = new_new_n16221__ & new_new_n16223__;
  assign new_new_n16225__ = new_new_n11010__ & ~new_new_n11055__;
  assign new_new_n16226__ = new_new_n11021__ & new_new_n11033__;
  assign new_new_n16227__ = ~new_new_n16225__ & new_new_n16226__;
  assign ys__n4791 = ~new_new_n11036__ & ~new_new_n16227__;
  assign ys__n4793 = ~new_new_n11026__ & ~new_new_n11036__;
  assign new_new_n16230__ = ~ys__n574 & ~ys__n4791;
  assign new_new_n16231__ = ~ys__n4793 & new_new_n16230__;
  assign ys__n4798 = ys__n576 | ~new_new_n16231__;
  assign ys__n18166 = ys__n402 & ~ys__n4566;
  assign new_new_n16234__ = ~ys__n164 & ~ys__n398;
  assign new_new_n16235__ = ~new_new_n14001__ & new_new_n16234__;
  assign new_new_n16236__ = ~ys__n18166 & new_new_n16235__;
  assign ys__n4817 = ys__n18166 | new_new_n16236__;
  assign new_new_n16238__ = ~ys__n164 & ys__n4826;
  assign new_new_n16239__ = ~new_new_n13941__ & ~new_new_n16238__;
  assign new_new_n16240__ = ~ys__n398 & ~new_new_n16239__;
  assign new_new_n16241__ = ~new_new_n14001__ & new_new_n16240__;
  assign ys__n4818 = ~ys__n18166 & new_new_n16241__;
  assign new_new_n16243__ = ys__n164 & ys__n4826;
  assign new_new_n16244__ = ~ys__n4832 & new_new_n16243__;
  assign new_new_n16245__ = ys__n4832 & ~new_new_n16243__;
  assign new_new_n16246__ = ~new_new_n16244__ & ~new_new_n16245__;
  assign new_new_n16247__ = ~ys__n398 & ~new_new_n14001__;
  assign new_new_n16248__ = ~new_new_n16246__ & new_new_n16247__;
  assign ys__n4820 = ~ys__n18166 & new_new_n16248__;
  assign new_new_n16250__ = ys__n4832 & new_new_n16243__;
  assign new_new_n16251__ = ~ys__n4833 & new_new_n16250__;
  assign new_new_n16252__ = ys__n4833 & ~new_new_n16250__;
  assign new_new_n16253__ = ~new_new_n16251__ & ~new_new_n16252__;
  assign new_new_n16254__ = new_new_n16247__ & ~new_new_n16253__;
  assign ys__n4821 = ~ys__n18166 & new_new_n16254__;
  assign new_new_n16256__ = ys__n4832 & ys__n4833;
  assign new_new_n16257__ = new_new_n16243__ & new_new_n16256__;
  assign new_new_n16258__ = ~ys__n354 & new_new_n16257__;
  assign new_new_n16259__ = ys__n354 & ~new_new_n16257__;
  assign new_new_n16260__ = ~new_new_n16258__ & ~new_new_n16259__;
  assign new_new_n16261__ = new_new_n16247__ & ~new_new_n16260__;
  assign ys__n4824 = ~ys__n18166 & new_new_n16261__;
  assign new_new_n16263__ = ~ys__n4818 & ~ys__n4820;
  assign new_new_n16264__ = ~ys__n4821 & ~ys__n4824;
  assign new_new_n16265__ = new_new_n16263__ & new_new_n16264__;
  assign ys__n4825 = ys__n4817 | ~new_new_n16265__;
  assign new_new_n16267__ = ~new_new_n12343__ & ~new_new_n12347__;
  assign new_new_n16268__ = ~new_new_n12350__ & new_new_n16267__;
  assign ys__n4839 = ys__n4836 & new_new_n16268__;
  assign ys__n4840 = ys__n4837 & new_new_n16268__;
  assign new_new_n16271__ = ys__n47661 & ~new_new_n10820__;
  assign new_new_n16272__ = ys__n23269 & ~new_new_n11180__;
  assign new_new_n16273__ = new_new_n10820__ & new_new_n16272__;
  assign ys__n12455 = new_new_n16271__ | new_new_n16273__;
  assign new_new_n16275__ = ys__n47662 & ~new_new_n10820__;
  assign new_new_n16276__ = ys__n23271 & ~new_new_n11180__;
  assign new_new_n16277__ = ys__n23272 & new_new_n11180__;
  assign new_new_n16278__ = ~new_new_n16276__ & ~new_new_n16277__;
  assign new_new_n16279__ = new_new_n10820__ & ~new_new_n16278__;
  assign ys__n12458 = new_new_n16275__ | new_new_n16279__;
  assign new_new_n16281__ = ys__n47663 & ~new_new_n10820__;
  assign new_new_n16282__ = ys__n23203 & ~new_new_n11180__;
  assign new_new_n16283__ = ys__n23274 & new_new_n11180__;
  assign new_new_n16284__ = ~new_new_n16282__ & ~new_new_n16283__;
  assign new_new_n16285__ = new_new_n10820__ & ~new_new_n16284__;
  assign ys__n12461 = new_new_n16281__ | new_new_n16285__;
  assign new_new_n16287__ = ys__n47664 & ~new_new_n10820__;
  assign new_new_n16288__ = ys__n23205 & ~new_new_n11180__;
  assign new_new_n16289__ = ys__n23276 & new_new_n11180__;
  assign new_new_n16290__ = ~new_new_n16288__ & ~new_new_n16289__;
  assign new_new_n16291__ = new_new_n10820__ & ~new_new_n16290__;
  assign ys__n12464 = new_new_n16287__ | new_new_n16291__;
  assign new_new_n16293__ = ys__n47665 & ~new_new_n10820__;
  assign new_new_n16294__ = ys__n23207 & ~new_new_n11180__;
  assign new_new_n16295__ = ys__n23278 & new_new_n11180__;
  assign new_new_n16296__ = ~new_new_n16294__ & ~new_new_n16295__;
  assign new_new_n16297__ = new_new_n10820__ & ~new_new_n16296__;
  assign ys__n12467 = new_new_n16293__ | new_new_n16297__;
  assign new_new_n16299__ = ys__n47666 & ~new_new_n10820__;
  assign new_new_n16300__ = ys__n23209 & ~new_new_n11180__;
  assign new_new_n16301__ = ys__n23280 & new_new_n11180__;
  assign new_new_n16302__ = ~new_new_n16300__ & ~new_new_n16301__;
  assign new_new_n16303__ = new_new_n10820__ & ~new_new_n16302__;
  assign ys__n12470 = new_new_n16299__ | new_new_n16303__;
  assign new_new_n16305__ = ys__n47667 & ~new_new_n10820__;
  assign new_new_n16306__ = ys__n23211 & ~new_new_n11180__;
  assign new_new_n16307__ = ys__n23282 & new_new_n11180__;
  assign new_new_n16308__ = ~new_new_n16306__ & ~new_new_n16307__;
  assign new_new_n16309__ = new_new_n10820__ & ~new_new_n16308__;
  assign ys__n12473 = new_new_n16305__ | new_new_n16309__;
  assign new_new_n16311__ = ys__n47668 & ~new_new_n10820__;
  assign new_new_n16312__ = ys__n23213 & ~new_new_n11180__;
  assign new_new_n16313__ = ys__n23284 & new_new_n11180__;
  assign new_new_n16314__ = ~new_new_n16312__ & ~new_new_n16313__;
  assign new_new_n16315__ = new_new_n10820__ & ~new_new_n16314__;
  assign ys__n12476 = new_new_n16311__ | new_new_n16315__;
  assign new_new_n16317__ = ys__n47669 & ~new_new_n10820__;
  assign new_new_n16318__ = ys__n23215 & ~new_new_n11180__;
  assign new_new_n16319__ = ys__n23286 & new_new_n11180__;
  assign new_new_n16320__ = ~new_new_n16318__ & ~new_new_n16319__;
  assign new_new_n16321__ = new_new_n10820__ & ~new_new_n16320__;
  assign ys__n12479 = new_new_n16317__ | new_new_n16321__;
  assign new_new_n16323__ = ys__n47670 & ~new_new_n10820__;
  assign new_new_n16324__ = ys__n23217 & ~new_new_n11180__;
  assign new_new_n16325__ = ys__n23288 & new_new_n11180__;
  assign new_new_n16326__ = ~new_new_n16324__ & ~new_new_n16325__;
  assign new_new_n16327__ = new_new_n10820__ & ~new_new_n16326__;
  assign ys__n12482 = new_new_n16323__ | new_new_n16327__;
  assign new_new_n16329__ = ys__n47671 & ~new_new_n10820__;
  assign new_new_n16330__ = ys__n23219 & ~new_new_n11180__;
  assign new_new_n16331__ = ys__n23290 & new_new_n11180__;
  assign new_new_n16332__ = ~new_new_n16330__ & ~new_new_n16331__;
  assign new_new_n16333__ = new_new_n10820__ & ~new_new_n16332__;
  assign ys__n12485 = new_new_n16329__ | new_new_n16333__;
  assign new_new_n16335__ = ys__n47672 & ~new_new_n10820__;
  assign new_new_n16336__ = ys__n23221 & ~new_new_n11180__;
  assign new_new_n16337__ = ys__n23292 & new_new_n11180__;
  assign new_new_n16338__ = ~new_new_n16336__ & ~new_new_n16337__;
  assign new_new_n16339__ = new_new_n10820__ & ~new_new_n16338__;
  assign ys__n12488 = new_new_n16335__ | new_new_n16339__;
  assign new_new_n16341__ = ys__n47673 & ~new_new_n10820__;
  assign new_new_n16342__ = ys__n23223 & ~new_new_n11180__;
  assign new_new_n16343__ = ys__n23294 & new_new_n11180__;
  assign new_new_n16344__ = ~new_new_n16342__ & ~new_new_n16343__;
  assign new_new_n16345__ = new_new_n10820__ & ~new_new_n16344__;
  assign ys__n12491 = new_new_n16341__ | new_new_n16345__;
  assign new_new_n16347__ = ys__n47674 & ~new_new_n10820__;
  assign new_new_n16348__ = ys__n23225 & ~new_new_n11180__;
  assign new_new_n16349__ = ys__n23296 & new_new_n11180__;
  assign new_new_n16350__ = ~new_new_n16348__ & ~new_new_n16349__;
  assign new_new_n16351__ = new_new_n10820__ & ~new_new_n16350__;
  assign ys__n12494 = new_new_n16347__ | new_new_n16351__;
  assign new_new_n16353__ = ys__n47675 & ~new_new_n10820__;
  assign new_new_n16354__ = ys__n23227 & ~new_new_n11180__;
  assign new_new_n16355__ = ys__n23298 & new_new_n11180__;
  assign new_new_n16356__ = ~new_new_n16354__ & ~new_new_n16355__;
  assign new_new_n16357__ = new_new_n10820__ & ~new_new_n16356__;
  assign ys__n12497 = new_new_n16353__ | new_new_n16357__;
  assign new_new_n16359__ = ys__n47676 & ~new_new_n10820__;
  assign new_new_n16360__ = ys__n23229 & ~new_new_n11180__;
  assign new_new_n16361__ = ys__n23300 & new_new_n11180__;
  assign new_new_n16362__ = ~new_new_n16360__ & ~new_new_n16361__;
  assign new_new_n16363__ = new_new_n10820__ & ~new_new_n16362__;
  assign ys__n12500 = new_new_n16359__ | new_new_n16363__;
  assign new_new_n16365__ = ys__n47677 & ~new_new_n10820__;
  assign new_new_n16366__ = ys__n23231 & ~new_new_n11180__;
  assign new_new_n16367__ = ys__n23302 & new_new_n11180__;
  assign new_new_n16368__ = ~new_new_n16366__ & ~new_new_n16367__;
  assign new_new_n16369__ = new_new_n10820__ & ~new_new_n16368__;
  assign ys__n12503 = new_new_n16365__ | new_new_n16369__;
  assign new_new_n16371__ = ys__n47678 & ~new_new_n10820__;
  assign new_new_n16372__ = ys__n23233 & ~new_new_n11180__;
  assign new_new_n16373__ = ys__n23304 & new_new_n11180__;
  assign new_new_n16374__ = ~new_new_n16372__ & ~new_new_n16373__;
  assign new_new_n16375__ = new_new_n10820__ & ~new_new_n16374__;
  assign ys__n12506 = new_new_n16371__ | new_new_n16375__;
  assign new_new_n16377__ = ys__n47679 & ~new_new_n10820__;
  assign new_new_n16378__ = ys__n23235 & ~new_new_n11180__;
  assign new_new_n16379__ = ys__n23306 & new_new_n11180__;
  assign new_new_n16380__ = ~new_new_n16378__ & ~new_new_n16379__;
  assign new_new_n16381__ = new_new_n10820__ & ~new_new_n16380__;
  assign ys__n12509 = new_new_n16377__ | new_new_n16381__;
  assign new_new_n16383__ = ys__n47680 & ~new_new_n10820__;
  assign new_new_n16384__ = ys__n23237 & ~new_new_n11180__;
  assign new_new_n16385__ = ys__n23308 & new_new_n11180__;
  assign new_new_n16386__ = ~new_new_n16384__ & ~new_new_n16385__;
  assign new_new_n16387__ = new_new_n10820__ & ~new_new_n16386__;
  assign ys__n12512 = new_new_n16383__ | new_new_n16387__;
  assign new_new_n16389__ = ys__n47681 & ~new_new_n10820__;
  assign new_new_n16390__ = ys__n23239 & ~new_new_n11180__;
  assign new_new_n16391__ = ys__n23310 & new_new_n11180__;
  assign new_new_n16392__ = ~new_new_n16390__ & ~new_new_n16391__;
  assign new_new_n16393__ = new_new_n10820__ & ~new_new_n16392__;
  assign ys__n12515 = new_new_n16389__ | new_new_n16393__;
  assign new_new_n16395__ = ys__n47682 & ~new_new_n10820__;
  assign new_new_n16396__ = ys__n23241 & ~new_new_n11180__;
  assign new_new_n16397__ = ys__n23312 & new_new_n11180__;
  assign new_new_n16398__ = ~new_new_n16396__ & ~new_new_n16397__;
  assign new_new_n16399__ = new_new_n10820__ & ~new_new_n16398__;
  assign ys__n12518 = new_new_n16395__ | new_new_n16399__;
  assign new_new_n16401__ = ys__n47683 & ~new_new_n10820__;
  assign new_new_n16402__ = ys__n23243 & ~new_new_n11180__;
  assign new_new_n16403__ = ys__n23314 & new_new_n11180__;
  assign new_new_n16404__ = ~new_new_n16402__ & ~new_new_n16403__;
  assign new_new_n16405__ = new_new_n10820__ & ~new_new_n16404__;
  assign ys__n12521 = new_new_n16401__ | new_new_n16405__;
  assign new_new_n16407__ = ys__n47684 & ~new_new_n10820__;
  assign new_new_n16408__ = ys__n23245 & ~new_new_n11180__;
  assign new_new_n16409__ = ys__n23316 & new_new_n11180__;
  assign new_new_n16410__ = ~new_new_n16408__ & ~new_new_n16409__;
  assign new_new_n16411__ = new_new_n10820__ & ~new_new_n16410__;
  assign ys__n12524 = new_new_n16407__ | new_new_n16411__;
  assign new_new_n16413__ = ys__n47685 & ~new_new_n10820__;
  assign new_new_n16414__ = ys__n23247 & ~new_new_n11180__;
  assign new_new_n16415__ = ys__n23318 & new_new_n11180__;
  assign new_new_n16416__ = ~new_new_n16414__ & ~new_new_n16415__;
  assign new_new_n16417__ = new_new_n10820__ & ~new_new_n16416__;
  assign ys__n12527 = new_new_n16413__ | new_new_n16417__;
  assign new_new_n16419__ = ys__n47686 & ~new_new_n10820__;
  assign new_new_n16420__ = ys__n23249 & ~new_new_n11180__;
  assign new_new_n16421__ = ys__n23320 & new_new_n11180__;
  assign new_new_n16422__ = ~new_new_n16420__ & ~new_new_n16421__;
  assign new_new_n16423__ = new_new_n10820__ & ~new_new_n16422__;
  assign ys__n12530 = new_new_n16419__ | new_new_n16423__;
  assign new_new_n16425__ = ys__n47687 & ~new_new_n10820__;
  assign new_new_n16426__ = ys__n23251 & ~new_new_n11180__;
  assign new_new_n16427__ = ys__n23322 & new_new_n11180__;
  assign new_new_n16428__ = ~new_new_n16426__ & ~new_new_n16427__;
  assign new_new_n16429__ = new_new_n10820__ & ~new_new_n16428__;
  assign ys__n12533 = new_new_n16425__ | new_new_n16429__;
  assign new_new_n16431__ = ys__n47688 & ~new_new_n10820__;
  assign new_new_n16432__ = ys__n23253 & ~new_new_n11180__;
  assign new_new_n16433__ = ys__n23324 & new_new_n11180__;
  assign new_new_n16434__ = ~new_new_n16432__ & ~new_new_n16433__;
  assign new_new_n16435__ = new_new_n10820__ & ~new_new_n16434__;
  assign ys__n12536 = new_new_n16431__ | new_new_n16435__;
  assign new_new_n16437__ = ys__n47689 & ~new_new_n10820__;
  assign new_new_n16438__ = ys__n23255 & ~new_new_n11180__;
  assign new_new_n16439__ = ys__n23326 & new_new_n11180__;
  assign new_new_n16440__ = ~new_new_n16438__ & ~new_new_n16439__;
  assign new_new_n16441__ = new_new_n10820__ & ~new_new_n16440__;
  assign ys__n12539 = new_new_n16437__ | new_new_n16441__;
  assign new_new_n16443__ = ys__n47690 & ~new_new_n10820__;
  assign new_new_n16444__ = ys__n23257 & ~new_new_n11180__;
  assign new_new_n16445__ = ~new_new_n11182__ & ~new_new_n16444__;
  assign new_new_n16446__ = new_new_n10820__ & ~new_new_n16445__;
  assign ys__n12542 = new_new_n16443__ | new_new_n16446__;
  assign new_new_n16448__ = ys__n47691 & ~new_new_n10820__;
  assign new_new_n16449__ = ys__n23259 & ~new_new_n11180__;
  assign new_new_n16450__ = ~new_new_n15985__ & ~new_new_n16449__;
  assign new_new_n16451__ = new_new_n10820__ & ~new_new_n16450__;
  assign ys__n12545 = new_new_n16448__ | new_new_n16451__;
  assign new_new_n16453__ = ys__n38311 & ~new_new_n10820__;
  assign new_new_n16454__ = ys__n23261 & ~new_new_n11180__;
  assign new_new_n16455__ = ~new_new_n11656__ & ~new_new_n16454__;
  assign new_new_n16456__ = new_new_n10820__ & ~new_new_n16455__;
  assign ys__n12548 = new_new_n16453__ | new_new_n16456__;
  assign new_new_n16458__ = ys__n30223 & new_new_n12152__;
  assign ys__n16188 = new_new_n12428__ | new_new_n16458__;
  assign new_new_n16460__ = ys__n740 & new_new_n12186__;
  assign new_new_n16461__ = new_new_n12188__ & ys__n3039;
  assign ys__n16412 = new_new_n16460__ | new_new_n16461__;
  assign new_new_n16463__ = new_new_n12188__ & ~ys__n3039;
  assign new_new_n16464__ = ys__n23850 & new_new_n12183__;
  assign ys__n16415 = new_new_n16463__ | new_new_n16464__;
  assign new_new_n16466__ = ys__n30223 & new_new_n12163__;
  assign ys__n16424 = new_new_n12450__ | new_new_n16466__;
  assign new_new_n16468__ = ys__n740 & new_new_n12175__;
  assign new_new_n16469__ = new_new_n12177__ & ys__n3039;
  assign ys__n16706 = new_new_n16468__ | new_new_n16469__;
  assign new_new_n16471__ = new_new_n12177__ & ~ys__n3039;
  assign new_new_n16472__ = ys__n23850 & new_new_n12172__;
  assign ys__n16709 = new_new_n16471__ | new_new_n16472__;
  assign new_new_n16474__ = ys__n30223 & new_new_n12196__;
  assign ys__n16718 = new_new_n12458__ | new_new_n16474__;
  assign new_new_n16476__ = ys__n740 & new_new_n12208__;
  assign new_new_n16477__ = new_new_n12210__ & ys__n3039;
  assign ys__n17692 = new_new_n16476__ | new_new_n16477__;
  assign new_new_n16479__ = new_new_n12210__ & ~ys__n3039;
  assign new_new_n16480__ = ys__n23850 & new_new_n12205__;
  assign ys__n17697 = new_new_n16479__ | new_new_n16480__;
  assign new_new_n16482__ = ys__n414 & ys__n728;
  assign new_new_n16483__ = ys__n724 & ys__n726;
  assign new_new_n16484__ = new_new_n16482__ & new_new_n16483__;
  assign new_new_n16485__ = ys__n718 & ys__n720;
  assign new_new_n16486__ = ys__n722 & new_new_n16485__;
  assign ys__n18007 = new_new_n16484__ & new_new_n16486__;
  assign new_new_n16488__ = ys__n714 & ys__n716;
  assign ys__n18009 = ~ys__n4615 & new_new_n16488__;
  assign new_new_n16490__ = ys__n312 & ys__n622;
  assign new_new_n16491__ = ys__n618 & ys__n620;
  assign new_new_n16492__ = new_new_n16490__ & new_new_n16491__;
  assign new_new_n16493__ = ys__n612 & ys__n614;
  assign new_new_n16494__ = ys__n616 & new_new_n16493__;
  assign ys__n18015 = new_new_n16492__ & new_new_n16494__;
  assign new_new_n16496__ = ys__n456 & ys__n710;
  assign new_new_n16497__ = ys__n706 & ys__n708;
  assign new_new_n16498__ = new_new_n16496__ & new_new_n16497__;
  assign new_new_n16499__ = ys__n700 & ys__n702;
  assign new_new_n16500__ = ys__n704 & new_new_n16499__;
  assign ys__n18019 = new_new_n16498__ & new_new_n16500__;
  assign new_new_n16502__ = ys__n574 & ~ys__n4791;
  assign new_new_n16503__ = ~ys__n4793 & new_new_n16502__;
  assign ys__n18028 = ys__n576 & new_new_n16503__;
  assign new_new_n16505__ = ~ys__n628 & ~ys__n794;
  assign new_new_n16506__ = ~ys__n786 & ~ys__n792;
  assign new_new_n16507__ = ~ys__n788 & new_new_n16506__;
  assign new_new_n16508__ = ys__n630 & new_new_n16507__;
  assign new_new_n16509__ = new_new_n16505__ & new_new_n16508__;
  assign new_new_n16510__ = ~ys__n790 & new_new_n16509__;
  assign new_new_n16511__ = ~ys__n630 & ~ys__n790;
  assign new_new_n16512__ = ~ys__n794 & new_new_n16507__;
  assign new_new_n16513__ = ys__n628 & new_new_n16512__;
  assign new_new_n16514__ = new_new_n16511__ & new_new_n16513__;
  assign ys__n18078 = new_new_n16510__ | new_new_n16514__;
  assign new_new_n16516__ = ys__n1301 & ~new_new_n11727__;
  assign new_new_n16517__ = ys__n816 & new_new_n11727__;
  assign new_new_n16518__ = ~new_new_n16516__ & ~new_new_n16517__;
  assign ys__n18080 = ~new_new_n11731__ & ~new_new_n16518__;
  assign new_new_n16520__ = new_new_n16505__ & new_new_n16511__;
  assign new_new_n16521__ = ~ys__n786 & ~ys__n788;
  assign new_new_n16522__ = ys__n792 & new_new_n16521__;
  assign new_new_n16523__ = new_new_n16520__ & new_new_n16522__;
  assign new_new_n16524__ = ys__n18080 & new_new_n16523__;
  assign new_new_n16525__ = ys__n794 & new_new_n16507__;
  assign new_new_n16526__ = ~ys__n628 & new_new_n16525__;
  assign new_new_n16527__ = new_new_n16511__ & new_new_n16526__;
  assign new_new_n16528__ = ~ys__n18078 & ~new_new_n16527__;
  assign ys__n18082 = new_new_n16524__ | ~new_new_n16528__;
  assign new_new_n16530__ = ~new_new_n16510__ & ~new_new_n16527__;
  assign new_new_n16531__ = ~new_new_n16523__ & new_new_n16530__;
  assign new_new_n16532__ = ~ys__n18080 & ~new_new_n16531__;
  assign new_new_n16533__ = ys__n786 & ~ys__n788;
  assign new_new_n16534__ = ~ys__n792 & new_new_n16533__;
  assign new_new_n16535__ = new_new_n16520__ & new_new_n16534__;
  assign ys__n18089 = new_new_n16514__ | new_new_n16535__;
  assign ys__n18087 = new_new_n16532__ | ys__n18089;
  assign new_new_n16538__ = ~ys__n630 & new_new_n16507__;
  assign new_new_n16539__ = new_new_n16505__ & new_new_n16538__;
  assign new_new_n16540__ = ys__n790 & new_new_n16539__;
  assign new_new_n16541__ = ys__n788 & new_new_n16506__;
  assign new_new_n16542__ = new_new_n16520__ & new_new_n16541__;
  assign ys__n18088 = ~new_new_n16540__ & ~new_new_n16542__;
  assign ys__n18125 = ys__n1094 | ys__n1088;
  assign ys__n24256 = ys__n30219 & ~ys__n4566;
  assign new_new_n16546__ = ~ys__n846 & new_new_n10609__;
  assign new_new_n16547__ = new_new_n12226__ & new_new_n16546__;
  assign new_new_n16548__ = new_new_n11042__ & new_new_n16547__;
  assign ys__n18227 = ys__n4176 | ~new_new_n16548__;
  assign new_new_n16550__ = ys__n24256 & ~ys__n18227;
  assign new_new_n16551__ = ys__n18149 & ~ys__n4566;
  assign new_new_n16552__ = ys__n18227 & new_new_n16551__;
  assign ys__n18128 = new_new_n16550__ | new_new_n16552__;
  assign new_new_n16554__ = ~ys__n4566 & new_new_n16548__;
  assign new_new_n16555__ = ys__n4696 & new_new_n16554__;
  assign new_new_n16556__ = ~ys__n33509 & ~ys__n4566;
  assign new_new_n16557__ = ys__n18150 & ys__n18137;
  assign new_new_n16558__ = new_new_n16548__ & new_new_n16557__;
  assign new_new_n16559__ = ys__n38776 & ys__n38777;
  assign new_new_n16560__ = new_new_n16558__ & new_new_n16559__;
  assign new_new_n16561__ = new_new_n16556__ & new_new_n16560__;
  assign new_new_n16562__ = new_new_n16555__ & new_new_n16561__;
  assign new_new_n16563__ = new_new_n16558__ & ~new_new_n16559__;
  assign new_new_n16564__ = ~ys__n33511 & new_new_n16556__;
  assign new_new_n16565__ = new_new_n16563__ & new_new_n16564__;
  assign new_new_n16566__ = new_new_n16555__ & new_new_n16565__;
  assign ys__n33515 = ~new_new_n16562__ & ~new_new_n16566__;
  assign new_new_n16568__ = ~ys__n1156 & ys__n1157;
  assign new_new_n16569__ = ~ys__n1156 & ~new_new_n16568__;
  assign new_new_n16570__ = ~ys__n1154 & ~new_new_n16569__;
  assign new_new_n16571__ = ys__n1154 & new_new_n16548__;
  assign new_new_n16572__ = ~new_new_n16570__ & ~new_new_n16571__;
  assign new_new_n16573__ = ~ys__n1153 & ~new_new_n16572__;
  assign new_new_n16574__ = ~ys__n18149 & ~ys__n33532;
  assign new_new_n16575__ = ~ys__n4566 & new_new_n16574__;
  assign new_new_n16576__ = new_new_n16555__ & new_new_n16575__;
  assign new_new_n16577__ = ys__n1153 & ~new_new_n16576__;
  assign new_new_n16578__ = ~new_new_n16573__ & ~new_new_n16577__;
  assign new_new_n16579__ = ~ys__n1151 & ~new_new_n16578__;
  assign new_new_n16580__ = ys__n18150 & new_new_n16555__;
  assign new_new_n16581__ = ~ys__n4566 & new_new_n16580__;
  assign new_new_n16582__ = new_new_n11042__ & new_new_n11046__;
  assign new_new_n16583__ = ys__n1119 & ~new_new_n16582__;
  assign new_new_n16584__ = ~ys__n33491 & ys__n33493;
  assign new_new_n16585__ = ys__n1088 & new_new_n16584__;
  assign new_new_n16586__ = new_new_n16582__ & new_new_n16585__;
  assign new_new_n16587__ = ~ys__n4566 & new_new_n16586__;
  assign new_new_n16588__ = ~ys__n4696 & new_new_n16587__;
  assign new_new_n16589__ = ~new_new_n16583__ & ~new_new_n16588__;
  assign new_new_n16590__ = ys__n24464 & ~new_new_n16582__;
  assign new_new_n16591__ = ys__n4696 & new_new_n16587__;
  assign new_new_n16592__ = ~new_new_n16590__ & ~new_new_n16591__;
  assign new_new_n16593__ = ys__n24590 & new_new_n16222__;
  assign new_new_n16594__ = ys__n1151 & ~new_new_n16593__;
  assign new_new_n16595__ = new_new_n16592__ & new_new_n16594__;
  assign new_new_n16596__ = new_new_n16589__ & new_new_n16595__;
  assign new_new_n16597__ = ~new_new_n16581__ & new_new_n16596__;
  assign new_new_n16598__ = ~new_new_n16579__ & ~new_new_n16597__;
  assign new_new_n16599__ = ~ys__n140 & ~new_new_n16598__;
  assign ys__n18133 = ys__n140 | new_new_n16599__;
  assign new_new_n16601__ = ~ys__n1151 & ys__n1153;
  assign new_new_n16602__ = ~ys__n33532 & new_new_n16601__;
  assign new_new_n16603__ = ~ys__n4566 & new_new_n16602__;
  assign new_new_n16604__ = new_new_n16580__ & new_new_n16603__;
  assign new_new_n16605__ = ys__n1151 & new_new_n16581__;
  assign new_new_n16606__ = ~new_new_n16604__ & ~new_new_n16605__;
  assign ys__n18134 = ~ys__n140 & ~new_new_n16606__;
  assign new_new_n16608__ = ~ys__n18133 & ~ys__n18134;
  assign new_new_n16609__ = ys__n23335 & ys__n27855;
  assign new_new_n16610__ = new_new_n10770__ & new_new_n16609__;
  assign new_new_n16611__ = ~new_new_n10770__ & ~new_new_n16609__;
  assign new_new_n16612__ = ~new_new_n16610__ & ~new_new_n16611__;
  assign new_new_n16613__ = ~new_new_n10767__ & new_new_n16612__;
  assign new_new_n16614__ = new_new_n10767__ & new_new_n16612__;
  assign new_new_n16615__ = ~new_new_n16613__ & ~new_new_n16614__;
  assign new_new_n16616__ = ~new_new_n10767__ & ~new_new_n16612__;
  assign new_new_n16617__ = new_new_n10767__ & ~new_new_n16612__;
  assign new_new_n16618__ = ~new_new_n16616__ & ~new_new_n16617__;
  assign new_new_n16619__ = new_new_n16615__ & new_new_n16618__;
  assign new_new_n16620__ = ~ys__n1509 & ys__n1511;
  assign new_new_n16621__ = ~new_new_n16619__ & new_new_n16620__;
  assign new_new_n16622__ = ys__n1509 & ~new_new_n16615__;
  assign new_new_n16623__ = ~new_new_n16619__ & new_new_n16622__;
  assign new_new_n16624__ = ~new_new_n16621__ & ~new_new_n16623__;
  assign new_new_n16625__ = ~ys__n1508 & ~new_new_n16624__;
  assign new_new_n16626__ = ys__n1508 & new_new_n16614__;
  assign new_new_n16627__ = ~new_new_n16619__ & new_new_n16626__;
  assign ys__n20045 = new_new_n16625__ | new_new_n16627__;
  assign new_new_n16629__ = ys__n1509 & ~new_new_n16618__;
  assign new_new_n16630__ = ~new_new_n16619__ & new_new_n16629__;
  assign new_new_n16631__ = ~new_new_n16621__ & ~new_new_n16630__;
  assign new_new_n16632__ = ~ys__n1508 & ~new_new_n16631__;
  assign new_new_n16633__ = ys__n1508 & new_new_n16617__;
  assign new_new_n16634__ = ~new_new_n16619__ & new_new_n16633__;
  assign ys__n20040 = new_new_n16632__ | new_new_n16634__;
  assign ys__n33521 = ~ys__n20045 | ~ys__n20040;
  assign new_new_n16637__ = ys__n30216 & ys__n33521;
  assign new_new_n16638__ = ~ys__n18128 & ~new_new_n16637__;
  assign new_new_n16639__ = ~ys__n33515 & ~new_new_n16638__;
  assign ys__n18136 = ~new_new_n16608__ & new_new_n16639__;
  assign new_new_n16641__ = ~ys__n17878 & ~ys__n17879;
  assign new_new_n16642__ = ~ys__n17881 & ~ys__n17882;
  assign new_new_n16643__ = new_new_n16641__ & new_new_n16642__;
  assign new_new_n16644__ = ~ys__n17872 & ~ys__n17873;
  assign new_new_n16645__ = ~ys__n17875 & ~ys__n17876;
  assign new_new_n16646__ = new_new_n16644__ & new_new_n16645__;
  assign new_new_n16647__ = new_new_n16643__ & new_new_n16646__;
  assign new_new_n16648__ = ~ys__n17890 & ~ys__n17891;
  assign new_new_n16649__ = ~ys__n17893 & ~ys__n17894;
  assign new_new_n16650__ = new_new_n16648__ & new_new_n16649__;
  assign new_new_n16651__ = ~ys__n17884 & ~ys__n17885;
  assign new_new_n16652__ = ~ys__n17887 & ~ys__n17888;
  assign new_new_n16653__ = new_new_n16651__ & new_new_n16652__;
  assign new_new_n16654__ = new_new_n16650__ & new_new_n16653__;
  assign new_new_n16655__ = new_new_n16647__ & new_new_n16654__;
  assign new_new_n16656__ = ~ys__n17827 & ~ys__n17828;
  assign new_new_n16657__ = ~ys__n17830 & ~ys__n17831;
  assign new_new_n16658__ = new_new_n16656__ & new_new_n16657__;
  assign new_new_n16659__ = ~ys__n17833 & ~ys__n17834;
  assign new_new_n16660__ = ~ys__n17836 & ~ys__n17837;
  assign new_new_n16661__ = new_new_n16659__ & new_new_n16660__;
  assign new_new_n16662__ = new_new_n16658__ & new_new_n16661__;
  assign new_new_n16663__ = ~ys__n17866 & ~ys__n17867;
  assign new_new_n16664__ = ~ys__n17869 & ~ys__n17870;
  assign new_new_n16665__ = new_new_n16663__ & new_new_n16664__;
  assign new_new_n16666__ = ~ys__n17845 & ~ys__n17846;
  assign new_new_n16667__ = ~ys__n17848 & ~ys__n17849;
  assign new_new_n16668__ = new_new_n16666__ & new_new_n16667__;
  assign new_new_n16669__ = new_new_n16665__ & new_new_n16668__;
  assign new_new_n16670__ = new_new_n16662__ & new_new_n16669__;
  assign new_new_n16671__ = new_new_n16655__ & new_new_n16670__;
  assign new_new_n16672__ = ~ys__n17803 & ~ys__n17804;
  assign new_new_n16673__ = ~ys__n17806 & ~ys__n17807;
  assign new_new_n16674__ = new_new_n16672__ & new_new_n16673__;
  assign new_new_n16675__ = ~ys__n17809 & ~ys__n17810;
  assign new_new_n16676__ = ~ys__n17812 & ~ys__n17813;
  assign new_new_n16677__ = new_new_n16675__ & new_new_n16676__;
  assign new_new_n16678__ = new_new_n16674__ & new_new_n16677__;
  assign new_new_n16679__ = ~ys__n17815 & ~ys__n17816;
  assign new_new_n16680__ = ~ys__n17818 & ~ys__n17819;
  assign new_new_n16681__ = new_new_n16679__ & new_new_n16680__;
  assign new_new_n16682__ = ~ys__n17821 & ~ys__n17822;
  assign new_new_n16683__ = ~ys__n17824 & ~ys__n17825;
  assign new_new_n16684__ = new_new_n16682__ & new_new_n16683__;
  assign new_new_n16685__ = new_new_n16681__ & new_new_n16684__;
  assign new_new_n16686__ = new_new_n16678__ & new_new_n16685__;
  assign new_new_n16687__ = ~ys__n17902 & ~ys__n17903;
  assign new_new_n16688__ = ~ys__n17905 & ~ys__n17906;
  assign new_new_n16689__ = new_new_n16687__ & new_new_n16688__;
  assign new_new_n16690__ = ~ys__n17896 & ~ys__n17897;
  assign new_new_n16691__ = ~ys__n17899 & ~ys__n17900;
  assign new_new_n16692__ = new_new_n16690__ & new_new_n16691__;
  assign new_new_n16693__ = new_new_n16689__ & new_new_n16692__;
  assign new_new_n16694__ = ~ys__n17839 & ~ys__n17840;
  assign new_new_n16695__ = ~ys__n17842 & ~ys__n17843;
  assign new_new_n16696__ = new_new_n16694__ & new_new_n16695__;
  assign new_new_n16697__ = ~ys__n17908 & ~ys__n17909;
  assign new_new_n16698__ = ~ys__n17911 & ~ys__n17912;
  assign new_new_n16699__ = new_new_n16697__ & new_new_n16698__;
  assign new_new_n16700__ = new_new_n16696__ & new_new_n16699__;
  assign new_new_n16701__ = new_new_n16693__ & new_new_n16700__;
  assign new_new_n16702__ = new_new_n16686__ & new_new_n16701__;
  assign new_new_n16703__ = new_new_n16671__ & new_new_n16702__;
  assign ys__n30330 = ys__n17912 & ~ys__n18156;
  assign new_new_n16705__ = ~ys__n404 & ys__n30330;
  assign new_new_n16706__ = ys__n404 & ~ys__n30330;
  assign new_new_n16707__ = ~new_new_n16705__ & ~new_new_n16706__;
  assign ys__n18154 = new_new_n16703__ | ~new_new_n16707__;
  assign ys__n18165 = ys__n948 & ~new_new_n16268__;
  assign new_new_n16710__ = ~ys__n326 & ys__n332;
  assign new_new_n16711__ = new_new_n12322__ & new_new_n16710__;
  assign new_new_n16712__ = ~ys__n336 & new_new_n16711__;
  assign new_new_n16713__ = new_new_n12320__ & new_new_n16710__;
  assign new_new_n16714__ = ~ys__n336 & new_new_n16713__;
  assign new_new_n16715__ = ~new_new_n16712__ & ~new_new_n16714__;
  assign ys__n18169 = ys__n598 & ~new_new_n16715__;
  assign new_new_n16717__ = ys__n26279 & ~ys__n18169;
  assign new_new_n16718__ = ys__n26437 & ~ys__n30941;
  assign new_new_n16719__ = ys__n18169 & new_new_n16718__;
  assign ys__n18170 = new_new_n16717__ | new_new_n16719__;
  assign new_new_n16721__ = new_new_n12313__ & new_new_n16710__;
  assign new_new_n16722__ = ~ys__n336 & new_new_n16721__;
  assign new_new_n16723__ = ~new_new_n16712__ & ~new_new_n16722__;
  assign new_new_n16724__ = ys__n598 & ys__n18173;
  assign ys__n18174 = ~new_new_n16723__ & new_new_n16724__;
  assign new_new_n16726__ = new_new_n12316__ & new_new_n16710__;
  assign new_new_n16727__ = ~ys__n336 & new_new_n16726__;
  assign new_new_n16728__ = ~new_new_n16712__ & ~new_new_n16727__;
  assign ys__n18176 = new_new_n16724__ & ~new_new_n16728__;
  assign ys__n18178 = ~ys__n18208 & new_new_n14022__;
  assign new_new_n16731__ = ~ys__n1508 & ~ys__n1509;
  assign new_new_n16732__ = ~ys__n1511 & new_new_n16731__;
  assign new_new_n16733__ = ys__n20035 & new_new_n16732__;
  assign new_new_n16734__ = ys__n23326 & ys__n28027;
  assign new_new_n16735__ = ~new_new_n10742__ & ~new_new_n10745__;
  assign new_new_n16736__ = ys__n23320 & ys__n28024;
  assign new_new_n16737__ = ys__n23318 & ys__n28023;
  assign new_new_n16738__ = ~new_new_n10738__ & new_new_n16737__;
  assign new_new_n16739__ = ~new_new_n16736__ & ~new_new_n16738__;
  assign new_new_n16740__ = new_new_n16735__ & ~new_new_n16739__;
  assign new_new_n16741__ = ys__n23324 & ys__n28026;
  assign new_new_n16742__ = ys__n23322 & ys__n28025;
  assign new_new_n16743__ = ~new_new_n10745__ & new_new_n16742__;
  assign new_new_n16744__ = ~new_new_n16741__ & ~new_new_n16743__;
  assign new_new_n16745__ = ~new_new_n16740__ & new_new_n16744__;
  assign new_new_n16746__ = ~new_new_n10735__ & ~new_new_n10738__;
  assign new_new_n16747__ = new_new_n16735__ & new_new_n16746__;
  assign new_new_n16748__ = ~new_new_n10696__ & ~new_new_n10699__;
  assign new_new_n16749__ = ~new_new_n10689__ & ~new_new_n10692__;
  assign new_new_n16750__ = new_new_n16748__ & new_new_n16749__;
  assign new_new_n16751__ = ~new_new_n10711__ & ~new_new_n10714__;
  assign new_new_n16752__ = ys__n23304 & ys__n28016;
  assign new_new_n16753__ = ys__n23302 & ys__n28015;
  assign new_new_n16754__ = ~new_new_n10707__ & new_new_n16753__;
  assign new_new_n16755__ = ~new_new_n16752__ & ~new_new_n16754__;
  assign new_new_n16756__ = new_new_n16751__ & ~new_new_n16755__;
  assign new_new_n16757__ = ys__n23308 & ys__n28018;
  assign new_new_n16758__ = ys__n23306 & ys__n28017;
  assign new_new_n16759__ = ~new_new_n10714__ & new_new_n16758__;
  assign new_new_n16760__ = ~new_new_n16757__ & ~new_new_n16759__;
  assign new_new_n16761__ = ~new_new_n16756__ & new_new_n16760__;
  assign new_new_n16762__ = new_new_n16750__ & ~new_new_n16761__;
  assign new_new_n16763__ = ys__n23312 & ys__n28020;
  assign new_new_n16764__ = ys__n23310 & ys__n28019;
  assign new_new_n16765__ = ~new_new_n10692__ & new_new_n16764__;
  assign new_new_n16766__ = ~new_new_n16763__ & ~new_new_n16765__;
  assign new_new_n16767__ = new_new_n16748__ & ~new_new_n16766__;
  assign new_new_n16768__ = ys__n23316 & ys__n28022;
  assign new_new_n16769__ = ys__n23314 & ys__n28021;
  assign new_new_n16770__ = ~new_new_n10699__ & new_new_n16769__;
  assign new_new_n16771__ = ~new_new_n16768__ & ~new_new_n16770__;
  assign new_new_n16772__ = ~new_new_n16767__ & new_new_n16771__;
  assign new_new_n16773__ = ~new_new_n16762__ & new_new_n16772__;
  assign new_new_n16774__ = ~new_new_n10704__ & ~new_new_n10707__;
  assign new_new_n16775__ = new_new_n16751__ & new_new_n16774__;
  assign new_new_n16776__ = new_new_n16750__ & new_new_n16775__;
  assign new_new_n16777__ = ys__n23272 & ys__n27857;
  assign new_new_n16778__ = ~new_new_n10770__ & new_new_n16609__;
  assign new_new_n16779__ = ~new_new_n16777__ & ~new_new_n16778__;
  assign new_new_n16780__ = ~new_new_n10774__ & ~new_new_n10777__;
  assign new_new_n16781__ = ~new_new_n16779__ & new_new_n16780__;
  assign new_new_n16782__ = ys__n23276 & ys__n27861;
  assign new_new_n16783__ = ys__n23274 & ys__n27859;
  assign new_new_n16784__ = ~new_new_n10777__ & new_new_n16783__;
  assign new_new_n16785__ = ~new_new_n16782__ & ~new_new_n16784__;
  assign new_new_n16786__ = ~new_new_n16781__ & new_new_n16785__;
  assign new_new_n16787__ = ~new_new_n10759__ & ~new_new_n10762__;
  assign new_new_n16788__ = ~new_new_n10752__ & ~new_new_n10755__;
  assign new_new_n16789__ = new_new_n16787__ & new_new_n16788__;
  assign new_new_n16790__ = ~new_new_n16786__ & new_new_n16789__;
  assign new_new_n16791__ = ys__n23280 & ys__n27865;
  assign new_new_n16792__ = ys__n23278 & ys__n27863;
  assign new_new_n16793__ = ~new_new_n10755__ & new_new_n16792__;
  assign new_new_n16794__ = ~new_new_n16791__ & ~new_new_n16793__;
  assign new_new_n16795__ = new_new_n16787__ & ~new_new_n16794__;
  assign new_new_n16796__ = ys__n23284 & ys__n27869;
  assign new_new_n16797__ = ys__n23282 & ys__n27867;
  assign new_new_n16798__ = ~new_new_n10762__ & new_new_n16797__;
  assign new_new_n16799__ = ~new_new_n16796__ & ~new_new_n16798__;
  assign new_new_n16800__ = ~new_new_n16795__ & new_new_n16799__;
  assign new_new_n16801__ = ~new_new_n16790__ & new_new_n16800__;
  assign new_new_n16802__ = ~new_new_n10790__ & ~new_new_n10793__;
  assign new_new_n16803__ = ~new_new_n10783__ & ~new_new_n10786__;
  assign new_new_n16804__ = new_new_n16802__ & new_new_n16803__;
  assign new_new_n16805__ = ~new_new_n10805__ & ~new_new_n10808__;
  assign new_new_n16806__ = ~new_new_n10798__ & ~new_new_n10801__;
  assign new_new_n16807__ = new_new_n16805__ & new_new_n16806__;
  assign new_new_n16808__ = new_new_n16804__ & new_new_n16807__;
  assign new_new_n16809__ = ~new_new_n16801__ & new_new_n16808__;
  assign new_new_n16810__ = ys__n23288 & ys__n27873;
  assign new_new_n16811__ = ys__n23286 & ys__n27871;
  assign new_new_n16812__ = ~new_new_n10801__ & new_new_n16811__;
  assign new_new_n16813__ = ~new_new_n16810__ & ~new_new_n16812__;
  assign new_new_n16814__ = new_new_n16805__ & ~new_new_n16813__;
  assign new_new_n16815__ = ys__n23292 & ys__n27877;
  assign new_new_n16816__ = ys__n23290 & ys__n27875;
  assign new_new_n16817__ = ~new_new_n10808__ & new_new_n16816__;
  assign new_new_n16818__ = ~new_new_n16815__ & ~new_new_n16817__;
  assign new_new_n16819__ = ~new_new_n16814__ & new_new_n16818__;
  assign new_new_n16820__ = new_new_n16804__ & ~new_new_n16819__;
  assign new_new_n16821__ = ys__n23296 & ys__n27881;
  assign new_new_n16822__ = ys__n23294 & ys__n27879;
  assign new_new_n16823__ = ~new_new_n10786__ & new_new_n16822__;
  assign new_new_n16824__ = ~new_new_n16821__ & ~new_new_n16823__;
  assign new_new_n16825__ = new_new_n16802__ & ~new_new_n16824__;
  assign new_new_n16826__ = ys__n23300 & ys__n27885;
  assign new_new_n16827__ = ys__n23298 & ys__n27883;
  assign new_new_n16828__ = ~new_new_n10793__ & new_new_n16827__;
  assign new_new_n16829__ = ~new_new_n16826__ & ~new_new_n16828__;
  assign new_new_n16830__ = ~new_new_n16825__ & new_new_n16829__;
  assign new_new_n16831__ = ~new_new_n16820__ & new_new_n16830__;
  assign new_new_n16832__ = ~new_new_n16809__ & new_new_n16831__;
  assign new_new_n16833__ = new_new_n16776__ & ~new_new_n16832__;
  assign new_new_n16834__ = new_new_n16773__ & ~new_new_n16833__;
  assign new_new_n16835__ = new_new_n16747__ & ~new_new_n16834__;
  assign new_new_n16836__ = new_new_n16745__ & ~new_new_n16835__;
  assign new_new_n16837__ = ~new_new_n10720__ & ~new_new_n16836__;
  assign new_new_n16838__ = ~new_new_n16734__ & ~new_new_n16837__;
  assign new_new_n16839__ = new_new_n10723__ & ~new_new_n16838__;
  assign new_new_n16840__ = ~new_new_n10723__ & new_new_n16838__;
  assign new_new_n16841__ = ~new_new_n16839__ & ~new_new_n16840__;
  assign new_new_n16842__ = ~new_new_n16732__ & ~new_new_n16841__;
  assign ys__n18214 = new_new_n16733__ | new_new_n16842__;
  assign new_new_n16844__ = ys__n23328 & ys__n28028;
  assign new_new_n16845__ = ~new_new_n10723__ & new_new_n16734__;
  assign new_new_n16846__ = ~new_new_n16844__ & ~new_new_n16845__;
  assign new_new_n16847__ = ~new_new_n10720__ & ~new_new_n10723__;
  assign new_new_n16848__ = ~new_new_n16836__ & new_new_n16847__;
  assign new_new_n16849__ = new_new_n16846__ & ~new_new_n16848__;
  assign new_new_n16850__ = new_new_n10727__ & ~new_new_n16849__;
  assign new_new_n16851__ = ~new_new_n10727__ & new_new_n16849__;
  assign new_new_n16852__ = ~new_new_n16850__ & ~new_new_n16851__;
  assign new_new_n16853__ = ~new_new_n16732__ & ~new_new_n16852__;
  assign ys__n18216 = new_new_n16733__ | new_new_n16853__;
  assign ys__n18217 = ys__n874 & ys__n18216;
  assign new_new_n16856__ = ys__n23330 & ys__n28029;
  assign new_new_n16857__ = ~new_new_n10727__ & ~new_new_n16849__;
  assign new_new_n16858__ = ~new_new_n16856__ & ~new_new_n16857__;
  assign new_new_n16859__ = new_new_n10730__ & ~new_new_n16858__;
  assign new_new_n16860__ = ~new_new_n10730__ & new_new_n16858__;
  assign new_new_n16861__ = ~new_new_n16859__ & ~new_new_n16860__;
  assign new_new_n16862__ = ~new_new_n16732__ & ~new_new_n16861__;
  assign ys__n18218 = new_new_n16733__ | new_new_n16862__;
  assign ys__n18241 = ~ys__n33548 & ys__n4764;
  assign new_new_n16865__ = ys__n18242 & ~ys__n18241;
  assign new_new_n16866__ = ys__n98 & ys__n18241;
  assign new_new_n16867__ = ~new_new_n16865__ & ~new_new_n16866__;
  assign ys__n18223 = ys__n874 & ~new_new_n16867__;
  assign new_new_n16869__ = ~ys__n18227 & ys__n18214;
  assign new_new_n16870__ = ys__n18226 & ys__n18227;
  assign new_new_n16871__ = ~new_new_n16869__ & ~new_new_n16870__;
  assign new_new_n16872__ = ys__n874 & ~new_new_n16871__;
  assign new_new_n16873__ = ~ys__n18227 & ys__n18218;
  assign new_new_n16874__ = ys__n18231 & ys__n18227;
  assign new_new_n16875__ = ~new_new_n16873__ & ~new_new_n16874__;
  assign new_new_n16876__ = ys__n874 & ~new_new_n16875__;
  assign new_new_n16877__ = new_new_n16872__ & ~new_new_n16876__;
  assign new_new_n16878__ = ~ys__n18227 & ys__n18216;
  assign new_new_n16879__ = ys__n18229 & ys__n18227;
  assign new_new_n16880__ = ~new_new_n16878__ & ~new_new_n16879__;
  assign ys__n18238 = ys__n874 & ~new_new_n16880__;
  assign new_new_n16882__ = new_new_n16872__ & ys__n18238;
  assign new_new_n16883__ = new_new_n16876__ & new_new_n16882__;
  assign ys__n18236 = new_new_n16877__ | new_new_n16883__;
  assign new_new_n16885__ = ~new_new_n16876__ & ~ys__n18238;
  assign new_new_n16886__ = new_new_n16876__ & ys__n18238;
  assign ys__n18239 = new_new_n16885__ | new_new_n16886__;
  assign new_new_n16888__ = ys__n29886 & ~new_new_n10603__;
  assign new_new_n16889__ = ~new_new_n10601__ & new_new_n16888__;
  assign new_new_n16890__ = ~ys__n23764 & new_new_n16889__;
  assign new_new_n16891__ = ys__n29902 & ~new_new_n10603__;
  assign new_new_n16892__ = ~new_new_n10601__ & new_new_n16891__;
  assign new_new_n16893__ = ~ys__n22466 & new_new_n16892__;
  assign new_new_n16894__ = ys__n22466 & new_new_n16889__;
  assign new_new_n16895__ = ~new_new_n16893__ & ~new_new_n16894__;
  assign new_new_n16896__ = ys__n23764 & ~new_new_n16895__;
  assign new_new_n16897__ = ~new_new_n16890__ & ~new_new_n16896__;
  assign ys__n25388 = new_new_n10866__ & ~new_new_n16897__;
  assign new_new_n16899__ = ~ys__n19256 & ys__n25388;
  assign new_new_n16900__ = ys__n530 & ys__n19256;
  assign new_new_n16901__ = ~new_new_n16899__ & ~new_new_n16900__;
  assign ys__n18251 = ys__n874 & ~new_new_n16901__;
  assign new_new_n16903__ = ys__n29893 & ~new_new_n10603__;
  assign new_new_n16904__ = ~new_new_n10601__ & new_new_n16903__;
  assign new_new_n16905__ = ~ys__n23764 & new_new_n16904__;
  assign new_new_n16906__ = ys__n29909 & ~new_new_n10603__;
  assign new_new_n16907__ = ~new_new_n10601__ & new_new_n16906__;
  assign new_new_n16908__ = ~ys__n22466 & new_new_n16907__;
  assign new_new_n16909__ = ys__n22466 & new_new_n16904__;
  assign new_new_n16910__ = ~new_new_n16908__ & ~new_new_n16909__;
  assign new_new_n16911__ = ys__n23764 & ~new_new_n16910__;
  assign new_new_n16912__ = ~new_new_n16905__ & ~new_new_n16911__;
  assign ys__n25432 = new_new_n10866__ & ~new_new_n16912__;
  assign new_new_n16914__ = ~ys__n19256 & ys__n25432;
  assign new_new_n16915__ = ys__n640 & ys__n19256;
  assign new_new_n16916__ = ~new_new_n16914__ & ~new_new_n16915__;
  assign ys__n18360 = ~ys__n874 | new_new_n16916__;
  assign new_new_n16918__ = ~new_new_n12143__ & ys__n18360;
  assign ys__n18268 = new_new_n12127__ & new_new_n16918__;
  assign ys__n18273 = ys__n18271 | ys__n4414;
  assign new_new_n16921__ = ~ys__n846 & ~ys__n4185;
  assign new_new_n16922__ = ~ys__n4625 & new_new_n16921__;
  assign new_new_n16923__ = new_new_n11041__ & new_new_n16922__;
  assign new_new_n16924__ = new_new_n12227__ & new_new_n16923__;
  assign new_new_n16925__ = ~ys__n4613 & new_new_n16924__;
  assign ys__n18303 = ys__n38522 | new_new_n16925__;
  assign new_new_n16927__ = ~ys__n18317 & ~ys__n33300;
  assign new_new_n16928__ = ys__n37692 & new_new_n16927__;
  assign new_new_n16929__ = ys__n3214 & ys__n33311;
  assign new_new_n16930__ = ~new_new_n12098__ & new_new_n16929__;
  assign new_new_n16931__ = ~ys__n37692 & ~new_new_n16930__;
  assign new_new_n16932__ = ys__n18317 & ~new_new_n16931__;
  assign ys__n18321 = new_new_n16928__ | new_new_n16932__;
  assign new_new_n16934__ = ys__n863 & ~new_new_n12108__;
  assign new_new_n16935__ = ys__n842 & new_new_n12108__;
  assign ys__n18329 = new_new_n16934__ | new_new_n16935__;
  assign new_new_n16937__ = ys__n844 & ys__n863;
  assign new_new_n16938__ = ~new_new_n12108__ & new_new_n16937__;
  assign new_new_n16939__ = ys__n840 & new_new_n12108__;
  assign ys__n18331 = new_new_n16938__ | new_new_n16939__;
  assign new_new_n16941__ = ys__n842 & ys__n863;
  assign new_new_n16942__ = ~new_new_n12108__ & new_new_n16941__;
  assign new_new_n16943__ = ys__n838 & new_new_n12108__;
  assign ys__n18333 = new_new_n16942__ | new_new_n16943__;
  assign new_new_n16945__ = ys__n840 & ys__n863;
  assign new_new_n16946__ = ~new_new_n12108__ & new_new_n16945__;
  assign new_new_n16947__ = ys__n836 & new_new_n12108__;
  assign ys__n18335 = new_new_n16946__ | new_new_n16947__;
  assign new_new_n16949__ = ys__n838 & ys__n863;
  assign new_new_n16950__ = ~new_new_n12108__ & new_new_n16949__;
  assign new_new_n16951__ = ys__n834 & new_new_n12108__;
  assign ys__n18337 = new_new_n16950__ | new_new_n16951__;
  assign new_new_n16953__ = ys__n836 & ys__n863;
  assign new_new_n16954__ = ~new_new_n12108__ & new_new_n16953__;
  assign new_new_n16955__ = ys__n832 & new_new_n12108__;
  assign ys__n18339 = new_new_n16954__ | new_new_n16955__;
  assign new_new_n16957__ = ys__n834 & ys__n863;
  assign new_new_n16958__ = ~new_new_n12108__ & new_new_n16957__;
  assign new_new_n16959__ = ys__n830 & new_new_n12108__;
  assign ys__n18341 = new_new_n16958__ | new_new_n16959__;
  assign new_new_n16961__ = ys__n832 & ys__n863;
  assign new_new_n16962__ = ~new_new_n12108__ & new_new_n16961__;
  assign new_new_n16963__ = ys__n858 & new_new_n12108__;
  assign ys__n18343 = new_new_n16962__ | new_new_n16963__;
  assign new_new_n16965__ = ys__n830 & ys__n863;
  assign new_new_n16966__ = ~new_new_n12108__ & new_new_n16965__;
  assign new_new_n16967__ = ys__n856 & new_new_n12108__;
  assign ys__n18345 = new_new_n16966__ | new_new_n16967__;
  assign new_new_n16969__ = ys__n858 & ys__n863;
  assign new_new_n16970__ = ~new_new_n12108__ & new_new_n16969__;
  assign new_new_n16971__ = ys__n854 & new_new_n12108__;
  assign ys__n18347 = new_new_n16970__ | new_new_n16971__;
  assign new_new_n16973__ = ys__n856 & ys__n863;
  assign new_new_n16974__ = ~new_new_n12108__ & new_new_n16973__;
  assign new_new_n16975__ = ys__n852 & new_new_n12108__;
  assign ys__n18349 = new_new_n16974__ | new_new_n16975__;
  assign new_new_n16977__ = ys__n854 & ys__n863;
  assign new_new_n16978__ = ~new_new_n12108__ & new_new_n16977__;
  assign new_new_n16979__ = ys__n850 & new_new_n12108__;
  assign ys__n18351 = new_new_n16978__ | new_new_n16979__;
  assign new_new_n16981__ = ys__n852 & ys__n863;
  assign new_new_n16982__ = ~new_new_n12108__ & new_new_n16981__;
  assign new_new_n16983__ = ys__n848 & new_new_n12108__;
  assign ys__n18353 = new_new_n16982__ | new_new_n16983__;
  assign new_new_n16985__ = ys__n850 & ys__n863;
  assign new_new_n16986__ = ~new_new_n12108__ & new_new_n16985__;
  assign new_new_n16987__ = ys__n846 & new_new_n12108__;
  assign ys__n18355 = new_new_n16986__ | new_new_n16987__;
  assign new_new_n16989__ = ys__n848 & ys__n863;
  assign new_new_n16990__ = ~new_new_n12108__ & new_new_n16989__;
  assign new_new_n16991__ = ys__n116 & new_new_n12108__;
  assign ys__n18357 = new_new_n16990__ | new_new_n16991__;
  assign new_new_n16993__ = ys__n18378 & ~ys__n18078;
  assign new_new_n16994__ = ~ys__n18393 & ys__n18544;
  assign new_new_n16995__ = ys__n19156 & ys__n18287;
  assign new_new_n16996__ = ~ys__n18284 & new_new_n16995__;
  assign new_new_n16997__ = ys__n18749 & ~new_new_n11122__;
  assign new_new_n16998__ = ~ys__n33552 & ~new_new_n11121__;
  assign new_new_n16999__ = ~ys__n18759 & ~new_new_n16998__;
  assign new_new_n17000__ = ~ys__n38894 & ~new_new_n16999__;
  assign new_new_n17001__ = ~ys__n38861 & ~new_new_n16999__;
  assign new_new_n17002__ = ~new_new_n17000__ & ~new_new_n17001__;
  assign new_new_n17003__ = ~ys__n38893 & ~new_new_n16999__;
  assign new_new_n17004__ = ~ys__n38862 & ~new_new_n16999__;
  assign new_new_n17005__ = new_new_n17003__ & new_new_n17004__;
  assign new_new_n17006__ = new_new_n17002__ & new_new_n17005__;
  assign new_new_n17007__ = ~new_new_n17003__ & ~new_new_n17004__;
  assign new_new_n17008__ = new_new_n17002__ & new_new_n17007__;
  assign new_new_n17009__ = new_new_n17000__ & new_new_n17001__;
  assign new_new_n17010__ = new_new_n17007__ & new_new_n17009__;
  assign new_new_n17011__ = ~new_new_n17008__ & ~new_new_n17010__;
  assign ys__n18750 = new_new_n17006__ | ~new_new_n17011__;
  assign new_new_n17013__ = new_new_n11122__ & ys__n18750;
  assign ys__n18751 = new_new_n16997__ | new_new_n17013__;
  assign new_new_n17015__ = ys__n18284 & ys__n18751;
  assign new_new_n17016__ = ~new_new_n16996__ & ~new_new_n17015__;
  assign new_new_n17017__ = ~ys__n18281 & ~new_new_n17016__;
  assign new_new_n17018__ = ~ys__n18281 & ~new_new_n17017__;
  assign new_new_n17019__ = ~ys__n18278 & ~new_new_n17018__;
  assign new_new_n17020__ = ~ys__n35049 & ys__n46214;
  assign new_new_n17021__ = ys__n30957 & ~new_new_n17020__;
  assign new_new_n17022__ = ys__n26557 & ~ys__n26558;
  assign new_new_n17023__ = ~ys__n26557 & ys__n26558;
  assign new_new_n17024__ = ~new_new_n17022__ & ~new_new_n17023__;
  assign new_new_n17025__ = new_new_n17020__ & ~new_new_n17024__;
  assign ys__n19149 = new_new_n17021__ | new_new_n17025__;
  assign new_new_n17027__ = ys__n18278 & ys__n19149;
  assign ys__n18545 = new_new_n17019__ | new_new_n17027__;
  assign new_new_n17029__ = ys__n18393 & ys__n18545;
  assign new_new_n17030__ = ~new_new_n16994__ & ~new_new_n17029__;
  assign new_new_n17031__ = ys__n18078 & ~new_new_n17030__;
  assign ys__n18380 = new_new_n16993__ | new_new_n17031__;
  assign new_new_n17033__ = ys__n18381 & ~ys__n18078;
  assign new_new_n17034__ = ~ys__n18393 & ys__n18546;
  assign new_new_n17035__ = ys__n19157 & ys__n18287;
  assign new_new_n17036__ = ~ys__n18284 & new_new_n17035__;
  assign new_new_n17037__ = ys__n18752 & ~new_new_n11122__;
  assign ys__n18753 = new_new_n17008__ & ys__n18750;
  assign new_new_n17039__ = new_new_n11122__ & ys__n18753;
  assign ys__n18754 = new_new_n17037__ | new_new_n17039__;
  assign new_new_n17041__ = ys__n18284 & ys__n18754;
  assign new_new_n17042__ = ~new_new_n17036__ & ~new_new_n17041__;
  assign new_new_n17043__ = ~ys__n18281 & ~new_new_n17042__;
  assign new_new_n17044__ = ~ys__n18281 & ~new_new_n17043__;
  assign new_new_n17045__ = ~ys__n18278 & ~new_new_n17044__;
  assign new_new_n17046__ = ys__n30960 & ~new_new_n17020__;
  assign new_new_n17047__ = ys__n26558 & new_new_n17020__;
  assign ys__n19151 = new_new_n17046__ | new_new_n17047__;
  assign new_new_n17049__ = ys__n18278 & ys__n19151;
  assign ys__n18547 = new_new_n17045__ | new_new_n17049__;
  assign new_new_n17051__ = ys__n18393 & ys__n18547;
  assign new_new_n17052__ = ~new_new_n17034__ & ~new_new_n17051__;
  assign new_new_n17053__ = ys__n18078 & ~new_new_n17052__;
  assign ys__n18383 = new_new_n17033__ | new_new_n17053__;
  assign new_new_n17055__ = ys__n18384 & ~ys__n18078;
  assign new_new_n17056__ = ys__n18208 & ~ys__n18393;
  assign new_new_n17057__ = ys__n18284 & ~ys__n18281;
  assign new_new_n17058__ = ~ys__n18281 & ~new_new_n17057__;
  assign new_new_n17059__ = ~ys__n18278 & ~new_new_n17058__;
  assign new_new_n17060__ = ys__n30961 & ~new_new_n17020__;
  assign new_new_n17061__ = ys__n26559 & new_new_n17020__;
  assign ys__n19159 = new_new_n17060__ | new_new_n17061__;
  assign new_new_n17063__ = ys__n18278 & ys__n19159;
  assign ys__n18555 = new_new_n17059__ | new_new_n17063__;
  assign new_new_n17065__ = ys__n18393 & ys__n18555;
  assign new_new_n17066__ = ~new_new_n17056__ & ~new_new_n17065__;
  assign new_new_n17067__ = ys__n18078 & ~new_new_n17066__;
  assign ys__n33324 = ~new_new_n17055__ & ~new_new_n17067__;
  assign new_new_n17069__ = ys__n18389 & ~ys__n18078;
  assign new_new_n17070__ = ~ys__n18393 & ys__n18556;
  assign new_new_n17071__ = ys__n18755 & ~new_new_n11122__;
  assign new_new_n17072__ = ~ys__n38864 & ~new_new_n11115__;
  assign new_new_n17073__ = ~ys__n24675 & ~ys__n18759;
  assign new_new_n17074__ = ~new_new_n17072__ & new_new_n17073__;
  assign new_new_n17075__ = new_new_n11122__ & new_new_n17074__;
  assign ys__n18757 = new_new_n17071__ | new_new_n17075__;
  assign new_new_n17077__ = ~ys__n18281 & ys__n18757;
  assign new_new_n17078__ = ys__n18284 & new_new_n17077__;
  assign new_new_n17079__ = ys__n18647 & ~new_new_n11125__;
  assign new_new_n17080__ = ys__n96 & ~ys__n98;
  assign new_new_n17081__ = ys__n100 & new_new_n17080__;
  assign new_new_n17082__ = ys__n78 & ys__n96;
  assign new_new_n17083__ = ys__n98 & ys__n100;
  assign new_new_n17084__ = new_new_n17082__ & new_new_n17083__;
  assign new_new_n17085__ = ys__n70 & ys__n72;
  assign new_new_n17086__ = ys__n74 & ys__n76;
  assign new_new_n17087__ = new_new_n17085__ & new_new_n17086__;
  assign new_new_n17088__ = new_new_n17084__ & new_new_n17087__;
  assign new_new_n17089__ = ~new_new_n17081__ & ~new_new_n17088__;
  assign new_new_n17090__ = new_new_n11125__ & ~new_new_n17089__;
  assign ys__n18649 = new_new_n17079__ | new_new_n17090__;
  assign new_new_n17092__ = ys__n18281 & ~ys__n18649;
  assign new_new_n17093__ = ~new_new_n17078__ & ~new_new_n17092__;
  assign ys__n18557 = ~ys__n18278 & ~new_new_n17093__;
  assign new_new_n17095__ = ys__n18393 & ys__n18557;
  assign new_new_n17096__ = ~new_new_n17070__ & ~new_new_n17095__;
  assign new_new_n17097__ = ys__n18078 & ~new_new_n17096__;
  assign ys__n33317 = ~new_new_n17069__ & ~new_new_n17097__;
  assign new_new_n17099__ = ys__n18956 & ys__n18287;
  assign new_new_n17100__ = ~ys__n18284 & new_new_n17099__;
  assign new_new_n17101__ = ys__n24615 & ~ys__n4764;
  assign new_new_n17102__ = ys__n24616 & ys__n4764;
  assign ys__n18764 = new_new_n17101__ | new_new_n17102__;
  assign new_new_n17104__ = ~ys__n18071 & ys__n18764;
  assign new_new_n17105__ = ys__n18071 & ys__n18765;
  assign new_new_n17106__ = ~new_new_n17104__ & ~new_new_n17105__;
  assign new_new_n17107__ = ~new_new_n11122__ & ~new_new_n17106__;
  assign new_new_n17108__ = ys__n24616 & ~ys__n24675;
  assign new_new_n17109__ = ys__n24674 & ys__n24675;
  assign new_new_n17110__ = ~new_new_n17108__ & ~new_new_n17109__;
  assign ys__n18654 = ~new_new_n16999__ & ~new_new_n17110__;
  assign new_new_n17112__ = new_new_n11122__ & ys__n18654;
  assign ys__n18655 = new_new_n17107__ | new_new_n17112__;
  assign new_new_n17114__ = ys__n18284 & ys__n18655;
  assign new_new_n17115__ = ~new_new_n17100__ & ~new_new_n17114__;
  assign new_new_n17116__ = ~ys__n18281 & ~new_new_n17115__;
  assign ys__n18559 = ys__n18558 & ~new_new_n11125__;
  assign new_new_n17118__ = ys__n18281 & ys__n18559;
  assign new_new_n17119__ = ~new_new_n17116__ & ~new_new_n17118__;
  assign new_new_n17120__ = ~ys__n18278 & ~new_new_n17119__;
  assign new_new_n17121__ = ys__n18829 & ys__n18278;
  assign ys__n18392 = new_new_n17120__ | new_new_n17121__;
  assign new_new_n17123__ = ys__n6112 & ~ys__n18393;
  assign new_new_n17124__ = ys__n18393 & ys__n18392;
  assign ys__n18394 = new_new_n17123__ | new_new_n17124__;
  assign new_new_n17126__ = ys__n18957 & ys__n18287;
  assign new_new_n17127__ = ~ys__n18284 & new_new_n17126__;
  assign new_new_n17128__ = ys__n24617 & ~ys__n4764;
  assign new_new_n17129__ = ys__n24618 & ys__n4764;
  assign ys__n18766 = new_new_n17128__ | new_new_n17129__;
  assign new_new_n17131__ = ~ys__n18071 & ys__n18766;
  assign new_new_n17132__ = ys__n18071 & ys__n18767;
  assign new_new_n17133__ = ~new_new_n17131__ & ~new_new_n17132__;
  assign new_new_n17134__ = ~new_new_n11122__ & ~new_new_n17133__;
  assign new_new_n17135__ = ys__n24618 & ~ys__n24675;
  assign new_new_n17136__ = ys__n24675 & ys__n24677;
  assign new_new_n17137__ = ~new_new_n17135__ & ~new_new_n17136__;
  assign ys__n18657 = ~new_new_n16999__ & ~new_new_n17137__;
  assign new_new_n17139__ = new_new_n11122__ & ys__n18657;
  assign ys__n18658 = new_new_n17134__ | new_new_n17139__;
  assign new_new_n17141__ = ys__n18284 & ys__n18658;
  assign new_new_n17142__ = ~new_new_n17127__ & ~new_new_n17141__;
  assign new_new_n17143__ = ~ys__n18281 & ~new_new_n17142__;
  assign ys__n18561 = ys__n18560 & ~new_new_n11125__;
  assign new_new_n17145__ = ys__n18281 & ys__n18561;
  assign new_new_n17146__ = ~new_new_n17143__ & ~new_new_n17145__;
  assign new_new_n17147__ = ~ys__n18278 & ~new_new_n17146__;
  assign new_new_n17148__ = ys__n18831 & ys__n18278;
  assign ys__n18395 = new_new_n17147__ | new_new_n17148__;
  assign new_new_n17150__ = ys__n6113 & ~ys__n18393;
  assign new_new_n17151__ = ys__n18393 & ys__n18395;
  assign ys__n18396 = new_new_n17150__ | new_new_n17151__;
  assign new_new_n17153__ = ys__n18958 & ys__n18287;
  assign new_new_n17154__ = ~ys__n18284 & new_new_n17153__;
  assign new_new_n17155__ = ys__n24619 & ~ys__n4764;
  assign new_new_n17156__ = ys__n24620 & ys__n4764;
  assign ys__n18768 = new_new_n17155__ | new_new_n17156__;
  assign new_new_n17158__ = ~ys__n18071 & ys__n18768;
  assign new_new_n17159__ = ys__n18071 & ys__n18769;
  assign new_new_n17160__ = ~new_new_n17158__ & ~new_new_n17159__;
  assign new_new_n17161__ = ~new_new_n11122__ & ~new_new_n17160__;
  assign new_new_n17162__ = ys__n24620 & ~ys__n24675;
  assign new_new_n17163__ = ys__n24675 & ys__n24679;
  assign new_new_n17164__ = ~new_new_n17162__ & ~new_new_n17163__;
  assign new_new_n17165__ = ys__n24107 & new_new_n17074__;
  assign ys__n18660 = ~new_new_n17164__ & ~new_new_n17165__;
  assign new_new_n17167__ = new_new_n11122__ & ys__n18660;
  assign ys__n18661 = new_new_n17161__ | new_new_n17167__;
  assign new_new_n17169__ = ys__n18284 & ys__n18661;
  assign new_new_n17170__ = ~new_new_n17154__ & ~new_new_n17169__;
  assign new_new_n17171__ = ~ys__n18281 & ~new_new_n17170__;
  assign new_new_n17172__ = ys__n18562 & ~new_new_n11125__;
  assign new_new_n17173__ = ys__n24107 & new_new_n17089__;
  assign new_new_n17174__ = ys__n38896 & new_new_n11125__;
  assign new_new_n17175__ = ~new_new_n17173__ & new_new_n17174__;
  assign ys__n18564 = new_new_n17172__ | new_new_n17175__;
  assign new_new_n17177__ = ys__n18281 & ys__n18564;
  assign new_new_n17178__ = ~new_new_n17171__ & ~new_new_n17177__;
  assign new_new_n17179__ = ~ys__n18278 & ~new_new_n17178__;
  assign new_new_n17180__ = ys__n18833 & ys__n18278;
  assign ys__n18397 = new_new_n17179__ | new_new_n17180__;
  assign new_new_n17182__ = ys__n172 & ~ys__n18393;
  assign new_new_n17183__ = ys__n18393 & ys__n18397;
  assign ys__n18398 = new_new_n17182__ | new_new_n17183__;
  assign new_new_n17185__ = ys__n18959 & ys__n18287;
  assign new_new_n17186__ = ~ys__n18284 & new_new_n17185__;
  assign new_new_n17187__ = ys__n24621 & ~ys__n4764;
  assign new_new_n17188__ = ys__n24622 & ys__n4764;
  assign ys__n18770 = new_new_n17187__ | new_new_n17188__;
  assign new_new_n17190__ = ~ys__n18071 & ys__n18770;
  assign new_new_n17191__ = ys__n18071 & ys__n18771;
  assign new_new_n17192__ = ~new_new_n17190__ & ~new_new_n17191__;
  assign new_new_n17193__ = ~new_new_n11122__ & ~new_new_n17192__;
  assign new_new_n17194__ = ys__n24622 & ~ys__n24675;
  assign new_new_n17195__ = ys__n24675 & ys__n24681;
  assign new_new_n17196__ = ~new_new_n17194__ & ~new_new_n17195__;
  assign ys__n18663 = ~new_new_n17165__ & ~new_new_n17196__;
  assign new_new_n17198__ = new_new_n11122__ & ys__n18663;
  assign ys__n18664 = new_new_n17193__ | new_new_n17198__;
  assign new_new_n17200__ = ys__n18284 & ys__n18664;
  assign new_new_n17201__ = ~new_new_n17186__ & ~new_new_n17200__;
  assign new_new_n17202__ = ~ys__n18281 & ~new_new_n17201__;
  assign new_new_n17203__ = ys__n18565 & ~new_new_n11125__;
  assign new_new_n17204__ = ys__n38897 & new_new_n11125__;
  assign new_new_n17205__ = ~new_new_n17173__ & new_new_n17204__;
  assign ys__n18567 = new_new_n17203__ | new_new_n17205__;
  assign new_new_n17207__ = ys__n18281 & ys__n18567;
  assign new_new_n17208__ = ~new_new_n17202__ & ~new_new_n17207__;
  assign new_new_n17209__ = ~ys__n18278 & ~new_new_n17208__;
  assign new_new_n17210__ = ys__n18835 & ys__n18278;
  assign ys__n18399 = new_new_n17209__ | new_new_n17210__;
  assign new_new_n17212__ = ys__n338 & ~ys__n18393;
  assign new_new_n17213__ = ys__n18393 & ys__n18399;
  assign ys__n18400 = new_new_n17212__ | new_new_n17213__;
  assign new_new_n17215__ = ys__n18960 & ys__n18287;
  assign new_new_n17216__ = ~ys__n18284 & new_new_n17215__;
  assign new_new_n17217__ = ys__n24623 & ~ys__n4764;
  assign new_new_n17218__ = ys__n24624 & ys__n4764;
  assign ys__n18772 = new_new_n17217__ | new_new_n17218__;
  assign new_new_n17220__ = ~ys__n18071 & ys__n18772;
  assign new_new_n17221__ = ys__n18071 & ys__n18773;
  assign new_new_n17222__ = ~new_new_n17220__ & ~new_new_n17221__;
  assign new_new_n17223__ = ~new_new_n11122__ & ~new_new_n17222__;
  assign new_new_n17224__ = ys__n24624 & ~ys__n24675;
  assign new_new_n17225__ = ys__n24675 & ys__n24683;
  assign ys__n18666 = new_new_n17224__ | new_new_n17225__;
  assign new_new_n17227__ = new_new_n11122__ & ys__n18666;
  assign ys__n18667 = new_new_n17223__ | new_new_n17227__;
  assign new_new_n17229__ = ys__n18284 & ys__n18667;
  assign new_new_n17230__ = ~new_new_n17216__ & ~new_new_n17229__;
  assign new_new_n17231__ = ~ys__n18281 & ~new_new_n17230__;
  assign new_new_n17232__ = ys__n18568 & ~new_new_n11125__;
  assign new_new_n17233__ = ys__n18569 & new_new_n11125__;
  assign ys__n18570 = new_new_n17232__ | new_new_n17233__;
  assign new_new_n17235__ = ys__n18281 & ys__n18570;
  assign new_new_n17236__ = ~new_new_n17231__ & ~new_new_n17235__;
  assign new_new_n17237__ = ~ys__n18278 & ~new_new_n17236__;
  assign new_new_n17238__ = ys__n18837 & ys__n18278;
  assign ys__n18401 = new_new_n17237__ | new_new_n17238__;
  assign new_new_n17240__ = ys__n22 & ~ys__n18393;
  assign new_new_n17241__ = ys__n18393 & ys__n18401;
  assign ys__n18402 = new_new_n17240__ | new_new_n17241__;
  assign new_new_n17243__ = ys__n18961 & ys__n18287;
  assign new_new_n17244__ = ~ys__n18284 & new_new_n17243__;
  assign new_new_n17245__ = ys__n24625 & ~ys__n4764;
  assign new_new_n17246__ = ys__n24626 & ys__n4764;
  assign ys__n18774 = new_new_n17245__ | new_new_n17246__;
  assign new_new_n17248__ = ~ys__n18071 & ys__n18774;
  assign new_new_n17249__ = ys__n18071 & ys__n18775;
  assign new_new_n17250__ = ~new_new_n17248__ & ~new_new_n17249__;
  assign new_new_n17251__ = ~new_new_n11122__ & ~new_new_n17250__;
  assign new_new_n17252__ = ys__n24626 & ~ys__n24675;
  assign new_new_n17253__ = ys__n24675 & ys__n24684;
  assign ys__n18669 = new_new_n17252__ | new_new_n17253__;
  assign new_new_n17255__ = new_new_n11122__ & ys__n18669;
  assign ys__n18670 = new_new_n17251__ | new_new_n17255__;
  assign new_new_n17257__ = ys__n18284 & ys__n18670;
  assign new_new_n17258__ = ~new_new_n17244__ & ~new_new_n17257__;
  assign new_new_n17259__ = ~ys__n18281 & ~new_new_n17258__;
  assign new_new_n17260__ = ys__n18571 & ~new_new_n11125__;
  assign new_new_n17261__ = ys__n18572 & new_new_n11125__;
  assign ys__n18573 = new_new_n17260__ | new_new_n17261__;
  assign new_new_n17263__ = ys__n18281 & ys__n18573;
  assign new_new_n17264__ = ~new_new_n17259__ & ~new_new_n17263__;
  assign new_new_n17265__ = ~ys__n18278 & ~new_new_n17264__;
  assign new_new_n17266__ = ys__n18839 & ys__n18278;
  assign ys__n18403 = new_new_n17265__ | new_new_n17266__;
  assign new_new_n17268__ = ys__n316 & ~ys__n18393;
  assign new_new_n17269__ = ys__n18393 & ys__n18403;
  assign ys__n18404 = new_new_n17268__ | new_new_n17269__;
  assign new_new_n17271__ = ys__n18962 & ys__n18287;
  assign new_new_n17272__ = ~ys__n18284 & new_new_n17271__;
  assign new_new_n17273__ = ys__n24627 & ~ys__n4764;
  assign new_new_n17274__ = ys__n24628 & ys__n4764;
  assign ys__n18776 = new_new_n17273__ | new_new_n17274__;
  assign new_new_n17276__ = ~ys__n18071 & ys__n18776;
  assign new_new_n17277__ = ys__n18071 & ys__n18777;
  assign new_new_n17278__ = ~new_new_n17276__ & ~new_new_n17277__;
  assign new_new_n17279__ = ~new_new_n11122__ & ~new_new_n17278__;
  assign new_new_n17280__ = ys__n24628 & ~ys__n24675;
  assign new_new_n17281__ = ys__n24675 & ys__n24685;
  assign ys__n18672 = new_new_n17280__ | new_new_n17281__;
  assign new_new_n17283__ = new_new_n11122__ & ys__n18672;
  assign ys__n18673 = new_new_n17279__ | new_new_n17283__;
  assign new_new_n17285__ = ys__n18284 & ys__n18673;
  assign new_new_n17286__ = ~new_new_n17272__ & ~new_new_n17285__;
  assign new_new_n17287__ = ~ys__n18281 & ~new_new_n17286__;
  assign new_new_n17288__ = ys__n18574 & ~new_new_n11125__;
  assign new_new_n17289__ = ys__n18575 & new_new_n11125__;
  assign ys__n18576 = new_new_n17288__ | new_new_n17289__;
  assign new_new_n17291__ = ys__n18281 & ys__n18576;
  assign new_new_n17292__ = ~new_new_n17287__ & ~new_new_n17291__;
  assign new_new_n17293__ = ~ys__n18278 & ~new_new_n17292__;
  assign new_new_n17294__ = ys__n18841 & ys__n18278;
  assign ys__n18405 = new_new_n17293__ | new_new_n17294__;
  assign new_new_n17296__ = ys__n6115 & ~ys__n18393;
  assign new_new_n17297__ = ys__n18393 & ys__n18405;
  assign ys__n18406 = new_new_n17296__ | new_new_n17297__;
  assign new_new_n17299__ = ys__n18963 & ys__n18287;
  assign new_new_n17300__ = ~ys__n18284 & new_new_n17299__;
  assign new_new_n17301__ = ys__n24629 & ~ys__n4764;
  assign new_new_n17302__ = ys__n24630 & ys__n4764;
  assign ys__n18778 = new_new_n17301__ | new_new_n17302__;
  assign new_new_n17304__ = ~ys__n18071 & ys__n18778;
  assign new_new_n17305__ = ys__n18071 & ys__n18779;
  assign new_new_n17306__ = ~new_new_n17304__ & ~new_new_n17305__;
  assign new_new_n17307__ = ~new_new_n11122__ & ~new_new_n17306__;
  assign new_new_n17308__ = ys__n24630 & ~ys__n24675;
  assign new_new_n17309__ = ys__n24675 & ys__n24686;
  assign ys__n18675 = new_new_n17308__ | new_new_n17309__;
  assign new_new_n17311__ = new_new_n11122__ & ys__n18675;
  assign ys__n18676 = new_new_n17307__ | new_new_n17311__;
  assign new_new_n17313__ = ys__n18284 & ys__n18676;
  assign new_new_n17314__ = ~new_new_n17300__ & ~new_new_n17313__;
  assign new_new_n17315__ = ~ys__n18281 & ~new_new_n17314__;
  assign new_new_n17316__ = ys__n18577 & ~new_new_n11125__;
  assign new_new_n17317__ = ys__n18578 & new_new_n11125__;
  assign ys__n18579 = new_new_n17316__ | new_new_n17317__;
  assign new_new_n17319__ = ys__n18281 & ys__n18579;
  assign new_new_n17320__ = ~new_new_n17315__ & ~new_new_n17319__;
  assign new_new_n17321__ = ~ys__n18278 & ~new_new_n17320__;
  assign new_new_n17322__ = ys__n18843 & ys__n18278;
  assign ys__n18407 = new_new_n17321__ | new_new_n17322__;
  assign new_new_n17324__ = ys__n44 & ~ys__n18393;
  assign new_new_n17325__ = ys__n18393 & ys__n18407;
  assign ys__n18408 = new_new_n17324__ | new_new_n17325__;
  assign new_new_n17327__ = ys__n18964 & ys__n18287;
  assign new_new_n17328__ = ~ys__n18284 & new_new_n17327__;
  assign new_new_n17329__ = ys__n24631 & ~ys__n4764;
  assign new_new_n17330__ = ys__n24632 & ys__n4764;
  assign ys__n18780 = new_new_n17329__ | new_new_n17330__;
  assign new_new_n17332__ = ~ys__n18071 & ys__n18780;
  assign new_new_n17333__ = ys__n18071 & ys__n18781;
  assign new_new_n17334__ = ~new_new_n17332__ & ~new_new_n17333__;
  assign new_new_n17335__ = ~new_new_n11122__ & ~new_new_n17334__;
  assign new_new_n17336__ = ys__n24632 & ~ys__n24675;
  assign new_new_n17337__ = ys__n24675 & ys__n24687;
  assign ys__n18678 = new_new_n17336__ | new_new_n17337__;
  assign new_new_n17339__ = new_new_n11122__ & ys__n18678;
  assign ys__n18679 = new_new_n17335__ | new_new_n17339__;
  assign new_new_n17341__ = ys__n18284 & ys__n18679;
  assign new_new_n17342__ = ~new_new_n17328__ & ~new_new_n17341__;
  assign new_new_n17343__ = ~ys__n18281 & ~new_new_n17342__;
  assign new_new_n17344__ = ys__n18580 & ~new_new_n11125__;
  assign new_new_n17345__ = ys__n18581 & new_new_n11125__;
  assign ys__n18582 = new_new_n17344__ | new_new_n17345__;
  assign new_new_n17347__ = ys__n18281 & ys__n18582;
  assign new_new_n17348__ = ~new_new_n17343__ & ~new_new_n17347__;
  assign new_new_n17349__ = ~ys__n18278 & ~new_new_n17348__;
  assign new_new_n17350__ = ys__n18845 & ys__n18278;
  assign ys__n18409 = new_new_n17349__ | new_new_n17350__;
  assign new_new_n17352__ = ys__n340 & ~ys__n18393;
  assign new_new_n17353__ = ys__n18393 & ys__n18409;
  assign ys__n18410 = new_new_n17352__ | new_new_n17353__;
  assign new_new_n17355__ = ys__n18965 & ys__n18287;
  assign new_new_n17356__ = ~ys__n18284 & new_new_n17355__;
  assign new_new_n17357__ = ys__n24633 & ~ys__n4764;
  assign new_new_n17358__ = ys__n24634 & ys__n4764;
  assign ys__n18782 = new_new_n17357__ | new_new_n17358__;
  assign new_new_n17360__ = ~ys__n18071 & ys__n18782;
  assign new_new_n17361__ = ys__n18071 & ys__n18783;
  assign new_new_n17362__ = ~new_new_n17360__ & ~new_new_n17361__;
  assign new_new_n17363__ = ~new_new_n11122__ & ~new_new_n17362__;
  assign new_new_n17364__ = ys__n24634 & ~ys__n24675;
  assign new_new_n17365__ = ys__n24675 & ys__n24688;
  assign ys__n18681 = new_new_n17364__ | new_new_n17365__;
  assign new_new_n17367__ = new_new_n11122__ & ys__n18681;
  assign ys__n18682 = new_new_n17363__ | new_new_n17367__;
  assign new_new_n17369__ = ys__n18284 & ys__n18682;
  assign new_new_n17370__ = ~new_new_n17356__ & ~new_new_n17369__;
  assign new_new_n17371__ = ~ys__n18281 & ~new_new_n17370__;
  assign new_new_n17372__ = ys__n18583 & ~new_new_n11125__;
  assign new_new_n17373__ = ys__n18584 & new_new_n11125__;
  assign ys__n18585 = new_new_n17372__ | new_new_n17373__;
  assign new_new_n17375__ = ys__n18281 & ys__n18585;
  assign new_new_n17376__ = ~new_new_n17371__ & ~new_new_n17375__;
  assign new_new_n17377__ = ~ys__n18278 & ~new_new_n17376__;
  assign new_new_n17378__ = ys__n18847 & ys__n18278;
  assign ys__n18411 = new_new_n17377__ | new_new_n17378__;
  assign new_new_n17380__ = ys__n46 & ~ys__n18393;
  assign new_new_n17381__ = ys__n18393 & ys__n18411;
  assign ys__n18412 = new_new_n17380__ | new_new_n17381__;
  assign new_new_n17383__ = ys__n18966 & ys__n18287;
  assign new_new_n17384__ = ~ys__n18284 & new_new_n17383__;
  assign new_new_n17385__ = ys__n24635 & ~ys__n4764;
  assign new_new_n17386__ = ys__n24636 & ys__n4764;
  assign ys__n18784 = new_new_n17385__ | new_new_n17386__;
  assign new_new_n17388__ = ~ys__n18071 & ys__n18784;
  assign new_new_n17389__ = ys__n18071 & ys__n18785;
  assign new_new_n17390__ = ~new_new_n17388__ & ~new_new_n17389__;
  assign new_new_n17391__ = ~new_new_n11122__ & ~new_new_n17390__;
  assign new_new_n17392__ = ys__n24636 & ~ys__n24675;
  assign new_new_n17393__ = ys__n24675 & ys__n24689;
  assign ys__n18684 = new_new_n17392__ | new_new_n17393__;
  assign new_new_n17395__ = new_new_n11122__ & ys__n18684;
  assign ys__n18685 = new_new_n17391__ | new_new_n17395__;
  assign new_new_n17397__ = ys__n18284 & ys__n18685;
  assign new_new_n17398__ = ~new_new_n17384__ & ~new_new_n17397__;
  assign new_new_n17399__ = ~ys__n18281 & ~new_new_n17398__;
  assign new_new_n17400__ = ys__n18586 & ~new_new_n11125__;
  assign new_new_n17401__ = ys__n18587 & new_new_n11125__;
  assign ys__n18588 = new_new_n17400__ | new_new_n17401__;
  assign new_new_n17403__ = ys__n18281 & ys__n18588;
  assign new_new_n17404__ = ~new_new_n17399__ & ~new_new_n17403__;
  assign new_new_n17405__ = ~ys__n18278 & ~new_new_n17404__;
  assign new_new_n17406__ = ys__n18849 & ys__n18278;
  assign ys__n18413 = new_new_n17405__ | new_new_n17406__;
  assign new_new_n17408__ = ys__n6118 & ~ys__n18393;
  assign new_new_n17409__ = ys__n18393 & ys__n18413;
  assign ys__n18414 = new_new_n17408__ | new_new_n17409__;
  assign new_new_n17411__ = ys__n18967 & ys__n18287;
  assign new_new_n17412__ = ~ys__n18284 & new_new_n17411__;
  assign new_new_n17413__ = ys__n24637 & ~ys__n4764;
  assign new_new_n17414__ = ys__n24638 & ys__n4764;
  assign ys__n18786 = new_new_n17413__ | new_new_n17414__;
  assign new_new_n17416__ = ~ys__n18071 & ys__n18786;
  assign new_new_n17417__ = ys__n18071 & ys__n18787;
  assign new_new_n17418__ = ~new_new_n17416__ & ~new_new_n17417__;
  assign new_new_n17419__ = ~new_new_n11122__ & ~new_new_n17418__;
  assign new_new_n17420__ = ys__n24638 & ~ys__n24675;
  assign new_new_n17421__ = ys__n24675 & ys__n24690;
  assign ys__n18687 = new_new_n17420__ | new_new_n17421__;
  assign new_new_n17423__ = new_new_n11122__ & ys__n18687;
  assign ys__n18688 = new_new_n17419__ | new_new_n17423__;
  assign new_new_n17425__ = ys__n18284 & ys__n18688;
  assign new_new_n17426__ = ~new_new_n17412__ & ~new_new_n17425__;
  assign new_new_n17427__ = ~ys__n18281 & ~new_new_n17426__;
  assign new_new_n17428__ = ys__n18589 & ~new_new_n11125__;
  assign new_new_n17429__ = ys__n18590 & new_new_n11125__;
  assign ys__n18591 = new_new_n17428__ | new_new_n17429__;
  assign new_new_n17431__ = ys__n18281 & ys__n18591;
  assign new_new_n17432__ = ~new_new_n17427__ & ~new_new_n17431__;
  assign new_new_n17433__ = ~ys__n18278 & ~new_new_n17432__;
  assign new_new_n17434__ = ys__n18851 & ys__n18278;
  assign ys__n18415 = new_new_n17433__ | new_new_n17434__;
  assign new_new_n17436__ = ys__n6119 & ~ys__n18393;
  assign new_new_n17437__ = ys__n18393 & ys__n18415;
  assign ys__n18416 = new_new_n17436__ | new_new_n17437__;
  assign new_new_n17439__ = ys__n18968 & ys__n18287;
  assign new_new_n17440__ = ~ys__n18284 & new_new_n17439__;
  assign new_new_n17441__ = ys__n24639 & ~ys__n4764;
  assign new_new_n17442__ = ys__n24640 & ys__n4764;
  assign ys__n18788 = new_new_n17441__ | new_new_n17442__;
  assign new_new_n17444__ = ~ys__n18071 & ys__n18788;
  assign new_new_n17445__ = ys__n18071 & ys__n18789;
  assign new_new_n17446__ = ~new_new_n17444__ & ~new_new_n17445__;
  assign new_new_n17447__ = ~new_new_n11122__ & ~new_new_n17446__;
  assign new_new_n17448__ = ys__n24640 & ~ys__n24675;
  assign new_new_n17449__ = ys__n24675 & ys__n24691;
  assign ys__n18690 = new_new_n17448__ | new_new_n17449__;
  assign new_new_n17451__ = new_new_n11122__ & ys__n18690;
  assign ys__n18691 = new_new_n17447__ | new_new_n17451__;
  assign new_new_n17453__ = ys__n18284 & ys__n18691;
  assign new_new_n17454__ = ~new_new_n17440__ & ~new_new_n17453__;
  assign new_new_n17455__ = ~ys__n18281 & ~new_new_n17454__;
  assign new_new_n17456__ = ys__n18592 & ~new_new_n11125__;
  assign new_new_n17457__ = ys__n18593 & new_new_n11125__;
  assign ys__n18594 = new_new_n17456__ | new_new_n17457__;
  assign new_new_n17459__ = ys__n18281 & ys__n18594;
  assign new_new_n17460__ = ~new_new_n17455__ & ~new_new_n17459__;
  assign new_new_n17461__ = ~ys__n18278 & ~new_new_n17460__;
  assign new_new_n17462__ = ys__n18853 & ys__n18278;
  assign ys__n18417 = new_new_n17461__ | new_new_n17462__;
  assign new_new_n17464__ = ys__n6120 & ~ys__n18393;
  assign new_new_n17465__ = ys__n18393 & ys__n18417;
  assign ys__n18418 = new_new_n17464__ | new_new_n17465__;
  assign new_new_n17467__ = ys__n18969 & ys__n18287;
  assign new_new_n17468__ = ~ys__n18284 & new_new_n17467__;
  assign new_new_n17469__ = ys__n24641 & ~ys__n4764;
  assign new_new_n17470__ = ys__n24642 & ys__n4764;
  assign ys__n18790 = new_new_n17469__ | new_new_n17470__;
  assign new_new_n17472__ = ~ys__n18071 & ys__n18790;
  assign new_new_n17473__ = ys__n18071 & ys__n18791;
  assign new_new_n17474__ = ~new_new_n17472__ & ~new_new_n17473__;
  assign new_new_n17475__ = ~new_new_n11122__ & ~new_new_n17474__;
  assign new_new_n17476__ = ys__n24642 & ~ys__n24675;
  assign new_new_n17477__ = ys__n24675 & ys__n24692;
  assign ys__n18693 = new_new_n17476__ | new_new_n17477__;
  assign new_new_n17479__ = new_new_n11122__ & ys__n18693;
  assign ys__n18694 = new_new_n17475__ | new_new_n17479__;
  assign new_new_n17481__ = ys__n18284 & ys__n18694;
  assign new_new_n17482__ = ~new_new_n17468__ & ~new_new_n17481__;
  assign new_new_n17483__ = ~ys__n18281 & ~new_new_n17482__;
  assign new_new_n17484__ = ys__n18595 & ~new_new_n11125__;
  assign new_new_n17485__ = ys__n18596 & new_new_n11125__;
  assign ys__n18597 = new_new_n17484__ | new_new_n17485__;
  assign new_new_n17487__ = ys__n18281 & ys__n18597;
  assign new_new_n17488__ = ~new_new_n17483__ & ~new_new_n17487__;
  assign new_new_n17489__ = ~ys__n18278 & ~new_new_n17488__;
  assign new_new_n17490__ = ys__n18855 & ys__n18278;
  assign ys__n18419 = new_new_n17489__ | new_new_n17490__;
  assign new_new_n17492__ = ys__n6121 & ~ys__n18393;
  assign new_new_n17493__ = ys__n18393 & ys__n18419;
  assign ys__n18420 = new_new_n17492__ | new_new_n17493__;
  assign new_new_n17495__ = ys__n18970 & ys__n18287;
  assign new_new_n17496__ = ~ys__n18284 & new_new_n17495__;
  assign new_new_n17497__ = ys__n24643 & ~ys__n4764;
  assign new_new_n17498__ = ys__n24644 & ys__n4764;
  assign ys__n18792 = new_new_n17497__ | new_new_n17498__;
  assign new_new_n17500__ = ~ys__n18071 & ys__n18792;
  assign new_new_n17501__ = ys__n18071 & ys__n18793;
  assign new_new_n17502__ = ~new_new_n17500__ & ~new_new_n17501__;
  assign new_new_n17503__ = ~new_new_n11122__ & ~new_new_n17502__;
  assign new_new_n17504__ = ys__n24644 & ~ys__n24675;
  assign new_new_n17505__ = ys__n24675 & ys__n24693;
  assign ys__n18696 = new_new_n17504__ | new_new_n17505__;
  assign new_new_n17507__ = new_new_n11122__ & ys__n18696;
  assign ys__n18697 = new_new_n17503__ | new_new_n17507__;
  assign new_new_n17509__ = ys__n18284 & ys__n18697;
  assign new_new_n17510__ = ~new_new_n17496__ & ~new_new_n17509__;
  assign new_new_n17511__ = ~ys__n18281 & ~new_new_n17510__;
  assign new_new_n17512__ = ys__n18598 & ~new_new_n11125__;
  assign new_new_n17513__ = ys__n18599 & new_new_n11125__;
  assign ys__n18600 = new_new_n17512__ | new_new_n17513__;
  assign new_new_n17515__ = ys__n18281 & ys__n18600;
  assign new_new_n17516__ = ~new_new_n17511__ & ~new_new_n17515__;
  assign new_new_n17517__ = ~ys__n18278 & ~new_new_n17516__;
  assign new_new_n17518__ = ys__n18857 & ys__n18278;
  assign ys__n18421 = new_new_n17517__ | new_new_n17518__;
  assign new_new_n17520__ = ys__n6123 & ~ys__n18393;
  assign new_new_n17521__ = ys__n18393 & ys__n18421;
  assign ys__n18422 = new_new_n17520__ | new_new_n17521__;
  assign new_new_n17523__ = ys__n18971 & ys__n18287;
  assign new_new_n17524__ = ~ys__n18284 & new_new_n17523__;
  assign new_new_n17525__ = ys__n24645 & ~ys__n4764;
  assign new_new_n17526__ = ys__n24646 & ys__n4764;
  assign ys__n18794 = new_new_n17525__ | new_new_n17526__;
  assign new_new_n17528__ = ~ys__n18071 & ys__n18794;
  assign new_new_n17529__ = ys__n18071 & ys__n18795;
  assign new_new_n17530__ = ~new_new_n17528__ & ~new_new_n17529__;
  assign new_new_n17531__ = ~new_new_n11122__ & ~new_new_n17530__;
  assign new_new_n17532__ = ys__n24646 & ~ys__n24675;
  assign new_new_n17533__ = ys__n24675 & ys__n24694;
  assign ys__n18699 = new_new_n17532__ | new_new_n17533__;
  assign new_new_n17535__ = new_new_n11122__ & ys__n18699;
  assign ys__n18700 = new_new_n17531__ | new_new_n17535__;
  assign new_new_n17537__ = ys__n18284 & ys__n18700;
  assign new_new_n17538__ = ~new_new_n17524__ & ~new_new_n17537__;
  assign new_new_n17539__ = ~ys__n18281 & ~new_new_n17538__;
  assign new_new_n17540__ = ys__n18601 & ~new_new_n11125__;
  assign new_new_n17541__ = ys__n18602 & new_new_n11125__;
  assign ys__n18603 = new_new_n17540__ | new_new_n17541__;
  assign new_new_n17543__ = ys__n18281 & ys__n18603;
  assign new_new_n17544__ = ~new_new_n17539__ & ~new_new_n17543__;
  assign new_new_n17545__ = ~ys__n18278 & ~new_new_n17544__;
  assign new_new_n17546__ = ys__n18859 & ys__n18278;
  assign ys__n18423 = new_new_n17545__ | new_new_n17546__;
  assign new_new_n17548__ = ys__n6124 & ~ys__n18393;
  assign new_new_n17549__ = ys__n18393 & ys__n18423;
  assign ys__n18424 = new_new_n17548__ | new_new_n17549__;
  assign new_new_n17551__ = ys__n18972 & ys__n18287;
  assign new_new_n17552__ = ~ys__n18284 & new_new_n17551__;
  assign new_new_n17553__ = ys__n24647 & ~ys__n4764;
  assign new_new_n17554__ = ys__n24648 & ys__n4764;
  assign ys__n18796 = new_new_n17553__ | new_new_n17554__;
  assign new_new_n17556__ = ~ys__n18071 & ys__n18796;
  assign new_new_n17557__ = ys__n18071 & ys__n18797;
  assign new_new_n17558__ = ~new_new_n17556__ & ~new_new_n17557__;
  assign new_new_n17559__ = ~new_new_n11122__ & ~new_new_n17558__;
  assign new_new_n17560__ = ys__n24648 & ~ys__n24675;
  assign new_new_n17561__ = ys__n24675 & ys__n24695;
  assign ys__n18702 = new_new_n17560__ | new_new_n17561__;
  assign new_new_n17563__ = new_new_n11122__ & ys__n18702;
  assign ys__n18703 = new_new_n17559__ | new_new_n17563__;
  assign new_new_n17565__ = ys__n18284 & ys__n18703;
  assign new_new_n17566__ = ~new_new_n17552__ & ~new_new_n17565__;
  assign new_new_n17567__ = ~ys__n18281 & ~new_new_n17566__;
  assign new_new_n17568__ = ys__n18604 & ~new_new_n11125__;
  assign new_new_n17569__ = ys__n18605 & new_new_n11125__;
  assign ys__n18606 = new_new_n17568__ | new_new_n17569__;
  assign new_new_n17571__ = ys__n18281 & ys__n18606;
  assign new_new_n17572__ = ~new_new_n17567__ & ~new_new_n17571__;
  assign new_new_n17573__ = ~ys__n18278 & ~new_new_n17572__;
  assign new_new_n17574__ = ys__n18861 & ys__n18278;
  assign ys__n18425 = new_new_n17573__ | new_new_n17574__;
  assign new_new_n17576__ = ys__n6126 & ~ys__n18393;
  assign new_new_n17577__ = ys__n18393 & ys__n18425;
  assign ys__n18426 = new_new_n17576__ | new_new_n17577__;
  assign new_new_n17579__ = ys__n18973 & ys__n18287;
  assign new_new_n17580__ = ~ys__n18284 & new_new_n17579__;
  assign new_new_n17581__ = ys__n24649 & ~ys__n4764;
  assign new_new_n17582__ = ys__n24650 & ys__n4764;
  assign ys__n18798 = new_new_n17581__ | new_new_n17582__;
  assign new_new_n17584__ = ~ys__n18071 & ys__n18798;
  assign new_new_n17585__ = ys__n18071 & ys__n18799;
  assign new_new_n17586__ = ~new_new_n17584__ & ~new_new_n17585__;
  assign new_new_n17587__ = ~new_new_n11122__ & ~new_new_n17586__;
  assign new_new_n17588__ = ys__n24650 & ~ys__n24675;
  assign new_new_n17589__ = ys__n24675 & ys__n24696;
  assign ys__n18705 = new_new_n17588__ | new_new_n17589__;
  assign new_new_n17591__ = new_new_n11122__ & ys__n18705;
  assign ys__n18706 = new_new_n17587__ | new_new_n17591__;
  assign new_new_n17593__ = ys__n18284 & ys__n18706;
  assign new_new_n17594__ = ~new_new_n17580__ & ~new_new_n17593__;
  assign new_new_n17595__ = ~ys__n18281 & ~new_new_n17594__;
  assign new_new_n17596__ = ys__n18607 & ~new_new_n11125__;
  assign new_new_n17597__ = ys__n18608 & new_new_n11125__;
  assign ys__n18609 = new_new_n17596__ | new_new_n17597__;
  assign new_new_n17599__ = ys__n18281 & ys__n18609;
  assign new_new_n17600__ = ~new_new_n17595__ & ~new_new_n17599__;
  assign new_new_n17601__ = ~ys__n18278 & ~new_new_n17600__;
  assign new_new_n17602__ = ys__n18863 & ys__n18278;
  assign ys__n18427 = new_new_n17601__ | new_new_n17602__;
  assign new_new_n17604__ = ys__n6127 & ~ys__n18393;
  assign new_new_n17605__ = ys__n18393 & ys__n18427;
  assign ys__n18428 = new_new_n17604__ | new_new_n17605__;
  assign new_new_n17607__ = ys__n18974 & ys__n18287;
  assign new_new_n17608__ = ~ys__n18284 & new_new_n17607__;
  assign new_new_n17609__ = ys__n24651 & ~ys__n4764;
  assign new_new_n17610__ = ys__n24652 & ys__n4764;
  assign ys__n18800 = new_new_n17609__ | new_new_n17610__;
  assign new_new_n17612__ = ~ys__n18071 & ys__n18800;
  assign new_new_n17613__ = ys__n18071 & ys__n18801;
  assign new_new_n17614__ = ~new_new_n17612__ & ~new_new_n17613__;
  assign new_new_n17615__ = ~new_new_n11122__ & ~new_new_n17614__;
  assign new_new_n17616__ = ys__n24652 & ~ys__n24675;
  assign new_new_n17617__ = ys__n24675 & ys__n24697;
  assign ys__n18708 = new_new_n17616__ | new_new_n17617__;
  assign new_new_n17619__ = new_new_n11122__ & ys__n18708;
  assign ys__n18709 = new_new_n17615__ | new_new_n17619__;
  assign new_new_n17621__ = ys__n18284 & ys__n18709;
  assign new_new_n17622__ = ~new_new_n17608__ & ~new_new_n17621__;
  assign new_new_n17623__ = ~ys__n18281 & ~new_new_n17622__;
  assign new_new_n17624__ = ys__n18610 & ~new_new_n11125__;
  assign new_new_n17625__ = ys__n18611 & new_new_n11125__;
  assign ys__n18612 = new_new_n17624__ | new_new_n17625__;
  assign new_new_n17627__ = ys__n18281 & ys__n18612;
  assign new_new_n17628__ = ~new_new_n17623__ & ~new_new_n17627__;
  assign new_new_n17629__ = ~ys__n18278 & ~new_new_n17628__;
  assign new_new_n17630__ = ys__n18865 & ys__n18278;
  assign ys__n18429 = new_new_n17629__ | new_new_n17630__;
  assign new_new_n17632__ = ys__n6129 & ~ys__n18393;
  assign new_new_n17633__ = ys__n18393 & ys__n18429;
  assign ys__n18430 = new_new_n17632__ | new_new_n17633__;
  assign new_new_n17635__ = ys__n18975 & ys__n18287;
  assign new_new_n17636__ = ~ys__n18284 & new_new_n17635__;
  assign new_new_n17637__ = ys__n24653 & ~ys__n4764;
  assign new_new_n17638__ = ys__n24654 & ys__n4764;
  assign ys__n18802 = new_new_n17637__ | new_new_n17638__;
  assign new_new_n17640__ = ~ys__n18071 & ys__n18802;
  assign new_new_n17641__ = ys__n18071 & ys__n18803;
  assign new_new_n17642__ = ~new_new_n17640__ & ~new_new_n17641__;
  assign new_new_n17643__ = ~new_new_n11122__ & ~new_new_n17642__;
  assign new_new_n17644__ = ys__n24654 & ~ys__n24675;
  assign new_new_n17645__ = ys__n24675 & ys__n24698;
  assign ys__n18711 = new_new_n17644__ | new_new_n17645__;
  assign new_new_n17647__ = new_new_n11122__ & ys__n18711;
  assign ys__n18712 = new_new_n17643__ | new_new_n17647__;
  assign new_new_n17649__ = ys__n18284 & ys__n18712;
  assign new_new_n17650__ = ~new_new_n17636__ & ~new_new_n17649__;
  assign new_new_n17651__ = ~ys__n18281 & ~new_new_n17650__;
  assign new_new_n17652__ = ys__n18613 & ~new_new_n11125__;
  assign new_new_n17653__ = ys__n18614 & new_new_n11125__;
  assign ys__n18615 = new_new_n17652__ | new_new_n17653__;
  assign new_new_n17655__ = ys__n18281 & ys__n18615;
  assign new_new_n17656__ = ~new_new_n17651__ & ~new_new_n17655__;
  assign new_new_n17657__ = ~ys__n18278 & ~new_new_n17656__;
  assign new_new_n17658__ = ys__n18867 & ys__n18278;
  assign ys__n18431 = new_new_n17657__ | new_new_n17658__;
  assign new_new_n17660__ = ys__n6130 & ~ys__n18393;
  assign new_new_n17661__ = ys__n18393 & ys__n18431;
  assign ys__n18432 = new_new_n17660__ | new_new_n17661__;
  assign new_new_n17663__ = ys__n18976 & ys__n18287;
  assign new_new_n17664__ = ~ys__n18284 & new_new_n17663__;
  assign new_new_n17665__ = ys__n24655 & ~ys__n4764;
  assign new_new_n17666__ = ys__n24656 & ys__n4764;
  assign ys__n18804 = new_new_n17665__ | new_new_n17666__;
  assign new_new_n17668__ = ~ys__n18071 & ys__n18804;
  assign new_new_n17669__ = ys__n18071 & ys__n18805;
  assign new_new_n17670__ = ~new_new_n17668__ & ~new_new_n17669__;
  assign new_new_n17671__ = ~new_new_n11122__ & ~new_new_n17670__;
  assign new_new_n17672__ = ys__n24656 & ~ys__n24675;
  assign new_new_n17673__ = ys__n24675 & ys__n24699;
  assign ys__n18714 = new_new_n17672__ | new_new_n17673__;
  assign new_new_n17675__ = new_new_n11122__ & ys__n18714;
  assign ys__n18715 = new_new_n17671__ | new_new_n17675__;
  assign new_new_n17677__ = ys__n18284 & ys__n18715;
  assign new_new_n17678__ = ~new_new_n17664__ & ~new_new_n17677__;
  assign new_new_n17679__ = ~ys__n18281 & ~new_new_n17678__;
  assign new_new_n17680__ = ys__n18616 & ~new_new_n11125__;
  assign new_new_n17681__ = ys__n18617 & new_new_n11125__;
  assign ys__n18618 = new_new_n17680__ | new_new_n17681__;
  assign new_new_n17683__ = ys__n18281 & ys__n18618;
  assign new_new_n17684__ = ~new_new_n17679__ & ~new_new_n17683__;
  assign new_new_n17685__ = ~ys__n18278 & ~new_new_n17684__;
  assign new_new_n17686__ = ys__n18869 & ys__n18278;
  assign ys__n18433 = new_new_n17685__ | new_new_n17686__;
  assign new_new_n17688__ = ys__n42 & ~ys__n18393;
  assign new_new_n17689__ = ys__n18393 & ys__n18433;
  assign ys__n18434 = new_new_n17688__ | new_new_n17689__;
  assign new_new_n17691__ = ys__n40 & ~ys__n18393;
  assign new_new_n17692__ = ys__n18393 & ys__n806;
  assign ys__n18435 = new_new_n17691__ | new_new_n17692__;
  assign new_new_n17694__ = ys__n6133 & ~ys__n18393;
  assign new_new_n17695__ = ys__n18393 & ys__n3250;
  assign ys__n18436 = new_new_n17694__ | new_new_n17695__;
  assign new_new_n17697__ = ys__n6134 & ~ys__n18393;
  assign new_new_n17698__ = ys__n18393 & ys__n3252;
  assign ys__n18437 = new_new_n17697__ | new_new_n17698__;
  assign new_new_n17700__ = ys__n38 & ~ys__n18393;
  assign new_new_n17701__ = ys__n18393 & ys__n804;
  assign ys__n18438 = new_new_n17700__ | new_new_n17701__;
  assign new_new_n17703__ = ys__n36 & ~ys__n18393;
  assign new_new_n17704__ = ys__n18393 & ys__n802;
  assign ys__n18439 = new_new_n17703__ | new_new_n17704__;
  assign new_new_n17706__ = ys__n34 & ~ys__n18393;
  assign new_new_n17707__ = ys__n18393 & ys__n800;
  assign ys__n18440 = new_new_n17706__ | new_new_n17707__;
  assign new_new_n17709__ = ys__n32 & ~ys__n18393;
  assign new_new_n17710__ = ys__n18393 & ys__n798;
  assign ys__n18441 = new_new_n17709__ | new_new_n17710__;
  assign new_new_n17712__ = ys__n30 & ~ys__n18393;
  assign new_new_n17713__ = ys__n18393 & ys__n796;
  assign ys__n18442 = new_new_n17712__ | new_new_n17713__;
  assign new_new_n17715__ = ys__n28 & ~ys__n18393;
  assign new_new_n17716__ = ys__n18393 & ys__n810;
  assign ys__n18443 = new_new_n17715__ | new_new_n17716__;
  assign new_new_n17718__ = ys__n26 & ~ys__n18393;
  assign new_new_n17719__ = ys__n18393 & ys__n808;
  assign ys__n18444 = new_new_n17718__ | new_new_n17719__;
  assign new_new_n17721__ = ys__n24 & ~ys__n18393;
  assign new_new_n17722__ = ys__n18393 & ys__n812;
  assign ys__n18445 = new_new_n17721__ | new_new_n17722__;
  assign new_new_n17724__ = ys__n19116 & ~ys__n18281;
  assign new_new_n17725__ = ~ys__n18278 & new_new_n17724__;
  assign new_new_n17726__ = ys__n18287 & new_new_n17725__;
  assign new_new_n17727__ = ~ys__n18284 & new_new_n17726__;
  assign new_new_n17728__ = ys__n18989 & ys__n18278;
  assign ys__n18449 = new_new_n17727__ | new_new_n17728__;
  assign new_new_n17730__ = ~ys__n18393 & ys__n18448;
  assign new_new_n17731__ = ys__n18393 & ys__n18449;
  assign ys__n18450 = new_new_n17730__ | new_new_n17731__;
  assign new_new_n17733__ = ys__n19117 & ~ys__n18281;
  assign new_new_n17734__ = ~ys__n18278 & new_new_n17733__;
  assign new_new_n17735__ = ys__n18287 & new_new_n17734__;
  assign new_new_n17736__ = ~ys__n18284 & new_new_n17735__;
  assign new_new_n17737__ = ys__n18991 & ys__n18278;
  assign ys__n18452 = new_new_n17736__ | new_new_n17737__;
  assign new_new_n17739__ = ~ys__n18393 & ys__n18451;
  assign new_new_n17740__ = ys__n18393 & ys__n18452;
  assign ys__n18453 = new_new_n17739__ | new_new_n17740__;
  assign new_new_n17742__ = ys__n19118 & ~ys__n18281;
  assign new_new_n17743__ = ~ys__n18278 & new_new_n17742__;
  assign new_new_n17744__ = ys__n18287 & new_new_n17743__;
  assign new_new_n17745__ = ~ys__n18284 & new_new_n17744__;
  assign new_new_n17746__ = ys__n18993 & ys__n18278;
  assign ys__n18455 = new_new_n17745__ | new_new_n17746__;
  assign new_new_n17748__ = ~ys__n18393 & ys__n18454;
  assign new_new_n17749__ = ys__n18393 & ys__n18455;
  assign ys__n18456 = new_new_n17748__ | new_new_n17749__;
  assign new_new_n17751__ = ys__n19119 & ~ys__n18281;
  assign new_new_n17752__ = ~ys__n18278 & new_new_n17751__;
  assign new_new_n17753__ = ys__n18287 & new_new_n17752__;
  assign new_new_n17754__ = ~ys__n18284 & new_new_n17753__;
  assign new_new_n17755__ = ys__n18995 & ys__n18278;
  assign ys__n18458 = new_new_n17754__ | new_new_n17755__;
  assign new_new_n17757__ = ~ys__n18393 & ys__n18457;
  assign new_new_n17758__ = ys__n18393 & ys__n18458;
  assign ys__n18459 = new_new_n17757__ | new_new_n17758__;
  assign new_new_n17760__ = ys__n19120 & ~ys__n18281;
  assign new_new_n17761__ = ~ys__n18278 & new_new_n17760__;
  assign new_new_n17762__ = ys__n18287 & new_new_n17761__;
  assign new_new_n17763__ = ~ys__n18284 & new_new_n17762__;
  assign new_new_n17764__ = ys__n18997 & ys__n18278;
  assign ys__n18461 = new_new_n17763__ | new_new_n17764__;
  assign new_new_n17766__ = ~ys__n18393 & ys__n18460;
  assign new_new_n17767__ = ys__n18393 & ys__n18461;
  assign ys__n18462 = new_new_n17766__ | new_new_n17767__;
  assign new_new_n17769__ = ys__n19121 & ~ys__n18281;
  assign new_new_n17770__ = ~ys__n18278 & new_new_n17769__;
  assign new_new_n17771__ = ys__n18287 & new_new_n17770__;
  assign new_new_n17772__ = ~ys__n18284 & new_new_n17771__;
  assign new_new_n17773__ = ys__n18999 & ys__n18278;
  assign ys__n18464 = new_new_n17772__ | new_new_n17773__;
  assign new_new_n17775__ = ~ys__n18393 & ys__n18463;
  assign new_new_n17776__ = ys__n18393 & ys__n18464;
  assign ys__n18465 = new_new_n17775__ | new_new_n17776__;
  assign new_new_n17778__ = ys__n19122 & ~ys__n18281;
  assign new_new_n17779__ = ~ys__n18278 & new_new_n17778__;
  assign new_new_n17780__ = ys__n18287 & new_new_n17779__;
  assign new_new_n17781__ = ~ys__n18284 & new_new_n17780__;
  assign new_new_n17782__ = ys__n19001 & ys__n18278;
  assign ys__n18467 = new_new_n17781__ | new_new_n17782__;
  assign new_new_n17784__ = ~ys__n18393 & ys__n18466;
  assign new_new_n17785__ = ys__n18393 & ys__n18467;
  assign ys__n18468 = new_new_n17784__ | new_new_n17785__;
  assign new_new_n17787__ = ys__n19123 & ~ys__n18281;
  assign new_new_n17788__ = ~ys__n18278 & new_new_n17787__;
  assign new_new_n17789__ = ys__n18287 & new_new_n17788__;
  assign new_new_n17790__ = ~ys__n18284 & new_new_n17789__;
  assign new_new_n17791__ = ys__n19003 & ys__n18278;
  assign ys__n18470 = new_new_n17790__ | new_new_n17791__;
  assign new_new_n17793__ = ~ys__n18393 & ys__n18469;
  assign new_new_n17794__ = ys__n18393 & ys__n18470;
  assign ys__n18471 = new_new_n17793__ | new_new_n17794__;
  assign new_new_n17796__ = ys__n19124 & ~ys__n18281;
  assign new_new_n17797__ = ~ys__n18278 & new_new_n17796__;
  assign new_new_n17798__ = ys__n18287 & new_new_n17797__;
  assign new_new_n17799__ = ~ys__n18284 & new_new_n17798__;
  assign new_new_n17800__ = ys__n19005 & ys__n18278;
  assign ys__n18473 = new_new_n17799__ | new_new_n17800__;
  assign new_new_n17802__ = ~ys__n18393 & ys__n18472;
  assign new_new_n17803__ = ys__n18393 & ys__n18473;
  assign ys__n18474 = new_new_n17802__ | new_new_n17803__;
  assign new_new_n17805__ = ys__n19125 & ~ys__n18281;
  assign new_new_n17806__ = ~ys__n18278 & new_new_n17805__;
  assign new_new_n17807__ = ys__n18287 & new_new_n17806__;
  assign new_new_n17808__ = ~ys__n18284 & new_new_n17807__;
  assign new_new_n17809__ = ys__n19007 & ys__n18278;
  assign ys__n18476 = new_new_n17808__ | new_new_n17809__;
  assign new_new_n17811__ = ~ys__n18393 & ys__n18475;
  assign new_new_n17812__ = ys__n18393 & ys__n18476;
  assign ys__n18477 = new_new_n17811__ | new_new_n17812__;
  assign new_new_n17814__ = ys__n19126 & ~ys__n18281;
  assign new_new_n17815__ = ~ys__n18278 & new_new_n17814__;
  assign new_new_n17816__ = ys__n18287 & new_new_n17815__;
  assign new_new_n17817__ = ~ys__n18284 & new_new_n17816__;
  assign new_new_n17818__ = ys__n19009 & ys__n18278;
  assign ys__n18479 = new_new_n17817__ | new_new_n17818__;
  assign new_new_n17820__ = ~ys__n18393 & ys__n18478;
  assign new_new_n17821__ = ys__n18393 & ys__n18479;
  assign ys__n18480 = new_new_n17820__ | new_new_n17821__;
  assign new_new_n17823__ = ys__n19127 & ~ys__n18281;
  assign new_new_n17824__ = ~ys__n18278 & new_new_n17823__;
  assign new_new_n17825__ = ys__n18287 & new_new_n17824__;
  assign new_new_n17826__ = ~ys__n18284 & new_new_n17825__;
  assign new_new_n17827__ = ys__n19011 & ys__n18278;
  assign ys__n18482 = new_new_n17826__ | new_new_n17827__;
  assign new_new_n17829__ = ~ys__n18393 & ys__n18481;
  assign new_new_n17830__ = ys__n18393 & ys__n18482;
  assign ys__n18483 = new_new_n17829__ | new_new_n17830__;
  assign new_new_n17832__ = ys__n19128 & ~ys__n18281;
  assign new_new_n17833__ = ~ys__n18278 & new_new_n17832__;
  assign new_new_n17834__ = ys__n18287 & new_new_n17833__;
  assign new_new_n17835__ = ~ys__n18284 & new_new_n17834__;
  assign new_new_n17836__ = ys__n19013 & ys__n18278;
  assign ys__n18485 = new_new_n17835__ | new_new_n17836__;
  assign new_new_n17838__ = ~ys__n18393 & ys__n18484;
  assign new_new_n17839__ = ys__n18393 & ys__n18485;
  assign ys__n18486 = new_new_n17838__ | new_new_n17839__;
  assign new_new_n17841__ = ys__n19129 & ~ys__n18281;
  assign new_new_n17842__ = ~ys__n18278 & new_new_n17841__;
  assign new_new_n17843__ = ys__n18287 & new_new_n17842__;
  assign new_new_n17844__ = ~ys__n18284 & new_new_n17843__;
  assign new_new_n17845__ = ys__n19015 & ys__n18278;
  assign ys__n18488 = new_new_n17844__ | new_new_n17845__;
  assign new_new_n17847__ = ~ys__n18393 & ys__n18487;
  assign new_new_n17848__ = ys__n18393 & ys__n18488;
  assign ys__n18489 = new_new_n17847__ | new_new_n17848__;
  assign new_new_n17850__ = ys__n19130 & ~ys__n18281;
  assign new_new_n17851__ = ~ys__n18278 & new_new_n17850__;
  assign new_new_n17852__ = ys__n18287 & new_new_n17851__;
  assign new_new_n17853__ = ~ys__n18284 & new_new_n17852__;
  assign new_new_n17854__ = ys__n19017 & ys__n18278;
  assign ys__n18491 = new_new_n17853__ | new_new_n17854__;
  assign new_new_n17856__ = ~ys__n18393 & ys__n18490;
  assign new_new_n17857__ = ys__n18393 & ys__n18491;
  assign ys__n18492 = new_new_n17856__ | new_new_n17857__;
  assign new_new_n17859__ = ys__n19131 & ~ys__n18281;
  assign new_new_n17860__ = ~ys__n18278 & new_new_n17859__;
  assign new_new_n17861__ = ys__n18287 & new_new_n17860__;
  assign new_new_n17862__ = ~ys__n18284 & new_new_n17861__;
  assign new_new_n17863__ = ys__n19019 & ys__n18278;
  assign ys__n18494 = new_new_n17862__ | new_new_n17863__;
  assign new_new_n17865__ = ~ys__n18393 & ys__n18493;
  assign new_new_n17866__ = ys__n18393 & ys__n18494;
  assign ys__n18495 = new_new_n17865__ | new_new_n17866__;
  assign new_new_n17868__ = ys__n19132 & ~ys__n18281;
  assign new_new_n17869__ = ~ys__n18278 & new_new_n17868__;
  assign new_new_n17870__ = ys__n18287 & new_new_n17869__;
  assign new_new_n17871__ = ~ys__n18284 & new_new_n17870__;
  assign new_new_n17872__ = ys__n19021 & ys__n18278;
  assign ys__n18497 = new_new_n17871__ | new_new_n17872__;
  assign new_new_n17874__ = ~ys__n18393 & ys__n18496;
  assign new_new_n17875__ = ys__n18393 & ys__n18497;
  assign ys__n18498 = new_new_n17874__ | new_new_n17875__;
  assign new_new_n17877__ = ys__n19133 & ~ys__n18281;
  assign new_new_n17878__ = ~ys__n18278 & new_new_n17877__;
  assign new_new_n17879__ = ys__n18287 & new_new_n17878__;
  assign new_new_n17880__ = ~ys__n18284 & new_new_n17879__;
  assign new_new_n17881__ = ys__n19023 & ys__n18278;
  assign ys__n18500 = new_new_n17880__ | new_new_n17881__;
  assign new_new_n17883__ = ~ys__n18393 & ys__n18499;
  assign new_new_n17884__ = ys__n18393 & ys__n18500;
  assign ys__n18501 = new_new_n17883__ | new_new_n17884__;
  assign new_new_n17886__ = ys__n19134 & ~ys__n18281;
  assign new_new_n17887__ = ~ys__n18278 & new_new_n17886__;
  assign new_new_n17888__ = ys__n18287 & new_new_n17887__;
  assign new_new_n17889__ = ~ys__n18284 & new_new_n17888__;
  assign new_new_n17890__ = ys__n19025 & ys__n18278;
  assign ys__n18503 = new_new_n17889__ | new_new_n17890__;
  assign new_new_n17892__ = ~ys__n18393 & ys__n18502;
  assign new_new_n17893__ = ys__n18393 & ys__n18503;
  assign ys__n18504 = new_new_n17892__ | new_new_n17893__;
  assign new_new_n17895__ = ys__n19135 & ~ys__n18281;
  assign new_new_n17896__ = ~ys__n18278 & new_new_n17895__;
  assign new_new_n17897__ = ys__n18287 & new_new_n17896__;
  assign new_new_n17898__ = ~ys__n18284 & new_new_n17897__;
  assign new_new_n17899__ = ys__n19027 & ys__n18278;
  assign ys__n18506 = new_new_n17898__ | new_new_n17899__;
  assign new_new_n17901__ = ~ys__n18393 & ys__n18505;
  assign new_new_n17902__ = ys__n18393 & ys__n18506;
  assign ys__n18507 = new_new_n17901__ | new_new_n17902__;
  assign new_new_n17904__ = ys__n19136 & ~ys__n18281;
  assign new_new_n17905__ = ~ys__n18278 & new_new_n17904__;
  assign new_new_n17906__ = ys__n18287 & new_new_n17905__;
  assign new_new_n17907__ = ~ys__n18284 & new_new_n17906__;
  assign new_new_n17908__ = ys__n19029 & ys__n18278;
  assign ys__n18509 = new_new_n17907__ | new_new_n17908__;
  assign new_new_n17910__ = ~ys__n18393 & ys__n18508;
  assign new_new_n17911__ = ys__n18393 & ys__n18509;
  assign ys__n18510 = new_new_n17910__ | new_new_n17911__;
  assign new_new_n17913__ = ys__n19137 & ~ys__n18281;
  assign new_new_n17914__ = ~ys__n18278 & new_new_n17913__;
  assign new_new_n17915__ = ys__n18287 & new_new_n17914__;
  assign new_new_n17916__ = ~ys__n18284 & new_new_n17915__;
  assign new_new_n17917__ = ys__n19031 & ys__n18278;
  assign ys__n18512 = new_new_n17916__ | new_new_n17917__;
  assign new_new_n17919__ = ~ys__n18393 & ys__n18511;
  assign new_new_n17920__ = ys__n18393 & ys__n18512;
  assign ys__n18513 = new_new_n17919__ | new_new_n17920__;
  assign new_new_n17922__ = ys__n19138 & ~ys__n18281;
  assign new_new_n17923__ = ~ys__n18278 & new_new_n17922__;
  assign new_new_n17924__ = ys__n18287 & new_new_n17923__;
  assign new_new_n17925__ = ~ys__n18284 & new_new_n17924__;
  assign new_new_n17926__ = ys__n19033 & ys__n18278;
  assign ys__n18515 = new_new_n17925__ | new_new_n17926__;
  assign new_new_n17928__ = ~ys__n18393 & ys__n18514;
  assign new_new_n17929__ = ys__n18393 & ys__n18515;
  assign ys__n18516 = new_new_n17928__ | new_new_n17929__;
  assign new_new_n17931__ = ys__n19139 & ~ys__n18281;
  assign new_new_n17932__ = ~ys__n18278 & new_new_n17931__;
  assign new_new_n17933__ = ys__n18287 & new_new_n17932__;
  assign new_new_n17934__ = ~ys__n18284 & new_new_n17933__;
  assign new_new_n17935__ = ys__n19035 & ys__n18278;
  assign ys__n18518 = new_new_n17934__ | new_new_n17935__;
  assign new_new_n17937__ = ~ys__n18393 & ys__n18517;
  assign new_new_n17938__ = ys__n18393 & ys__n18518;
  assign ys__n18519 = new_new_n17937__ | new_new_n17938__;
  assign new_new_n17940__ = ys__n19140 & ~ys__n18281;
  assign new_new_n17941__ = ~ys__n18278 & new_new_n17940__;
  assign new_new_n17942__ = ys__n18287 & new_new_n17941__;
  assign new_new_n17943__ = ~ys__n18284 & new_new_n17942__;
  assign new_new_n17944__ = ys__n19037 & ys__n18278;
  assign ys__n18521 = new_new_n17943__ | new_new_n17944__;
  assign new_new_n17946__ = ~ys__n18393 & ys__n18520;
  assign new_new_n17947__ = ys__n18393 & ys__n18521;
  assign ys__n18522 = new_new_n17946__ | new_new_n17947__;
  assign new_new_n17949__ = ys__n19141 & ~ys__n18281;
  assign new_new_n17950__ = ~ys__n18278 & new_new_n17949__;
  assign new_new_n17951__ = ys__n18287 & new_new_n17950__;
  assign new_new_n17952__ = ~ys__n18284 & new_new_n17951__;
  assign new_new_n17953__ = ys__n19039 & ys__n18278;
  assign ys__n18524 = new_new_n17952__ | new_new_n17953__;
  assign new_new_n17955__ = ~ys__n18393 & ys__n18523;
  assign new_new_n17956__ = ys__n18393 & ys__n18524;
  assign ys__n18525 = new_new_n17955__ | new_new_n17956__;
  assign new_new_n17958__ = ys__n19142 & ~ys__n18281;
  assign new_new_n17959__ = ~ys__n18278 & new_new_n17958__;
  assign new_new_n17960__ = ys__n18287 & new_new_n17959__;
  assign new_new_n17961__ = ~ys__n18284 & new_new_n17960__;
  assign new_new_n17962__ = ys__n19041 & ys__n18278;
  assign ys__n18527 = new_new_n17961__ | new_new_n17962__;
  assign new_new_n17964__ = ~ys__n18393 & ys__n18526;
  assign new_new_n17965__ = ys__n18393 & ys__n18527;
  assign ys__n18528 = new_new_n17964__ | new_new_n17965__;
  assign new_new_n17967__ = ys__n19143 & ~ys__n18281;
  assign new_new_n17968__ = ~ys__n18278 & new_new_n17967__;
  assign new_new_n17969__ = ys__n18287 & new_new_n17968__;
  assign new_new_n17970__ = ~ys__n18284 & new_new_n17969__;
  assign new_new_n17971__ = ys__n19043 & ys__n18278;
  assign ys__n18530 = new_new_n17970__ | new_new_n17971__;
  assign new_new_n17973__ = ~ys__n18393 & ys__n18529;
  assign new_new_n17974__ = ys__n18393 & ys__n18530;
  assign ys__n18531 = new_new_n17973__ | new_new_n17974__;
  assign new_new_n17976__ = ys__n19144 & ~ys__n18281;
  assign new_new_n17977__ = ~ys__n18278 & new_new_n17976__;
  assign new_new_n17978__ = ys__n18287 & new_new_n17977__;
  assign new_new_n17979__ = ~ys__n18284 & new_new_n17978__;
  assign new_new_n17980__ = ys__n19045 & ys__n18278;
  assign ys__n18533 = new_new_n17979__ | new_new_n17980__;
  assign new_new_n17982__ = ~ys__n18393 & ys__n18532;
  assign new_new_n17983__ = ys__n18393 & ys__n18533;
  assign ys__n18534 = new_new_n17982__ | new_new_n17983__;
  assign new_new_n17985__ = ys__n19145 & ~ys__n18281;
  assign new_new_n17986__ = ~ys__n18278 & new_new_n17985__;
  assign new_new_n17987__ = ys__n18287 & new_new_n17986__;
  assign new_new_n17988__ = ~ys__n18284 & new_new_n17987__;
  assign new_new_n17989__ = ys__n19047 & ys__n18278;
  assign ys__n18536 = new_new_n17988__ | new_new_n17989__;
  assign new_new_n17991__ = ~ys__n18393 & ys__n18535;
  assign new_new_n17992__ = ys__n18393 & ys__n18536;
  assign ys__n18537 = new_new_n17991__ | new_new_n17992__;
  assign new_new_n17994__ = ys__n19146 & ~ys__n18281;
  assign new_new_n17995__ = ~ys__n18278 & new_new_n17994__;
  assign new_new_n17996__ = ys__n18287 & new_new_n17995__;
  assign new_new_n17997__ = ~ys__n18284 & new_new_n17996__;
  assign new_new_n17998__ = ys__n19049 & ys__n18278;
  assign ys__n18539 = new_new_n17997__ | new_new_n17998__;
  assign new_new_n18000__ = ~ys__n18393 & ys__n18538;
  assign new_new_n18001__ = ys__n18393 & ys__n18539;
  assign ys__n18540 = new_new_n18000__ | new_new_n18001__;
  assign new_new_n18003__ = ys__n19147 & ~ys__n18281;
  assign new_new_n18004__ = ~ys__n18278 & new_new_n18003__;
  assign new_new_n18005__ = ys__n18287 & new_new_n18004__;
  assign new_new_n18006__ = ~ys__n18284 & new_new_n18005__;
  assign new_new_n18007__ = ys__n19051 & ys__n18278;
  assign ys__n18542 = new_new_n18006__ | new_new_n18007__;
  assign new_new_n18009__ = ~ys__n18393 & ys__n18541;
  assign new_new_n18010__ = ys__n18393 & ys__n18542;
  assign ys__n18543 = new_new_n18009__ | new_new_n18010__;
  assign new_new_n18012__ = ys__n18281 & ~ys__n18278;
  assign ys__n18548 = ys__n18278 | new_new_n18012__;
  assign new_new_n18014__ = ys__n18065 & ~ys__n18393;
  assign new_new_n18015__ = ys__n18393 & ys__n18548;
  assign ys__n18549 = new_new_n18014__ | new_new_n18015__;
  assign new_new_n18017__ = ys__n19166 & ys__n18287;
  assign new_new_n18018__ = ~ys__n18284 & new_new_n18017__;
  assign new_new_n18019__ = ys__n18758 & ~new_new_n11122__;
  assign new_new_n18020__ = ys__n18759 & new_new_n11122__;
  assign ys__n18760 = new_new_n18019__ | new_new_n18020__;
  assign new_new_n18022__ = ys__n18284 & ys__n18760;
  assign new_new_n18023__ = ~new_new_n18018__ & ~new_new_n18022__;
  assign new_new_n18024__ = ~ys__n18281 & ~new_new_n18023__;
  assign new_new_n18025__ = ys__n18281 & ys__n18649;
  assign new_new_n18026__ = ~new_new_n18024__ & ~new_new_n18025__;
  assign ys__n18550 = ~ys__n18278 & ~new_new_n18026__;
  assign new_new_n18028__ = ys__n18059 & ~ys__n18393;
  assign new_new_n18029__ = ys__n18393 & ys__n18550;
  assign ys__n18551 = new_new_n18028__ | new_new_n18029__;
  assign ys__n19183 = ~new_new_n12143__ & ~ys__n18360;
  assign new_new_n18032__ = ~new_new_n12143__ & ~ys__n19183;
  assign new_new_n18033__ = new_new_n12070__ & ~new_new_n12127__;
  assign new_new_n18034__ = ~new_new_n18032__ & new_new_n18033__;
  assign new_new_n18035__ = new_new_n12070__ & ~new_new_n18034__;
  assign new_new_n18036__ = ~ys__n2 & ~new_new_n18035__;
  assign new_new_n18037__ = ~new_new_n12070__ & new_new_n12143__;
  assign new_new_n18038__ = new_new_n12143__ & ys__n18360;
  assign new_new_n18039__ = new_new_n12143__ & ~new_new_n18038__;
  assign new_new_n18040__ = new_new_n12127__ & ~new_new_n18039__;
  assign new_new_n18041__ = new_new_n12127__ & ~new_new_n18040__;
  assign new_new_n18042__ = new_new_n12070__ & ~new_new_n18041__;
  assign new_new_n18043__ = ~new_new_n18037__ & ~new_new_n18042__;
  assign new_new_n18044__ = ys__n2 & ~new_new_n18043__;
  assign ys__n18553 = new_new_n18036__ | new_new_n18044__;
  assign new_new_n18046__ = ys__n18277 & ~ys__n18393;
  assign new_new_n18047__ = ys__n18393 & ys__n18278;
  assign ys__n18554 = new_new_n18046__ | new_new_n18047__;
  assign new_new_n18049__ = ys__n18650 & ~new_new_n11125__;
  assign new_new_n18050__ = ys__n18651 & new_new_n11125__;
  assign ys__n18652 = new_new_n18049__ | new_new_n18050__;
  assign new_new_n18052__ = ys__n18761 & ~new_new_n11122__;
  assign new_new_n18053__ = ys__n18762 & new_new_n11122__;
  assign ys__n18763 = new_new_n18052__ | new_new_n18053__;
  assign new_new_n18055__ = ys__n124 & ~ys__n18303;
  assign new_new_n18056__ = ys__n4615 & ys__n18303;
  assign new_new_n18057__ = ~new_new_n18055__ & ~new_new_n18056__;
  assign ys__n19173 = ys__n874 & ~new_new_n18057__;
  assign new_new_n18059__ = ys__n126 & ~ys__n18303;
  assign new_new_n18060__ = ys__n714 & ys__n18303;
  assign new_new_n18061__ = ~new_new_n18059__ & ~new_new_n18060__;
  assign new_new_n18062__ = ys__n874 & ~new_new_n18061__;
  assign new_new_n18063__ = ys__n122 & ~ys__n18303;
  assign new_new_n18064__ = ys__n716 & ys__n18303;
  assign new_new_n18065__ = ~new_new_n18063__ & ~new_new_n18064__;
  assign new_new_n18066__ = ys__n874 & ~new_new_n18065__;
  assign new_new_n18067__ = new_new_n18062__ & ~new_new_n18066__;
  assign new_new_n18068__ = ys__n19173 & new_new_n18062__;
  assign new_new_n18069__ = new_new_n18066__ & new_new_n18068__;
  assign ys__n19177 = new_new_n18067__ | new_new_n18069__;
  assign new_new_n18071__ = ~ys__n19173 & ~new_new_n18066__;
  assign new_new_n18072__ = ys__n19173 & new_new_n18066__;
  assign ys__n19178 = new_new_n18071__ | new_new_n18072__;
  assign new_new_n18074__ = ys__n826 & new_new_n11727__;
  assign new_new_n18075__ = ~new_new_n11731__ & new_new_n18074__;
  assign new_new_n18076__ = ys__n822 & new_new_n11731__;
  assign ys__n19227 = new_new_n18075__ | new_new_n18076__;
  assign new_new_n18078__ = ys__n824 & new_new_n11727__;
  assign new_new_n18079__ = ~new_new_n11731__ & new_new_n18078__;
  assign new_new_n18080__ = ys__n820 & new_new_n11731__;
  assign ys__n19229 = new_new_n18079__ | new_new_n18080__;
  assign new_new_n18082__ = ys__n822 & new_new_n11727__;
  assign new_new_n18083__ = ~new_new_n11731__ & new_new_n18082__;
  assign new_new_n18084__ = ys__n818 & new_new_n11731__;
  assign ys__n19231 = new_new_n18083__ | new_new_n18084__;
  assign new_new_n18086__ = ys__n820 & new_new_n11727__;
  assign new_new_n18087__ = ~new_new_n11731__ & new_new_n18086__;
  assign new_new_n18088__ = ys__n816 & new_new_n11731__;
  assign ys__n19233 = new_new_n18087__ | new_new_n18088__;
  assign new_new_n18090__ = ys__n818 & new_new_n11727__;
  assign new_new_n18091__ = ~new_new_n11731__ & new_new_n18090__;
  assign new_new_n18092__ = ys__n1301 & new_new_n11731__;
  assign ys__n19235 = new_new_n18091__ | new_new_n18092__;
  assign new_new_n18094__ = ~ys__n27737 & ys__n732;
  assign new_new_n18095__ = new_new_n11726__ & new_new_n18094__;
  assign new_new_n18096__ = ~ys__n730 & new_new_n18095__;
  assign new_new_n18097__ = ~ys__n27737 & ~new_new_n11726__;
  assign new_new_n18098__ = ys__n4603 & new_new_n18097__;
  assign ys__n19239 = new_new_n18096__ | new_new_n18098__;
  assign new_new_n18100__ = ys__n19245 & ~ys__n19251;
  assign new_new_n18101__ = ~new_new_n10860__ & ~new_new_n18100__;
  assign new_new_n18102__ = ~ys__n19253 & ~new_new_n18101__;
  assign ys__n19254 = new_new_n10858__ | new_new_n18102__;
  assign new_new_n18104__ = ys__n19251 & new_new_n10834__;
  assign ys__n19257 = new_new_n10872__ | new_new_n18104__;
  assign new_new_n18106__ = ys__n140 & ~ys__n19259;
  assign new_new_n18107__ = ys__n19259 & ~ys__n19261;
  assign new_new_n18108__ = ~new_new_n18106__ & ~new_new_n18107__;
  assign new_new_n18109__ = ~ys__n19263 & ~new_new_n18108__;
  assign new_new_n18110__ = ys__n19263 & ys__n3039;
  assign ys__n19264 = new_new_n18109__ | new_new_n18110__;
  assign new_new_n18112__ = ys__n19259 & ys__n19261;
  assign new_new_n18113__ = ~ys__n19263 & new_new_n18112__;
  assign new_new_n18114__ = ys__n19263 & ~ys__n3039;
  assign ys__n19266 = new_new_n18113__ | new_new_n18114__;
  assign new_new_n18116__ = ~ys__n1505 & ~ys__n1506;
  assign new_new_n18117__ = ys__n19843 & ys__n19844;
  assign new_new_n18118__ = new_new_n18116__ & new_new_n18117__;
  assign new_new_n18119__ = ys__n23335 & ys__n27857;
  assign new_new_n18120__ = ~new_new_n10765__ & ~new_new_n18119__;
  assign new_new_n18121__ = ~ys__n23272 & ~new_new_n18120__;
  assign new_new_n18122__ = ~ys__n23335 & ys__n27859;
  assign new_new_n18123__ = ys__n23335 & ys__n27861;
  assign new_new_n18124__ = ~new_new_n18122__ & ~new_new_n18123__;
  assign new_new_n18125__ = ys__n23272 & ~new_new_n18124__;
  assign new_new_n18126__ = ~new_new_n18121__ & ~new_new_n18125__;
  assign new_new_n18127__ = ~ys__n23274 & ~new_new_n18126__;
  assign new_new_n18128__ = ~ys__n23335 & ys__n27863;
  assign new_new_n18129__ = ys__n23335 & ys__n27865;
  assign new_new_n18130__ = ~new_new_n18128__ & ~new_new_n18129__;
  assign new_new_n18131__ = ~ys__n23272 & ~new_new_n18130__;
  assign new_new_n18132__ = ~ys__n23335 & ys__n27867;
  assign new_new_n18133__ = ys__n23335 & ys__n27869;
  assign new_new_n18134__ = ~new_new_n18132__ & ~new_new_n18133__;
  assign new_new_n18135__ = ys__n23272 & ~new_new_n18134__;
  assign new_new_n18136__ = ~new_new_n18131__ & ~new_new_n18135__;
  assign new_new_n18137__ = ys__n23274 & ~new_new_n18136__;
  assign new_new_n18138__ = ~new_new_n18127__ & ~new_new_n18137__;
  assign new_new_n18139__ = ~ys__n23276 & ~new_new_n18138__;
  assign new_new_n18140__ = ~ys__n23335 & ys__n27871;
  assign new_new_n18141__ = ys__n23335 & ys__n27873;
  assign new_new_n18142__ = ~new_new_n18140__ & ~new_new_n18141__;
  assign new_new_n18143__ = ~ys__n23272 & ~new_new_n18142__;
  assign new_new_n18144__ = ~ys__n23335 & ys__n27875;
  assign new_new_n18145__ = ys__n23335 & ys__n27877;
  assign new_new_n18146__ = ~new_new_n18144__ & ~new_new_n18145__;
  assign new_new_n18147__ = ys__n23272 & ~new_new_n18146__;
  assign new_new_n18148__ = ~new_new_n18143__ & ~new_new_n18147__;
  assign new_new_n18149__ = ~ys__n23274 & ~new_new_n18148__;
  assign new_new_n18150__ = ~ys__n23335 & ys__n27879;
  assign new_new_n18151__ = ys__n23335 & ys__n27881;
  assign new_new_n18152__ = ~new_new_n18150__ & ~new_new_n18151__;
  assign new_new_n18153__ = ~ys__n23272 & ~new_new_n18152__;
  assign new_new_n18154__ = ~ys__n23335 & ys__n27883;
  assign new_new_n18155__ = ys__n23335 & ys__n27885;
  assign new_new_n18156__ = ~new_new_n18154__ & ~new_new_n18155__;
  assign new_new_n18157__ = ys__n23272 & ~new_new_n18156__;
  assign new_new_n18158__ = ~new_new_n18153__ & ~new_new_n18157__;
  assign new_new_n18159__ = ys__n23274 & ~new_new_n18158__;
  assign new_new_n18160__ = ~new_new_n18149__ & ~new_new_n18159__;
  assign new_new_n18161__ = ys__n23276 & ~new_new_n18160__;
  assign new_new_n18162__ = ~new_new_n18139__ & ~new_new_n18161__;
  assign new_new_n18163__ = ~ys__n23278 & ~new_new_n18162__;
  assign new_new_n18164__ = ~ys__n23335 & ys__n28015;
  assign new_new_n18165__ = ys__n23335 & ys__n28016;
  assign new_new_n18166__ = ~new_new_n18164__ & ~new_new_n18165__;
  assign new_new_n18167__ = ~ys__n23272 & ~new_new_n18166__;
  assign new_new_n18168__ = ~ys__n23335 & ys__n28017;
  assign new_new_n18169__ = ys__n23335 & ys__n28018;
  assign new_new_n18170__ = ~new_new_n18168__ & ~new_new_n18169__;
  assign new_new_n18171__ = ys__n23272 & ~new_new_n18170__;
  assign new_new_n18172__ = ~new_new_n18167__ & ~new_new_n18171__;
  assign new_new_n18173__ = ~ys__n23274 & ~new_new_n18172__;
  assign new_new_n18174__ = ~ys__n23335 & ys__n28019;
  assign new_new_n18175__ = ys__n23335 & ys__n28020;
  assign new_new_n18176__ = ~new_new_n18174__ & ~new_new_n18175__;
  assign new_new_n18177__ = ~ys__n23272 & ~new_new_n18176__;
  assign new_new_n18178__ = ~ys__n23335 & ys__n28021;
  assign new_new_n18179__ = ys__n23335 & ys__n28022;
  assign new_new_n18180__ = ~new_new_n18178__ & ~new_new_n18179__;
  assign new_new_n18181__ = ys__n23272 & ~new_new_n18180__;
  assign new_new_n18182__ = ~new_new_n18177__ & ~new_new_n18181__;
  assign new_new_n18183__ = ys__n23274 & ~new_new_n18182__;
  assign new_new_n18184__ = ~new_new_n18173__ & ~new_new_n18183__;
  assign new_new_n18185__ = ~ys__n23276 & ~new_new_n18184__;
  assign new_new_n18186__ = ~ys__n23335 & ys__n28023;
  assign new_new_n18187__ = ys__n23335 & ys__n28024;
  assign new_new_n18188__ = ~new_new_n18186__ & ~new_new_n18187__;
  assign new_new_n18189__ = ~ys__n23272 & ~new_new_n18188__;
  assign new_new_n18190__ = ~ys__n23335 & ys__n28025;
  assign new_new_n18191__ = ys__n23335 & ys__n28026;
  assign new_new_n18192__ = ~new_new_n18190__ & ~new_new_n18191__;
  assign new_new_n18193__ = ys__n23272 & ~new_new_n18192__;
  assign new_new_n18194__ = ~new_new_n18189__ & ~new_new_n18193__;
  assign new_new_n18195__ = ~ys__n23274 & ~new_new_n18194__;
  assign new_new_n18196__ = ~ys__n23335 & ys__n28027;
  assign new_new_n18197__ = ys__n23335 & ys__n28028;
  assign new_new_n18198__ = ~new_new_n18196__ & ~new_new_n18197__;
  assign new_new_n18199__ = ~ys__n23272 & ~new_new_n18198__;
  assign new_new_n18200__ = ~ys__n23335 & ys__n28029;
  assign new_new_n18201__ = ys__n23335 & ys__n28030;
  assign new_new_n18202__ = ~new_new_n18200__ & ~new_new_n18201__;
  assign new_new_n18203__ = ys__n23272 & ~new_new_n18202__;
  assign new_new_n18204__ = ~new_new_n18199__ & ~new_new_n18203__;
  assign new_new_n18205__ = ys__n23274 & ~new_new_n18204__;
  assign new_new_n18206__ = ~new_new_n18195__ & ~new_new_n18205__;
  assign new_new_n18207__ = ys__n23276 & ~new_new_n18206__;
  assign new_new_n18208__ = ~new_new_n18185__ & ~new_new_n18207__;
  assign new_new_n18209__ = ys__n23278 & ~new_new_n18208__;
  assign new_new_n18210__ = ~new_new_n18163__ & ~new_new_n18209__;
  assign new_new_n18211__ = ~new_new_n18116__ & ~new_new_n18210__;
  assign new_new_n18212__ = ~new_new_n18118__ & ~new_new_n18211__;
  assign new_new_n18213__ = ~ys__n1502 & ~ys__n1503;
  assign new_new_n18214__ = ~new_new_n18212__ & new_new_n18213__;
  assign new_new_n18215__ = ~ys__n23272 & new_new_n10765__;
  assign new_new_n18216__ = ~ys__n23274 & new_new_n18215__;
  assign new_new_n18217__ = ~ys__n23276 & new_new_n18216__;
  assign new_new_n18218__ = ys__n1502 & ~ys__n23278;
  assign new_new_n18219__ = ~new_new_n18213__ & new_new_n18218__;
  assign new_new_n18220__ = new_new_n18217__ & new_new_n18219__;
  assign new_new_n18221__ = ~new_new_n18214__ & ~new_new_n18220__;
  assign new_new_n18222__ = ~ys__n1495 & ~ys__n1496;
  assign new_new_n18223__ = ~ys__n1498 & ~ys__n1499;
  assign new_new_n18224__ = new_new_n18222__ & new_new_n18223__;
  assign new_new_n18225__ = ~new_new_n18221__ & new_new_n18224__;
  assign new_new_n18226__ = ~ys__n1498 & ys__n1499;
  assign new_new_n18227__ = ~new_new_n10767__ & new_new_n18226__;
  assign new_new_n18228__ = ~ys__n23335 & ~ys__n27855;
  assign new_new_n18229__ = ys__n1498 & new_new_n18228__;
  assign new_new_n18230__ = ~new_new_n18227__ & ~new_new_n18229__;
  assign new_new_n18231__ = ~ys__n1496 & ~new_new_n18230__;
  assign new_new_n18232__ = ys__n1496 & ~new_new_n18228__;
  assign new_new_n18233__ = ~new_new_n18231__ & ~new_new_n18232__;
  assign new_new_n18234__ = ~ys__n1495 & ~new_new_n18233__;
  assign new_new_n18235__ = ys__n1495 & new_new_n16609__;
  assign new_new_n18236__ = ~new_new_n18234__ & ~new_new_n18235__;
  assign new_new_n18237__ = ~new_new_n18224__ & ~new_new_n18236__;
  assign new_new_n18238__ = ~new_new_n18225__ & ~new_new_n18237__;
  assign new_new_n18239__ = ~ys__n1492 & ~ys__n1493;
  assign new_new_n18240__ = ~new_new_n18238__ & new_new_n18239__;
  assign new_new_n18241__ = ~ys__n1492 & ys__n23332;
  assign new_new_n18242__ = ~ys__n1492 & ys__n28030;
  assign new_new_n18243__ = ~new_new_n18241__ & ~new_new_n18242__;
  assign new_new_n18244__ = new_new_n18241__ & new_new_n18242__;
  assign new_new_n18245__ = ~new_new_n18243__ & ~new_new_n18244__;
  assign new_new_n18246__ = ~ys__n23272 & ~ys__n27857;
  assign new_new_n18247__ = ~new_new_n16777__ & ~new_new_n18246__;
  assign new_new_n18248__ = ~new_new_n16609__ & ~new_new_n18228__;
  assign new_new_n18249__ = ~new_new_n10766__ & new_new_n18248__;
  assign new_new_n18250__ = ~new_new_n18247__ & ~new_new_n18249__;
  assign new_new_n18251__ = ~new_new_n10769__ & ~new_new_n18250__;
  assign new_new_n18252__ = ~ys__n23276 & ~ys__n27861;
  assign new_new_n18253__ = ~new_new_n16782__ & ~new_new_n18252__;
  assign new_new_n18254__ = ~ys__n23274 & ~ys__n27859;
  assign new_new_n18255__ = ~new_new_n16783__ & ~new_new_n18254__;
  assign new_new_n18256__ = ~new_new_n18253__ & ~new_new_n18255__;
  assign new_new_n18257__ = ~new_new_n18251__ & new_new_n18256__;
  assign new_new_n18258__ = new_new_n10773__ & ~new_new_n18253__;
  assign new_new_n18259__ = ~new_new_n10776__ & ~new_new_n18258__;
  assign new_new_n18260__ = ~new_new_n18257__ & new_new_n18259__;
  assign new_new_n18261__ = ~ys__n23284 & ~ys__n27869;
  assign new_new_n18262__ = ~new_new_n16796__ & ~new_new_n18261__;
  assign new_new_n18263__ = ~ys__n23282 & ~ys__n27867;
  assign new_new_n18264__ = ~new_new_n16797__ & ~new_new_n18263__;
  assign new_new_n18265__ = ~new_new_n18262__ & ~new_new_n18264__;
  assign new_new_n18266__ = ~ys__n23280 & ~ys__n27865;
  assign new_new_n18267__ = ~new_new_n16791__ & ~new_new_n18266__;
  assign new_new_n18268__ = ~ys__n23278 & ~ys__n27863;
  assign new_new_n18269__ = ~new_new_n16792__ & ~new_new_n18268__;
  assign new_new_n18270__ = ~new_new_n18267__ & ~new_new_n18269__;
  assign new_new_n18271__ = new_new_n18265__ & new_new_n18270__;
  assign new_new_n18272__ = ~new_new_n18260__ & new_new_n18271__;
  assign new_new_n18273__ = new_new_n10751__ & ~new_new_n18267__;
  assign new_new_n18274__ = ~new_new_n10754__ & ~new_new_n18273__;
  assign new_new_n18275__ = new_new_n18265__ & ~new_new_n18274__;
  assign new_new_n18276__ = new_new_n10758__ & ~new_new_n18262__;
  assign new_new_n18277__ = ~new_new_n10761__ & ~new_new_n18276__;
  assign new_new_n18278__ = ~new_new_n18275__ & new_new_n18277__;
  assign new_new_n18279__ = ~new_new_n18272__ & new_new_n18278__;
  assign new_new_n18280__ = ~ys__n23300 & ~ys__n27885;
  assign new_new_n18281__ = ~new_new_n16826__ & ~new_new_n18280__;
  assign new_new_n18282__ = ~ys__n23298 & ~ys__n27883;
  assign new_new_n18283__ = ~new_new_n16827__ & ~new_new_n18282__;
  assign new_new_n18284__ = ~new_new_n18281__ & ~new_new_n18283__;
  assign new_new_n18285__ = ~ys__n23296 & ~ys__n27881;
  assign new_new_n18286__ = ~new_new_n16821__ & ~new_new_n18285__;
  assign new_new_n18287__ = ~ys__n23294 & ~ys__n27879;
  assign new_new_n18288__ = ~new_new_n16822__ & ~new_new_n18287__;
  assign new_new_n18289__ = ~new_new_n18286__ & ~new_new_n18288__;
  assign new_new_n18290__ = new_new_n18284__ & new_new_n18289__;
  assign new_new_n18291__ = ~ys__n23292 & ~ys__n27877;
  assign new_new_n18292__ = ~new_new_n16815__ & ~new_new_n18291__;
  assign new_new_n18293__ = ~ys__n23290 & ~ys__n27875;
  assign new_new_n18294__ = ~new_new_n16816__ & ~new_new_n18293__;
  assign new_new_n18295__ = ~new_new_n18292__ & ~new_new_n18294__;
  assign new_new_n18296__ = ~ys__n23288 & ~ys__n27873;
  assign new_new_n18297__ = ~new_new_n16810__ & ~new_new_n18296__;
  assign new_new_n18298__ = ~ys__n23286 & ~ys__n27871;
  assign new_new_n18299__ = ~new_new_n16811__ & ~new_new_n18298__;
  assign new_new_n18300__ = ~new_new_n18297__ & ~new_new_n18299__;
  assign new_new_n18301__ = new_new_n18295__ & new_new_n18300__;
  assign new_new_n18302__ = new_new_n18290__ & new_new_n18301__;
  assign new_new_n18303__ = ~new_new_n18279__ & new_new_n18302__;
  assign new_new_n18304__ = new_new_n10797__ & ~new_new_n18297__;
  assign new_new_n18305__ = ~new_new_n10800__ & ~new_new_n18304__;
  assign new_new_n18306__ = new_new_n18295__ & ~new_new_n18305__;
  assign new_new_n18307__ = new_new_n10804__ & ~new_new_n18292__;
  assign new_new_n18308__ = ~new_new_n10807__ & ~new_new_n18307__;
  assign new_new_n18309__ = ~new_new_n18306__ & new_new_n18308__;
  assign new_new_n18310__ = new_new_n18290__ & ~new_new_n18309__;
  assign new_new_n18311__ = new_new_n10782__ & ~new_new_n18286__;
  assign new_new_n18312__ = ~new_new_n10785__ & ~new_new_n18311__;
  assign new_new_n18313__ = new_new_n18284__ & ~new_new_n18312__;
  assign new_new_n18314__ = new_new_n10789__ & ~new_new_n18281__;
  assign new_new_n18315__ = ~new_new_n10792__ & ~new_new_n18314__;
  assign new_new_n18316__ = ~new_new_n18313__ & new_new_n18315__;
  assign new_new_n18317__ = ~new_new_n18310__ & new_new_n18316__;
  assign new_new_n18318__ = ~new_new_n18303__ & new_new_n18317__;
  assign new_new_n18319__ = ~ys__n23332 & ~ys__n28030;
  assign new_new_n18320__ = ys__n23332 & ys__n28030;
  assign new_new_n18321__ = ~new_new_n18319__ & ~new_new_n18320__;
  assign new_new_n18322__ = ~ys__n23330 & ~ys__n28029;
  assign new_new_n18323__ = ~new_new_n16856__ & ~new_new_n18322__;
  assign new_new_n18324__ = ~new_new_n18321__ & ~new_new_n18323__;
  assign new_new_n18325__ = ~ys__n23328 & ~ys__n28028;
  assign new_new_n18326__ = ~new_new_n16844__ & ~new_new_n18325__;
  assign new_new_n18327__ = ~ys__n23326 & ~ys__n28027;
  assign new_new_n18328__ = ~new_new_n16734__ & ~new_new_n18327__;
  assign new_new_n18329__ = ~new_new_n18326__ & ~new_new_n18328__;
  assign new_new_n18330__ = new_new_n18324__ & new_new_n18329__;
  assign new_new_n18331__ = ~ys__n23324 & ~ys__n28026;
  assign new_new_n18332__ = ~new_new_n16741__ & ~new_new_n18331__;
  assign new_new_n18333__ = ~ys__n23322 & ~ys__n28025;
  assign new_new_n18334__ = ~new_new_n16742__ & ~new_new_n18333__;
  assign new_new_n18335__ = ~new_new_n18332__ & ~new_new_n18334__;
  assign new_new_n18336__ = ~ys__n23320 & ~ys__n28024;
  assign new_new_n18337__ = ~new_new_n16736__ & ~new_new_n18336__;
  assign new_new_n18338__ = ~ys__n23318 & ~ys__n28023;
  assign new_new_n18339__ = ~new_new_n16737__ & ~new_new_n18338__;
  assign new_new_n18340__ = ~new_new_n18337__ & ~new_new_n18339__;
  assign new_new_n18341__ = new_new_n18335__ & new_new_n18340__;
  assign new_new_n18342__ = new_new_n18330__ & new_new_n18341__;
  assign new_new_n18343__ = ~ys__n23316 & ~ys__n28022;
  assign new_new_n18344__ = ~new_new_n16768__ & ~new_new_n18343__;
  assign new_new_n18345__ = ~ys__n23314 & ~ys__n28021;
  assign new_new_n18346__ = ~new_new_n16769__ & ~new_new_n18345__;
  assign new_new_n18347__ = ~new_new_n18344__ & ~new_new_n18346__;
  assign new_new_n18348__ = ~ys__n23312 & ~ys__n28020;
  assign new_new_n18349__ = ~new_new_n16763__ & ~new_new_n18348__;
  assign new_new_n18350__ = ~ys__n23310 & ~ys__n28019;
  assign new_new_n18351__ = ~new_new_n16764__ & ~new_new_n18350__;
  assign new_new_n18352__ = ~new_new_n18349__ & ~new_new_n18351__;
  assign new_new_n18353__ = new_new_n18347__ & new_new_n18352__;
  assign new_new_n18354__ = ~ys__n23308 & ~ys__n28018;
  assign new_new_n18355__ = ~new_new_n16757__ & ~new_new_n18354__;
  assign new_new_n18356__ = ~ys__n23306 & ~ys__n28017;
  assign new_new_n18357__ = ~new_new_n16758__ & ~new_new_n18356__;
  assign new_new_n18358__ = ~new_new_n18355__ & ~new_new_n18357__;
  assign new_new_n18359__ = ~ys__n23304 & ~ys__n28016;
  assign new_new_n18360__ = ~new_new_n16752__ & ~new_new_n18359__;
  assign new_new_n18361__ = ~ys__n23302 & ~ys__n28015;
  assign new_new_n18362__ = ~new_new_n16753__ & ~new_new_n18361__;
  assign new_new_n18363__ = ~new_new_n18360__ & ~new_new_n18362__;
  assign new_new_n18364__ = new_new_n18358__ & new_new_n18363__;
  assign new_new_n18365__ = new_new_n18353__ & new_new_n18364__;
  assign new_new_n18366__ = new_new_n18342__ & new_new_n18365__;
  assign new_new_n18367__ = ~new_new_n18318__ & new_new_n18366__;
  assign new_new_n18368__ = new_new_n10703__ & ~new_new_n18360__;
  assign new_new_n18369__ = ~new_new_n10706__ & ~new_new_n18368__;
  assign new_new_n18370__ = new_new_n18358__ & ~new_new_n18369__;
  assign new_new_n18371__ = new_new_n10710__ & ~new_new_n18355__;
  assign new_new_n18372__ = ~new_new_n10713__ & ~new_new_n18371__;
  assign new_new_n18373__ = ~new_new_n18370__ & new_new_n18372__;
  assign new_new_n18374__ = new_new_n18353__ & ~new_new_n18373__;
  assign new_new_n18375__ = new_new_n10688__ & ~new_new_n18349__;
  assign new_new_n18376__ = ~new_new_n10691__ & ~new_new_n18375__;
  assign new_new_n18377__ = new_new_n18347__ & ~new_new_n18376__;
  assign new_new_n18378__ = new_new_n10695__ & ~new_new_n18344__;
  assign new_new_n18379__ = ~new_new_n10698__ & ~new_new_n18378__;
  assign new_new_n18380__ = ~new_new_n18377__ & new_new_n18379__;
  assign new_new_n18381__ = ~new_new_n18374__ & new_new_n18380__;
  assign new_new_n18382__ = new_new_n18342__ & ~new_new_n18381__;
  assign new_new_n18383__ = new_new_n10734__ & ~new_new_n18337__;
  assign new_new_n18384__ = ~new_new_n10737__ & ~new_new_n18383__;
  assign new_new_n18385__ = new_new_n18335__ & ~new_new_n18384__;
  assign new_new_n18386__ = new_new_n10741__ & ~new_new_n18332__;
  assign new_new_n18387__ = ~new_new_n10744__ & ~new_new_n18386__;
  assign new_new_n18388__ = ~new_new_n18385__ & new_new_n18387__;
  assign new_new_n18389__ = new_new_n18330__ & ~new_new_n18388__;
  assign new_new_n18390__ = new_new_n10719__ & ~new_new_n18326__;
  assign new_new_n18391__ = ~new_new_n10722__ & ~new_new_n18390__;
  assign new_new_n18392__ = new_new_n18324__ & ~new_new_n18391__;
  assign new_new_n18393__ = new_new_n10726__ & ~new_new_n18321__;
  assign new_new_n18394__ = ~new_new_n10729__ & ~new_new_n18393__;
  assign new_new_n18395__ = ~new_new_n18392__ & new_new_n18394__;
  assign new_new_n18396__ = ~new_new_n18389__ & new_new_n18395__;
  assign new_new_n18397__ = ~new_new_n18382__ & new_new_n18396__;
  assign new_new_n18398__ = ~new_new_n18367__ & new_new_n18397__;
  assign new_new_n18399__ = new_new_n18245__ & ~new_new_n18398__;
  assign new_new_n18400__ = ~new_new_n18245__ & new_new_n18398__;
  assign new_new_n18401__ = ~new_new_n18399__ & ~new_new_n18400__;
  assign new_new_n18402__ = ~ys__n1489 & ~new_new_n18401__;
  assign new_new_n18403__ = ~new_new_n18241__ & new_new_n18242__;
  assign new_new_n18404__ = new_new_n18241__ & ~new_new_n18242__;
  assign new_new_n18405__ = ~new_new_n18403__ & ~new_new_n18404__;
  assign new_new_n18406__ = ~new_new_n10727__ & ~new_new_n10730__;
  assign new_new_n18407__ = new_new_n16847__ & new_new_n18406__;
  assign new_new_n18408__ = new_new_n16747__ & new_new_n18407__;
  assign new_new_n18409__ = new_new_n16776__ & new_new_n18408__;
  assign new_new_n18410__ = ~new_new_n16832__ & new_new_n18409__;
  assign new_new_n18411__ = ~new_new_n16773__ & new_new_n18408__;
  assign new_new_n18412__ = ~new_new_n16745__ & new_new_n18407__;
  assign new_new_n18413__ = ~new_new_n16846__ & new_new_n18406__;
  assign new_new_n18414__ = ~new_new_n10730__ & new_new_n16856__;
  assign new_new_n18415__ = ~new_new_n18320__ & ~new_new_n18414__;
  assign new_new_n18416__ = ~new_new_n18413__ & new_new_n18415__;
  assign new_new_n18417__ = ~new_new_n18412__ & new_new_n18416__;
  assign new_new_n18418__ = ~new_new_n18411__ & new_new_n18417__;
  assign new_new_n18419__ = ~new_new_n18410__ & new_new_n18418__;
  assign new_new_n18420__ = new_new_n18405__ & ~new_new_n18419__;
  assign new_new_n18421__ = ~new_new_n18405__ & new_new_n18419__;
  assign new_new_n18422__ = ~new_new_n18420__ & ~new_new_n18421__;
  assign new_new_n18423__ = ys__n1489 & ~new_new_n18422__;
  assign new_new_n18424__ = ~new_new_n18402__ & ~new_new_n18423__;
  assign new_new_n18425__ = ~new_new_n18239__ & ~new_new_n18424__;
  assign new_new_n18426__ = ~new_new_n18240__ & ~new_new_n18425__;
  assign new_new_n18427__ = ~ys__n1489 & ~ys__n1490;
  assign new_new_n18428__ = ~new_new_n18426__ & new_new_n18427__;
  assign new_new_n18429__ = ~ys__n1489 & new_new_n18248__;
  assign new_new_n18430__ = ys__n1489 & ~new_new_n10767__;
  assign new_new_n18431__ = ~new_new_n18429__ & ~new_new_n18430__;
  assign new_new_n18432__ = ~new_new_n18427__ & ~new_new_n18431__;
  assign new_new_n18433__ = ~new_new_n18428__ & ~new_new_n18432__;
  assign new_new_n18434__ = ~ys__n19973 & ~new_new_n18433__;
  assign new_new_n18435__ = ys__n19972 & ys__n19973;
  assign new_new_n18436__ = ~new_new_n18434__ & ~new_new_n18435__;
  assign new_new_n18437__ = ~ys__n352 & ~new_new_n18436__;
  assign new_new_n18438__ = ~ys__n220 & ys__n47026;
  assign new_new_n18439__ = ys__n222 & ys__n248;
  assign new_new_n18440__ = new_new_n18438__ & new_new_n18439__;
  assign new_new_n18441__ = ys__n222 & ~ys__n248;
  assign new_new_n18442__ = ~ys__n220 & ys__n47074;
  assign new_new_n18443__ = new_new_n18441__ & new_new_n18442__;
  assign new_new_n18444__ = ~ys__n222 & ys__n248;
  assign new_new_n18445__ = ~ys__n220 & ys__n47010;
  assign new_new_n18446__ = new_new_n18444__ & new_new_n18445__;
  assign new_new_n18447__ = ~new_new_n18443__ & ~new_new_n18446__;
  assign new_new_n18448__ = ~new_new_n18440__ & new_new_n18447__;
  assign new_new_n18449__ = ~new_new_n18441__ & ~new_new_n18444__;
  assign new_new_n18450__ = ~ys__n222 & ~ys__n248;
  assign new_new_n18451__ = ~new_new_n18439__ & ~new_new_n18450__;
  assign new_new_n18452__ = new_new_n18449__ & new_new_n18451__;
  assign new_new_n18453__ = ys__n352 & ~new_new_n18452__;
  assign new_new_n18454__ = ~new_new_n18448__ & new_new_n18453__;
  assign ys__n19878 = new_new_n18437__ | new_new_n18454__;
  assign new_new_n18456__ = ys__n19844 & ys__n19845;
  assign new_new_n18457__ = new_new_n18116__ & new_new_n18456__;
  assign new_new_n18458__ = ~ys__n23335 & ys__n27857;
  assign new_new_n18459__ = ys__n23335 & ys__n27859;
  assign new_new_n18460__ = ~new_new_n18458__ & ~new_new_n18459__;
  assign new_new_n18461__ = ~ys__n23272 & ~new_new_n18460__;
  assign new_new_n18462__ = ~ys__n23335 & ys__n27861;
  assign new_new_n18463__ = ys__n23335 & ys__n27863;
  assign new_new_n18464__ = ~new_new_n18462__ & ~new_new_n18463__;
  assign new_new_n18465__ = ys__n23272 & ~new_new_n18464__;
  assign new_new_n18466__ = ~new_new_n18461__ & ~new_new_n18465__;
  assign new_new_n18467__ = ~ys__n23274 & ~new_new_n18466__;
  assign new_new_n18468__ = ~ys__n23335 & ys__n27865;
  assign new_new_n18469__ = ys__n23335 & ys__n27867;
  assign new_new_n18470__ = ~new_new_n18468__ & ~new_new_n18469__;
  assign new_new_n18471__ = ~ys__n23272 & ~new_new_n18470__;
  assign new_new_n18472__ = ~ys__n23335 & ys__n27869;
  assign new_new_n18473__ = ys__n23335 & ys__n27871;
  assign new_new_n18474__ = ~new_new_n18472__ & ~new_new_n18473__;
  assign new_new_n18475__ = ys__n23272 & ~new_new_n18474__;
  assign new_new_n18476__ = ~new_new_n18471__ & ~new_new_n18475__;
  assign new_new_n18477__ = ys__n23274 & ~new_new_n18476__;
  assign new_new_n18478__ = ~new_new_n18467__ & ~new_new_n18477__;
  assign new_new_n18479__ = ~ys__n23276 & ~new_new_n18478__;
  assign new_new_n18480__ = ~ys__n23335 & ys__n27873;
  assign new_new_n18481__ = ys__n23335 & ys__n27875;
  assign new_new_n18482__ = ~new_new_n18480__ & ~new_new_n18481__;
  assign new_new_n18483__ = ~ys__n23272 & ~new_new_n18482__;
  assign new_new_n18484__ = ~ys__n23335 & ys__n27877;
  assign new_new_n18485__ = ys__n23335 & ys__n27879;
  assign new_new_n18486__ = ~new_new_n18484__ & ~new_new_n18485__;
  assign new_new_n18487__ = ys__n23272 & ~new_new_n18486__;
  assign new_new_n18488__ = ~new_new_n18483__ & ~new_new_n18487__;
  assign new_new_n18489__ = ~ys__n23274 & ~new_new_n18488__;
  assign new_new_n18490__ = ~ys__n23335 & ys__n27881;
  assign new_new_n18491__ = ys__n23335 & ys__n27883;
  assign new_new_n18492__ = ~new_new_n18490__ & ~new_new_n18491__;
  assign new_new_n18493__ = ~ys__n23272 & ~new_new_n18492__;
  assign new_new_n18494__ = ~ys__n23335 & ys__n27885;
  assign new_new_n18495__ = ys__n23335 & ys__n28015;
  assign new_new_n18496__ = ~new_new_n18494__ & ~new_new_n18495__;
  assign new_new_n18497__ = ys__n23272 & ~new_new_n18496__;
  assign new_new_n18498__ = ~new_new_n18493__ & ~new_new_n18497__;
  assign new_new_n18499__ = ys__n23274 & ~new_new_n18498__;
  assign new_new_n18500__ = ~new_new_n18489__ & ~new_new_n18499__;
  assign new_new_n18501__ = ys__n23276 & ~new_new_n18500__;
  assign new_new_n18502__ = ~new_new_n18479__ & ~new_new_n18501__;
  assign new_new_n18503__ = ~ys__n23278 & ~new_new_n18502__;
  assign new_new_n18504__ = ~ys__n23335 & ys__n28016;
  assign new_new_n18505__ = ys__n23335 & ys__n28017;
  assign new_new_n18506__ = ~new_new_n18504__ & ~new_new_n18505__;
  assign new_new_n18507__ = ~ys__n23272 & ~new_new_n18506__;
  assign new_new_n18508__ = ~ys__n23335 & ys__n28018;
  assign new_new_n18509__ = ys__n23335 & ys__n28019;
  assign new_new_n18510__ = ~new_new_n18508__ & ~new_new_n18509__;
  assign new_new_n18511__ = ys__n23272 & ~new_new_n18510__;
  assign new_new_n18512__ = ~new_new_n18507__ & ~new_new_n18511__;
  assign new_new_n18513__ = ~ys__n23274 & ~new_new_n18512__;
  assign new_new_n18514__ = ~ys__n23335 & ys__n28020;
  assign new_new_n18515__ = ys__n23335 & ys__n28021;
  assign new_new_n18516__ = ~new_new_n18514__ & ~new_new_n18515__;
  assign new_new_n18517__ = ~ys__n23272 & ~new_new_n18516__;
  assign new_new_n18518__ = ~ys__n23335 & ys__n28022;
  assign new_new_n18519__ = ys__n23335 & ys__n28023;
  assign new_new_n18520__ = ~new_new_n18518__ & ~new_new_n18519__;
  assign new_new_n18521__ = ys__n23272 & ~new_new_n18520__;
  assign new_new_n18522__ = ~new_new_n18517__ & ~new_new_n18521__;
  assign new_new_n18523__ = ys__n23274 & ~new_new_n18522__;
  assign new_new_n18524__ = ~new_new_n18513__ & ~new_new_n18523__;
  assign new_new_n18525__ = ~ys__n23276 & ~new_new_n18524__;
  assign new_new_n18526__ = ~ys__n23335 & ys__n28024;
  assign new_new_n18527__ = ys__n23335 & ys__n28025;
  assign new_new_n18528__ = ~new_new_n18526__ & ~new_new_n18527__;
  assign new_new_n18529__ = ~ys__n23272 & ~new_new_n18528__;
  assign new_new_n18530__ = ~ys__n23335 & ys__n28026;
  assign new_new_n18531__ = ys__n23335 & ys__n28027;
  assign new_new_n18532__ = ~new_new_n18530__ & ~new_new_n18531__;
  assign new_new_n18533__ = ys__n23272 & ~new_new_n18532__;
  assign new_new_n18534__ = ~new_new_n18529__ & ~new_new_n18533__;
  assign new_new_n18535__ = ~ys__n23274 & ~new_new_n18534__;
  assign new_new_n18536__ = ~ys__n23335 & ys__n28028;
  assign new_new_n18537__ = ys__n23335 & ys__n28029;
  assign new_new_n18538__ = ~new_new_n18536__ & ~new_new_n18537__;
  assign new_new_n18539__ = ~ys__n23272 & ~new_new_n18538__;
  assign new_new_n18540__ = ys__n23272 & ys__n28030;
  assign new_new_n18541__ = ~new_new_n18539__ & ~new_new_n18540__;
  assign new_new_n18542__ = ys__n23274 & ~new_new_n18541__;
  assign new_new_n18543__ = ~new_new_n18535__ & ~new_new_n18542__;
  assign new_new_n18544__ = ys__n23276 & ~new_new_n18543__;
  assign new_new_n18545__ = ~new_new_n18525__ & ~new_new_n18544__;
  assign new_new_n18546__ = ys__n23278 & ~new_new_n18545__;
  assign new_new_n18547__ = ~new_new_n18503__ & ~new_new_n18546__;
  assign new_new_n18548__ = ~ys__n1505 & ~new_new_n18547__;
  assign new_new_n18549__ = ~ys__n23335 & ys__n28030;
  assign new_new_n18550__ = ys__n23272 & new_new_n18549__;
  assign new_new_n18551__ = ~new_new_n18539__ & ~new_new_n18550__;
  assign new_new_n18552__ = ys__n23274 & ~new_new_n18551__;
  assign new_new_n18553__ = ~new_new_n18535__ & ~new_new_n18552__;
  assign new_new_n18554__ = ys__n23276 & ~new_new_n18553__;
  assign new_new_n18555__ = ~new_new_n18525__ & ~new_new_n18554__;
  assign new_new_n18556__ = ys__n23278 & ~new_new_n18555__;
  assign new_new_n18557__ = ~new_new_n18503__ & ~new_new_n18556__;
  assign new_new_n18558__ = ys__n1505 & ~new_new_n18557__;
  assign new_new_n18559__ = ~new_new_n18548__ & ~new_new_n18558__;
  assign new_new_n18560__ = ~new_new_n18116__ & ~new_new_n18559__;
  assign new_new_n18561__ = ~new_new_n18457__ & ~new_new_n18560__;
  assign new_new_n18562__ = new_new_n18213__ & ~new_new_n18561__;
  assign new_new_n18563__ = ~new_new_n16609__ & ~new_new_n18458__;
  assign new_new_n18564__ = ~ys__n23272 & ~new_new_n18563__;
  assign new_new_n18565__ = ~ys__n23274 & new_new_n18564__;
  assign new_new_n18566__ = ~ys__n23276 & new_new_n18565__;
  assign new_new_n18567__ = new_new_n18219__ & new_new_n18566__;
  assign new_new_n18568__ = ~new_new_n18562__ & ~new_new_n18567__;
  assign new_new_n18569__ = new_new_n18224__ & ~new_new_n18568__;
  assign new_new_n18570__ = ~new_new_n10770__ & new_new_n18226__;
  assign new_new_n18571__ = ys__n1498 & new_new_n18246__;
  assign new_new_n18572__ = ~new_new_n18570__ & ~new_new_n18571__;
  assign new_new_n18573__ = ~ys__n1496 & ~new_new_n18572__;
  assign new_new_n18574__ = ys__n1496 & ~new_new_n18246__;
  assign new_new_n18575__ = ~new_new_n18573__ & ~new_new_n18574__;
  assign new_new_n18576__ = ~ys__n1495 & ~new_new_n18575__;
  assign new_new_n18577__ = ys__n1495 & new_new_n16777__;
  assign new_new_n18578__ = ~new_new_n18576__ & ~new_new_n18577__;
  assign new_new_n18579__ = ~new_new_n18224__ & ~new_new_n18578__;
  assign new_new_n18580__ = ~new_new_n18569__ & ~new_new_n18579__;
  assign new_new_n18581__ = new_new_n18239__ & new_new_n18427__;
  assign new_new_n18582__ = ~new_new_n18580__ & new_new_n18581__;
  assign new_new_n18583__ = new_new_n18247__ & ~new_new_n18249__;
  assign new_new_n18584__ = ~new_new_n18247__ & new_new_n18249__;
  assign new_new_n18585__ = ~new_new_n18583__ & ~new_new_n18584__;
  assign new_new_n18586__ = ~ys__n1489 & ~new_new_n18585__;
  assign new_new_n18587__ = ys__n1489 & ~new_new_n16612__;
  assign new_new_n18588__ = ~new_new_n18586__ & ~new_new_n18587__;
  assign new_new_n18589__ = ~new_new_n18427__ & ~new_new_n18588__;
  assign new_new_n18590__ = ~new_new_n18582__ & ~new_new_n18589__;
  assign new_new_n18591__ = ~ys__n19973 & ~new_new_n18590__;
  assign new_new_n18592__ = ys__n19973 & ys__n19974;
  assign new_new_n18593__ = ~new_new_n18591__ & ~new_new_n18592__;
  assign new_new_n18594__ = ~ys__n352 & ~new_new_n18593__;
  assign new_new_n18595__ = ~ys__n220 & ys__n47027;
  assign new_new_n18596__ = new_new_n18439__ & new_new_n18595__;
  assign new_new_n18597__ = ~ys__n220 & ys__n47075;
  assign new_new_n18598__ = new_new_n18441__ & new_new_n18597__;
  assign new_new_n18599__ = ~ys__n220 & ys__n47011;
  assign new_new_n18600__ = new_new_n18444__ & new_new_n18599__;
  assign new_new_n18601__ = ~new_new_n18598__ & ~new_new_n18600__;
  assign new_new_n18602__ = ~new_new_n18596__ & new_new_n18601__;
  assign new_new_n18603__ = new_new_n18453__ & ~new_new_n18602__;
  assign ys__n19881 = new_new_n18594__ | new_new_n18603__;
  assign new_new_n18605__ = ys__n19844 & ys__n19846;
  assign new_new_n18606__ = new_new_n18116__ & new_new_n18605__;
  assign new_new_n18607__ = ~ys__n23272 & ~new_new_n18124__;
  assign new_new_n18608__ = ys__n23272 & ~new_new_n18130__;
  assign new_new_n18609__ = ~new_new_n18607__ & ~new_new_n18608__;
  assign new_new_n18610__ = ~ys__n23274 & ~new_new_n18609__;
  assign new_new_n18611__ = ~ys__n23272 & ~new_new_n18134__;
  assign new_new_n18612__ = ys__n23272 & ~new_new_n18142__;
  assign new_new_n18613__ = ~new_new_n18611__ & ~new_new_n18612__;
  assign new_new_n18614__ = ys__n23274 & ~new_new_n18613__;
  assign new_new_n18615__ = ~new_new_n18610__ & ~new_new_n18614__;
  assign new_new_n18616__ = ~ys__n23276 & ~new_new_n18615__;
  assign new_new_n18617__ = ~ys__n23272 & ~new_new_n18146__;
  assign new_new_n18618__ = ys__n23272 & ~new_new_n18152__;
  assign new_new_n18619__ = ~new_new_n18617__ & ~new_new_n18618__;
  assign new_new_n18620__ = ~ys__n23274 & ~new_new_n18619__;
  assign new_new_n18621__ = ~ys__n23272 & ~new_new_n18156__;
  assign new_new_n18622__ = ys__n23272 & ~new_new_n18166__;
  assign new_new_n18623__ = ~new_new_n18621__ & ~new_new_n18622__;
  assign new_new_n18624__ = ys__n23274 & ~new_new_n18623__;
  assign new_new_n18625__ = ~new_new_n18620__ & ~new_new_n18624__;
  assign new_new_n18626__ = ys__n23276 & ~new_new_n18625__;
  assign new_new_n18627__ = ~new_new_n18616__ & ~new_new_n18626__;
  assign new_new_n18628__ = ~ys__n23278 & ~new_new_n18627__;
  assign new_new_n18629__ = ~ys__n23272 & ~new_new_n18170__;
  assign new_new_n18630__ = ys__n23272 & ~new_new_n18176__;
  assign new_new_n18631__ = ~new_new_n18629__ & ~new_new_n18630__;
  assign new_new_n18632__ = ~ys__n23274 & ~new_new_n18631__;
  assign new_new_n18633__ = ~ys__n23272 & ~new_new_n18180__;
  assign new_new_n18634__ = ys__n23272 & ~new_new_n18188__;
  assign new_new_n18635__ = ~new_new_n18633__ & ~new_new_n18634__;
  assign new_new_n18636__ = ys__n23274 & ~new_new_n18635__;
  assign new_new_n18637__ = ~new_new_n18632__ & ~new_new_n18636__;
  assign new_new_n18638__ = ~ys__n23276 & ~new_new_n18637__;
  assign new_new_n18639__ = ~ys__n23272 & ~new_new_n18192__;
  assign new_new_n18640__ = ys__n23272 & ~new_new_n18198__;
  assign new_new_n18641__ = ~new_new_n18639__ & ~new_new_n18640__;
  assign new_new_n18642__ = ~ys__n23274 & ~new_new_n18641__;
  assign new_new_n18643__ = ~ys__n23272 & ~new_new_n18202__;
  assign new_new_n18644__ = ~new_new_n18540__ & ~new_new_n18643__;
  assign new_new_n18645__ = ys__n23274 & ~new_new_n18644__;
  assign new_new_n18646__ = ~new_new_n18642__ & ~new_new_n18645__;
  assign new_new_n18647__ = ys__n23276 & ~new_new_n18646__;
  assign new_new_n18648__ = ~new_new_n18638__ & ~new_new_n18647__;
  assign new_new_n18649__ = ys__n23278 & ~new_new_n18648__;
  assign new_new_n18650__ = ~new_new_n18628__ & ~new_new_n18649__;
  assign new_new_n18651__ = ~ys__n1505 & ~new_new_n18650__;
  assign new_new_n18652__ = ys__n23274 & new_new_n18643__;
  assign new_new_n18653__ = ~new_new_n18642__ & ~new_new_n18652__;
  assign new_new_n18654__ = ys__n23276 & ~new_new_n18653__;
  assign new_new_n18655__ = ~new_new_n18638__ & ~new_new_n18654__;
  assign new_new_n18656__ = ys__n23278 & ~new_new_n18655__;
  assign new_new_n18657__ = ~new_new_n18628__ & ~new_new_n18656__;
  assign new_new_n18658__ = ys__n1505 & ~new_new_n18657__;
  assign new_new_n18659__ = ~new_new_n18651__ & ~new_new_n18658__;
  assign new_new_n18660__ = ~new_new_n18116__ & ~new_new_n18659__;
  assign new_new_n18661__ = ~new_new_n18606__ & ~new_new_n18660__;
  assign new_new_n18662__ = new_new_n18213__ & ~new_new_n18661__;
  assign new_new_n18663__ = ~new_new_n18119__ & ~new_new_n18122__;
  assign new_new_n18664__ = ~ys__n23272 & ~new_new_n18663__;
  assign new_new_n18665__ = ys__n23272 & new_new_n10765__;
  assign new_new_n18666__ = ~new_new_n18664__ & ~new_new_n18665__;
  assign new_new_n18667__ = ~ys__n23274 & ~new_new_n18666__;
  assign new_new_n18668__ = ~ys__n23276 & new_new_n18667__;
  assign new_new_n18669__ = new_new_n18219__ & new_new_n18668__;
  assign new_new_n18670__ = ~new_new_n18662__ & ~new_new_n18669__;
  assign new_new_n18671__ = new_new_n18224__ & ~new_new_n18670__;
  assign new_new_n18672__ = ~new_new_n10774__ & new_new_n18226__;
  assign new_new_n18673__ = ys__n1498 & new_new_n18254__;
  assign new_new_n18674__ = ~new_new_n18672__ & ~new_new_n18673__;
  assign new_new_n18675__ = ~ys__n1496 & ~new_new_n18674__;
  assign new_new_n18676__ = ys__n1496 & ~new_new_n18254__;
  assign new_new_n18677__ = ~new_new_n18675__ & ~new_new_n18676__;
  assign new_new_n18678__ = ~ys__n1495 & ~new_new_n18677__;
  assign new_new_n18679__ = ys__n1495 & new_new_n16783__;
  assign new_new_n18680__ = ~new_new_n18678__ & ~new_new_n18679__;
  assign new_new_n18681__ = ~new_new_n18224__ & ~new_new_n18680__;
  assign new_new_n18682__ = ~new_new_n18671__ & ~new_new_n18681__;
  assign new_new_n18683__ = new_new_n18581__ & ~new_new_n18682__;
  assign new_new_n18684__ = ~new_new_n18251__ & new_new_n18255__;
  assign new_new_n18685__ = new_new_n18251__ & ~new_new_n18255__;
  assign new_new_n18686__ = ~new_new_n18684__ & ~new_new_n18685__;
  assign new_new_n18687__ = ~ys__n1489 & ~new_new_n18686__;
  assign new_new_n18688__ = new_new_n10774__ & ~new_new_n16779__;
  assign new_new_n18689__ = ~new_new_n10774__ & new_new_n16779__;
  assign new_new_n18690__ = ~new_new_n18688__ & ~new_new_n18689__;
  assign new_new_n18691__ = ys__n1489 & ~new_new_n18690__;
  assign new_new_n18692__ = ~new_new_n18687__ & ~new_new_n18691__;
  assign new_new_n18693__ = ~new_new_n18427__ & ~new_new_n18692__;
  assign new_new_n18694__ = ~new_new_n18683__ & ~new_new_n18693__;
  assign new_new_n18695__ = ~ys__n19973 & ~new_new_n18694__;
  assign new_new_n18696__ = ys__n19973 & ys__n19975;
  assign new_new_n18697__ = ~new_new_n18695__ & ~new_new_n18696__;
  assign new_new_n18698__ = ~ys__n352 & ~new_new_n18697__;
  assign new_new_n18699__ = ~ys__n220 & ys__n47028;
  assign new_new_n18700__ = new_new_n18439__ & new_new_n18699__;
  assign new_new_n18701__ = ~ys__n220 & ys__n47076;
  assign new_new_n18702__ = new_new_n18441__ & new_new_n18701__;
  assign new_new_n18703__ = ~ys__n220 & ys__n47012;
  assign new_new_n18704__ = new_new_n18444__ & new_new_n18703__;
  assign new_new_n18705__ = ~new_new_n18702__ & ~new_new_n18704__;
  assign new_new_n18706__ = ~new_new_n18700__ & new_new_n18705__;
  assign new_new_n18707__ = new_new_n18453__ & ~new_new_n18706__;
  assign ys__n19884 = new_new_n18698__ | new_new_n18707__;
  assign new_new_n18709__ = ys__n19844 & ys__n19847;
  assign new_new_n18710__ = new_new_n18116__ & new_new_n18709__;
  assign new_new_n18711__ = ~ys__n23272 & ~new_new_n18464__;
  assign new_new_n18712__ = ys__n23272 & ~new_new_n18470__;
  assign new_new_n18713__ = ~new_new_n18711__ & ~new_new_n18712__;
  assign new_new_n18714__ = ~ys__n23274 & ~new_new_n18713__;
  assign new_new_n18715__ = ~ys__n23272 & ~new_new_n18474__;
  assign new_new_n18716__ = ys__n23272 & ~new_new_n18482__;
  assign new_new_n18717__ = ~new_new_n18715__ & ~new_new_n18716__;
  assign new_new_n18718__ = ys__n23274 & ~new_new_n18717__;
  assign new_new_n18719__ = ~new_new_n18714__ & ~new_new_n18718__;
  assign new_new_n18720__ = ~ys__n23276 & ~new_new_n18719__;
  assign new_new_n18721__ = ~ys__n23272 & ~new_new_n18486__;
  assign new_new_n18722__ = ys__n23272 & ~new_new_n18492__;
  assign new_new_n18723__ = ~new_new_n18721__ & ~new_new_n18722__;
  assign new_new_n18724__ = ~ys__n23274 & ~new_new_n18723__;
  assign new_new_n18725__ = ~ys__n23272 & ~new_new_n18496__;
  assign new_new_n18726__ = ys__n23272 & ~new_new_n18506__;
  assign new_new_n18727__ = ~new_new_n18725__ & ~new_new_n18726__;
  assign new_new_n18728__ = ys__n23274 & ~new_new_n18727__;
  assign new_new_n18729__ = ~new_new_n18724__ & ~new_new_n18728__;
  assign new_new_n18730__ = ys__n23276 & ~new_new_n18729__;
  assign new_new_n18731__ = ~new_new_n18720__ & ~new_new_n18730__;
  assign new_new_n18732__ = ~ys__n23278 & ~new_new_n18731__;
  assign new_new_n18733__ = ~ys__n23272 & ~new_new_n18510__;
  assign new_new_n18734__ = ys__n23272 & ~new_new_n18516__;
  assign new_new_n18735__ = ~new_new_n18733__ & ~new_new_n18734__;
  assign new_new_n18736__ = ~ys__n23274 & ~new_new_n18735__;
  assign new_new_n18737__ = ~ys__n23272 & ~new_new_n18520__;
  assign new_new_n18738__ = ys__n23272 & ~new_new_n18528__;
  assign new_new_n18739__ = ~new_new_n18737__ & ~new_new_n18738__;
  assign new_new_n18740__ = ys__n23274 & ~new_new_n18739__;
  assign new_new_n18741__ = ~new_new_n18736__ & ~new_new_n18740__;
  assign new_new_n18742__ = ~ys__n23276 & ~new_new_n18741__;
  assign new_new_n18743__ = ~ys__n23272 & ~new_new_n18532__;
  assign new_new_n18744__ = ys__n23272 & ~new_new_n18538__;
  assign new_new_n18745__ = ~new_new_n18743__ & ~new_new_n18744__;
  assign new_new_n18746__ = ~ys__n23274 & ~new_new_n18745__;
  assign new_new_n18747__ = ys__n23274 & ys__n28030;
  assign new_new_n18748__ = ~new_new_n18746__ & ~new_new_n18747__;
  assign new_new_n18749__ = ys__n23276 & ~new_new_n18748__;
  assign new_new_n18750__ = ~new_new_n18742__ & ~new_new_n18749__;
  assign new_new_n18751__ = ys__n23278 & ~new_new_n18750__;
  assign new_new_n18752__ = ~new_new_n18732__ & ~new_new_n18751__;
  assign new_new_n18753__ = ~ys__n1505 & ~new_new_n18752__;
  assign new_new_n18754__ = ~ys__n23272 & new_new_n18549__;
  assign new_new_n18755__ = ys__n23274 & new_new_n18754__;
  assign new_new_n18756__ = ~new_new_n18746__ & ~new_new_n18755__;
  assign new_new_n18757__ = ys__n23276 & ~new_new_n18756__;
  assign new_new_n18758__ = ~new_new_n18742__ & ~new_new_n18757__;
  assign new_new_n18759__ = ys__n23278 & ~new_new_n18758__;
  assign new_new_n18760__ = ~new_new_n18732__ & ~new_new_n18759__;
  assign new_new_n18761__ = ys__n1505 & ~new_new_n18760__;
  assign new_new_n18762__ = ~new_new_n18753__ & ~new_new_n18761__;
  assign new_new_n18763__ = ~new_new_n18116__ & ~new_new_n18762__;
  assign new_new_n18764__ = ~new_new_n18710__ & ~new_new_n18763__;
  assign new_new_n18765__ = new_new_n18213__ & ~new_new_n18764__;
  assign new_new_n18766__ = ~new_new_n18459__ & ~new_new_n18462__;
  assign new_new_n18767__ = ~ys__n23272 & ~new_new_n18766__;
  assign new_new_n18768__ = ys__n23272 & ~new_new_n18563__;
  assign new_new_n18769__ = ~new_new_n18767__ & ~new_new_n18768__;
  assign new_new_n18770__ = ~ys__n23274 & ~new_new_n18769__;
  assign new_new_n18771__ = ~ys__n23276 & new_new_n18770__;
  assign new_new_n18772__ = new_new_n18219__ & new_new_n18771__;
  assign new_new_n18773__ = ~new_new_n18765__ & ~new_new_n18772__;
  assign new_new_n18774__ = new_new_n18224__ & ~new_new_n18773__;
  assign new_new_n18775__ = ~new_new_n10777__ & new_new_n18226__;
  assign new_new_n18776__ = ys__n1498 & new_new_n18252__;
  assign new_new_n18777__ = ~new_new_n18775__ & ~new_new_n18776__;
  assign new_new_n18778__ = ~ys__n1496 & ~new_new_n18777__;
  assign new_new_n18779__ = ys__n1496 & ~new_new_n18252__;
  assign new_new_n18780__ = ~new_new_n18778__ & ~new_new_n18779__;
  assign new_new_n18781__ = ~ys__n1495 & ~new_new_n18780__;
  assign new_new_n18782__ = ys__n1495 & new_new_n16782__;
  assign new_new_n18783__ = ~new_new_n18781__ & ~new_new_n18782__;
  assign new_new_n18784__ = ~new_new_n18224__ & ~new_new_n18783__;
  assign new_new_n18785__ = ~new_new_n18774__ & ~new_new_n18784__;
  assign new_new_n18786__ = new_new_n18581__ & ~new_new_n18785__;
  assign new_new_n18787__ = ~new_new_n18251__ & ~new_new_n18255__;
  assign new_new_n18788__ = ~new_new_n10773__ & ~new_new_n18787__;
  assign new_new_n18789__ = new_new_n18253__ & ~new_new_n18788__;
  assign new_new_n18790__ = ~new_new_n18253__ & new_new_n18788__;
  assign new_new_n18791__ = ~new_new_n18789__ & ~new_new_n18790__;
  assign new_new_n18792__ = ~ys__n1489 & ~new_new_n18791__;
  assign new_new_n18793__ = ~new_new_n10774__ & ~new_new_n16779__;
  assign new_new_n18794__ = ~new_new_n16783__ & ~new_new_n18793__;
  assign new_new_n18795__ = new_new_n10777__ & ~new_new_n18794__;
  assign new_new_n18796__ = ~new_new_n10777__ & new_new_n18794__;
  assign new_new_n18797__ = ~new_new_n18795__ & ~new_new_n18796__;
  assign new_new_n18798__ = ys__n1489 & ~new_new_n18797__;
  assign new_new_n18799__ = ~new_new_n18792__ & ~new_new_n18798__;
  assign new_new_n18800__ = ~new_new_n18427__ & ~new_new_n18799__;
  assign new_new_n18801__ = ~new_new_n18786__ & ~new_new_n18800__;
  assign new_new_n18802__ = ~ys__n19973 & ~new_new_n18801__;
  assign new_new_n18803__ = ys__n19973 & ys__n19976;
  assign new_new_n18804__ = ~new_new_n18802__ & ~new_new_n18803__;
  assign new_new_n18805__ = ~ys__n352 & ~new_new_n18804__;
  assign new_new_n18806__ = ~ys__n220 & ys__n47029;
  assign new_new_n18807__ = new_new_n18439__ & new_new_n18806__;
  assign new_new_n18808__ = ~ys__n220 & ys__n47077;
  assign new_new_n18809__ = new_new_n18441__ & new_new_n18808__;
  assign new_new_n18810__ = ~ys__n220 & ys__n47013;
  assign new_new_n18811__ = new_new_n18444__ & new_new_n18810__;
  assign new_new_n18812__ = ~new_new_n18809__ & ~new_new_n18811__;
  assign new_new_n18813__ = ~new_new_n18807__ & new_new_n18812__;
  assign new_new_n18814__ = new_new_n18453__ & ~new_new_n18813__;
  assign ys__n19887 = new_new_n18805__ | new_new_n18814__;
  assign new_new_n18816__ = ys__n19844 & ys__n19848;
  assign new_new_n18817__ = new_new_n18116__ & new_new_n18816__;
  assign new_new_n18818__ = ~ys__n23274 & ~new_new_n18136__;
  assign new_new_n18819__ = ys__n23274 & ~new_new_n18148__;
  assign new_new_n18820__ = ~new_new_n18818__ & ~new_new_n18819__;
  assign new_new_n18821__ = ~ys__n23276 & ~new_new_n18820__;
  assign new_new_n18822__ = ~ys__n23274 & ~new_new_n18158__;
  assign new_new_n18823__ = ys__n23274 & ~new_new_n18172__;
  assign new_new_n18824__ = ~new_new_n18822__ & ~new_new_n18823__;
  assign new_new_n18825__ = ys__n23276 & ~new_new_n18824__;
  assign new_new_n18826__ = ~new_new_n18821__ & ~new_new_n18825__;
  assign new_new_n18827__ = ~ys__n23278 & ~new_new_n18826__;
  assign new_new_n18828__ = ~ys__n23274 & ~new_new_n18182__;
  assign new_new_n18829__ = ys__n23274 & ~new_new_n18194__;
  assign new_new_n18830__ = ~new_new_n18828__ & ~new_new_n18829__;
  assign new_new_n18831__ = ~ys__n23276 & ~new_new_n18830__;
  assign new_new_n18832__ = ~ys__n23274 & ~new_new_n18204__;
  assign new_new_n18833__ = ~new_new_n18747__ & ~new_new_n18832__;
  assign new_new_n18834__ = ys__n23276 & ~new_new_n18833__;
  assign new_new_n18835__ = ~new_new_n18831__ & ~new_new_n18834__;
  assign new_new_n18836__ = ys__n23278 & ~new_new_n18835__;
  assign new_new_n18837__ = ~new_new_n18827__ & ~new_new_n18836__;
  assign new_new_n18838__ = ~ys__n1505 & ~new_new_n18837__;
  assign new_new_n18839__ = ys__n23276 & new_new_n18832__;
  assign new_new_n18840__ = ~new_new_n18831__ & ~new_new_n18839__;
  assign new_new_n18841__ = ys__n23278 & ~new_new_n18840__;
  assign new_new_n18842__ = ~new_new_n18827__ & ~new_new_n18841__;
  assign new_new_n18843__ = ys__n1505 & ~new_new_n18842__;
  assign new_new_n18844__ = ~new_new_n18838__ & ~new_new_n18843__;
  assign new_new_n18845__ = ~new_new_n18116__ & ~new_new_n18844__;
  assign new_new_n18846__ = ~new_new_n18817__ & ~new_new_n18845__;
  assign new_new_n18847__ = new_new_n18213__ & ~new_new_n18846__;
  assign new_new_n18848__ = ~new_new_n18123__ & ~new_new_n18128__;
  assign new_new_n18849__ = ~ys__n23272 & ~new_new_n18848__;
  assign new_new_n18850__ = ys__n23272 & ~new_new_n18663__;
  assign new_new_n18851__ = ~new_new_n18849__ & ~new_new_n18850__;
  assign new_new_n18852__ = ~ys__n23274 & ~new_new_n18851__;
  assign new_new_n18853__ = ys__n23274 & new_new_n18215__;
  assign new_new_n18854__ = ~new_new_n18852__ & ~new_new_n18853__;
  assign new_new_n18855__ = ~ys__n23276 & ~new_new_n18854__;
  assign new_new_n18856__ = new_new_n18219__ & new_new_n18855__;
  assign new_new_n18857__ = ~new_new_n18847__ & ~new_new_n18856__;
  assign new_new_n18858__ = new_new_n18224__ & ~new_new_n18857__;
  assign new_new_n18859__ = ~new_new_n10752__ & new_new_n18226__;
  assign new_new_n18860__ = ys__n1498 & new_new_n18268__;
  assign new_new_n18861__ = ~new_new_n18859__ & ~new_new_n18860__;
  assign new_new_n18862__ = ~ys__n1496 & ~new_new_n18861__;
  assign new_new_n18863__ = ys__n1496 & ~new_new_n18268__;
  assign new_new_n18864__ = ~new_new_n18862__ & ~new_new_n18863__;
  assign new_new_n18865__ = ~ys__n1495 & ~new_new_n18864__;
  assign new_new_n18866__ = ys__n1495 & new_new_n16792__;
  assign new_new_n18867__ = ~new_new_n18865__ & ~new_new_n18866__;
  assign new_new_n18868__ = ~new_new_n18224__ & ~new_new_n18867__;
  assign new_new_n18869__ = ~new_new_n18858__ & ~new_new_n18868__;
  assign new_new_n18870__ = new_new_n18581__ & ~new_new_n18869__;
  assign new_new_n18871__ = ~new_new_n18260__ & new_new_n18269__;
  assign new_new_n18872__ = new_new_n18260__ & ~new_new_n18269__;
  assign new_new_n18873__ = ~new_new_n18871__ & ~new_new_n18872__;
  assign new_new_n18874__ = ~ys__n1489 & ~new_new_n18873__;
  assign new_new_n18875__ = new_new_n10752__ & ~new_new_n16786__;
  assign new_new_n18876__ = ~new_new_n10752__ & new_new_n16786__;
  assign new_new_n18877__ = ~new_new_n18875__ & ~new_new_n18876__;
  assign new_new_n18878__ = ys__n1489 & ~new_new_n18877__;
  assign new_new_n18879__ = ~new_new_n18874__ & ~new_new_n18878__;
  assign new_new_n18880__ = ~new_new_n18427__ & ~new_new_n18879__;
  assign new_new_n18881__ = ~new_new_n18870__ & ~new_new_n18880__;
  assign new_new_n18882__ = ~ys__n19973 & ~new_new_n18881__;
  assign new_new_n18883__ = ys__n19973 & ys__n19977;
  assign new_new_n18884__ = ~new_new_n18882__ & ~new_new_n18883__;
  assign new_new_n18885__ = ~ys__n352 & ~new_new_n18884__;
  assign new_new_n18886__ = ~ys__n220 & ys__n47030;
  assign new_new_n18887__ = new_new_n18439__ & new_new_n18886__;
  assign new_new_n18888__ = ~ys__n220 & ys__n47078;
  assign new_new_n18889__ = new_new_n18441__ & new_new_n18888__;
  assign new_new_n18890__ = ~ys__n220 & ys__n47014;
  assign new_new_n18891__ = new_new_n18444__ & new_new_n18890__;
  assign new_new_n18892__ = ~new_new_n18889__ & ~new_new_n18891__;
  assign new_new_n18893__ = ~new_new_n18887__ & new_new_n18892__;
  assign new_new_n18894__ = new_new_n18453__ & ~new_new_n18893__;
  assign ys__n19890 = new_new_n18885__ | new_new_n18894__;
  assign new_new_n18896__ = ys__n19844 & ys__n19849;
  assign new_new_n18897__ = new_new_n18116__ & new_new_n18896__;
  assign new_new_n18898__ = ~ys__n23274 & ~new_new_n18476__;
  assign new_new_n18899__ = ys__n23274 & ~new_new_n18488__;
  assign new_new_n18900__ = ~new_new_n18898__ & ~new_new_n18899__;
  assign new_new_n18901__ = ~ys__n23276 & ~new_new_n18900__;
  assign new_new_n18902__ = ~ys__n23274 & ~new_new_n18498__;
  assign new_new_n18903__ = ys__n23274 & ~new_new_n18512__;
  assign new_new_n18904__ = ~new_new_n18902__ & ~new_new_n18903__;
  assign new_new_n18905__ = ys__n23276 & ~new_new_n18904__;
  assign new_new_n18906__ = ~new_new_n18901__ & ~new_new_n18905__;
  assign new_new_n18907__ = ~ys__n23278 & ~new_new_n18906__;
  assign new_new_n18908__ = ~ys__n23274 & ~new_new_n18522__;
  assign new_new_n18909__ = ys__n23274 & ~new_new_n18534__;
  assign new_new_n18910__ = ~new_new_n18908__ & ~new_new_n18909__;
  assign new_new_n18911__ = ~ys__n23276 & ~new_new_n18910__;
  assign new_new_n18912__ = ~ys__n23274 & ~new_new_n18541__;
  assign new_new_n18913__ = ~new_new_n18747__ & ~new_new_n18912__;
  assign new_new_n18914__ = ys__n23276 & ~new_new_n18913__;
  assign new_new_n18915__ = ~new_new_n18911__ & ~new_new_n18914__;
  assign new_new_n18916__ = ys__n23278 & ~new_new_n18915__;
  assign new_new_n18917__ = ~new_new_n18907__ & ~new_new_n18916__;
  assign new_new_n18918__ = ~ys__n1505 & ~new_new_n18917__;
  assign new_new_n18919__ = ~ys__n23274 & ~new_new_n18551__;
  assign new_new_n18920__ = ys__n23276 & new_new_n18919__;
  assign new_new_n18921__ = ~new_new_n18911__ & ~new_new_n18920__;
  assign new_new_n18922__ = ys__n23278 & ~new_new_n18921__;
  assign new_new_n18923__ = ~new_new_n18907__ & ~new_new_n18922__;
  assign new_new_n18924__ = ys__n1505 & ~new_new_n18923__;
  assign new_new_n18925__ = ~new_new_n18918__ & ~new_new_n18924__;
  assign new_new_n18926__ = ~new_new_n18116__ & ~new_new_n18925__;
  assign new_new_n18927__ = ~new_new_n18897__ & ~new_new_n18926__;
  assign new_new_n18928__ = new_new_n18213__ & ~new_new_n18927__;
  assign new_new_n18929__ = ~new_new_n18463__ & ~new_new_n18468__;
  assign new_new_n18930__ = ~ys__n23272 & ~new_new_n18929__;
  assign new_new_n18931__ = ys__n23272 & ~new_new_n18766__;
  assign new_new_n18932__ = ~new_new_n18930__ & ~new_new_n18931__;
  assign new_new_n18933__ = ~ys__n23274 & ~new_new_n18932__;
  assign new_new_n18934__ = ys__n23274 & new_new_n18564__;
  assign new_new_n18935__ = ~new_new_n18933__ & ~new_new_n18934__;
  assign new_new_n18936__ = ~ys__n23276 & ~new_new_n18935__;
  assign new_new_n18937__ = new_new_n18219__ & new_new_n18936__;
  assign new_new_n18938__ = ~new_new_n18928__ & ~new_new_n18937__;
  assign new_new_n18939__ = new_new_n18224__ & ~new_new_n18938__;
  assign new_new_n18940__ = ~new_new_n10755__ & new_new_n18226__;
  assign new_new_n18941__ = ys__n1498 & new_new_n18266__;
  assign new_new_n18942__ = ~new_new_n18940__ & ~new_new_n18941__;
  assign new_new_n18943__ = ~ys__n1496 & ~new_new_n18942__;
  assign new_new_n18944__ = ys__n1496 & ~new_new_n18266__;
  assign new_new_n18945__ = ~new_new_n18943__ & ~new_new_n18944__;
  assign new_new_n18946__ = ~ys__n1495 & ~new_new_n18945__;
  assign new_new_n18947__ = ys__n1495 & new_new_n16791__;
  assign new_new_n18948__ = ~new_new_n18946__ & ~new_new_n18947__;
  assign new_new_n18949__ = ~new_new_n18224__ & ~new_new_n18948__;
  assign new_new_n18950__ = ~new_new_n18939__ & ~new_new_n18949__;
  assign new_new_n18951__ = new_new_n18581__ & ~new_new_n18950__;
  assign new_new_n18952__ = ~new_new_n18260__ & ~new_new_n18269__;
  assign new_new_n18953__ = ~new_new_n10751__ & ~new_new_n18952__;
  assign new_new_n18954__ = new_new_n18267__ & ~new_new_n18953__;
  assign new_new_n18955__ = ~new_new_n18267__ & new_new_n18953__;
  assign new_new_n18956__ = ~new_new_n18954__ & ~new_new_n18955__;
  assign new_new_n18957__ = ~ys__n1489 & ~new_new_n18956__;
  assign new_new_n18958__ = ~new_new_n10752__ & ~new_new_n16786__;
  assign new_new_n18959__ = ~new_new_n16792__ & ~new_new_n18958__;
  assign new_new_n18960__ = new_new_n10755__ & ~new_new_n18959__;
  assign new_new_n18961__ = ~new_new_n10755__ & new_new_n18959__;
  assign new_new_n18962__ = ~new_new_n18960__ & ~new_new_n18961__;
  assign new_new_n18963__ = ys__n1489 & ~new_new_n18962__;
  assign new_new_n18964__ = ~new_new_n18957__ & ~new_new_n18963__;
  assign new_new_n18965__ = ~new_new_n18427__ & ~new_new_n18964__;
  assign new_new_n18966__ = ~new_new_n18951__ & ~new_new_n18965__;
  assign new_new_n18967__ = ~ys__n19973 & ~new_new_n18966__;
  assign new_new_n18968__ = ys__n19973 & ys__n19978;
  assign new_new_n18969__ = ~new_new_n18967__ & ~new_new_n18968__;
  assign new_new_n18970__ = ~ys__n352 & ~new_new_n18969__;
  assign new_new_n18971__ = ~ys__n220 & ys__n47031;
  assign new_new_n18972__ = new_new_n18439__ & new_new_n18971__;
  assign new_new_n18973__ = ~ys__n220 & ys__n47079;
  assign new_new_n18974__ = new_new_n18441__ & new_new_n18973__;
  assign new_new_n18975__ = ~ys__n220 & ys__n47015;
  assign new_new_n18976__ = new_new_n18444__ & new_new_n18975__;
  assign new_new_n18977__ = ~new_new_n18974__ & ~new_new_n18976__;
  assign new_new_n18978__ = ~new_new_n18972__ & new_new_n18977__;
  assign new_new_n18979__ = new_new_n18453__ & ~new_new_n18978__;
  assign ys__n19893 = new_new_n18970__ | new_new_n18979__;
  assign new_new_n18981__ = ys__n19844 & ys__n19850;
  assign new_new_n18982__ = new_new_n18116__ & new_new_n18981__;
  assign new_new_n18983__ = ~ys__n23274 & ~new_new_n18613__;
  assign new_new_n18984__ = ys__n23274 & ~new_new_n18619__;
  assign new_new_n18985__ = ~new_new_n18983__ & ~new_new_n18984__;
  assign new_new_n18986__ = ~ys__n23276 & ~new_new_n18985__;
  assign new_new_n18987__ = ~ys__n23274 & ~new_new_n18623__;
  assign new_new_n18988__ = ys__n23274 & ~new_new_n18631__;
  assign new_new_n18989__ = ~new_new_n18987__ & ~new_new_n18988__;
  assign new_new_n18990__ = ys__n23276 & ~new_new_n18989__;
  assign new_new_n18991__ = ~new_new_n18986__ & ~new_new_n18990__;
  assign new_new_n18992__ = ~ys__n23278 & ~new_new_n18991__;
  assign new_new_n18993__ = ~ys__n23274 & ~new_new_n18635__;
  assign new_new_n18994__ = ys__n23274 & ~new_new_n18641__;
  assign new_new_n18995__ = ~new_new_n18993__ & ~new_new_n18994__;
  assign new_new_n18996__ = ~ys__n23276 & ~new_new_n18995__;
  assign new_new_n18997__ = ~ys__n23274 & ~new_new_n18644__;
  assign new_new_n18998__ = ~new_new_n18747__ & ~new_new_n18997__;
  assign new_new_n18999__ = ys__n23276 & ~new_new_n18998__;
  assign new_new_n19000__ = ~new_new_n18996__ & ~new_new_n18999__;
  assign new_new_n19001__ = ys__n23278 & ~new_new_n19000__;
  assign new_new_n19002__ = ~new_new_n18992__ & ~new_new_n19001__;
  assign new_new_n19003__ = ~ys__n1505 & ~new_new_n19002__;
  assign new_new_n19004__ = ~ys__n23274 & new_new_n18643__;
  assign new_new_n19005__ = ys__n23276 & new_new_n19004__;
  assign new_new_n19006__ = ~new_new_n18996__ & ~new_new_n19005__;
  assign new_new_n19007__ = ys__n23278 & ~new_new_n19006__;
  assign new_new_n19008__ = ~new_new_n18992__ & ~new_new_n19007__;
  assign new_new_n19009__ = ys__n1505 & ~new_new_n19008__;
  assign new_new_n19010__ = ~new_new_n19003__ & ~new_new_n19009__;
  assign new_new_n19011__ = ~new_new_n18116__ & ~new_new_n19010__;
  assign new_new_n19012__ = ~new_new_n18982__ & ~new_new_n19011__;
  assign new_new_n19013__ = new_new_n18213__ & ~new_new_n19012__;
  assign new_new_n19014__ = ~new_new_n18129__ & ~new_new_n18132__;
  assign new_new_n19015__ = ~ys__n23272 & ~new_new_n19014__;
  assign new_new_n19016__ = ys__n23272 & ~new_new_n18848__;
  assign new_new_n19017__ = ~new_new_n19015__ & ~new_new_n19016__;
  assign new_new_n19018__ = ~ys__n23274 & ~new_new_n19017__;
  assign new_new_n19019__ = ys__n23274 & ~new_new_n18666__;
  assign new_new_n19020__ = ~new_new_n19018__ & ~new_new_n19019__;
  assign new_new_n19021__ = ~ys__n23276 & ~new_new_n19020__;
  assign new_new_n19022__ = new_new_n18219__ & new_new_n19021__;
  assign new_new_n19023__ = ~new_new_n19013__ & ~new_new_n19022__;
  assign new_new_n19024__ = new_new_n18224__ & ~new_new_n19023__;
  assign new_new_n19025__ = ~new_new_n10759__ & new_new_n18226__;
  assign new_new_n19026__ = ys__n1498 & new_new_n18263__;
  assign new_new_n19027__ = ~new_new_n19025__ & ~new_new_n19026__;
  assign new_new_n19028__ = ~ys__n1496 & ~new_new_n19027__;
  assign new_new_n19029__ = ys__n1496 & ~new_new_n18263__;
  assign new_new_n19030__ = ~new_new_n19028__ & ~new_new_n19029__;
  assign new_new_n19031__ = ~ys__n1495 & ~new_new_n19030__;
  assign new_new_n19032__ = ys__n1495 & new_new_n16797__;
  assign new_new_n19033__ = ~new_new_n19031__ & ~new_new_n19032__;
  assign new_new_n19034__ = ~new_new_n18224__ & ~new_new_n19033__;
  assign new_new_n19035__ = ~new_new_n19024__ & ~new_new_n19034__;
  assign new_new_n19036__ = new_new_n18581__ & ~new_new_n19035__;
  assign new_new_n19037__ = ~new_new_n18260__ & new_new_n18270__;
  assign new_new_n19038__ = new_new_n18274__ & ~new_new_n19037__;
  assign new_new_n19039__ = new_new_n18264__ & ~new_new_n19038__;
  assign new_new_n19040__ = ~new_new_n18264__ & new_new_n19038__;
  assign new_new_n19041__ = ~new_new_n19039__ & ~new_new_n19040__;
  assign new_new_n19042__ = ~ys__n1489 & ~new_new_n19041__;
  assign new_new_n19043__ = ~new_new_n16786__ & new_new_n16788__;
  assign new_new_n19044__ = new_new_n16794__ & ~new_new_n19043__;
  assign new_new_n19045__ = new_new_n10759__ & ~new_new_n19044__;
  assign new_new_n19046__ = ~new_new_n10759__ & new_new_n19044__;
  assign new_new_n19047__ = ~new_new_n19045__ & ~new_new_n19046__;
  assign new_new_n19048__ = ys__n1489 & ~new_new_n19047__;
  assign new_new_n19049__ = ~new_new_n19042__ & ~new_new_n19048__;
  assign new_new_n19050__ = ~new_new_n18427__ & ~new_new_n19049__;
  assign new_new_n19051__ = ~new_new_n19036__ & ~new_new_n19050__;
  assign new_new_n19052__ = ~ys__n19973 & ~new_new_n19051__;
  assign new_new_n19053__ = ys__n19973 & ys__n19979;
  assign new_new_n19054__ = ~new_new_n19052__ & ~new_new_n19053__;
  assign new_new_n19055__ = ~ys__n352 & ~new_new_n19054__;
  assign new_new_n19056__ = ~ys__n220 & ys__n47032;
  assign new_new_n19057__ = new_new_n18439__ & new_new_n19056__;
  assign new_new_n19058__ = ~ys__n220 & ys__n47080;
  assign new_new_n19059__ = new_new_n18441__ & new_new_n19058__;
  assign new_new_n19060__ = ~ys__n220 & ys__n47016;
  assign new_new_n19061__ = new_new_n18444__ & new_new_n19060__;
  assign new_new_n19062__ = ~new_new_n19059__ & ~new_new_n19061__;
  assign new_new_n19063__ = ~new_new_n19057__ & new_new_n19062__;
  assign new_new_n19064__ = new_new_n18453__ & ~new_new_n19063__;
  assign ys__n19896 = new_new_n19055__ | new_new_n19064__;
  assign new_new_n19066__ = ys__n19844 & ys__n19851;
  assign new_new_n19067__ = new_new_n18116__ & new_new_n19066__;
  assign new_new_n19068__ = ~ys__n23274 & ~new_new_n18717__;
  assign new_new_n19069__ = ys__n23274 & ~new_new_n18723__;
  assign new_new_n19070__ = ~new_new_n19068__ & ~new_new_n19069__;
  assign new_new_n19071__ = ~ys__n23276 & ~new_new_n19070__;
  assign new_new_n19072__ = ~ys__n23274 & ~new_new_n18727__;
  assign new_new_n19073__ = ys__n23274 & ~new_new_n18735__;
  assign new_new_n19074__ = ~new_new_n19072__ & ~new_new_n19073__;
  assign new_new_n19075__ = ys__n23276 & ~new_new_n19074__;
  assign new_new_n19076__ = ~new_new_n19071__ & ~new_new_n19075__;
  assign new_new_n19077__ = ~ys__n23278 & ~new_new_n19076__;
  assign new_new_n19078__ = ~ys__n23274 & ~new_new_n18739__;
  assign new_new_n19079__ = ys__n23274 & ~new_new_n18745__;
  assign new_new_n19080__ = ~new_new_n19078__ & ~new_new_n19079__;
  assign new_new_n19081__ = ~ys__n23276 & ~new_new_n19080__;
  assign new_new_n19082__ = ys__n23276 & ys__n28030;
  assign new_new_n19083__ = ~new_new_n19081__ & ~new_new_n19082__;
  assign new_new_n19084__ = ys__n23278 & ~new_new_n19083__;
  assign new_new_n19085__ = ~new_new_n19077__ & ~new_new_n19084__;
  assign new_new_n19086__ = ~ys__n1505 & ~new_new_n19085__;
  assign new_new_n19087__ = ~ys__n23274 & new_new_n18754__;
  assign new_new_n19088__ = ys__n23276 & new_new_n19087__;
  assign new_new_n19089__ = ~new_new_n19081__ & ~new_new_n19088__;
  assign new_new_n19090__ = ys__n23278 & ~new_new_n19089__;
  assign new_new_n19091__ = ~new_new_n19077__ & ~new_new_n19090__;
  assign new_new_n19092__ = ys__n1505 & ~new_new_n19091__;
  assign new_new_n19093__ = ~new_new_n19086__ & ~new_new_n19092__;
  assign new_new_n19094__ = ~new_new_n18116__ & ~new_new_n19093__;
  assign new_new_n19095__ = ~new_new_n19067__ & ~new_new_n19094__;
  assign new_new_n19096__ = new_new_n18213__ & ~new_new_n19095__;
  assign new_new_n19097__ = ~new_new_n18469__ & ~new_new_n18472__;
  assign new_new_n19098__ = ~ys__n23272 & ~new_new_n19097__;
  assign new_new_n19099__ = ys__n23272 & ~new_new_n18929__;
  assign new_new_n19100__ = ~new_new_n19098__ & ~new_new_n19099__;
  assign new_new_n19101__ = ~ys__n23274 & ~new_new_n19100__;
  assign new_new_n19102__ = ys__n23274 & ~new_new_n18769__;
  assign new_new_n19103__ = ~new_new_n19101__ & ~new_new_n19102__;
  assign new_new_n19104__ = ~ys__n23276 & ~new_new_n19103__;
  assign new_new_n19105__ = new_new_n18219__ & new_new_n19104__;
  assign new_new_n19106__ = ~new_new_n19096__ & ~new_new_n19105__;
  assign new_new_n19107__ = new_new_n18224__ & ~new_new_n19106__;
  assign new_new_n19108__ = ~new_new_n10762__ & new_new_n18226__;
  assign new_new_n19109__ = ys__n1498 & new_new_n18261__;
  assign new_new_n19110__ = ~new_new_n19108__ & ~new_new_n19109__;
  assign new_new_n19111__ = ~ys__n1496 & ~new_new_n19110__;
  assign new_new_n19112__ = ys__n1496 & ~new_new_n18261__;
  assign new_new_n19113__ = ~new_new_n19111__ & ~new_new_n19112__;
  assign new_new_n19114__ = ~ys__n1495 & ~new_new_n19113__;
  assign new_new_n19115__ = ys__n1495 & new_new_n16796__;
  assign new_new_n19116__ = ~new_new_n19114__ & ~new_new_n19115__;
  assign new_new_n19117__ = ~new_new_n18224__ & ~new_new_n19116__;
  assign new_new_n19118__ = ~new_new_n19107__ & ~new_new_n19117__;
  assign new_new_n19119__ = new_new_n18581__ & ~new_new_n19118__;
  assign new_new_n19120__ = ~new_new_n18264__ & ~new_new_n19038__;
  assign new_new_n19121__ = ~new_new_n10758__ & ~new_new_n19120__;
  assign new_new_n19122__ = new_new_n18262__ & ~new_new_n19121__;
  assign new_new_n19123__ = ~new_new_n18262__ & new_new_n19121__;
  assign new_new_n19124__ = ~new_new_n19122__ & ~new_new_n19123__;
  assign new_new_n19125__ = ~ys__n1489 & ~new_new_n19124__;
  assign new_new_n19126__ = ~new_new_n10759__ & ~new_new_n19044__;
  assign new_new_n19127__ = ~new_new_n16797__ & ~new_new_n19126__;
  assign new_new_n19128__ = new_new_n10762__ & ~new_new_n19127__;
  assign new_new_n19129__ = ~new_new_n10762__ & new_new_n19127__;
  assign new_new_n19130__ = ~new_new_n19128__ & ~new_new_n19129__;
  assign new_new_n19131__ = ys__n1489 & ~new_new_n19130__;
  assign new_new_n19132__ = ~new_new_n19125__ & ~new_new_n19131__;
  assign new_new_n19133__ = ~new_new_n18427__ & ~new_new_n19132__;
  assign new_new_n19134__ = ~new_new_n19119__ & ~new_new_n19133__;
  assign new_new_n19135__ = ~ys__n19973 & ~new_new_n19134__;
  assign new_new_n19136__ = ys__n19973 & ys__n19980;
  assign new_new_n19137__ = ~new_new_n19135__ & ~new_new_n19136__;
  assign new_new_n19138__ = ~ys__n352 & ~new_new_n19137__;
  assign new_new_n19139__ = ~ys__n220 & ys__n47033;
  assign new_new_n19140__ = new_new_n18439__ & new_new_n19139__;
  assign new_new_n19141__ = ~ys__n220 & ys__n47081;
  assign new_new_n19142__ = new_new_n18441__ & new_new_n19141__;
  assign new_new_n19143__ = ~ys__n220 & ys__n47017;
  assign new_new_n19144__ = new_new_n18444__ & new_new_n19143__;
  assign new_new_n19145__ = ~new_new_n19142__ & ~new_new_n19144__;
  assign new_new_n19146__ = ~new_new_n19140__ & new_new_n19145__;
  assign new_new_n19147__ = new_new_n18453__ & ~new_new_n19146__;
  assign ys__n19899 = new_new_n19138__ | new_new_n19147__;
  assign new_new_n19149__ = ys__n19844 & ys__n19852;
  assign new_new_n19150__ = new_new_n18116__ & new_new_n19149__;
  assign new_new_n19151__ = ~ys__n23276 & ~new_new_n18160__;
  assign new_new_n19152__ = ys__n23276 & ~new_new_n18184__;
  assign new_new_n19153__ = ~new_new_n19151__ & ~new_new_n19152__;
  assign new_new_n19154__ = ~ys__n23278 & ~new_new_n19153__;
  assign new_new_n19155__ = ~ys__n23276 & ~new_new_n18206__;
  assign new_new_n19156__ = ~new_new_n19082__ & ~new_new_n19155__;
  assign new_new_n19157__ = ys__n23278 & ~new_new_n19156__;
  assign new_new_n19158__ = ~new_new_n19154__ & ~new_new_n19157__;
  assign new_new_n19159__ = ~ys__n1505 & ~new_new_n19158__;
  assign new_new_n19160__ = ys__n23278 & new_new_n19155__;
  assign new_new_n19161__ = ~new_new_n19154__ & ~new_new_n19160__;
  assign new_new_n19162__ = ys__n1505 & ~new_new_n19161__;
  assign new_new_n19163__ = ~new_new_n19159__ & ~new_new_n19162__;
  assign new_new_n19164__ = ~new_new_n18116__ & ~new_new_n19163__;
  assign new_new_n19165__ = ~new_new_n19150__ & ~new_new_n19164__;
  assign new_new_n19166__ = new_new_n18213__ & ~new_new_n19165__;
  assign new_new_n19167__ = ~new_new_n18133__ & ~new_new_n18140__;
  assign new_new_n19168__ = ~ys__n23272 & ~new_new_n19167__;
  assign new_new_n19169__ = ys__n23272 & ~new_new_n19014__;
  assign new_new_n19170__ = ~new_new_n19168__ & ~new_new_n19169__;
  assign new_new_n19171__ = ~ys__n23274 & ~new_new_n19170__;
  assign new_new_n19172__ = ys__n23274 & ~new_new_n18851__;
  assign new_new_n19173__ = ~new_new_n19171__ & ~new_new_n19172__;
  assign new_new_n19174__ = ~ys__n23276 & ~new_new_n19173__;
  assign new_new_n19175__ = ys__n23276 & new_new_n18216__;
  assign new_new_n19176__ = ~new_new_n19174__ & ~new_new_n19175__;
  assign new_new_n19177__ = new_new_n18219__ & ~new_new_n19176__;
  assign new_new_n19178__ = ~new_new_n19166__ & ~new_new_n19177__;
  assign new_new_n19179__ = new_new_n18224__ & ~new_new_n19178__;
  assign new_new_n19180__ = ~new_new_n10798__ & new_new_n18226__;
  assign new_new_n19181__ = ys__n1498 & new_new_n18298__;
  assign new_new_n19182__ = ~new_new_n19180__ & ~new_new_n19181__;
  assign new_new_n19183__ = ~ys__n1496 & ~new_new_n19182__;
  assign new_new_n19184__ = ys__n1496 & ~new_new_n18298__;
  assign new_new_n19185__ = ~new_new_n19183__ & ~new_new_n19184__;
  assign new_new_n19186__ = ~ys__n1495 & ~new_new_n19185__;
  assign new_new_n19187__ = ys__n1495 & new_new_n16811__;
  assign new_new_n19188__ = ~new_new_n19186__ & ~new_new_n19187__;
  assign new_new_n19189__ = ~new_new_n18224__ & ~new_new_n19188__;
  assign new_new_n19190__ = ~new_new_n19179__ & ~new_new_n19189__;
  assign new_new_n19191__ = new_new_n18581__ & ~new_new_n19190__;
  assign new_new_n19192__ = ~new_new_n18279__ & new_new_n18299__;
  assign new_new_n19193__ = new_new_n18279__ & ~new_new_n18299__;
  assign new_new_n19194__ = ~new_new_n19192__ & ~new_new_n19193__;
  assign new_new_n19195__ = ~ys__n1489 & ~new_new_n19194__;
  assign new_new_n19196__ = new_new_n10798__ & ~new_new_n16801__;
  assign new_new_n19197__ = ~new_new_n10798__ & new_new_n16801__;
  assign new_new_n19198__ = ~new_new_n19196__ & ~new_new_n19197__;
  assign new_new_n19199__ = ys__n1489 & ~new_new_n19198__;
  assign new_new_n19200__ = ~new_new_n19195__ & ~new_new_n19199__;
  assign new_new_n19201__ = ~new_new_n18427__ & ~new_new_n19200__;
  assign new_new_n19202__ = ~new_new_n19191__ & ~new_new_n19201__;
  assign new_new_n19203__ = ~ys__n19973 & ~new_new_n19202__;
  assign new_new_n19204__ = ys__n19973 & ys__n19981;
  assign new_new_n19205__ = ~new_new_n19203__ & ~new_new_n19204__;
  assign new_new_n19206__ = ~ys__n352 & ~new_new_n19205__;
  assign new_new_n19207__ = ~ys__n220 & ys__n47034;
  assign new_new_n19208__ = new_new_n18439__ & new_new_n19207__;
  assign new_new_n19209__ = ~ys__n220 & ys__n47082;
  assign new_new_n19210__ = new_new_n18441__ & new_new_n19209__;
  assign new_new_n19211__ = ~ys__n220 & ys__n47018;
  assign new_new_n19212__ = new_new_n18444__ & new_new_n19211__;
  assign new_new_n19213__ = ~new_new_n19210__ & ~new_new_n19212__;
  assign new_new_n19214__ = ~new_new_n19208__ & new_new_n19213__;
  assign new_new_n19215__ = new_new_n18453__ & ~new_new_n19214__;
  assign ys__n19902 = new_new_n19206__ | new_new_n19215__;
  assign new_new_n19217__ = ys__n19844 & ys__n19853;
  assign new_new_n19218__ = new_new_n18116__ & new_new_n19217__;
  assign new_new_n19219__ = ~ys__n23276 & ~new_new_n18500__;
  assign new_new_n19220__ = ys__n23276 & ~new_new_n18524__;
  assign new_new_n19221__ = ~new_new_n19219__ & ~new_new_n19220__;
  assign new_new_n19222__ = ~ys__n23278 & ~new_new_n19221__;
  assign new_new_n19223__ = ~ys__n23276 & ~new_new_n18543__;
  assign new_new_n19224__ = ~new_new_n19082__ & ~new_new_n19223__;
  assign new_new_n19225__ = ys__n23278 & ~new_new_n19224__;
  assign new_new_n19226__ = ~new_new_n19222__ & ~new_new_n19225__;
  assign new_new_n19227__ = ~ys__n1505 & ~new_new_n19226__;
  assign new_new_n19228__ = ~ys__n23276 & ~new_new_n18553__;
  assign new_new_n19229__ = ys__n23278 & new_new_n19228__;
  assign new_new_n19230__ = ~new_new_n19222__ & ~new_new_n19229__;
  assign new_new_n19231__ = ys__n1505 & ~new_new_n19230__;
  assign new_new_n19232__ = ~new_new_n19227__ & ~new_new_n19231__;
  assign new_new_n19233__ = ~new_new_n18116__ & ~new_new_n19232__;
  assign new_new_n19234__ = ~new_new_n19218__ & ~new_new_n19233__;
  assign new_new_n19235__ = new_new_n18213__ & ~new_new_n19234__;
  assign new_new_n19236__ = ~new_new_n18473__ & ~new_new_n18480__;
  assign new_new_n19237__ = ~ys__n23272 & ~new_new_n19236__;
  assign new_new_n19238__ = ys__n23272 & ~new_new_n19097__;
  assign new_new_n19239__ = ~new_new_n19237__ & ~new_new_n19238__;
  assign new_new_n19240__ = ~ys__n23274 & ~new_new_n19239__;
  assign new_new_n19241__ = ys__n23274 & ~new_new_n18932__;
  assign new_new_n19242__ = ~new_new_n19240__ & ~new_new_n19241__;
  assign new_new_n19243__ = ~ys__n23276 & ~new_new_n19242__;
  assign new_new_n19244__ = ys__n23276 & new_new_n18565__;
  assign new_new_n19245__ = ~new_new_n19243__ & ~new_new_n19244__;
  assign new_new_n19246__ = new_new_n18219__ & ~new_new_n19245__;
  assign new_new_n19247__ = ~new_new_n19235__ & ~new_new_n19246__;
  assign new_new_n19248__ = new_new_n18224__ & ~new_new_n19247__;
  assign new_new_n19249__ = ~new_new_n10801__ & new_new_n18226__;
  assign new_new_n19250__ = ys__n1498 & new_new_n18296__;
  assign new_new_n19251__ = ~new_new_n19249__ & ~new_new_n19250__;
  assign new_new_n19252__ = ~ys__n1496 & ~new_new_n19251__;
  assign new_new_n19253__ = ys__n1496 & ~new_new_n18296__;
  assign new_new_n19254__ = ~new_new_n19252__ & ~new_new_n19253__;
  assign new_new_n19255__ = ~ys__n1495 & ~new_new_n19254__;
  assign new_new_n19256__ = ys__n1495 & new_new_n16810__;
  assign new_new_n19257__ = ~new_new_n19255__ & ~new_new_n19256__;
  assign new_new_n19258__ = ~new_new_n18224__ & ~new_new_n19257__;
  assign new_new_n19259__ = ~new_new_n19248__ & ~new_new_n19258__;
  assign new_new_n19260__ = new_new_n18581__ & ~new_new_n19259__;
  assign new_new_n19261__ = ~new_new_n18279__ & ~new_new_n18299__;
  assign new_new_n19262__ = ~new_new_n10797__ & ~new_new_n19261__;
  assign new_new_n19263__ = new_new_n18297__ & ~new_new_n19262__;
  assign new_new_n19264__ = ~new_new_n18297__ & new_new_n19262__;
  assign new_new_n19265__ = ~new_new_n19263__ & ~new_new_n19264__;
  assign new_new_n19266__ = ~ys__n1489 & ~new_new_n19265__;
  assign new_new_n19267__ = ~new_new_n10798__ & ~new_new_n16801__;
  assign new_new_n19268__ = ~new_new_n16811__ & ~new_new_n19267__;
  assign new_new_n19269__ = new_new_n10801__ & ~new_new_n19268__;
  assign new_new_n19270__ = ~new_new_n10801__ & new_new_n19268__;
  assign new_new_n19271__ = ~new_new_n19269__ & ~new_new_n19270__;
  assign new_new_n19272__ = ys__n1489 & ~new_new_n19271__;
  assign new_new_n19273__ = ~new_new_n19266__ & ~new_new_n19272__;
  assign new_new_n19274__ = ~new_new_n18427__ & ~new_new_n19273__;
  assign new_new_n19275__ = ~new_new_n19260__ & ~new_new_n19274__;
  assign new_new_n19276__ = ~ys__n19973 & ~new_new_n19275__;
  assign new_new_n19277__ = ys__n19973 & ys__n19982;
  assign new_new_n19278__ = ~new_new_n19276__ & ~new_new_n19277__;
  assign new_new_n19279__ = ~ys__n352 & ~new_new_n19278__;
  assign new_new_n19280__ = ~ys__n220 & ys__n47035;
  assign new_new_n19281__ = new_new_n18439__ & new_new_n19280__;
  assign new_new_n19282__ = ~ys__n220 & ys__n47083;
  assign new_new_n19283__ = new_new_n18441__ & new_new_n19282__;
  assign new_new_n19284__ = ~ys__n220 & ys__n47019;
  assign new_new_n19285__ = new_new_n18444__ & new_new_n19284__;
  assign new_new_n19286__ = ~new_new_n19283__ & ~new_new_n19285__;
  assign new_new_n19287__ = ~new_new_n19281__ & new_new_n19286__;
  assign new_new_n19288__ = new_new_n18453__ & ~new_new_n19287__;
  assign ys__n19905 = new_new_n19279__ | new_new_n19288__;
  assign new_new_n19290__ = ys__n19844 & ys__n19854;
  assign new_new_n19291__ = new_new_n18116__ & new_new_n19290__;
  assign new_new_n19292__ = ~ys__n23276 & ~new_new_n18625__;
  assign new_new_n19293__ = ys__n23276 & ~new_new_n18637__;
  assign new_new_n19294__ = ~new_new_n19292__ & ~new_new_n19293__;
  assign new_new_n19295__ = ~ys__n23278 & ~new_new_n19294__;
  assign new_new_n19296__ = ~ys__n23276 & ~new_new_n18646__;
  assign new_new_n19297__ = ~new_new_n19082__ & ~new_new_n19296__;
  assign new_new_n19298__ = ys__n23278 & ~new_new_n19297__;
  assign new_new_n19299__ = ~new_new_n19295__ & ~new_new_n19298__;
  assign new_new_n19300__ = ~ys__n1505 & ~new_new_n19299__;
  assign new_new_n19301__ = ~ys__n23276 & ~new_new_n18653__;
  assign new_new_n19302__ = ys__n23278 & new_new_n19301__;
  assign new_new_n19303__ = ~new_new_n19295__ & ~new_new_n19302__;
  assign new_new_n19304__ = ys__n1505 & ~new_new_n19303__;
  assign new_new_n19305__ = ~new_new_n19300__ & ~new_new_n19304__;
  assign new_new_n19306__ = ~new_new_n18116__ & ~new_new_n19305__;
  assign new_new_n19307__ = ~new_new_n19291__ & ~new_new_n19306__;
  assign new_new_n19308__ = new_new_n18213__ & ~new_new_n19307__;
  assign new_new_n19309__ = ~new_new_n18141__ & ~new_new_n18144__;
  assign new_new_n19310__ = ~ys__n23272 & ~new_new_n19309__;
  assign new_new_n19311__ = ys__n23272 & ~new_new_n19167__;
  assign new_new_n19312__ = ~new_new_n19310__ & ~new_new_n19311__;
  assign new_new_n19313__ = ~ys__n23274 & ~new_new_n19312__;
  assign new_new_n19314__ = ys__n23274 & ~new_new_n19017__;
  assign new_new_n19315__ = ~new_new_n19313__ & ~new_new_n19314__;
  assign new_new_n19316__ = ~ys__n23276 & ~new_new_n19315__;
  assign new_new_n19317__ = ys__n23276 & new_new_n18667__;
  assign new_new_n19318__ = ~new_new_n19316__ & ~new_new_n19317__;
  assign new_new_n19319__ = new_new_n18219__ & ~new_new_n19318__;
  assign new_new_n19320__ = ~new_new_n19308__ & ~new_new_n19319__;
  assign new_new_n19321__ = new_new_n18224__ & ~new_new_n19320__;
  assign new_new_n19322__ = ~new_new_n10805__ & new_new_n18226__;
  assign new_new_n19323__ = ys__n1498 & new_new_n18293__;
  assign new_new_n19324__ = ~new_new_n19322__ & ~new_new_n19323__;
  assign new_new_n19325__ = ~ys__n1496 & ~new_new_n19324__;
  assign new_new_n19326__ = ys__n1496 & ~new_new_n18293__;
  assign new_new_n19327__ = ~new_new_n19325__ & ~new_new_n19326__;
  assign new_new_n19328__ = ~ys__n1495 & ~new_new_n19327__;
  assign new_new_n19329__ = ys__n1495 & new_new_n16816__;
  assign new_new_n19330__ = ~new_new_n19328__ & ~new_new_n19329__;
  assign new_new_n19331__ = ~new_new_n18224__ & ~new_new_n19330__;
  assign new_new_n19332__ = ~new_new_n19321__ & ~new_new_n19331__;
  assign new_new_n19333__ = new_new_n18581__ & ~new_new_n19332__;
  assign new_new_n19334__ = ~new_new_n18279__ & new_new_n18300__;
  assign new_new_n19335__ = new_new_n18305__ & ~new_new_n19334__;
  assign new_new_n19336__ = new_new_n18294__ & ~new_new_n19335__;
  assign new_new_n19337__ = ~new_new_n18294__ & new_new_n19335__;
  assign new_new_n19338__ = ~new_new_n19336__ & ~new_new_n19337__;
  assign new_new_n19339__ = ~ys__n1489 & ~new_new_n19338__;
  assign new_new_n19340__ = ~new_new_n16801__ & new_new_n16806__;
  assign new_new_n19341__ = new_new_n16813__ & ~new_new_n19340__;
  assign new_new_n19342__ = new_new_n10805__ & ~new_new_n19341__;
  assign new_new_n19343__ = ~new_new_n10805__ & new_new_n19341__;
  assign new_new_n19344__ = ~new_new_n19342__ & ~new_new_n19343__;
  assign new_new_n19345__ = ys__n1489 & ~new_new_n19344__;
  assign new_new_n19346__ = ~new_new_n19339__ & ~new_new_n19345__;
  assign new_new_n19347__ = ~new_new_n18427__ & ~new_new_n19346__;
  assign new_new_n19348__ = ~new_new_n19333__ & ~new_new_n19347__;
  assign new_new_n19349__ = ~ys__n19973 & ~new_new_n19348__;
  assign new_new_n19350__ = ys__n19973 & ys__n19983;
  assign new_new_n19351__ = ~new_new_n19349__ & ~new_new_n19350__;
  assign new_new_n19352__ = ~ys__n352 & ~new_new_n19351__;
  assign new_new_n19353__ = ~ys__n220 & ys__n47036;
  assign new_new_n19354__ = new_new_n18439__ & new_new_n19353__;
  assign new_new_n19355__ = ~ys__n220 & ys__n47084;
  assign new_new_n19356__ = new_new_n18441__ & new_new_n19355__;
  assign new_new_n19357__ = ~ys__n220 & ys__n47020;
  assign new_new_n19358__ = new_new_n18444__ & new_new_n19357__;
  assign new_new_n19359__ = ~new_new_n19356__ & ~new_new_n19358__;
  assign new_new_n19360__ = ~new_new_n19354__ & new_new_n19359__;
  assign new_new_n19361__ = new_new_n18453__ & ~new_new_n19360__;
  assign ys__n19908 = new_new_n19352__ | new_new_n19361__;
  assign new_new_n19363__ = ys__n19844 & ys__n19855;
  assign new_new_n19364__ = new_new_n18116__ & new_new_n19363__;
  assign new_new_n19365__ = ~ys__n23276 & ~new_new_n18729__;
  assign new_new_n19366__ = ys__n23276 & ~new_new_n18741__;
  assign new_new_n19367__ = ~new_new_n19365__ & ~new_new_n19366__;
  assign new_new_n19368__ = ~ys__n23278 & ~new_new_n19367__;
  assign new_new_n19369__ = ~ys__n23276 & ~new_new_n18748__;
  assign new_new_n19370__ = ~new_new_n19082__ & ~new_new_n19369__;
  assign new_new_n19371__ = ys__n23278 & ~new_new_n19370__;
  assign new_new_n19372__ = ~new_new_n19368__ & ~new_new_n19371__;
  assign new_new_n19373__ = ~ys__n1505 & ~new_new_n19372__;
  assign new_new_n19374__ = ~ys__n23276 & ~new_new_n18756__;
  assign new_new_n19375__ = ys__n23278 & new_new_n19374__;
  assign new_new_n19376__ = ~new_new_n19368__ & ~new_new_n19375__;
  assign new_new_n19377__ = ys__n1505 & ~new_new_n19376__;
  assign new_new_n19378__ = ~new_new_n19373__ & ~new_new_n19377__;
  assign new_new_n19379__ = ~new_new_n18116__ & ~new_new_n19378__;
  assign new_new_n19380__ = ~new_new_n19364__ & ~new_new_n19379__;
  assign new_new_n19381__ = new_new_n18213__ & ~new_new_n19380__;
  assign new_new_n19382__ = ~new_new_n18481__ & ~new_new_n18484__;
  assign new_new_n19383__ = ~ys__n23272 & ~new_new_n19382__;
  assign new_new_n19384__ = ys__n23272 & ~new_new_n19236__;
  assign new_new_n19385__ = ~new_new_n19383__ & ~new_new_n19384__;
  assign new_new_n19386__ = ~ys__n23274 & ~new_new_n19385__;
  assign new_new_n19387__ = ys__n23274 & ~new_new_n19100__;
  assign new_new_n19388__ = ~new_new_n19386__ & ~new_new_n19387__;
  assign new_new_n19389__ = ~ys__n23276 & ~new_new_n19388__;
  assign new_new_n19390__ = ys__n23276 & new_new_n18770__;
  assign new_new_n19391__ = ~new_new_n19389__ & ~new_new_n19390__;
  assign new_new_n19392__ = new_new_n18219__ & ~new_new_n19391__;
  assign new_new_n19393__ = ~new_new_n19381__ & ~new_new_n19392__;
  assign new_new_n19394__ = new_new_n18224__ & ~new_new_n19393__;
  assign new_new_n19395__ = ~new_new_n10808__ & new_new_n18226__;
  assign new_new_n19396__ = ys__n1498 & new_new_n18291__;
  assign new_new_n19397__ = ~new_new_n19395__ & ~new_new_n19396__;
  assign new_new_n19398__ = ~ys__n1496 & ~new_new_n19397__;
  assign new_new_n19399__ = ys__n1496 & ~new_new_n18291__;
  assign new_new_n19400__ = ~new_new_n19398__ & ~new_new_n19399__;
  assign new_new_n19401__ = ~ys__n1495 & ~new_new_n19400__;
  assign new_new_n19402__ = ys__n1495 & new_new_n16815__;
  assign new_new_n19403__ = ~new_new_n19401__ & ~new_new_n19402__;
  assign new_new_n19404__ = ~new_new_n18224__ & ~new_new_n19403__;
  assign new_new_n19405__ = ~new_new_n19394__ & ~new_new_n19404__;
  assign new_new_n19406__ = new_new_n18581__ & ~new_new_n19405__;
  assign new_new_n19407__ = ~new_new_n18294__ & ~new_new_n19335__;
  assign new_new_n19408__ = ~new_new_n10804__ & ~new_new_n19407__;
  assign new_new_n19409__ = new_new_n18292__ & ~new_new_n19408__;
  assign new_new_n19410__ = ~new_new_n18292__ & new_new_n19408__;
  assign new_new_n19411__ = ~new_new_n19409__ & ~new_new_n19410__;
  assign new_new_n19412__ = ~ys__n1489 & ~new_new_n19411__;
  assign new_new_n19413__ = ~new_new_n10805__ & ~new_new_n19341__;
  assign new_new_n19414__ = ~new_new_n16816__ & ~new_new_n19413__;
  assign new_new_n19415__ = new_new_n10808__ & ~new_new_n19414__;
  assign new_new_n19416__ = ~new_new_n10808__ & new_new_n19414__;
  assign new_new_n19417__ = ~new_new_n19415__ & ~new_new_n19416__;
  assign new_new_n19418__ = ys__n1489 & ~new_new_n19417__;
  assign new_new_n19419__ = ~new_new_n19412__ & ~new_new_n19418__;
  assign new_new_n19420__ = ~new_new_n18427__ & ~new_new_n19419__;
  assign new_new_n19421__ = ~new_new_n19406__ & ~new_new_n19420__;
  assign new_new_n19422__ = ~ys__n19973 & ~new_new_n19421__;
  assign new_new_n19423__ = ys__n19973 & ys__n19984;
  assign new_new_n19424__ = ~new_new_n19422__ & ~new_new_n19423__;
  assign new_new_n19425__ = ~ys__n352 & ~new_new_n19424__;
  assign new_new_n19426__ = ~ys__n220 & ys__n47037;
  assign new_new_n19427__ = new_new_n18439__ & new_new_n19426__;
  assign new_new_n19428__ = ~ys__n220 & ys__n47085;
  assign new_new_n19429__ = new_new_n18441__ & new_new_n19428__;
  assign new_new_n19430__ = ~ys__n220 & ys__n47021;
  assign new_new_n19431__ = new_new_n18444__ & new_new_n19430__;
  assign new_new_n19432__ = ~new_new_n19429__ & ~new_new_n19431__;
  assign new_new_n19433__ = ~new_new_n19427__ & new_new_n19432__;
  assign new_new_n19434__ = new_new_n18453__ & ~new_new_n19433__;
  assign ys__n19911 = new_new_n19425__ | new_new_n19434__;
  assign new_new_n19436__ = ys__n19844 & ys__n19856;
  assign new_new_n19437__ = new_new_n18116__ & new_new_n19436__;
  assign new_new_n19438__ = ~ys__n23276 & ~new_new_n18824__;
  assign new_new_n19439__ = ys__n23276 & ~new_new_n18830__;
  assign new_new_n19440__ = ~new_new_n19438__ & ~new_new_n19439__;
  assign new_new_n19441__ = ~ys__n23278 & ~new_new_n19440__;
  assign new_new_n19442__ = ~ys__n23276 & ~new_new_n18833__;
  assign new_new_n19443__ = ~new_new_n19082__ & ~new_new_n19442__;
  assign new_new_n19444__ = ys__n23278 & ~new_new_n19443__;
  assign new_new_n19445__ = ~new_new_n19441__ & ~new_new_n19444__;
  assign new_new_n19446__ = ~ys__n1505 & ~new_new_n19445__;
  assign new_new_n19447__ = ~ys__n23276 & new_new_n18832__;
  assign new_new_n19448__ = ys__n23278 & new_new_n19447__;
  assign new_new_n19449__ = ~new_new_n19441__ & ~new_new_n19448__;
  assign new_new_n19450__ = ys__n1505 & ~new_new_n19449__;
  assign new_new_n19451__ = ~new_new_n19446__ & ~new_new_n19450__;
  assign new_new_n19452__ = ~new_new_n18116__ & ~new_new_n19451__;
  assign new_new_n19453__ = ~new_new_n19437__ & ~new_new_n19452__;
  assign new_new_n19454__ = new_new_n18213__ & ~new_new_n19453__;
  assign new_new_n19455__ = ~new_new_n18145__ & ~new_new_n18150__;
  assign new_new_n19456__ = ~ys__n23272 & ~new_new_n19455__;
  assign new_new_n19457__ = ys__n23272 & ~new_new_n19309__;
  assign new_new_n19458__ = ~new_new_n19456__ & ~new_new_n19457__;
  assign new_new_n19459__ = ~ys__n23274 & ~new_new_n19458__;
  assign new_new_n19460__ = ys__n23274 & ~new_new_n19170__;
  assign new_new_n19461__ = ~new_new_n19459__ & ~new_new_n19460__;
  assign new_new_n19462__ = ~ys__n23276 & ~new_new_n19461__;
  assign new_new_n19463__ = ys__n23276 & ~new_new_n18854__;
  assign new_new_n19464__ = ~new_new_n19462__ & ~new_new_n19463__;
  assign new_new_n19465__ = new_new_n18219__ & ~new_new_n19464__;
  assign new_new_n19466__ = ~new_new_n19454__ & ~new_new_n19465__;
  assign new_new_n19467__ = new_new_n18224__ & ~new_new_n19466__;
  assign new_new_n19468__ = ~new_new_n10783__ & new_new_n18226__;
  assign new_new_n19469__ = ys__n1498 & new_new_n18287__;
  assign new_new_n19470__ = ~new_new_n19468__ & ~new_new_n19469__;
  assign new_new_n19471__ = ~ys__n1496 & ~new_new_n19470__;
  assign new_new_n19472__ = ys__n1496 & ~new_new_n18287__;
  assign new_new_n19473__ = ~new_new_n19471__ & ~new_new_n19472__;
  assign new_new_n19474__ = ~ys__n1495 & ~new_new_n19473__;
  assign new_new_n19475__ = ys__n1495 & new_new_n16822__;
  assign new_new_n19476__ = ~new_new_n19474__ & ~new_new_n19475__;
  assign new_new_n19477__ = ~new_new_n18224__ & ~new_new_n19476__;
  assign new_new_n19478__ = ~new_new_n19467__ & ~new_new_n19477__;
  assign new_new_n19479__ = new_new_n18581__ & ~new_new_n19478__;
  assign new_new_n19480__ = ~new_new_n18279__ & new_new_n18301__;
  assign new_new_n19481__ = new_new_n18309__ & ~new_new_n19480__;
  assign new_new_n19482__ = new_new_n18288__ & ~new_new_n19481__;
  assign new_new_n19483__ = ~new_new_n18288__ & new_new_n19481__;
  assign new_new_n19484__ = ~new_new_n19482__ & ~new_new_n19483__;
  assign new_new_n19485__ = ~ys__n1489 & ~new_new_n19484__;
  assign new_new_n19486__ = ~new_new_n16801__ & new_new_n16807__;
  assign new_new_n19487__ = new_new_n16819__ & ~new_new_n19486__;
  assign new_new_n19488__ = new_new_n10783__ & ~new_new_n19487__;
  assign new_new_n19489__ = ~new_new_n10783__ & new_new_n19487__;
  assign new_new_n19490__ = ~new_new_n19488__ & ~new_new_n19489__;
  assign new_new_n19491__ = ys__n1489 & ~new_new_n19490__;
  assign new_new_n19492__ = ~new_new_n19485__ & ~new_new_n19491__;
  assign new_new_n19493__ = ~new_new_n18427__ & ~new_new_n19492__;
  assign new_new_n19494__ = ~new_new_n19479__ & ~new_new_n19493__;
  assign new_new_n19495__ = ~ys__n19973 & ~new_new_n19494__;
  assign new_new_n19496__ = ys__n19973 & ys__n19985;
  assign new_new_n19497__ = ~new_new_n19495__ & ~new_new_n19496__;
  assign new_new_n19498__ = ~ys__n352 & ~new_new_n19497__;
  assign new_new_n19499__ = ~ys__n220 & ys__n47038;
  assign new_new_n19500__ = new_new_n18439__ & new_new_n19499__;
  assign new_new_n19501__ = ~ys__n220 & ys__n47086;
  assign new_new_n19502__ = new_new_n18441__ & new_new_n19501__;
  assign new_new_n19503__ = ~ys__n220 & ys__n47022;
  assign new_new_n19504__ = new_new_n18444__ & new_new_n19503__;
  assign new_new_n19505__ = ~new_new_n19502__ & ~new_new_n19504__;
  assign new_new_n19506__ = ~new_new_n19500__ & new_new_n19505__;
  assign new_new_n19507__ = new_new_n18453__ & ~new_new_n19506__;
  assign ys__n19914 = new_new_n19498__ | new_new_n19507__;
  assign new_new_n19509__ = ys__n19844 & ys__n19857;
  assign new_new_n19510__ = new_new_n18116__ & new_new_n19509__;
  assign new_new_n19511__ = ~ys__n23276 & ~new_new_n18904__;
  assign new_new_n19512__ = ys__n23276 & ~new_new_n18910__;
  assign new_new_n19513__ = ~new_new_n19511__ & ~new_new_n19512__;
  assign new_new_n19514__ = ~ys__n23278 & ~new_new_n19513__;
  assign new_new_n19515__ = ~ys__n23276 & ~new_new_n18913__;
  assign new_new_n19516__ = ~new_new_n19082__ & ~new_new_n19515__;
  assign new_new_n19517__ = ys__n23278 & ~new_new_n19516__;
  assign new_new_n19518__ = ~new_new_n19514__ & ~new_new_n19517__;
  assign new_new_n19519__ = ~ys__n1505 & ~new_new_n19518__;
  assign new_new_n19520__ = ~ys__n23276 & new_new_n18919__;
  assign new_new_n19521__ = ys__n23278 & new_new_n19520__;
  assign new_new_n19522__ = ~new_new_n19514__ & ~new_new_n19521__;
  assign new_new_n19523__ = ys__n1505 & ~new_new_n19522__;
  assign new_new_n19524__ = ~new_new_n19519__ & ~new_new_n19523__;
  assign new_new_n19525__ = ~new_new_n18116__ & ~new_new_n19524__;
  assign new_new_n19526__ = ~new_new_n19510__ & ~new_new_n19525__;
  assign new_new_n19527__ = new_new_n18213__ & ~new_new_n19526__;
  assign new_new_n19528__ = ~new_new_n18485__ & ~new_new_n18490__;
  assign new_new_n19529__ = ~ys__n23272 & ~new_new_n19528__;
  assign new_new_n19530__ = ys__n23272 & ~new_new_n19382__;
  assign new_new_n19531__ = ~new_new_n19529__ & ~new_new_n19530__;
  assign new_new_n19532__ = ~ys__n23274 & ~new_new_n19531__;
  assign new_new_n19533__ = ys__n23274 & ~new_new_n19239__;
  assign new_new_n19534__ = ~new_new_n19532__ & ~new_new_n19533__;
  assign new_new_n19535__ = ~ys__n23276 & ~new_new_n19534__;
  assign new_new_n19536__ = ys__n23276 & ~new_new_n18935__;
  assign new_new_n19537__ = ~new_new_n19535__ & ~new_new_n19536__;
  assign new_new_n19538__ = new_new_n18219__ & ~new_new_n19537__;
  assign new_new_n19539__ = ~new_new_n19527__ & ~new_new_n19538__;
  assign new_new_n19540__ = new_new_n18224__ & ~new_new_n19539__;
  assign new_new_n19541__ = ~new_new_n10786__ & new_new_n18226__;
  assign new_new_n19542__ = ys__n1498 & new_new_n18285__;
  assign new_new_n19543__ = ~new_new_n19541__ & ~new_new_n19542__;
  assign new_new_n19544__ = ~ys__n1496 & ~new_new_n19543__;
  assign new_new_n19545__ = ys__n1496 & ~new_new_n18285__;
  assign new_new_n19546__ = ~new_new_n19544__ & ~new_new_n19545__;
  assign new_new_n19547__ = ~ys__n1495 & ~new_new_n19546__;
  assign new_new_n19548__ = ys__n1495 & new_new_n16821__;
  assign new_new_n19549__ = ~new_new_n19547__ & ~new_new_n19548__;
  assign new_new_n19550__ = ~new_new_n18224__ & ~new_new_n19549__;
  assign new_new_n19551__ = ~new_new_n19540__ & ~new_new_n19550__;
  assign new_new_n19552__ = new_new_n18581__ & ~new_new_n19551__;
  assign new_new_n19553__ = ~new_new_n18288__ & ~new_new_n19481__;
  assign new_new_n19554__ = ~new_new_n10782__ & ~new_new_n19553__;
  assign new_new_n19555__ = new_new_n18286__ & ~new_new_n19554__;
  assign new_new_n19556__ = ~new_new_n18286__ & new_new_n19554__;
  assign new_new_n19557__ = ~new_new_n19555__ & ~new_new_n19556__;
  assign new_new_n19558__ = ~ys__n1489 & ~new_new_n19557__;
  assign new_new_n19559__ = ~new_new_n10783__ & ~new_new_n19487__;
  assign new_new_n19560__ = ~new_new_n16822__ & ~new_new_n19559__;
  assign new_new_n19561__ = new_new_n10786__ & ~new_new_n19560__;
  assign new_new_n19562__ = ~new_new_n10786__ & new_new_n19560__;
  assign new_new_n19563__ = ~new_new_n19561__ & ~new_new_n19562__;
  assign new_new_n19564__ = ys__n1489 & ~new_new_n19563__;
  assign new_new_n19565__ = ~new_new_n19558__ & ~new_new_n19564__;
  assign new_new_n19566__ = ~new_new_n18427__ & ~new_new_n19565__;
  assign new_new_n19567__ = ~new_new_n19552__ & ~new_new_n19566__;
  assign new_new_n19568__ = ~ys__n19973 & ~new_new_n19567__;
  assign new_new_n19569__ = ys__n19973 & ys__n19986;
  assign new_new_n19570__ = ~new_new_n19568__ & ~new_new_n19569__;
  assign new_new_n19571__ = ~ys__n352 & ~new_new_n19570__;
  assign new_new_n19572__ = ~ys__n220 & ys__n47039;
  assign new_new_n19573__ = new_new_n18439__ & new_new_n19572__;
  assign new_new_n19574__ = ~ys__n220 & ys__n47087;
  assign new_new_n19575__ = new_new_n18441__ & new_new_n19574__;
  assign new_new_n19576__ = ~ys__n220 & ys__n47023;
  assign new_new_n19577__ = new_new_n18444__ & new_new_n19576__;
  assign new_new_n19578__ = ~new_new_n19575__ & ~new_new_n19577__;
  assign new_new_n19579__ = ~new_new_n19573__ & new_new_n19578__;
  assign new_new_n19580__ = new_new_n18453__ & ~new_new_n19579__;
  assign ys__n19917 = new_new_n19571__ | new_new_n19580__;
  assign new_new_n19582__ = ys__n19844 & ys__n19858;
  assign new_new_n19583__ = new_new_n18116__ & new_new_n19582__;
  assign new_new_n19584__ = ~ys__n23276 & ~new_new_n18989__;
  assign new_new_n19585__ = ys__n23276 & ~new_new_n18995__;
  assign new_new_n19586__ = ~new_new_n19584__ & ~new_new_n19585__;
  assign new_new_n19587__ = ~ys__n23278 & ~new_new_n19586__;
  assign new_new_n19588__ = ~ys__n23276 & ~new_new_n18998__;
  assign new_new_n19589__ = ~new_new_n19082__ & ~new_new_n19588__;
  assign new_new_n19590__ = ys__n23278 & ~new_new_n19589__;
  assign new_new_n19591__ = ~new_new_n19587__ & ~new_new_n19590__;
  assign new_new_n19592__ = ~ys__n1505 & ~new_new_n19591__;
  assign new_new_n19593__ = ~ys__n23276 & new_new_n19004__;
  assign new_new_n19594__ = ys__n23278 & new_new_n19593__;
  assign new_new_n19595__ = ~new_new_n19587__ & ~new_new_n19594__;
  assign new_new_n19596__ = ys__n1505 & ~new_new_n19595__;
  assign new_new_n19597__ = ~new_new_n19592__ & ~new_new_n19596__;
  assign new_new_n19598__ = ~new_new_n18116__ & ~new_new_n19597__;
  assign new_new_n19599__ = ~new_new_n19583__ & ~new_new_n19598__;
  assign new_new_n19600__ = new_new_n18213__ & ~new_new_n19599__;
  assign new_new_n19601__ = ~new_new_n18151__ & ~new_new_n18154__;
  assign new_new_n19602__ = ~ys__n23272 & ~new_new_n19601__;
  assign new_new_n19603__ = ys__n23272 & ~new_new_n19455__;
  assign new_new_n19604__ = ~new_new_n19602__ & ~new_new_n19603__;
  assign new_new_n19605__ = ~ys__n23274 & ~new_new_n19604__;
  assign new_new_n19606__ = ys__n23274 & ~new_new_n19312__;
  assign new_new_n19607__ = ~new_new_n19605__ & ~new_new_n19606__;
  assign new_new_n19608__ = ~ys__n23276 & ~new_new_n19607__;
  assign new_new_n19609__ = ys__n23276 & ~new_new_n19020__;
  assign new_new_n19610__ = ~new_new_n19608__ & ~new_new_n19609__;
  assign new_new_n19611__ = new_new_n18219__ & ~new_new_n19610__;
  assign new_new_n19612__ = ~new_new_n19600__ & ~new_new_n19611__;
  assign new_new_n19613__ = new_new_n18224__ & ~new_new_n19612__;
  assign new_new_n19614__ = ~new_new_n10790__ & new_new_n18226__;
  assign new_new_n19615__ = ys__n1498 & new_new_n18282__;
  assign new_new_n19616__ = ~new_new_n19614__ & ~new_new_n19615__;
  assign new_new_n19617__ = ~ys__n1496 & ~new_new_n19616__;
  assign new_new_n19618__ = ys__n1496 & ~new_new_n18282__;
  assign new_new_n19619__ = ~new_new_n19617__ & ~new_new_n19618__;
  assign new_new_n19620__ = ~ys__n1495 & ~new_new_n19619__;
  assign new_new_n19621__ = ys__n1495 & new_new_n16827__;
  assign new_new_n19622__ = ~new_new_n19620__ & ~new_new_n19621__;
  assign new_new_n19623__ = ~new_new_n18224__ & ~new_new_n19622__;
  assign new_new_n19624__ = ~new_new_n19613__ & ~new_new_n19623__;
  assign new_new_n19625__ = new_new_n18581__ & ~new_new_n19624__;
  assign new_new_n19626__ = new_new_n18289__ & ~new_new_n19481__;
  assign new_new_n19627__ = new_new_n18312__ & ~new_new_n19626__;
  assign new_new_n19628__ = new_new_n18283__ & ~new_new_n19627__;
  assign new_new_n19629__ = ~new_new_n18283__ & new_new_n19627__;
  assign new_new_n19630__ = ~new_new_n19628__ & ~new_new_n19629__;
  assign new_new_n19631__ = ~ys__n1489 & ~new_new_n19630__;
  assign new_new_n19632__ = new_new_n16803__ & ~new_new_n19487__;
  assign new_new_n19633__ = new_new_n16824__ & ~new_new_n19632__;
  assign new_new_n19634__ = new_new_n10790__ & ~new_new_n19633__;
  assign new_new_n19635__ = ~new_new_n10790__ & new_new_n19633__;
  assign new_new_n19636__ = ~new_new_n19634__ & ~new_new_n19635__;
  assign new_new_n19637__ = ys__n1489 & ~new_new_n19636__;
  assign new_new_n19638__ = ~new_new_n19631__ & ~new_new_n19637__;
  assign new_new_n19639__ = ~new_new_n18427__ & ~new_new_n19638__;
  assign new_new_n19640__ = ~new_new_n19625__ & ~new_new_n19639__;
  assign new_new_n19641__ = ~ys__n19973 & ~new_new_n19640__;
  assign new_new_n19642__ = ys__n19973 & ys__n19987;
  assign new_new_n19643__ = ~new_new_n19641__ & ~new_new_n19642__;
  assign new_new_n19644__ = ~ys__n352 & ~new_new_n19643__;
  assign new_new_n19645__ = ~ys__n220 & ys__n47040;
  assign new_new_n19646__ = new_new_n18439__ & new_new_n19645__;
  assign new_new_n19647__ = ~ys__n220 & ys__n47088;
  assign new_new_n19648__ = new_new_n18441__ & new_new_n19647__;
  assign new_new_n19649__ = ~ys__n220 & ys__n47024;
  assign new_new_n19650__ = new_new_n18444__ & new_new_n19649__;
  assign new_new_n19651__ = ~new_new_n19648__ & ~new_new_n19650__;
  assign new_new_n19652__ = ~new_new_n19646__ & new_new_n19651__;
  assign new_new_n19653__ = new_new_n18453__ & ~new_new_n19652__;
  assign ys__n19920 = new_new_n19644__ | new_new_n19653__;
  assign new_new_n19655__ = ys__n19844 & ys__n19859;
  assign new_new_n19656__ = new_new_n18116__ & new_new_n19655__;
  assign new_new_n19657__ = ~ys__n23276 & ~new_new_n19074__;
  assign new_new_n19658__ = ys__n23276 & ~new_new_n19080__;
  assign new_new_n19659__ = ~new_new_n19657__ & ~new_new_n19658__;
  assign new_new_n19660__ = ~ys__n23278 & ~new_new_n19659__;
  assign new_new_n19661__ = ys__n23278 & ys__n28030;
  assign new_new_n19662__ = ~new_new_n19660__ & ~new_new_n19661__;
  assign new_new_n19663__ = ~ys__n1505 & ~new_new_n19662__;
  assign new_new_n19664__ = ~ys__n23276 & new_new_n19087__;
  assign new_new_n19665__ = ys__n23278 & new_new_n19664__;
  assign new_new_n19666__ = ~new_new_n19660__ & ~new_new_n19665__;
  assign new_new_n19667__ = ys__n1505 & ~new_new_n19666__;
  assign new_new_n19668__ = ~new_new_n19663__ & ~new_new_n19667__;
  assign new_new_n19669__ = ~new_new_n18116__ & ~new_new_n19668__;
  assign new_new_n19670__ = ~new_new_n19656__ & ~new_new_n19669__;
  assign new_new_n19671__ = new_new_n18213__ & ~new_new_n19670__;
  assign new_new_n19672__ = ~new_new_n18491__ & ~new_new_n18494__;
  assign new_new_n19673__ = ~ys__n23272 & ~new_new_n19672__;
  assign new_new_n19674__ = ys__n23272 & ~new_new_n19528__;
  assign new_new_n19675__ = ~new_new_n19673__ & ~new_new_n19674__;
  assign new_new_n19676__ = ~ys__n23274 & ~new_new_n19675__;
  assign new_new_n19677__ = ys__n23274 & ~new_new_n19385__;
  assign new_new_n19678__ = ~new_new_n19676__ & ~new_new_n19677__;
  assign new_new_n19679__ = ~ys__n23276 & ~new_new_n19678__;
  assign new_new_n19680__ = ys__n23276 & ~new_new_n19103__;
  assign new_new_n19681__ = ~new_new_n19679__ & ~new_new_n19680__;
  assign new_new_n19682__ = new_new_n18219__ & ~new_new_n19681__;
  assign new_new_n19683__ = ~new_new_n19671__ & ~new_new_n19682__;
  assign new_new_n19684__ = new_new_n18224__ & ~new_new_n19683__;
  assign new_new_n19685__ = ~new_new_n10793__ & new_new_n18226__;
  assign new_new_n19686__ = ys__n1498 & new_new_n18280__;
  assign new_new_n19687__ = ~new_new_n19685__ & ~new_new_n19686__;
  assign new_new_n19688__ = ~ys__n1496 & ~new_new_n19687__;
  assign new_new_n19689__ = ys__n1496 & ~new_new_n18280__;
  assign new_new_n19690__ = ~new_new_n19688__ & ~new_new_n19689__;
  assign new_new_n19691__ = ~ys__n1495 & ~new_new_n19690__;
  assign new_new_n19692__ = ys__n1495 & new_new_n16826__;
  assign new_new_n19693__ = ~new_new_n19691__ & ~new_new_n19692__;
  assign new_new_n19694__ = ~new_new_n18224__ & ~new_new_n19693__;
  assign new_new_n19695__ = ~new_new_n19684__ & ~new_new_n19694__;
  assign new_new_n19696__ = new_new_n18581__ & ~new_new_n19695__;
  assign new_new_n19697__ = ~new_new_n18283__ & ~new_new_n19627__;
  assign new_new_n19698__ = ~new_new_n10789__ & ~new_new_n19697__;
  assign new_new_n19699__ = new_new_n18281__ & ~new_new_n19698__;
  assign new_new_n19700__ = ~new_new_n18281__ & new_new_n19698__;
  assign new_new_n19701__ = ~new_new_n19699__ & ~new_new_n19700__;
  assign new_new_n19702__ = ~ys__n1489 & ~new_new_n19701__;
  assign new_new_n19703__ = ~new_new_n10790__ & ~new_new_n19633__;
  assign new_new_n19704__ = ~new_new_n16827__ & ~new_new_n19703__;
  assign new_new_n19705__ = new_new_n10793__ & ~new_new_n19704__;
  assign new_new_n19706__ = ~new_new_n10793__ & new_new_n19704__;
  assign new_new_n19707__ = ~new_new_n19705__ & ~new_new_n19706__;
  assign new_new_n19708__ = ys__n1489 & ~new_new_n19707__;
  assign new_new_n19709__ = ~new_new_n19702__ & ~new_new_n19708__;
  assign new_new_n19710__ = ~new_new_n18427__ & ~new_new_n19709__;
  assign new_new_n19711__ = ~new_new_n19696__ & ~new_new_n19710__;
  assign new_new_n19712__ = ~ys__n19973 & ~new_new_n19711__;
  assign new_new_n19713__ = ys__n19973 & ys__n19988;
  assign new_new_n19714__ = ~new_new_n19712__ & ~new_new_n19713__;
  assign new_new_n19715__ = ~ys__n352 & ~new_new_n19714__;
  assign new_new_n19716__ = ~ys__n220 & ys__n47041;
  assign new_new_n19717__ = new_new_n18439__ & new_new_n19716__;
  assign new_new_n19718__ = ~ys__n220 & ys__n47089;
  assign new_new_n19719__ = new_new_n18441__ & new_new_n19718__;
  assign new_new_n19720__ = ~ys__n220 & ys__n47025;
  assign new_new_n19721__ = new_new_n18444__ & new_new_n19720__;
  assign new_new_n19722__ = ~new_new_n19719__ & ~new_new_n19721__;
  assign new_new_n19723__ = ~new_new_n19717__ & new_new_n19722__;
  assign new_new_n19724__ = new_new_n18453__ & ~new_new_n19723__;
  assign ys__n19923 = new_new_n19715__ | new_new_n19724__;
  assign new_new_n19726__ = ys__n19844 & ys__n19860;
  assign new_new_n19727__ = new_new_n18116__ & new_new_n19726__;
  assign new_new_n19728__ = ~ys__n23278 & ~new_new_n18208__;
  assign new_new_n19729__ = ~new_new_n19661__ & ~new_new_n19728__;
  assign new_new_n19730__ = ~ys__n1505 & ~new_new_n19729__;
  assign new_new_n19731__ = ys__n1505 & new_new_n19728__;
  assign new_new_n19732__ = ~new_new_n19730__ & ~new_new_n19731__;
  assign new_new_n19733__ = ~new_new_n18116__ & ~new_new_n19732__;
  assign new_new_n19734__ = ~new_new_n19727__ & ~new_new_n19733__;
  assign new_new_n19735__ = new_new_n18213__ & ~new_new_n19734__;
  assign new_new_n19736__ = ~ys__n1502 & ys__n27855;
  assign new_new_n19737__ = ~new_new_n18155__ & ~new_new_n18164__;
  assign new_new_n19738__ = ~ys__n23272 & ~new_new_n19737__;
  assign new_new_n19739__ = ys__n23272 & ~new_new_n19601__;
  assign new_new_n19740__ = ~new_new_n19738__ & ~new_new_n19739__;
  assign new_new_n19741__ = ~ys__n23274 & ~new_new_n19740__;
  assign new_new_n19742__ = ys__n23274 & ~new_new_n19458__;
  assign new_new_n19743__ = ~new_new_n19741__ & ~new_new_n19742__;
  assign new_new_n19744__ = ~ys__n23276 & ~new_new_n19743__;
  assign new_new_n19745__ = ys__n23276 & ~new_new_n19173__;
  assign new_new_n19746__ = ~new_new_n19744__ & ~new_new_n19745__;
  assign new_new_n19747__ = ~ys__n23278 & ~new_new_n19746__;
  assign new_new_n19748__ = ys__n23278 & new_new_n18217__;
  assign new_new_n19749__ = ~new_new_n19747__ & ~new_new_n19748__;
  assign new_new_n19750__ = ys__n1502 & ~new_new_n19749__;
  assign new_new_n19751__ = ~new_new_n19736__ & ~new_new_n19750__;
  assign new_new_n19752__ = ~new_new_n18213__ & ~new_new_n19751__;
  assign new_new_n19753__ = ~new_new_n19735__ & ~new_new_n19752__;
  assign new_new_n19754__ = new_new_n18224__ & ~new_new_n19753__;
  assign new_new_n19755__ = ~new_new_n10704__ & new_new_n18226__;
  assign new_new_n19756__ = ys__n1498 & new_new_n18361__;
  assign new_new_n19757__ = ~new_new_n19755__ & ~new_new_n19756__;
  assign new_new_n19758__ = ~ys__n1496 & ~new_new_n19757__;
  assign new_new_n19759__ = ys__n1496 & ~new_new_n18361__;
  assign new_new_n19760__ = ~new_new_n19758__ & ~new_new_n19759__;
  assign new_new_n19761__ = ~ys__n1495 & ~new_new_n19760__;
  assign new_new_n19762__ = ys__n1495 & new_new_n16753__;
  assign new_new_n19763__ = ~new_new_n19761__ & ~new_new_n19762__;
  assign new_new_n19764__ = ~new_new_n18224__ & ~new_new_n19763__;
  assign new_new_n19765__ = ~new_new_n19754__ & ~new_new_n19764__;
  assign new_new_n19766__ = new_new_n18581__ & ~new_new_n19765__;
  assign new_new_n19767__ = ~new_new_n18318__ & new_new_n18362__;
  assign new_new_n19768__ = new_new_n18318__ & ~new_new_n18362__;
  assign new_new_n19769__ = ~new_new_n19767__ & ~new_new_n19768__;
  assign new_new_n19770__ = ~ys__n1489 & ~new_new_n19769__;
  assign new_new_n19771__ = new_new_n10704__ & ~new_new_n16832__;
  assign new_new_n19772__ = ~new_new_n10704__ & new_new_n16832__;
  assign new_new_n19773__ = ~new_new_n19771__ & ~new_new_n19772__;
  assign new_new_n19774__ = ys__n1489 & ~new_new_n19773__;
  assign new_new_n19775__ = ~new_new_n19770__ & ~new_new_n19774__;
  assign new_new_n19776__ = ~new_new_n18427__ & ~new_new_n19775__;
  assign new_new_n19777__ = ~new_new_n19766__ & ~new_new_n19776__;
  assign new_new_n19778__ = ~ys__n19973 & ~new_new_n19777__;
  assign new_new_n19779__ = ys__n19973 & ys__n19989;
  assign new_new_n19780__ = ~new_new_n19778__ & ~new_new_n19779__;
  assign new_new_n19781__ = ~ys__n352 & ~new_new_n19780__;
  assign new_new_n19782__ = ~ys__n220 & ys__n47090;
  assign new_new_n19783__ = new_new_n18439__ & new_new_n19782__;
  assign new_new_n19784__ = new_new_n18441__ & new_new_n19782__;
  assign new_new_n19785__ = new_new_n18438__ & new_new_n18444__;
  assign new_new_n19786__ = ~new_new_n19784__ & ~new_new_n19785__;
  assign new_new_n19787__ = ~new_new_n19783__ & new_new_n19786__;
  assign new_new_n19788__ = new_new_n18453__ & ~new_new_n19787__;
  assign ys__n19926 = new_new_n19781__ | new_new_n19788__;
  assign new_new_n19790__ = ys__n19844 & ys__n19861;
  assign new_new_n19791__ = new_new_n18116__ & new_new_n19790__;
  assign new_new_n19792__ = ~ys__n23278 & ~new_new_n18545__;
  assign new_new_n19793__ = ~new_new_n19661__ & ~new_new_n19792__;
  assign new_new_n19794__ = ~ys__n1505 & ~new_new_n19793__;
  assign new_new_n19795__ = ys__n1505 & ~ys__n23278;
  assign new_new_n19796__ = ~new_new_n18555__ & new_new_n19795__;
  assign new_new_n19797__ = ~new_new_n19794__ & ~new_new_n19796__;
  assign new_new_n19798__ = ~new_new_n18116__ & ~new_new_n19797__;
  assign new_new_n19799__ = ~new_new_n19791__ & ~new_new_n19798__;
  assign new_new_n19800__ = new_new_n18213__ & ~new_new_n19799__;
  assign new_new_n19801__ = ~ys__n1502 & ys__n27857;
  assign new_new_n19802__ = ~new_new_n18495__ & ~new_new_n18504__;
  assign new_new_n19803__ = ~ys__n23272 & ~new_new_n19802__;
  assign new_new_n19804__ = ys__n23272 & ~new_new_n19672__;
  assign new_new_n19805__ = ~new_new_n19803__ & ~new_new_n19804__;
  assign new_new_n19806__ = ~ys__n23274 & ~new_new_n19805__;
  assign new_new_n19807__ = ys__n23274 & ~new_new_n19531__;
  assign new_new_n19808__ = ~new_new_n19806__ & ~new_new_n19807__;
  assign new_new_n19809__ = ~ys__n23276 & ~new_new_n19808__;
  assign new_new_n19810__ = ys__n23276 & ~new_new_n19242__;
  assign new_new_n19811__ = ~new_new_n19809__ & ~new_new_n19810__;
  assign new_new_n19812__ = ~ys__n23278 & ~new_new_n19811__;
  assign new_new_n19813__ = ys__n23278 & new_new_n18566__;
  assign new_new_n19814__ = ~new_new_n19812__ & ~new_new_n19813__;
  assign new_new_n19815__ = ys__n1502 & ~new_new_n19814__;
  assign new_new_n19816__ = ~new_new_n19801__ & ~new_new_n19815__;
  assign new_new_n19817__ = ~new_new_n18213__ & ~new_new_n19816__;
  assign new_new_n19818__ = ~new_new_n19800__ & ~new_new_n19817__;
  assign new_new_n19819__ = new_new_n18224__ & ~new_new_n19818__;
  assign new_new_n19820__ = ~new_new_n10707__ & new_new_n18226__;
  assign new_new_n19821__ = ys__n1498 & new_new_n18359__;
  assign new_new_n19822__ = ~new_new_n19820__ & ~new_new_n19821__;
  assign new_new_n19823__ = ~ys__n1496 & ~new_new_n19822__;
  assign new_new_n19824__ = ys__n1496 & ~new_new_n18359__;
  assign new_new_n19825__ = ~new_new_n19823__ & ~new_new_n19824__;
  assign new_new_n19826__ = ~ys__n1495 & ~new_new_n19825__;
  assign new_new_n19827__ = ys__n1495 & new_new_n16752__;
  assign new_new_n19828__ = ~new_new_n19826__ & ~new_new_n19827__;
  assign new_new_n19829__ = ~new_new_n18224__ & ~new_new_n19828__;
  assign new_new_n19830__ = ~new_new_n19819__ & ~new_new_n19829__;
  assign new_new_n19831__ = new_new_n18581__ & ~new_new_n19830__;
  assign new_new_n19832__ = ~new_new_n18318__ & ~new_new_n18362__;
  assign new_new_n19833__ = ~new_new_n10703__ & ~new_new_n19832__;
  assign new_new_n19834__ = new_new_n18360__ & ~new_new_n19833__;
  assign new_new_n19835__ = ~new_new_n18360__ & new_new_n19833__;
  assign new_new_n19836__ = ~new_new_n19834__ & ~new_new_n19835__;
  assign new_new_n19837__ = ~ys__n1489 & ~new_new_n19836__;
  assign new_new_n19838__ = ~new_new_n10704__ & ~new_new_n16832__;
  assign new_new_n19839__ = ~new_new_n16753__ & ~new_new_n19838__;
  assign new_new_n19840__ = new_new_n10707__ & ~new_new_n19839__;
  assign new_new_n19841__ = ~new_new_n10707__ & new_new_n19839__;
  assign new_new_n19842__ = ~new_new_n19840__ & ~new_new_n19841__;
  assign new_new_n19843__ = ys__n1489 & ~new_new_n19842__;
  assign new_new_n19844__ = ~new_new_n19837__ & ~new_new_n19843__;
  assign new_new_n19845__ = ~new_new_n18427__ & ~new_new_n19844__;
  assign new_new_n19846__ = ~new_new_n19831__ & ~new_new_n19845__;
  assign new_new_n19847__ = ~ys__n19973 & ~new_new_n19846__;
  assign new_new_n19848__ = ys__n19973 & ys__n19990;
  assign new_new_n19849__ = ~new_new_n19847__ & ~new_new_n19848__;
  assign new_new_n19850__ = ~ys__n352 & ~new_new_n19849__;
  assign new_new_n19851__ = ~ys__n220 & ys__n47091;
  assign new_new_n19852__ = new_new_n18439__ & new_new_n19851__;
  assign new_new_n19853__ = new_new_n18441__ & new_new_n19851__;
  assign new_new_n19854__ = new_new_n18444__ & new_new_n18595__;
  assign new_new_n19855__ = ~new_new_n19853__ & ~new_new_n19854__;
  assign new_new_n19856__ = ~new_new_n19852__ & new_new_n19855__;
  assign new_new_n19857__ = new_new_n18453__ & ~new_new_n19856__;
  assign ys__n19929 = new_new_n19850__ | new_new_n19857__;
  assign new_new_n19859__ = ys__n19844 & ys__n19862;
  assign new_new_n19860__ = new_new_n18116__ & new_new_n19859__;
  assign new_new_n19861__ = ~ys__n23278 & ~new_new_n18648__;
  assign new_new_n19862__ = ~new_new_n19661__ & ~new_new_n19861__;
  assign new_new_n19863__ = ~ys__n1505 & ~new_new_n19862__;
  assign new_new_n19864__ = ~new_new_n18655__ & new_new_n19795__;
  assign new_new_n19865__ = ~new_new_n19863__ & ~new_new_n19864__;
  assign new_new_n19866__ = ~new_new_n18116__ & ~new_new_n19865__;
  assign new_new_n19867__ = ~new_new_n19860__ & ~new_new_n19866__;
  assign new_new_n19868__ = new_new_n18213__ & ~new_new_n19867__;
  assign new_new_n19869__ = ~ys__n1502 & ys__n27859;
  assign new_new_n19870__ = ~new_new_n18165__ & ~new_new_n18168__;
  assign new_new_n19871__ = ~ys__n23272 & ~new_new_n19870__;
  assign new_new_n19872__ = ys__n23272 & ~new_new_n19737__;
  assign new_new_n19873__ = ~new_new_n19871__ & ~new_new_n19872__;
  assign new_new_n19874__ = ~ys__n23274 & ~new_new_n19873__;
  assign new_new_n19875__ = ys__n23274 & ~new_new_n19604__;
  assign new_new_n19876__ = ~new_new_n19874__ & ~new_new_n19875__;
  assign new_new_n19877__ = ~ys__n23276 & ~new_new_n19876__;
  assign new_new_n19878__ = ys__n23276 & ~new_new_n19315__;
  assign new_new_n19879__ = ~new_new_n19877__ & ~new_new_n19878__;
  assign new_new_n19880__ = ~ys__n23278 & ~new_new_n19879__;
  assign new_new_n19881__ = ys__n23278 & new_new_n18668__;
  assign new_new_n19882__ = ~new_new_n19880__ & ~new_new_n19881__;
  assign new_new_n19883__ = ys__n1502 & ~new_new_n19882__;
  assign new_new_n19884__ = ~new_new_n19869__ & ~new_new_n19883__;
  assign new_new_n19885__ = ~new_new_n18213__ & ~new_new_n19884__;
  assign new_new_n19886__ = ~new_new_n19868__ & ~new_new_n19885__;
  assign new_new_n19887__ = new_new_n18224__ & ~new_new_n19886__;
  assign new_new_n19888__ = ~new_new_n10711__ & new_new_n18226__;
  assign new_new_n19889__ = ys__n1498 & new_new_n18356__;
  assign new_new_n19890__ = ~new_new_n19888__ & ~new_new_n19889__;
  assign new_new_n19891__ = ~ys__n1496 & ~new_new_n19890__;
  assign new_new_n19892__ = ys__n1496 & ~new_new_n18356__;
  assign new_new_n19893__ = ~new_new_n19891__ & ~new_new_n19892__;
  assign new_new_n19894__ = ~ys__n1495 & ~new_new_n19893__;
  assign new_new_n19895__ = ys__n1495 & new_new_n16758__;
  assign new_new_n19896__ = ~new_new_n19894__ & ~new_new_n19895__;
  assign new_new_n19897__ = ~new_new_n18224__ & ~new_new_n19896__;
  assign new_new_n19898__ = ~new_new_n19887__ & ~new_new_n19897__;
  assign new_new_n19899__ = new_new_n18581__ & ~new_new_n19898__;
  assign new_new_n19900__ = ~new_new_n18318__ & new_new_n18363__;
  assign new_new_n19901__ = new_new_n18369__ & ~new_new_n19900__;
  assign new_new_n19902__ = new_new_n18357__ & ~new_new_n19901__;
  assign new_new_n19903__ = ~new_new_n18357__ & new_new_n19901__;
  assign new_new_n19904__ = ~new_new_n19902__ & ~new_new_n19903__;
  assign new_new_n19905__ = ~ys__n1489 & ~new_new_n19904__;
  assign new_new_n19906__ = new_new_n16774__ & ~new_new_n16832__;
  assign new_new_n19907__ = new_new_n16755__ & ~new_new_n19906__;
  assign new_new_n19908__ = new_new_n10711__ & ~new_new_n19907__;
  assign new_new_n19909__ = ~new_new_n10711__ & new_new_n19907__;
  assign new_new_n19910__ = ~new_new_n19908__ & ~new_new_n19909__;
  assign new_new_n19911__ = ys__n1489 & ~new_new_n19910__;
  assign new_new_n19912__ = ~new_new_n19905__ & ~new_new_n19911__;
  assign new_new_n19913__ = ~new_new_n18427__ & ~new_new_n19912__;
  assign new_new_n19914__ = ~new_new_n19899__ & ~new_new_n19913__;
  assign new_new_n19915__ = ~ys__n19973 & ~new_new_n19914__;
  assign new_new_n19916__ = ys__n19973 & ys__n19991;
  assign new_new_n19917__ = ~new_new_n19915__ & ~new_new_n19916__;
  assign new_new_n19918__ = ~ys__n352 & ~new_new_n19917__;
  assign new_new_n19919__ = ~ys__n220 & ys__n47092;
  assign new_new_n19920__ = new_new_n18439__ & new_new_n19919__;
  assign new_new_n19921__ = new_new_n18441__ & new_new_n19919__;
  assign new_new_n19922__ = new_new_n18444__ & new_new_n18699__;
  assign new_new_n19923__ = ~new_new_n19921__ & ~new_new_n19922__;
  assign new_new_n19924__ = ~new_new_n19920__ & new_new_n19923__;
  assign new_new_n19925__ = new_new_n18453__ & ~new_new_n19924__;
  assign ys__n19932 = new_new_n19918__ | new_new_n19925__;
  assign new_new_n19927__ = ys__n19844 & ys__n19863;
  assign new_new_n19928__ = new_new_n18116__ & new_new_n19927__;
  assign new_new_n19929__ = ~ys__n23278 & ~new_new_n18750__;
  assign new_new_n19930__ = ~new_new_n19661__ & ~new_new_n19929__;
  assign new_new_n19931__ = ~ys__n1505 & ~new_new_n19930__;
  assign new_new_n19932__ = ~new_new_n18758__ & new_new_n19795__;
  assign new_new_n19933__ = ~new_new_n19931__ & ~new_new_n19932__;
  assign new_new_n19934__ = ~new_new_n18116__ & ~new_new_n19933__;
  assign new_new_n19935__ = ~new_new_n19928__ & ~new_new_n19934__;
  assign new_new_n19936__ = new_new_n18213__ & ~new_new_n19935__;
  assign new_new_n19937__ = ~ys__n1502 & ys__n27861;
  assign new_new_n19938__ = ~new_new_n18505__ & ~new_new_n18508__;
  assign new_new_n19939__ = ~ys__n23272 & ~new_new_n19938__;
  assign new_new_n19940__ = ys__n23272 & ~new_new_n19802__;
  assign new_new_n19941__ = ~new_new_n19939__ & ~new_new_n19940__;
  assign new_new_n19942__ = ~ys__n23274 & ~new_new_n19941__;
  assign new_new_n19943__ = ys__n23274 & ~new_new_n19675__;
  assign new_new_n19944__ = ~new_new_n19942__ & ~new_new_n19943__;
  assign new_new_n19945__ = ~ys__n23276 & ~new_new_n19944__;
  assign new_new_n19946__ = ys__n23276 & ~new_new_n19388__;
  assign new_new_n19947__ = ~new_new_n19945__ & ~new_new_n19946__;
  assign new_new_n19948__ = ~ys__n23278 & ~new_new_n19947__;
  assign new_new_n19949__ = ys__n23278 & new_new_n18771__;
  assign new_new_n19950__ = ~new_new_n19948__ & ~new_new_n19949__;
  assign new_new_n19951__ = ys__n1502 & ~new_new_n19950__;
  assign new_new_n19952__ = ~new_new_n19937__ & ~new_new_n19951__;
  assign new_new_n19953__ = ~new_new_n18213__ & ~new_new_n19952__;
  assign new_new_n19954__ = ~new_new_n19936__ & ~new_new_n19953__;
  assign new_new_n19955__ = new_new_n18224__ & ~new_new_n19954__;
  assign new_new_n19956__ = ~new_new_n10714__ & new_new_n18226__;
  assign new_new_n19957__ = ys__n1498 & new_new_n18354__;
  assign new_new_n19958__ = ~new_new_n19956__ & ~new_new_n19957__;
  assign new_new_n19959__ = ~ys__n1496 & ~new_new_n19958__;
  assign new_new_n19960__ = ys__n1496 & ~new_new_n18354__;
  assign new_new_n19961__ = ~new_new_n19959__ & ~new_new_n19960__;
  assign new_new_n19962__ = ~ys__n1495 & ~new_new_n19961__;
  assign new_new_n19963__ = ys__n1495 & new_new_n16757__;
  assign new_new_n19964__ = ~new_new_n19962__ & ~new_new_n19963__;
  assign new_new_n19965__ = ~new_new_n18224__ & ~new_new_n19964__;
  assign new_new_n19966__ = ~new_new_n19955__ & ~new_new_n19965__;
  assign new_new_n19967__ = new_new_n18581__ & ~new_new_n19966__;
  assign new_new_n19968__ = ~new_new_n18357__ & ~new_new_n19901__;
  assign new_new_n19969__ = ~new_new_n10710__ & ~new_new_n19968__;
  assign new_new_n19970__ = new_new_n18355__ & ~new_new_n19969__;
  assign new_new_n19971__ = ~new_new_n18355__ & new_new_n19969__;
  assign new_new_n19972__ = ~new_new_n19970__ & ~new_new_n19971__;
  assign new_new_n19973__ = ~ys__n1489 & ~new_new_n19972__;
  assign new_new_n19974__ = ~new_new_n10711__ & ~new_new_n19907__;
  assign new_new_n19975__ = ~new_new_n16758__ & ~new_new_n19974__;
  assign new_new_n19976__ = new_new_n10714__ & ~new_new_n19975__;
  assign new_new_n19977__ = ~new_new_n10714__ & new_new_n19975__;
  assign new_new_n19978__ = ~new_new_n19976__ & ~new_new_n19977__;
  assign new_new_n19979__ = ys__n1489 & ~new_new_n19978__;
  assign new_new_n19980__ = ~new_new_n19973__ & ~new_new_n19979__;
  assign new_new_n19981__ = ~new_new_n18427__ & ~new_new_n19980__;
  assign new_new_n19982__ = ~new_new_n19967__ & ~new_new_n19981__;
  assign new_new_n19983__ = ~ys__n19973 & ~new_new_n19982__;
  assign new_new_n19984__ = ys__n19973 & ys__n19992;
  assign new_new_n19985__ = ~new_new_n19983__ & ~new_new_n19984__;
  assign new_new_n19986__ = ~ys__n352 & ~new_new_n19985__;
  assign new_new_n19987__ = ~ys__n220 & ys__n47093;
  assign new_new_n19988__ = new_new_n18439__ & new_new_n19987__;
  assign new_new_n19989__ = new_new_n18441__ & new_new_n19987__;
  assign new_new_n19990__ = new_new_n18444__ & new_new_n18806__;
  assign new_new_n19991__ = ~new_new_n19989__ & ~new_new_n19990__;
  assign new_new_n19992__ = ~new_new_n19988__ & new_new_n19991__;
  assign new_new_n19993__ = new_new_n18453__ & ~new_new_n19992__;
  assign ys__n19935 = new_new_n19986__ | new_new_n19993__;
  assign new_new_n19995__ = ys__n19844 & ys__n19864;
  assign new_new_n19996__ = new_new_n18116__ & new_new_n19995__;
  assign new_new_n19997__ = ~ys__n23278 & ~new_new_n18835__;
  assign new_new_n19998__ = ~new_new_n19661__ & ~new_new_n19997__;
  assign new_new_n19999__ = ~ys__n1505 & ~new_new_n19998__;
  assign new_new_n20000__ = ~new_new_n18840__ & new_new_n19795__;
  assign new_new_n20001__ = ~new_new_n19999__ & ~new_new_n20000__;
  assign new_new_n20002__ = ~new_new_n18116__ & ~new_new_n20001__;
  assign new_new_n20003__ = ~new_new_n19996__ & ~new_new_n20002__;
  assign new_new_n20004__ = new_new_n18213__ & ~new_new_n20003__;
  assign new_new_n20005__ = ~ys__n1502 & ys__n27863;
  assign new_new_n20006__ = ~new_new_n18169__ & ~new_new_n18174__;
  assign new_new_n20007__ = ~ys__n23272 & ~new_new_n20006__;
  assign new_new_n20008__ = ys__n23272 & ~new_new_n19870__;
  assign new_new_n20009__ = ~new_new_n20007__ & ~new_new_n20008__;
  assign new_new_n20010__ = ~ys__n23274 & ~new_new_n20009__;
  assign new_new_n20011__ = ys__n23274 & ~new_new_n19740__;
  assign new_new_n20012__ = ~new_new_n20010__ & ~new_new_n20011__;
  assign new_new_n20013__ = ~ys__n23276 & ~new_new_n20012__;
  assign new_new_n20014__ = ys__n23276 & ~new_new_n19461__;
  assign new_new_n20015__ = ~new_new_n20013__ & ~new_new_n20014__;
  assign new_new_n20016__ = ~ys__n23278 & ~new_new_n20015__;
  assign new_new_n20017__ = ys__n23278 & new_new_n18855__;
  assign new_new_n20018__ = ~new_new_n20016__ & ~new_new_n20017__;
  assign new_new_n20019__ = ys__n1502 & ~new_new_n20018__;
  assign new_new_n20020__ = ~new_new_n20005__ & ~new_new_n20019__;
  assign new_new_n20021__ = ~new_new_n18213__ & ~new_new_n20020__;
  assign new_new_n20022__ = ~new_new_n20004__ & ~new_new_n20021__;
  assign new_new_n20023__ = new_new_n18224__ & ~new_new_n20022__;
  assign new_new_n20024__ = ~new_new_n10689__ & new_new_n18226__;
  assign new_new_n20025__ = ys__n1498 & new_new_n18350__;
  assign new_new_n20026__ = ~new_new_n20024__ & ~new_new_n20025__;
  assign new_new_n20027__ = ~ys__n1496 & ~new_new_n20026__;
  assign new_new_n20028__ = ys__n1496 & ~new_new_n18350__;
  assign new_new_n20029__ = ~new_new_n20027__ & ~new_new_n20028__;
  assign new_new_n20030__ = ~ys__n1495 & ~new_new_n20029__;
  assign new_new_n20031__ = ys__n1495 & new_new_n16764__;
  assign new_new_n20032__ = ~new_new_n20030__ & ~new_new_n20031__;
  assign new_new_n20033__ = ~new_new_n18224__ & ~new_new_n20032__;
  assign new_new_n20034__ = ~new_new_n20023__ & ~new_new_n20033__;
  assign new_new_n20035__ = new_new_n18581__ & ~new_new_n20034__;
  assign new_new_n20036__ = ~new_new_n18318__ & new_new_n18364__;
  assign new_new_n20037__ = new_new_n18373__ & ~new_new_n20036__;
  assign new_new_n20038__ = new_new_n18351__ & ~new_new_n20037__;
  assign new_new_n20039__ = ~new_new_n18351__ & new_new_n20037__;
  assign new_new_n20040__ = ~new_new_n20038__ & ~new_new_n20039__;
  assign new_new_n20041__ = ~ys__n1489 & ~new_new_n20040__;
  assign new_new_n20042__ = new_new_n16775__ & ~new_new_n16832__;
  assign new_new_n20043__ = new_new_n16761__ & ~new_new_n20042__;
  assign new_new_n20044__ = new_new_n10689__ & ~new_new_n20043__;
  assign new_new_n20045__ = ~new_new_n10689__ & new_new_n20043__;
  assign new_new_n20046__ = ~new_new_n20044__ & ~new_new_n20045__;
  assign new_new_n20047__ = ys__n1489 & ~new_new_n20046__;
  assign new_new_n20048__ = ~new_new_n20041__ & ~new_new_n20047__;
  assign new_new_n20049__ = ~new_new_n18427__ & ~new_new_n20048__;
  assign new_new_n20050__ = ~new_new_n20035__ & ~new_new_n20049__;
  assign new_new_n20051__ = ~ys__n19973 & ~new_new_n20050__;
  assign new_new_n20052__ = ys__n19973 & ys__n19993;
  assign new_new_n20053__ = ~new_new_n20051__ & ~new_new_n20052__;
  assign new_new_n20054__ = ~ys__n352 & ~new_new_n20053__;
  assign new_new_n20055__ = ~ys__n220 & ys__n47094;
  assign new_new_n20056__ = new_new_n18439__ & new_new_n20055__;
  assign new_new_n20057__ = new_new_n18441__ & new_new_n20055__;
  assign new_new_n20058__ = new_new_n18444__ & new_new_n18886__;
  assign new_new_n20059__ = ~new_new_n20057__ & ~new_new_n20058__;
  assign new_new_n20060__ = ~new_new_n20056__ & new_new_n20059__;
  assign new_new_n20061__ = new_new_n18453__ & ~new_new_n20060__;
  assign ys__n19938 = new_new_n20054__ | new_new_n20061__;
  assign new_new_n20063__ = ys__n19844 & ys__n19865;
  assign new_new_n20064__ = new_new_n18116__ & new_new_n20063__;
  assign new_new_n20065__ = ~ys__n23278 & ~new_new_n18915__;
  assign new_new_n20066__ = ~new_new_n19661__ & ~new_new_n20065__;
  assign new_new_n20067__ = ~ys__n1505 & ~new_new_n20066__;
  assign new_new_n20068__ = ~new_new_n18921__ & new_new_n19795__;
  assign new_new_n20069__ = ~new_new_n20067__ & ~new_new_n20068__;
  assign new_new_n20070__ = ~new_new_n18116__ & ~new_new_n20069__;
  assign new_new_n20071__ = ~new_new_n20064__ & ~new_new_n20070__;
  assign new_new_n20072__ = new_new_n18213__ & ~new_new_n20071__;
  assign new_new_n20073__ = ~ys__n1502 & ys__n27865;
  assign new_new_n20074__ = ~new_new_n18509__ & ~new_new_n18514__;
  assign new_new_n20075__ = ~ys__n23272 & ~new_new_n20074__;
  assign new_new_n20076__ = ys__n23272 & ~new_new_n19938__;
  assign new_new_n20077__ = ~new_new_n20075__ & ~new_new_n20076__;
  assign new_new_n20078__ = ~ys__n23274 & ~new_new_n20077__;
  assign new_new_n20079__ = ys__n23274 & ~new_new_n19805__;
  assign new_new_n20080__ = ~new_new_n20078__ & ~new_new_n20079__;
  assign new_new_n20081__ = ~ys__n23276 & ~new_new_n20080__;
  assign new_new_n20082__ = ys__n23276 & ~new_new_n19534__;
  assign new_new_n20083__ = ~new_new_n20081__ & ~new_new_n20082__;
  assign new_new_n20084__ = ~ys__n23278 & ~new_new_n20083__;
  assign new_new_n20085__ = ys__n23278 & new_new_n18936__;
  assign new_new_n20086__ = ~new_new_n20084__ & ~new_new_n20085__;
  assign new_new_n20087__ = ys__n1502 & ~new_new_n20086__;
  assign new_new_n20088__ = ~new_new_n20073__ & ~new_new_n20087__;
  assign new_new_n20089__ = ~new_new_n18213__ & ~new_new_n20088__;
  assign new_new_n20090__ = ~new_new_n20072__ & ~new_new_n20089__;
  assign new_new_n20091__ = new_new_n18224__ & ~new_new_n20090__;
  assign new_new_n20092__ = ~new_new_n10692__ & new_new_n18226__;
  assign new_new_n20093__ = ys__n1498 & new_new_n18348__;
  assign new_new_n20094__ = ~new_new_n20092__ & ~new_new_n20093__;
  assign new_new_n20095__ = ~ys__n1496 & ~new_new_n20094__;
  assign new_new_n20096__ = ys__n1496 & ~new_new_n18348__;
  assign new_new_n20097__ = ~new_new_n20095__ & ~new_new_n20096__;
  assign new_new_n20098__ = ~ys__n1495 & ~new_new_n20097__;
  assign new_new_n20099__ = ys__n1495 & new_new_n16763__;
  assign new_new_n20100__ = ~new_new_n20098__ & ~new_new_n20099__;
  assign new_new_n20101__ = ~new_new_n18224__ & ~new_new_n20100__;
  assign new_new_n20102__ = ~new_new_n20091__ & ~new_new_n20101__;
  assign new_new_n20103__ = new_new_n18581__ & ~new_new_n20102__;
  assign new_new_n20104__ = ~new_new_n18351__ & ~new_new_n20037__;
  assign new_new_n20105__ = ~new_new_n10688__ & ~new_new_n20104__;
  assign new_new_n20106__ = new_new_n18349__ & ~new_new_n20105__;
  assign new_new_n20107__ = ~new_new_n18349__ & new_new_n20105__;
  assign new_new_n20108__ = ~new_new_n20106__ & ~new_new_n20107__;
  assign new_new_n20109__ = ~ys__n1489 & ~new_new_n20108__;
  assign new_new_n20110__ = ~new_new_n10689__ & ~new_new_n20043__;
  assign new_new_n20111__ = ~new_new_n16764__ & ~new_new_n20110__;
  assign new_new_n20112__ = new_new_n10692__ & ~new_new_n20111__;
  assign new_new_n20113__ = ~new_new_n10692__ & new_new_n20111__;
  assign new_new_n20114__ = ~new_new_n20112__ & ~new_new_n20113__;
  assign new_new_n20115__ = ys__n1489 & ~new_new_n20114__;
  assign new_new_n20116__ = ~new_new_n20109__ & ~new_new_n20115__;
  assign new_new_n20117__ = ~new_new_n18427__ & ~new_new_n20116__;
  assign new_new_n20118__ = ~new_new_n20103__ & ~new_new_n20117__;
  assign new_new_n20119__ = ~ys__n19973 & ~new_new_n20118__;
  assign new_new_n20120__ = ys__n19973 & ys__n19994;
  assign new_new_n20121__ = ~new_new_n20119__ & ~new_new_n20120__;
  assign new_new_n20122__ = ~ys__n352 & ~new_new_n20121__;
  assign new_new_n20123__ = ~ys__n220 & ys__n47095;
  assign new_new_n20124__ = new_new_n18439__ & new_new_n20123__;
  assign new_new_n20125__ = new_new_n18441__ & new_new_n20123__;
  assign new_new_n20126__ = new_new_n18444__ & new_new_n18971__;
  assign new_new_n20127__ = ~new_new_n20125__ & ~new_new_n20126__;
  assign new_new_n20128__ = ~new_new_n20124__ & new_new_n20127__;
  assign new_new_n20129__ = new_new_n18453__ & ~new_new_n20128__;
  assign ys__n19941 = new_new_n20122__ | new_new_n20129__;
  assign new_new_n20131__ = ys__n19844 & ys__n19866;
  assign new_new_n20132__ = new_new_n18116__ & new_new_n20131__;
  assign new_new_n20133__ = ~ys__n23278 & ~new_new_n19000__;
  assign new_new_n20134__ = ~new_new_n19661__ & ~new_new_n20133__;
  assign new_new_n20135__ = ~ys__n1505 & ~new_new_n20134__;
  assign new_new_n20136__ = ~new_new_n19006__ & new_new_n19795__;
  assign new_new_n20137__ = ~new_new_n20135__ & ~new_new_n20136__;
  assign new_new_n20138__ = ~new_new_n18116__ & ~new_new_n20137__;
  assign new_new_n20139__ = ~new_new_n20132__ & ~new_new_n20138__;
  assign new_new_n20140__ = new_new_n18213__ & ~new_new_n20139__;
  assign new_new_n20141__ = ~ys__n1502 & ys__n27867;
  assign new_new_n20142__ = ~new_new_n18175__ & ~new_new_n18178__;
  assign new_new_n20143__ = ~ys__n23272 & ~new_new_n20142__;
  assign new_new_n20144__ = ys__n23272 & ~new_new_n20006__;
  assign new_new_n20145__ = ~new_new_n20143__ & ~new_new_n20144__;
  assign new_new_n20146__ = ~ys__n23274 & ~new_new_n20145__;
  assign new_new_n20147__ = ys__n23274 & ~new_new_n19873__;
  assign new_new_n20148__ = ~new_new_n20146__ & ~new_new_n20147__;
  assign new_new_n20149__ = ~ys__n23276 & ~new_new_n20148__;
  assign new_new_n20150__ = ys__n23276 & ~new_new_n19607__;
  assign new_new_n20151__ = ~new_new_n20149__ & ~new_new_n20150__;
  assign new_new_n20152__ = ~ys__n23278 & ~new_new_n20151__;
  assign new_new_n20153__ = ys__n23278 & new_new_n19021__;
  assign new_new_n20154__ = ~new_new_n20152__ & ~new_new_n20153__;
  assign new_new_n20155__ = ys__n1502 & ~new_new_n20154__;
  assign new_new_n20156__ = ~new_new_n20141__ & ~new_new_n20155__;
  assign new_new_n20157__ = ~new_new_n18213__ & ~new_new_n20156__;
  assign new_new_n20158__ = ~new_new_n20140__ & ~new_new_n20157__;
  assign new_new_n20159__ = new_new_n18224__ & ~new_new_n20158__;
  assign new_new_n20160__ = ~new_new_n10696__ & new_new_n18226__;
  assign new_new_n20161__ = ys__n1498 & new_new_n18345__;
  assign new_new_n20162__ = ~new_new_n20160__ & ~new_new_n20161__;
  assign new_new_n20163__ = ~ys__n1496 & ~new_new_n20162__;
  assign new_new_n20164__ = ys__n1496 & ~new_new_n18345__;
  assign new_new_n20165__ = ~new_new_n20163__ & ~new_new_n20164__;
  assign new_new_n20166__ = ~ys__n1495 & ~new_new_n20165__;
  assign new_new_n20167__ = ys__n1495 & new_new_n16769__;
  assign new_new_n20168__ = ~new_new_n20166__ & ~new_new_n20167__;
  assign new_new_n20169__ = ~new_new_n18224__ & ~new_new_n20168__;
  assign new_new_n20170__ = ~new_new_n20159__ & ~new_new_n20169__;
  assign new_new_n20171__ = new_new_n18581__ & ~new_new_n20170__;
  assign new_new_n20172__ = new_new_n18352__ & ~new_new_n20037__;
  assign new_new_n20173__ = new_new_n18376__ & ~new_new_n20172__;
  assign new_new_n20174__ = new_new_n18346__ & ~new_new_n20173__;
  assign new_new_n20175__ = ~new_new_n18346__ & new_new_n20173__;
  assign new_new_n20176__ = ~new_new_n20174__ & ~new_new_n20175__;
  assign new_new_n20177__ = ~ys__n1489 & ~new_new_n20176__;
  assign new_new_n20178__ = new_new_n16749__ & ~new_new_n20043__;
  assign new_new_n20179__ = new_new_n16766__ & ~new_new_n20178__;
  assign new_new_n20180__ = new_new_n10696__ & ~new_new_n20179__;
  assign new_new_n20181__ = ~new_new_n10696__ & new_new_n20179__;
  assign new_new_n20182__ = ~new_new_n20180__ & ~new_new_n20181__;
  assign new_new_n20183__ = ys__n1489 & ~new_new_n20182__;
  assign new_new_n20184__ = ~new_new_n20177__ & ~new_new_n20183__;
  assign new_new_n20185__ = ~new_new_n18427__ & ~new_new_n20184__;
  assign new_new_n20186__ = ~new_new_n20171__ & ~new_new_n20185__;
  assign new_new_n20187__ = ~ys__n19973 & ~new_new_n20186__;
  assign new_new_n20188__ = ys__n19973 & ys__n19995;
  assign new_new_n20189__ = ~new_new_n20187__ & ~new_new_n20188__;
  assign new_new_n20190__ = ~ys__n352 & ~new_new_n20189__;
  assign new_new_n20191__ = ~ys__n220 & ys__n47096;
  assign new_new_n20192__ = new_new_n18439__ & new_new_n20191__;
  assign new_new_n20193__ = new_new_n18441__ & new_new_n20191__;
  assign new_new_n20194__ = new_new_n18444__ & new_new_n19056__;
  assign new_new_n20195__ = ~new_new_n20193__ & ~new_new_n20194__;
  assign new_new_n20196__ = ~new_new_n20192__ & new_new_n20195__;
  assign new_new_n20197__ = new_new_n18453__ & ~new_new_n20196__;
  assign ys__n19944 = new_new_n20190__ | new_new_n20197__;
  assign new_new_n20199__ = ys__n19844 & ys__n19867;
  assign new_new_n20200__ = new_new_n18116__ & new_new_n20199__;
  assign new_new_n20201__ = ~ys__n23278 & ~new_new_n19083__;
  assign new_new_n20202__ = ~new_new_n19661__ & ~new_new_n20201__;
  assign new_new_n20203__ = ~ys__n1505 & ~new_new_n20202__;
  assign new_new_n20204__ = ~new_new_n19089__ & new_new_n19795__;
  assign new_new_n20205__ = ~new_new_n20203__ & ~new_new_n20204__;
  assign new_new_n20206__ = ~new_new_n18116__ & ~new_new_n20205__;
  assign new_new_n20207__ = ~new_new_n20200__ & ~new_new_n20206__;
  assign new_new_n20208__ = new_new_n18213__ & ~new_new_n20207__;
  assign new_new_n20209__ = ~ys__n1502 & ys__n27869;
  assign new_new_n20210__ = ~new_new_n18515__ & ~new_new_n18518__;
  assign new_new_n20211__ = ~ys__n23272 & ~new_new_n20210__;
  assign new_new_n20212__ = ys__n23272 & ~new_new_n20074__;
  assign new_new_n20213__ = ~new_new_n20211__ & ~new_new_n20212__;
  assign new_new_n20214__ = ~ys__n23274 & ~new_new_n20213__;
  assign new_new_n20215__ = ys__n23274 & ~new_new_n19941__;
  assign new_new_n20216__ = ~new_new_n20214__ & ~new_new_n20215__;
  assign new_new_n20217__ = ~ys__n23276 & ~new_new_n20216__;
  assign new_new_n20218__ = ys__n23276 & ~new_new_n19678__;
  assign new_new_n20219__ = ~new_new_n20217__ & ~new_new_n20218__;
  assign new_new_n20220__ = ~ys__n23278 & ~new_new_n20219__;
  assign new_new_n20221__ = ys__n23278 & new_new_n19104__;
  assign new_new_n20222__ = ~new_new_n20220__ & ~new_new_n20221__;
  assign new_new_n20223__ = ys__n1502 & ~new_new_n20222__;
  assign new_new_n20224__ = ~new_new_n20209__ & ~new_new_n20223__;
  assign new_new_n20225__ = ~new_new_n18213__ & ~new_new_n20224__;
  assign new_new_n20226__ = ~new_new_n20208__ & ~new_new_n20225__;
  assign new_new_n20227__ = new_new_n18224__ & ~new_new_n20226__;
  assign new_new_n20228__ = ~new_new_n10699__ & new_new_n18226__;
  assign new_new_n20229__ = ys__n1498 & new_new_n18343__;
  assign new_new_n20230__ = ~new_new_n20228__ & ~new_new_n20229__;
  assign new_new_n20231__ = ~ys__n1496 & ~new_new_n20230__;
  assign new_new_n20232__ = ys__n1496 & ~new_new_n18343__;
  assign new_new_n20233__ = ~new_new_n20231__ & ~new_new_n20232__;
  assign new_new_n20234__ = ~ys__n1495 & ~new_new_n20233__;
  assign new_new_n20235__ = ys__n1495 & new_new_n16768__;
  assign new_new_n20236__ = ~new_new_n20234__ & ~new_new_n20235__;
  assign new_new_n20237__ = ~new_new_n18224__ & ~new_new_n20236__;
  assign new_new_n20238__ = ~new_new_n20227__ & ~new_new_n20237__;
  assign new_new_n20239__ = new_new_n18581__ & ~new_new_n20238__;
  assign new_new_n20240__ = ~new_new_n18346__ & ~new_new_n20173__;
  assign new_new_n20241__ = ~new_new_n10695__ & ~new_new_n20240__;
  assign new_new_n20242__ = new_new_n18344__ & ~new_new_n20241__;
  assign new_new_n20243__ = ~new_new_n18344__ & new_new_n20241__;
  assign new_new_n20244__ = ~new_new_n20242__ & ~new_new_n20243__;
  assign new_new_n20245__ = ~ys__n1489 & ~new_new_n20244__;
  assign new_new_n20246__ = ~new_new_n10696__ & ~new_new_n20179__;
  assign new_new_n20247__ = ~new_new_n16769__ & ~new_new_n20246__;
  assign new_new_n20248__ = new_new_n10699__ & ~new_new_n20247__;
  assign new_new_n20249__ = ~new_new_n10699__ & new_new_n20247__;
  assign new_new_n20250__ = ~new_new_n20248__ & ~new_new_n20249__;
  assign new_new_n20251__ = ys__n1489 & ~new_new_n20250__;
  assign new_new_n20252__ = ~new_new_n20245__ & ~new_new_n20251__;
  assign new_new_n20253__ = ~new_new_n18427__ & ~new_new_n20252__;
  assign new_new_n20254__ = ~new_new_n20239__ & ~new_new_n20253__;
  assign new_new_n20255__ = ~ys__n19973 & ~new_new_n20254__;
  assign new_new_n20256__ = ys__n19973 & ys__n19996;
  assign new_new_n20257__ = ~new_new_n20255__ & ~new_new_n20256__;
  assign new_new_n20258__ = ~ys__n352 & ~new_new_n20257__;
  assign new_new_n20259__ = ~ys__n220 & ys__n47097;
  assign new_new_n20260__ = new_new_n18439__ & new_new_n20259__;
  assign new_new_n20261__ = new_new_n18441__ & new_new_n20259__;
  assign new_new_n20262__ = new_new_n18444__ & new_new_n19139__;
  assign new_new_n20263__ = ~new_new_n20261__ & ~new_new_n20262__;
  assign new_new_n20264__ = ~new_new_n20260__ & new_new_n20263__;
  assign new_new_n20265__ = new_new_n18453__ & ~new_new_n20264__;
  assign ys__n19947 = new_new_n20258__ | new_new_n20265__;
  assign new_new_n20267__ = ys__n19844 & ys__n19868;
  assign new_new_n20268__ = new_new_n18116__ & new_new_n20267__;
  assign new_new_n20269__ = ~ys__n23278 & ~new_new_n19156__;
  assign new_new_n20270__ = ~new_new_n19661__ & ~new_new_n20269__;
  assign new_new_n20271__ = ~ys__n1505 & ~new_new_n20270__;
  assign new_new_n20272__ = new_new_n19155__ & new_new_n19795__;
  assign new_new_n20273__ = ~new_new_n20271__ & ~new_new_n20272__;
  assign new_new_n20274__ = ~new_new_n18116__ & ~new_new_n20273__;
  assign new_new_n20275__ = ~new_new_n20268__ & ~new_new_n20274__;
  assign new_new_n20276__ = new_new_n18213__ & ~new_new_n20275__;
  assign new_new_n20277__ = ~ys__n1502 & ys__n27871;
  assign new_new_n20278__ = ~new_new_n18179__ & ~new_new_n18186__;
  assign new_new_n20279__ = ~ys__n23272 & ~new_new_n20278__;
  assign new_new_n20280__ = ys__n23272 & ~new_new_n20142__;
  assign new_new_n20281__ = ~new_new_n20279__ & ~new_new_n20280__;
  assign new_new_n20282__ = ~ys__n23274 & ~new_new_n20281__;
  assign new_new_n20283__ = ys__n23274 & ~new_new_n20009__;
  assign new_new_n20284__ = ~new_new_n20282__ & ~new_new_n20283__;
  assign new_new_n20285__ = ~ys__n23276 & ~new_new_n20284__;
  assign new_new_n20286__ = ys__n23276 & ~new_new_n19743__;
  assign new_new_n20287__ = ~new_new_n20285__ & ~new_new_n20286__;
  assign new_new_n20288__ = ~ys__n23278 & ~new_new_n20287__;
  assign new_new_n20289__ = ys__n23278 & ~new_new_n19176__;
  assign new_new_n20290__ = ~new_new_n20288__ & ~new_new_n20289__;
  assign new_new_n20291__ = ys__n1502 & ~new_new_n20290__;
  assign new_new_n20292__ = ~new_new_n20277__ & ~new_new_n20291__;
  assign new_new_n20293__ = ~new_new_n18213__ & ~new_new_n20292__;
  assign new_new_n20294__ = ~new_new_n20276__ & ~new_new_n20293__;
  assign new_new_n20295__ = new_new_n18224__ & ~new_new_n20294__;
  assign new_new_n20296__ = ~new_new_n10735__ & new_new_n18226__;
  assign new_new_n20297__ = ys__n1498 & new_new_n18338__;
  assign new_new_n20298__ = ~new_new_n20296__ & ~new_new_n20297__;
  assign new_new_n20299__ = ~ys__n1496 & ~new_new_n20298__;
  assign new_new_n20300__ = ys__n1496 & ~new_new_n18338__;
  assign new_new_n20301__ = ~new_new_n20299__ & ~new_new_n20300__;
  assign new_new_n20302__ = ~ys__n1495 & ~new_new_n20301__;
  assign new_new_n20303__ = ys__n1495 & new_new_n16737__;
  assign new_new_n20304__ = ~new_new_n20302__ & ~new_new_n20303__;
  assign new_new_n20305__ = ~new_new_n18224__ & ~new_new_n20304__;
  assign new_new_n20306__ = ~new_new_n20295__ & ~new_new_n20305__;
  assign new_new_n20307__ = new_new_n18581__ & ~new_new_n20306__;
  assign new_new_n20308__ = ~new_new_n18318__ & new_new_n18365__;
  assign new_new_n20309__ = new_new_n18381__ & ~new_new_n20308__;
  assign new_new_n20310__ = new_new_n18339__ & ~new_new_n20309__;
  assign new_new_n20311__ = ~new_new_n18339__ & new_new_n20309__;
  assign new_new_n20312__ = ~new_new_n20310__ & ~new_new_n20311__;
  assign new_new_n20313__ = ~ys__n1489 & ~new_new_n20312__;
  assign new_new_n20314__ = new_new_n10735__ & ~new_new_n16834__;
  assign new_new_n20315__ = ~new_new_n10735__ & new_new_n16834__;
  assign new_new_n20316__ = ~new_new_n20314__ & ~new_new_n20315__;
  assign new_new_n20317__ = ys__n1489 & ~new_new_n20316__;
  assign new_new_n20318__ = ~new_new_n20313__ & ~new_new_n20317__;
  assign new_new_n20319__ = ~new_new_n18427__ & ~new_new_n20318__;
  assign new_new_n20320__ = ~new_new_n20307__ & ~new_new_n20319__;
  assign new_new_n20321__ = ~ys__n19973 & ~new_new_n20320__;
  assign new_new_n20322__ = ys__n19973 & ys__n19997;
  assign new_new_n20323__ = ~new_new_n20321__ & ~new_new_n20322__;
  assign new_new_n20324__ = ~ys__n352 & ~new_new_n20323__;
  assign new_new_n20325__ = ~ys__n220 & ys__n47098;
  assign new_new_n20326__ = new_new_n18439__ & new_new_n20325__;
  assign new_new_n20327__ = new_new_n18441__ & new_new_n20325__;
  assign new_new_n20328__ = new_new_n18444__ & new_new_n19207__;
  assign new_new_n20329__ = ~new_new_n20327__ & ~new_new_n20328__;
  assign new_new_n20330__ = ~new_new_n20326__ & new_new_n20329__;
  assign new_new_n20331__ = new_new_n18453__ & ~new_new_n20330__;
  assign ys__n19950 = new_new_n20324__ | new_new_n20331__;
  assign new_new_n20333__ = ys__n19844 & ys__n19869;
  assign new_new_n20334__ = new_new_n18116__ & new_new_n20333__;
  assign new_new_n20335__ = ~ys__n23278 & ~new_new_n19224__;
  assign new_new_n20336__ = ~new_new_n19661__ & ~new_new_n20335__;
  assign new_new_n20337__ = ~ys__n1505 & ~new_new_n20336__;
  assign new_new_n20338__ = new_new_n19228__ & new_new_n19795__;
  assign new_new_n20339__ = ~new_new_n20337__ & ~new_new_n20338__;
  assign new_new_n20340__ = ~new_new_n18116__ & ~new_new_n20339__;
  assign new_new_n20341__ = ~new_new_n20334__ & ~new_new_n20340__;
  assign new_new_n20342__ = new_new_n18213__ & ~new_new_n20341__;
  assign new_new_n20343__ = ~ys__n1502 & ys__n27873;
  assign new_new_n20344__ = ~new_new_n18519__ & ~new_new_n18526__;
  assign new_new_n20345__ = ~ys__n23272 & ~new_new_n20344__;
  assign new_new_n20346__ = ys__n23272 & ~new_new_n20210__;
  assign new_new_n20347__ = ~new_new_n20345__ & ~new_new_n20346__;
  assign new_new_n20348__ = ~ys__n23274 & ~new_new_n20347__;
  assign new_new_n20349__ = ys__n23274 & ~new_new_n20077__;
  assign new_new_n20350__ = ~new_new_n20348__ & ~new_new_n20349__;
  assign new_new_n20351__ = ~ys__n23276 & ~new_new_n20350__;
  assign new_new_n20352__ = ys__n23276 & ~new_new_n19808__;
  assign new_new_n20353__ = ~new_new_n20351__ & ~new_new_n20352__;
  assign new_new_n20354__ = ~ys__n23278 & ~new_new_n20353__;
  assign new_new_n20355__ = ys__n23278 & ~new_new_n19245__;
  assign new_new_n20356__ = ~new_new_n20354__ & ~new_new_n20355__;
  assign new_new_n20357__ = ys__n1502 & ~new_new_n20356__;
  assign new_new_n20358__ = ~new_new_n20343__ & ~new_new_n20357__;
  assign new_new_n20359__ = ~new_new_n18213__ & ~new_new_n20358__;
  assign new_new_n20360__ = ~new_new_n20342__ & ~new_new_n20359__;
  assign new_new_n20361__ = new_new_n18224__ & ~new_new_n20360__;
  assign new_new_n20362__ = ~new_new_n10738__ & new_new_n18226__;
  assign new_new_n20363__ = ys__n1498 & new_new_n18336__;
  assign new_new_n20364__ = ~new_new_n20362__ & ~new_new_n20363__;
  assign new_new_n20365__ = ~ys__n1496 & ~new_new_n20364__;
  assign new_new_n20366__ = ys__n1496 & ~new_new_n18336__;
  assign new_new_n20367__ = ~new_new_n20365__ & ~new_new_n20366__;
  assign new_new_n20368__ = ~ys__n1495 & ~new_new_n20367__;
  assign new_new_n20369__ = ys__n1495 & new_new_n16736__;
  assign new_new_n20370__ = ~new_new_n20368__ & ~new_new_n20369__;
  assign new_new_n20371__ = ~new_new_n18224__ & ~new_new_n20370__;
  assign new_new_n20372__ = ~new_new_n20361__ & ~new_new_n20371__;
  assign new_new_n20373__ = new_new_n18581__ & ~new_new_n20372__;
  assign new_new_n20374__ = ~new_new_n18339__ & ~new_new_n20309__;
  assign new_new_n20375__ = ~new_new_n10734__ & ~new_new_n20374__;
  assign new_new_n20376__ = new_new_n18337__ & ~new_new_n20375__;
  assign new_new_n20377__ = ~new_new_n18337__ & new_new_n20375__;
  assign new_new_n20378__ = ~new_new_n20376__ & ~new_new_n20377__;
  assign new_new_n20379__ = ~ys__n1489 & ~new_new_n20378__;
  assign new_new_n20380__ = ~new_new_n10735__ & ~new_new_n16834__;
  assign new_new_n20381__ = ~new_new_n16737__ & ~new_new_n20380__;
  assign new_new_n20382__ = new_new_n10738__ & ~new_new_n20381__;
  assign new_new_n20383__ = ~new_new_n10738__ & new_new_n20381__;
  assign new_new_n20384__ = ~new_new_n20382__ & ~new_new_n20383__;
  assign new_new_n20385__ = ys__n1489 & ~new_new_n20384__;
  assign new_new_n20386__ = ~new_new_n20379__ & ~new_new_n20385__;
  assign new_new_n20387__ = ~new_new_n18427__ & ~new_new_n20386__;
  assign new_new_n20388__ = ~new_new_n20373__ & ~new_new_n20387__;
  assign new_new_n20389__ = ~ys__n19973 & ~new_new_n20388__;
  assign new_new_n20390__ = ys__n19973 & ys__n19998;
  assign new_new_n20391__ = ~new_new_n20389__ & ~new_new_n20390__;
  assign new_new_n20392__ = ~ys__n352 & ~new_new_n20391__;
  assign new_new_n20393__ = ~ys__n220 & ys__n47099;
  assign new_new_n20394__ = new_new_n18439__ & new_new_n20393__;
  assign new_new_n20395__ = new_new_n18441__ & new_new_n20393__;
  assign new_new_n20396__ = new_new_n18444__ & new_new_n19280__;
  assign new_new_n20397__ = ~new_new_n20395__ & ~new_new_n20396__;
  assign new_new_n20398__ = ~new_new_n20394__ & new_new_n20397__;
  assign new_new_n20399__ = new_new_n18453__ & ~new_new_n20398__;
  assign ys__n19953 = new_new_n20392__ | new_new_n20399__;
  assign new_new_n20401__ = ys__n19844 & ys__n19870;
  assign new_new_n20402__ = new_new_n18116__ & new_new_n20401__;
  assign new_new_n20403__ = ~ys__n23278 & ~new_new_n19297__;
  assign new_new_n20404__ = ~new_new_n19661__ & ~new_new_n20403__;
  assign new_new_n20405__ = ~ys__n1505 & ~new_new_n20404__;
  assign new_new_n20406__ = new_new_n19301__ & new_new_n19795__;
  assign new_new_n20407__ = ~new_new_n20405__ & ~new_new_n20406__;
  assign new_new_n20408__ = ~new_new_n18116__ & ~new_new_n20407__;
  assign new_new_n20409__ = ~new_new_n20402__ & ~new_new_n20408__;
  assign new_new_n20410__ = new_new_n18213__ & ~new_new_n20409__;
  assign new_new_n20411__ = ~ys__n1502 & ys__n27875;
  assign new_new_n20412__ = ~new_new_n18187__ & ~new_new_n18190__;
  assign new_new_n20413__ = ~ys__n23272 & ~new_new_n20412__;
  assign new_new_n20414__ = ys__n23272 & ~new_new_n20278__;
  assign new_new_n20415__ = ~new_new_n20413__ & ~new_new_n20414__;
  assign new_new_n20416__ = ~ys__n23274 & ~new_new_n20415__;
  assign new_new_n20417__ = ys__n23274 & ~new_new_n20145__;
  assign new_new_n20418__ = ~new_new_n20416__ & ~new_new_n20417__;
  assign new_new_n20419__ = ~ys__n23276 & ~new_new_n20418__;
  assign new_new_n20420__ = ys__n23276 & ~new_new_n19876__;
  assign new_new_n20421__ = ~new_new_n20419__ & ~new_new_n20420__;
  assign new_new_n20422__ = ~ys__n23278 & ~new_new_n20421__;
  assign new_new_n20423__ = ys__n23278 & ~new_new_n19318__;
  assign new_new_n20424__ = ~new_new_n20422__ & ~new_new_n20423__;
  assign new_new_n20425__ = ys__n1502 & ~new_new_n20424__;
  assign new_new_n20426__ = ~new_new_n20411__ & ~new_new_n20425__;
  assign new_new_n20427__ = ~new_new_n18213__ & ~new_new_n20426__;
  assign new_new_n20428__ = ~new_new_n20410__ & ~new_new_n20427__;
  assign new_new_n20429__ = new_new_n18224__ & ~new_new_n20428__;
  assign new_new_n20430__ = ~new_new_n10742__ & new_new_n18226__;
  assign new_new_n20431__ = ys__n1498 & new_new_n18333__;
  assign new_new_n20432__ = ~new_new_n20430__ & ~new_new_n20431__;
  assign new_new_n20433__ = ~ys__n1496 & ~new_new_n20432__;
  assign new_new_n20434__ = ys__n1496 & ~new_new_n18333__;
  assign new_new_n20435__ = ~new_new_n20433__ & ~new_new_n20434__;
  assign new_new_n20436__ = ~ys__n1495 & ~new_new_n20435__;
  assign new_new_n20437__ = ys__n1495 & new_new_n16742__;
  assign new_new_n20438__ = ~new_new_n20436__ & ~new_new_n20437__;
  assign new_new_n20439__ = ~new_new_n18224__ & ~new_new_n20438__;
  assign new_new_n20440__ = ~new_new_n20429__ & ~new_new_n20439__;
  assign new_new_n20441__ = new_new_n18581__ & ~new_new_n20440__;
  assign new_new_n20442__ = new_new_n18340__ & ~new_new_n20309__;
  assign new_new_n20443__ = new_new_n18384__ & ~new_new_n20442__;
  assign new_new_n20444__ = new_new_n18334__ & ~new_new_n20443__;
  assign new_new_n20445__ = ~new_new_n18334__ & new_new_n20443__;
  assign new_new_n20446__ = ~new_new_n20444__ & ~new_new_n20445__;
  assign new_new_n20447__ = ~ys__n1489 & ~new_new_n20446__;
  assign new_new_n20448__ = new_new_n16746__ & ~new_new_n16834__;
  assign new_new_n20449__ = new_new_n16739__ & ~new_new_n20448__;
  assign new_new_n20450__ = new_new_n10742__ & ~new_new_n20449__;
  assign new_new_n20451__ = ~new_new_n10742__ & new_new_n20449__;
  assign new_new_n20452__ = ~new_new_n20450__ & ~new_new_n20451__;
  assign new_new_n20453__ = ys__n1489 & ~new_new_n20452__;
  assign new_new_n20454__ = ~new_new_n20447__ & ~new_new_n20453__;
  assign new_new_n20455__ = ~new_new_n18427__ & ~new_new_n20454__;
  assign new_new_n20456__ = ~new_new_n20441__ & ~new_new_n20455__;
  assign new_new_n20457__ = ~ys__n19973 & ~new_new_n20456__;
  assign new_new_n20458__ = ys__n19973 & ys__n19999;
  assign new_new_n20459__ = ~new_new_n20457__ & ~new_new_n20458__;
  assign new_new_n20460__ = ~ys__n352 & ~new_new_n20459__;
  assign new_new_n20461__ = ~ys__n220 & ys__n47100;
  assign new_new_n20462__ = new_new_n18439__ & new_new_n20461__;
  assign new_new_n20463__ = new_new_n18441__ & new_new_n20461__;
  assign new_new_n20464__ = new_new_n18444__ & new_new_n19353__;
  assign new_new_n20465__ = ~new_new_n20463__ & ~new_new_n20464__;
  assign new_new_n20466__ = ~new_new_n20462__ & new_new_n20465__;
  assign new_new_n20467__ = new_new_n18453__ & ~new_new_n20466__;
  assign ys__n19956 = new_new_n20460__ | new_new_n20467__;
  assign new_new_n20469__ = ys__n19844 & ys__n19871;
  assign new_new_n20470__ = new_new_n18116__ & new_new_n20469__;
  assign new_new_n20471__ = ~ys__n23278 & ~new_new_n19370__;
  assign new_new_n20472__ = ~new_new_n19661__ & ~new_new_n20471__;
  assign new_new_n20473__ = ~ys__n1505 & ~new_new_n20472__;
  assign new_new_n20474__ = new_new_n19374__ & new_new_n19795__;
  assign new_new_n20475__ = ~new_new_n20473__ & ~new_new_n20474__;
  assign new_new_n20476__ = ~new_new_n18116__ & ~new_new_n20475__;
  assign new_new_n20477__ = ~new_new_n20470__ & ~new_new_n20476__;
  assign new_new_n20478__ = new_new_n18213__ & ~new_new_n20477__;
  assign new_new_n20479__ = ~ys__n1502 & ys__n27877;
  assign new_new_n20480__ = ~new_new_n18527__ & ~new_new_n18530__;
  assign new_new_n20481__ = ~ys__n23272 & ~new_new_n20480__;
  assign new_new_n20482__ = ys__n23272 & ~new_new_n20344__;
  assign new_new_n20483__ = ~new_new_n20481__ & ~new_new_n20482__;
  assign new_new_n20484__ = ~ys__n23274 & ~new_new_n20483__;
  assign new_new_n20485__ = ys__n23274 & ~new_new_n20213__;
  assign new_new_n20486__ = ~new_new_n20484__ & ~new_new_n20485__;
  assign new_new_n20487__ = ~ys__n23276 & ~new_new_n20486__;
  assign new_new_n20488__ = ys__n23276 & ~new_new_n19944__;
  assign new_new_n20489__ = ~new_new_n20487__ & ~new_new_n20488__;
  assign new_new_n20490__ = ~ys__n23278 & ~new_new_n20489__;
  assign new_new_n20491__ = ys__n23278 & ~new_new_n19391__;
  assign new_new_n20492__ = ~new_new_n20490__ & ~new_new_n20491__;
  assign new_new_n20493__ = ys__n1502 & ~new_new_n20492__;
  assign new_new_n20494__ = ~new_new_n20479__ & ~new_new_n20493__;
  assign new_new_n20495__ = ~new_new_n18213__ & ~new_new_n20494__;
  assign new_new_n20496__ = ~new_new_n20478__ & ~new_new_n20495__;
  assign new_new_n20497__ = new_new_n18224__ & ~new_new_n20496__;
  assign new_new_n20498__ = ~new_new_n10745__ & new_new_n18226__;
  assign new_new_n20499__ = ys__n1498 & new_new_n18331__;
  assign new_new_n20500__ = ~new_new_n20498__ & ~new_new_n20499__;
  assign new_new_n20501__ = ~ys__n1496 & ~new_new_n20500__;
  assign new_new_n20502__ = ys__n1496 & ~new_new_n18331__;
  assign new_new_n20503__ = ~new_new_n20501__ & ~new_new_n20502__;
  assign new_new_n20504__ = ~ys__n1495 & ~new_new_n20503__;
  assign new_new_n20505__ = ys__n1495 & new_new_n16741__;
  assign new_new_n20506__ = ~new_new_n20504__ & ~new_new_n20505__;
  assign new_new_n20507__ = ~new_new_n18224__ & ~new_new_n20506__;
  assign new_new_n20508__ = ~new_new_n20497__ & ~new_new_n20507__;
  assign new_new_n20509__ = new_new_n18581__ & ~new_new_n20508__;
  assign new_new_n20510__ = ~new_new_n18334__ & ~new_new_n20443__;
  assign new_new_n20511__ = ~new_new_n10741__ & ~new_new_n20510__;
  assign new_new_n20512__ = new_new_n18332__ & ~new_new_n20511__;
  assign new_new_n20513__ = ~new_new_n18332__ & new_new_n20511__;
  assign new_new_n20514__ = ~new_new_n20512__ & ~new_new_n20513__;
  assign new_new_n20515__ = ~ys__n1489 & ~new_new_n20514__;
  assign new_new_n20516__ = ~new_new_n10742__ & ~new_new_n20449__;
  assign new_new_n20517__ = ~new_new_n16742__ & ~new_new_n20516__;
  assign new_new_n20518__ = new_new_n10745__ & ~new_new_n20517__;
  assign new_new_n20519__ = ~new_new_n10745__ & new_new_n20517__;
  assign new_new_n20520__ = ~new_new_n20518__ & ~new_new_n20519__;
  assign new_new_n20521__ = ys__n1489 & ~new_new_n20520__;
  assign new_new_n20522__ = ~new_new_n20515__ & ~new_new_n20521__;
  assign new_new_n20523__ = ~new_new_n18427__ & ~new_new_n20522__;
  assign new_new_n20524__ = ~new_new_n20509__ & ~new_new_n20523__;
  assign new_new_n20525__ = ~ys__n19973 & ~new_new_n20524__;
  assign new_new_n20526__ = ys__n19973 & ys__n20000;
  assign new_new_n20527__ = ~new_new_n20525__ & ~new_new_n20526__;
  assign new_new_n20528__ = ~ys__n352 & ~new_new_n20527__;
  assign new_new_n20529__ = ~ys__n220 & ys__n47101;
  assign new_new_n20530__ = new_new_n18439__ & new_new_n20529__;
  assign new_new_n20531__ = new_new_n18441__ & new_new_n20529__;
  assign new_new_n20532__ = new_new_n18444__ & new_new_n19426__;
  assign new_new_n20533__ = ~new_new_n20531__ & ~new_new_n20532__;
  assign new_new_n20534__ = ~new_new_n20530__ & new_new_n20533__;
  assign new_new_n20535__ = new_new_n18453__ & ~new_new_n20534__;
  assign ys__n19959 = new_new_n20528__ | new_new_n20535__;
  assign new_new_n20537__ = ys__n19844 & ys__n19872;
  assign new_new_n20538__ = new_new_n18116__ & new_new_n20537__;
  assign new_new_n20539__ = ~ys__n23278 & ~new_new_n19443__;
  assign new_new_n20540__ = ~new_new_n19661__ & ~new_new_n20539__;
  assign new_new_n20541__ = ~ys__n1505 & ~new_new_n20540__;
  assign new_new_n20542__ = new_new_n19447__ & new_new_n19795__;
  assign new_new_n20543__ = ~new_new_n20541__ & ~new_new_n20542__;
  assign new_new_n20544__ = ~new_new_n18116__ & ~new_new_n20543__;
  assign new_new_n20545__ = ~new_new_n20538__ & ~new_new_n20544__;
  assign new_new_n20546__ = new_new_n18213__ & ~new_new_n20545__;
  assign new_new_n20547__ = ~ys__n1502 & ys__n27879;
  assign new_new_n20548__ = ~new_new_n18191__ & ~new_new_n18196__;
  assign new_new_n20549__ = ~ys__n23272 & ~new_new_n20548__;
  assign new_new_n20550__ = ys__n23272 & ~new_new_n20412__;
  assign new_new_n20551__ = ~new_new_n20549__ & ~new_new_n20550__;
  assign new_new_n20552__ = ~ys__n23274 & ~new_new_n20551__;
  assign new_new_n20553__ = ys__n23274 & ~new_new_n20281__;
  assign new_new_n20554__ = ~new_new_n20552__ & ~new_new_n20553__;
  assign new_new_n20555__ = ~ys__n23276 & ~new_new_n20554__;
  assign new_new_n20556__ = ys__n23276 & ~new_new_n20012__;
  assign new_new_n20557__ = ~new_new_n20555__ & ~new_new_n20556__;
  assign new_new_n20558__ = ~ys__n23278 & ~new_new_n20557__;
  assign new_new_n20559__ = ys__n23278 & ~new_new_n19464__;
  assign new_new_n20560__ = ~new_new_n20558__ & ~new_new_n20559__;
  assign new_new_n20561__ = ys__n1502 & ~new_new_n20560__;
  assign new_new_n20562__ = ~new_new_n20547__ & ~new_new_n20561__;
  assign new_new_n20563__ = ~new_new_n18213__ & ~new_new_n20562__;
  assign new_new_n20564__ = ~new_new_n20546__ & ~new_new_n20563__;
  assign new_new_n20565__ = new_new_n18224__ & ~new_new_n20564__;
  assign new_new_n20566__ = ~new_new_n10720__ & new_new_n18226__;
  assign new_new_n20567__ = ys__n1498 & new_new_n18327__;
  assign new_new_n20568__ = ~new_new_n20566__ & ~new_new_n20567__;
  assign new_new_n20569__ = ~ys__n1496 & ~new_new_n20568__;
  assign new_new_n20570__ = ys__n1496 & ~new_new_n18327__;
  assign new_new_n20571__ = ~new_new_n20569__ & ~new_new_n20570__;
  assign new_new_n20572__ = ~ys__n1495 & ~new_new_n20571__;
  assign new_new_n20573__ = ys__n1495 & new_new_n16734__;
  assign new_new_n20574__ = ~new_new_n20572__ & ~new_new_n20573__;
  assign new_new_n20575__ = ~new_new_n18224__ & ~new_new_n20574__;
  assign new_new_n20576__ = ~new_new_n20565__ & ~new_new_n20575__;
  assign new_new_n20577__ = new_new_n18581__ & ~new_new_n20576__;
  assign new_new_n20578__ = new_new_n18341__ & ~new_new_n20309__;
  assign new_new_n20579__ = new_new_n18388__ & ~new_new_n20578__;
  assign new_new_n20580__ = new_new_n18328__ & ~new_new_n20579__;
  assign new_new_n20581__ = ~new_new_n18328__ & new_new_n20579__;
  assign new_new_n20582__ = ~new_new_n20580__ & ~new_new_n20581__;
  assign new_new_n20583__ = ~ys__n1489 & ~new_new_n20582__;
  assign new_new_n20584__ = new_new_n10720__ & ~new_new_n16836__;
  assign new_new_n20585__ = ~new_new_n10720__ & new_new_n16836__;
  assign new_new_n20586__ = ~new_new_n20584__ & ~new_new_n20585__;
  assign new_new_n20587__ = ys__n1489 & ~new_new_n20586__;
  assign new_new_n20588__ = ~new_new_n20583__ & ~new_new_n20587__;
  assign new_new_n20589__ = ~new_new_n18427__ & ~new_new_n20588__;
  assign new_new_n20590__ = ~new_new_n20577__ & ~new_new_n20589__;
  assign new_new_n20591__ = ~ys__n19973 & ~new_new_n20590__;
  assign new_new_n20592__ = ys__n19973 & ys__n20001;
  assign new_new_n20593__ = ~new_new_n20591__ & ~new_new_n20592__;
  assign new_new_n20594__ = ~ys__n352 & ~new_new_n20593__;
  assign new_new_n20595__ = ~ys__n220 & ys__n47102;
  assign new_new_n20596__ = new_new_n18439__ & new_new_n20595__;
  assign new_new_n20597__ = new_new_n18441__ & new_new_n20595__;
  assign new_new_n20598__ = new_new_n18444__ & new_new_n19499__;
  assign new_new_n20599__ = ~new_new_n20597__ & ~new_new_n20598__;
  assign new_new_n20600__ = ~new_new_n20596__ & new_new_n20599__;
  assign new_new_n20601__ = new_new_n18453__ & ~new_new_n20600__;
  assign ys__n19962 = new_new_n20594__ | new_new_n20601__;
  assign new_new_n20603__ = ys__n19844 & ys__n19873;
  assign new_new_n20604__ = new_new_n18116__ & new_new_n20603__;
  assign new_new_n20605__ = ~ys__n23278 & ~new_new_n19516__;
  assign new_new_n20606__ = ~new_new_n19661__ & ~new_new_n20605__;
  assign new_new_n20607__ = ~ys__n1505 & ~new_new_n20606__;
  assign new_new_n20608__ = new_new_n19520__ & new_new_n19795__;
  assign new_new_n20609__ = ~new_new_n20607__ & ~new_new_n20608__;
  assign new_new_n20610__ = ~new_new_n18116__ & ~new_new_n20609__;
  assign new_new_n20611__ = ~new_new_n20604__ & ~new_new_n20610__;
  assign new_new_n20612__ = new_new_n18213__ & ~new_new_n20611__;
  assign new_new_n20613__ = ~ys__n1502 & ys__n27881;
  assign new_new_n20614__ = ~new_new_n18531__ & ~new_new_n18536__;
  assign new_new_n20615__ = ~ys__n23272 & ~new_new_n20614__;
  assign new_new_n20616__ = ys__n23272 & ~new_new_n20480__;
  assign new_new_n20617__ = ~new_new_n20615__ & ~new_new_n20616__;
  assign new_new_n20618__ = ~ys__n23274 & ~new_new_n20617__;
  assign new_new_n20619__ = ys__n23274 & ~new_new_n20347__;
  assign new_new_n20620__ = ~new_new_n20618__ & ~new_new_n20619__;
  assign new_new_n20621__ = ~ys__n23276 & ~new_new_n20620__;
  assign new_new_n20622__ = ys__n23276 & ~new_new_n20080__;
  assign new_new_n20623__ = ~new_new_n20621__ & ~new_new_n20622__;
  assign new_new_n20624__ = ~ys__n23278 & ~new_new_n20623__;
  assign new_new_n20625__ = ys__n23278 & ~new_new_n19537__;
  assign new_new_n20626__ = ~new_new_n20624__ & ~new_new_n20625__;
  assign new_new_n20627__ = ys__n1502 & ~new_new_n20626__;
  assign new_new_n20628__ = ~new_new_n20613__ & ~new_new_n20627__;
  assign new_new_n20629__ = ~new_new_n18213__ & ~new_new_n20628__;
  assign new_new_n20630__ = ~new_new_n20612__ & ~new_new_n20629__;
  assign new_new_n20631__ = new_new_n18224__ & ~new_new_n20630__;
  assign new_new_n20632__ = ~new_new_n10723__ & new_new_n18226__;
  assign new_new_n20633__ = ys__n1498 & new_new_n18325__;
  assign new_new_n20634__ = ~new_new_n20632__ & ~new_new_n20633__;
  assign new_new_n20635__ = ~ys__n1496 & ~new_new_n20634__;
  assign new_new_n20636__ = ys__n1496 & ~new_new_n18325__;
  assign new_new_n20637__ = ~new_new_n20635__ & ~new_new_n20636__;
  assign new_new_n20638__ = ~ys__n1495 & ~new_new_n20637__;
  assign new_new_n20639__ = ys__n1495 & new_new_n16844__;
  assign new_new_n20640__ = ~new_new_n20638__ & ~new_new_n20639__;
  assign new_new_n20641__ = ~new_new_n18224__ & ~new_new_n20640__;
  assign new_new_n20642__ = ~new_new_n20631__ & ~new_new_n20641__;
  assign new_new_n20643__ = new_new_n18581__ & ~new_new_n20642__;
  assign new_new_n20644__ = ~new_new_n18328__ & ~new_new_n20579__;
  assign new_new_n20645__ = ~new_new_n10719__ & ~new_new_n20644__;
  assign new_new_n20646__ = new_new_n18326__ & ~new_new_n20645__;
  assign new_new_n20647__ = ~new_new_n18326__ & new_new_n20645__;
  assign new_new_n20648__ = ~new_new_n20646__ & ~new_new_n20647__;
  assign new_new_n20649__ = ~ys__n1489 & ~new_new_n20648__;
  assign new_new_n20650__ = ys__n1489 & ~new_new_n16841__;
  assign new_new_n20651__ = ~new_new_n20649__ & ~new_new_n20650__;
  assign new_new_n20652__ = ~new_new_n18427__ & ~new_new_n20651__;
  assign new_new_n20653__ = ~new_new_n20643__ & ~new_new_n20652__;
  assign new_new_n20654__ = ~ys__n19973 & ~new_new_n20653__;
  assign new_new_n20655__ = ys__n19973 & ys__n20002;
  assign new_new_n20656__ = ~new_new_n20654__ & ~new_new_n20655__;
  assign new_new_n20657__ = ~ys__n352 & ~new_new_n20656__;
  assign new_new_n20658__ = ~ys__n220 & ys__n47103;
  assign new_new_n20659__ = new_new_n18439__ & new_new_n20658__;
  assign new_new_n20660__ = new_new_n18441__ & new_new_n20658__;
  assign new_new_n20661__ = new_new_n18444__ & new_new_n19572__;
  assign new_new_n20662__ = ~new_new_n20660__ & ~new_new_n20661__;
  assign new_new_n20663__ = ~new_new_n20659__ & new_new_n20662__;
  assign new_new_n20664__ = new_new_n18453__ & ~new_new_n20663__;
  assign ys__n19965 = new_new_n20657__ | new_new_n20664__;
  assign new_new_n20666__ = ys__n19844 & ys__n19874;
  assign new_new_n20667__ = new_new_n18116__ & new_new_n20666__;
  assign new_new_n20668__ = ~ys__n23278 & ~new_new_n19589__;
  assign new_new_n20669__ = ~new_new_n19661__ & ~new_new_n20668__;
  assign new_new_n20670__ = ~ys__n1505 & ~new_new_n20669__;
  assign new_new_n20671__ = new_new_n19593__ & new_new_n19795__;
  assign new_new_n20672__ = ~new_new_n20670__ & ~new_new_n20671__;
  assign new_new_n20673__ = ~new_new_n18116__ & ~new_new_n20672__;
  assign new_new_n20674__ = ~new_new_n20667__ & ~new_new_n20673__;
  assign new_new_n20675__ = new_new_n18213__ & ~new_new_n20674__;
  assign new_new_n20676__ = ~ys__n1502 & ys__n27883;
  assign new_new_n20677__ = ~new_new_n18197__ & ~new_new_n18200__;
  assign new_new_n20678__ = ~ys__n23272 & ~new_new_n20677__;
  assign new_new_n20679__ = ys__n23272 & ~new_new_n20548__;
  assign new_new_n20680__ = ~new_new_n20678__ & ~new_new_n20679__;
  assign new_new_n20681__ = ~ys__n23274 & ~new_new_n20680__;
  assign new_new_n20682__ = ys__n23274 & ~new_new_n20415__;
  assign new_new_n20683__ = ~new_new_n20681__ & ~new_new_n20682__;
  assign new_new_n20684__ = ~ys__n23276 & ~new_new_n20683__;
  assign new_new_n20685__ = ys__n23276 & ~new_new_n20148__;
  assign new_new_n20686__ = ~new_new_n20684__ & ~new_new_n20685__;
  assign new_new_n20687__ = ~ys__n23278 & ~new_new_n20686__;
  assign new_new_n20688__ = ys__n23278 & ~new_new_n19610__;
  assign new_new_n20689__ = ~new_new_n20687__ & ~new_new_n20688__;
  assign new_new_n20690__ = ys__n1502 & ~new_new_n20689__;
  assign new_new_n20691__ = ~new_new_n20676__ & ~new_new_n20690__;
  assign new_new_n20692__ = ~new_new_n18213__ & ~new_new_n20691__;
  assign new_new_n20693__ = ~new_new_n20675__ & ~new_new_n20692__;
  assign new_new_n20694__ = new_new_n18224__ & ~new_new_n20693__;
  assign new_new_n20695__ = ~new_new_n10727__ & new_new_n18226__;
  assign new_new_n20696__ = ys__n1498 & new_new_n18322__;
  assign new_new_n20697__ = ~new_new_n20695__ & ~new_new_n20696__;
  assign new_new_n20698__ = ~ys__n1496 & ~new_new_n20697__;
  assign new_new_n20699__ = ys__n1496 & ~new_new_n18322__;
  assign new_new_n20700__ = ~new_new_n20698__ & ~new_new_n20699__;
  assign new_new_n20701__ = ~ys__n1495 & ~new_new_n20700__;
  assign new_new_n20702__ = ys__n1495 & new_new_n16856__;
  assign new_new_n20703__ = ~new_new_n20701__ & ~new_new_n20702__;
  assign new_new_n20704__ = ~new_new_n18224__ & ~new_new_n20703__;
  assign new_new_n20705__ = ~new_new_n20694__ & ~new_new_n20704__;
  assign new_new_n20706__ = new_new_n18581__ & ~new_new_n20705__;
  assign new_new_n20707__ = new_new_n18329__ & ~new_new_n20579__;
  assign new_new_n20708__ = new_new_n18391__ & ~new_new_n20707__;
  assign new_new_n20709__ = new_new_n18323__ & ~new_new_n20708__;
  assign new_new_n20710__ = ~new_new_n18323__ & new_new_n20708__;
  assign new_new_n20711__ = ~new_new_n20709__ & ~new_new_n20710__;
  assign new_new_n20712__ = ~ys__n1489 & ~new_new_n20711__;
  assign new_new_n20713__ = ys__n1489 & ~new_new_n16852__;
  assign new_new_n20714__ = ~new_new_n20712__ & ~new_new_n20713__;
  assign new_new_n20715__ = ~new_new_n18427__ & ~new_new_n20714__;
  assign new_new_n20716__ = ~new_new_n20706__ & ~new_new_n20715__;
  assign new_new_n20717__ = ~ys__n19973 & ~new_new_n20716__;
  assign new_new_n20718__ = ys__n19973 & ys__n20003;
  assign new_new_n20719__ = ~new_new_n20717__ & ~new_new_n20718__;
  assign new_new_n20720__ = ~ys__n352 & ~new_new_n20719__;
  assign new_new_n20721__ = ~ys__n220 & ys__n47104;
  assign new_new_n20722__ = new_new_n18439__ & new_new_n20721__;
  assign new_new_n20723__ = new_new_n18441__ & new_new_n20721__;
  assign new_new_n20724__ = new_new_n18444__ & new_new_n19645__;
  assign new_new_n20725__ = ~new_new_n20723__ & ~new_new_n20724__;
  assign new_new_n20726__ = ~new_new_n20722__ & new_new_n20725__;
  assign new_new_n20727__ = new_new_n18453__ & ~new_new_n20726__;
  assign ys__n19968 = new_new_n20720__ | new_new_n20727__;
  assign new_new_n20729__ = ys__n19844 & ys__n19875;
  assign new_new_n20730__ = new_new_n18116__ & new_new_n20729__;
  assign new_new_n20731__ = ~ys__n1505 & ys__n28030;
  assign new_new_n20732__ = new_new_n19664__ & new_new_n19795__;
  assign new_new_n20733__ = ~new_new_n20731__ & ~new_new_n20732__;
  assign new_new_n20734__ = ~new_new_n18116__ & ~new_new_n20733__;
  assign new_new_n20735__ = ~new_new_n20730__ & ~new_new_n20734__;
  assign new_new_n20736__ = new_new_n18213__ & ~new_new_n20735__;
  assign new_new_n20737__ = ~ys__n1502 & ys__n27885;
  assign new_new_n20738__ = ~new_new_n18537__ & ~new_new_n18549__;
  assign new_new_n20739__ = ~ys__n23272 & ~new_new_n20738__;
  assign new_new_n20740__ = ys__n23272 & ~new_new_n20614__;
  assign new_new_n20741__ = ~new_new_n20739__ & ~new_new_n20740__;
  assign new_new_n20742__ = ~ys__n23274 & ~new_new_n20741__;
  assign new_new_n20743__ = ys__n23274 & ~new_new_n20483__;
  assign new_new_n20744__ = ~new_new_n20742__ & ~new_new_n20743__;
  assign new_new_n20745__ = ~ys__n23276 & ~new_new_n20744__;
  assign new_new_n20746__ = ys__n23276 & ~new_new_n20216__;
  assign new_new_n20747__ = ~new_new_n20745__ & ~new_new_n20746__;
  assign new_new_n20748__ = ~ys__n23278 & ~new_new_n20747__;
  assign new_new_n20749__ = ys__n23278 & ~new_new_n19681__;
  assign new_new_n20750__ = ~new_new_n20748__ & ~new_new_n20749__;
  assign new_new_n20751__ = ys__n1502 & ~new_new_n20750__;
  assign new_new_n20752__ = ~new_new_n20737__ & ~new_new_n20751__;
  assign new_new_n20753__ = ~new_new_n18213__ & ~new_new_n20752__;
  assign new_new_n20754__ = ~new_new_n20736__ & ~new_new_n20753__;
  assign new_new_n20755__ = new_new_n18224__ & ~new_new_n20754__;
  assign new_new_n20756__ = ~new_new_n10730__ & new_new_n18226__;
  assign new_new_n20757__ = ys__n1498 & new_new_n18319__;
  assign new_new_n20758__ = ~new_new_n20756__ & ~new_new_n20757__;
  assign new_new_n20759__ = ~ys__n1496 & ~new_new_n20758__;
  assign new_new_n20760__ = ys__n1496 & ~new_new_n18319__;
  assign new_new_n20761__ = ~new_new_n20759__ & ~new_new_n20760__;
  assign new_new_n20762__ = ~ys__n1495 & ~new_new_n20761__;
  assign new_new_n20763__ = ys__n1495 & new_new_n18320__;
  assign new_new_n20764__ = ~new_new_n20762__ & ~new_new_n20763__;
  assign new_new_n20765__ = ~new_new_n18224__ & ~new_new_n20764__;
  assign new_new_n20766__ = ~new_new_n20755__ & ~new_new_n20765__;
  assign new_new_n20767__ = new_new_n18581__ & ~new_new_n20766__;
  assign new_new_n20768__ = ~new_new_n18323__ & ~new_new_n20708__;
  assign new_new_n20769__ = ~new_new_n10726__ & ~new_new_n20768__;
  assign new_new_n20770__ = new_new_n18321__ & ~new_new_n20769__;
  assign new_new_n20771__ = ~new_new_n18321__ & new_new_n20769__;
  assign new_new_n20772__ = ~new_new_n20770__ & ~new_new_n20771__;
  assign new_new_n20773__ = ~ys__n1489 & ~new_new_n20772__;
  assign new_new_n20774__ = ys__n1489 & ~new_new_n16861__;
  assign new_new_n20775__ = ~new_new_n20773__ & ~new_new_n20774__;
  assign new_new_n20776__ = ~new_new_n18427__ & ~new_new_n20775__;
  assign new_new_n20777__ = ~new_new_n20767__ & ~new_new_n20776__;
  assign new_new_n20778__ = ~ys__n19973 & ~new_new_n20777__;
  assign new_new_n20779__ = ys__n19973 & ys__n20004;
  assign new_new_n20780__ = ~new_new_n20778__ & ~new_new_n20779__;
  assign new_new_n20781__ = ~ys__n352 & ~new_new_n20780__;
  assign new_new_n20782__ = ~ys__n220 & ys__n47105;
  assign new_new_n20783__ = new_new_n18439__ & new_new_n20782__;
  assign new_new_n20784__ = new_new_n18441__ & new_new_n20782__;
  assign new_new_n20785__ = new_new_n18444__ & new_new_n19716__;
  assign new_new_n20786__ = ~new_new_n20784__ & ~new_new_n20785__;
  assign new_new_n20787__ = ~new_new_n20783__ & new_new_n20786__;
  assign new_new_n20788__ = new_new_n18453__ & ~new_new_n20787__;
  assign ys__n19971 = new_new_n20781__ | new_new_n20788__;
  assign new_new_n20790__ = ~new_new_n10767__ & ~new_new_n16732__;
  assign ys__n20006 = new_new_n16733__ | new_new_n20790__;
  assign new_new_n20792__ = ~new_new_n16612__ & ~new_new_n16732__;
  assign ys__n20007 = new_new_n16733__ | new_new_n20792__;
  assign new_new_n20794__ = ~new_new_n16732__ & ~new_new_n18690__;
  assign ys__n20008 = new_new_n16733__ | new_new_n20794__;
  assign new_new_n20796__ = ~new_new_n16732__ & ~new_new_n18797__;
  assign ys__n20009 = new_new_n16733__ | new_new_n20796__;
  assign new_new_n20798__ = ~new_new_n16732__ & ~new_new_n18877__;
  assign ys__n20010 = new_new_n16733__ | new_new_n20798__;
  assign new_new_n20800__ = ~new_new_n16732__ & ~new_new_n18962__;
  assign ys__n20011 = new_new_n16733__ | new_new_n20800__;
  assign new_new_n20802__ = ~new_new_n16732__ & ~new_new_n19047__;
  assign ys__n20012 = new_new_n16733__ | new_new_n20802__;
  assign new_new_n20804__ = ~new_new_n16732__ & ~new_new_n19130__;
  assign ys__n20013 = new_new_n16733__ | new_new_n20804__;
  assign new_new_n20806__ = ~new_new_n16732__ & ~new_new_n19198__;
  assign ys__n20014 = new_new_n16733__ | new_new_n20806__;
  assign new_new_n20808__ = ~new_new_n16732__ & ~new_new_n19271__;
  assign ys__n20015 = new_new_n16733__ | new_new_n20808__;
  assign new_new_n20810__ = ~new_new_n16732__ & ~new_new_n19344__;
  assign ys__n20016 = new_new_n16733__ | new_new_n20810__;
  assign new_new_n20812__ = ~new_new_n16732__ & ~new_new_n19417__;
  assign ys__n20017 = new_new_n16733__ | new_new_n20812__;
  assign new_new_n20814__ = ~new_new_n16732__ & ~new_new_n19490__;
  assign ys__n20018 = new_new_n16733__ | new_new_n20814__;
  assign new_new_n20816__ = ~new_new_n16732__ & ~new_new_n19563__;
  assign ys__n20019 = new_new_n16733__ | new_new_n20816__;
  assign new_new_n20818__ = ~new_new_n16732__ & ~new_new_n19636__;
  assign ys__n20020 = new_new_n16733__ | new_new_n20818__;
  assign new_new_n20820__ = ~new_new_n16732__ & ~new_new_n19707__;
  assign ys__n20021 = new_new_n16733__ | new_new_n20820__;
  assign new_new_n20822__ = ~new_new_n16732__ & ~new_new_n19773__;
  assign ys__n20022 = new_new_n16733__ | new_new_n20822__;
  assign new_new_n20824__ = ~new_new_n16732__ & ~new_new_n19842__;
  assign ys__n20023 = new_new_n16733__ | new_new_n20824__;
  assign new_new_n20826__ = ~new_new_n16732__ & ~new_new_n19910__;
  assign ys__n20024 = new_new_n16733__ | new_new_n20826__;
  assign new_new_n20828__ = ~new_new_n16732__ & ~new_new_n19978__;
  assign ys__n20025 = new_new_n16733__ | new_new_n20828__;
  assign new_new_n20830__ = ~new_new_n16732__ & ~new_new_n20046__;
  assign ys__n20026 = new_new_n16733__ | new_new_n20830__;
  assign new_new_n20832__ = ~new_new_n16732__ & ~new_new_n20114__;
  assign ys__n20027 = new_new_n16733__ | new_new_n20832__;
  assign new_new_n20834__ = ~new_new_n16732__ & ~new_new_n20182__;
  assign ys__n20028 = new_new_n16733__ | new_new_n20834__;
  assign new_new_n20836__ = ~new_new_n16732__ & ~new_new_n20250__;
  assign ys__n20029 = new_new_n16733__ | new_new_n20836__;
  assign new_new_n20838__ = ~new_new_n16732__ & ~new_new_n20316__;
  assign ys__n20030 = new_new_n16733__ | new_new_n20838__;
  assign new_new_n20840__ = ~new_new_n16732__ & ~new_new_n20384__;
  assign ys__n20031 = new_new_n16733__ | new_new_n20840__;
  assign new_new_n20842__ = ~new_new_n16732__ & ~new_new_n20452__;
  assign ys__n20032 = new_new_n16733__ | new_new_n20842__;
  assign new_new_n20844__ = ~new_new_n16732__ & ~new_new_n20520__;
  assign ys__n20033 = new_new_n16733__ | new_new_n20844__;
  assign new_new_n20846__ = ~new_new_n16732__ & ~new_new_n20586__;
  assign ys__n20034 = new_new_n16733__ | new_new_n20846__;
  assign new_new_n20848__ = ys__n1508 & new_new_n16616__;
  assign new_new_n20849__ = ~new_new_n16619__ & new_new_n20848__;
  assign ys__n20038 = new_new_n16632__ | new_new_n20849__;
  assign new_new_n20851__ = ys__n1508 & new_new_n16613__;
  assign new_new_n20852__ = ~new_new_n16619__ & new_new_n20851__;
  assign ys__n20043 = new_new_n16625__ | new_new_n20852__;
  assign new_new_n20854__ = ~new_new_n16613__ & ~new_new_n16616__;
  assign new_new_n20855__ = ~new_new_n16617__ & new_new_n20854__;
  assign new_new_n20856__ = ~new_new_n16614__ & new_new_n20855__;
  assign new_new_n20857__ = new_new_n16620__ & ~new_new_n20855__;
  assign new_new_n20858__ = ~new_new_n20856__ & new_new_n20857__;
  assign new_new_n20859__ = ~new_new_n16614__ & ~new_new_n16617__;
  assign new_new_n20860__ = new_new_n20854__ & new_new_n20859__;
  assign new_new_n20861__ = ys__n1509 & ~new_new_n20854__;
  assign new_new_n20862__ = ~new_new_n20860__ & new_new_n20861__;
  assign new_new_n20863__ = ~new_new_n20858__ & ~new_new_n20862__;
  assign ys__n20053 = ~ys__n1508 & ~new_new_n20863__;
  assign new_new_n20865__ = ~ys__n1511 & ys__n20035;
  assign new_new_n20866__ = ys__n20058 & new_new_n20865__;
  assign new_new_n20867__ = ys__n1511 & ys__n20058;
  assign new_new_n20868__ = ~new_new_n20866__ & ~new_new_n20867__;
  assign new_new_n20869__ = ~ys__n1509 & ~new_new_n20868__;
  assign new_new_n20870__ = ys__n1509 & ys__n20058;
  assign new_new_n20871__ = ~new_new_n20869__ & ~new_new_n20870__;
  assign new_new_n20872__ = ~ys__n1508 & ~new_new_n20871__;
  assign new_new_n20873__ = ys__n1508 & ys__n20058;
  assign ys__n20059 = new_new_n20872__ | new_new_n20873__;
  assign new_new_n20875__ = ys__n20061 & new_new_n20865__;
  assign new_new_n20876__ = ys__n1511 & ys__n20061;
  assign new_new_n20877__ = ~new_new_n20875__ & ~new_new_n20876__;
  assign new_new_n20878__ = ~ys__n1509 & ~new_new_n20877__;
  assign new_new_n20879__ = ys__n1509 & ys__n20061;
  assign new_new_n20880__ = ~new_new_n20878__ & ~new_new_n20879__;
  assign new_new_n20881__ = ~ys__n1508 & ~new_new_n20880__;
  assign new_new_n20882__ = ys__n1508 & ys__n20061;
  assign ys__n20062 = new_new_n20881__ | new_new_n20882__;
  assign new_new_n20884__ = ys__n20064 & new_new_n20865__;
  assign new_new_n20885__ = ys__n1511 & ys__n20064;
  assign new_new_n20886__ = ~new_new_n20884__ & ~new_new_n20885__;
  assign new_new_n20887__ = ~ys__n1509 & ~new_new_n20886__;
  assign new_new_n20888__ = ys__n1509 & ys__n20064;
  assign new_new_n20889__ = ~new_new_n20887__ & ~new_new_n20888__;
  assign new_new_n20890__ = ~ys__n1508 & ~new_new_n20889__;
  assign new_new_n20891__ = ys__n1508 & ys__n20064;
  assign ys__n20065 = new_new_n20890__ | new_new_n20891__;
  assign new_new_n20893__ = ys__n20067 & new_new_n20865__;
  assign new_new_n20894__ = ys__n1511 & ys__n20067;
  assign new_new_n20895__ = ~new_new_n20893__ & ~new_new_n20894__;
  assign new_new_n20896__ = ~ys__n1509 & ~new_new_n20895__;
  assign new_new_n20897__ = ys__n1509 & ys__n20067;
  assign new_new_n20898__ = ~new_new_n20896__ & ~new_new_n20897__;
  assign new_new_n20899__ = ~ys__n1508 & ~new_new_n20898__;
  assign new_new_n20900__ = ys__n1508 & ys__n20067;
  assign ys__n20068 = new_new_n20899__ | new_new_n20900__;
  assign new_new_n20902__ = ys__n20070 & new_new_n20865__;
  assign new_new_n20903__ = ys__n1511 & ys__n20070;
  assign new_new_n20904__ = ~new_new_n20902__ & ~new_new_n20903__;
  assign new_new_n20905__ = ~ys__n1509 & ~new_new_n20904__;
  assign new_new_n20906__ = ys__n1509 & ys__n20070;
  assign new_new_n20907__ = ~new_new_n20905__ & ~new_new_n20906__;
  assign new_new_n20908__ = ~ys__n1508 & ~new_new_n20907__;
  assign new_new_n20909__ = ys__n1508 & ys__n20070;
  assign ys__n20071 = new_new_n20908__ | new_new_n20909__;
  assign new_new_n20911__ = ys__n20073 & new_new_n20865__;
  assign new_new_n20912__ = ys__n1511 & ys__n20073;
  assign new_new_n20913__ = ~new_new_n20911__ & ~new_new_n20912__;
  assign new_new_n20914__ = ~ys__n1509 & ~new_new_n20913__;
  assign new_new_n20915__ = ys__n1509 & ys__n20073;
  assign new_new_n20916__ = ~new_new_n20914__ & ~new_new_n20915__;
  assign new_new_n20917__ = ~ys__n1508 & ~new_new_n20916__;
  assign new_new_n20918__ = ys__n1508 & ys__n20073;
  assign ys__n20074 = new_new_n20917__ | new_new_n20918__;
  assign new_new_n20920__ = ys__n20076 & new_new_n20865__;
  assign new_new_n20921__ = ys__n1511 & ys__n20076;
  assign new_new_n20922__ = ~new_new_n20920__ & ~new_new_n20921__;
  assign new_new_n20923__ = ~ys__n1509 & ~new_new_n20922__;
  assign new_new_n20924__ = ys__n1509 & ys__n20076;
  assign new_new_n20925__ = ~new_new_n20923__ & ~new_new_n20924__;
  assign new_new_n20926__ = ~ys__n1508 & ~new_new_n20925__;
  assign new_new_n20927__ = ys__n1508 & ys__n20076;
  assign ys__n20077 = new_new_n20926__ | new_new_n20927__;
  assign new_new_n20929__ = ys__n20079 & new_new_n20865__;
  assign new_new_n20930__ = ys__n1511 & ys__n20079;
  assign new_new_n20931__ = ~new_new_n20929__ & ~new_new_n20930__;
  assign new_new_n20932__ = ~ys__n1509 & ~new_new_n20931__;
  assign new_new_n20933__ = ys__n1509 & ys__n20079;
  assign new_new_n20934__ = ~new_new_n20932__ & ~new_new_n20933__;
  assign new_new_n20935__ = ~ys__n1508 & ~new_new_n20934__;
  assign new_new_n20936__ = ys__n1508 & ys__n20079;
  assign ys__n20080 = new_new_n20935__ | new_new_n20936__;
  assign new_new_n20938__ = ys__n20138 & new_new_n20865__;
  assign new_new_n20939__ = ys__n1511 & ys__n20138;
  assign new_new_n20940__ = ~new_new_n20938__ & ~new_new_n20939__;
  assign new_new_n20941__ = ~ys__n1509 & ~new_new_n20940__;
  assign new_new_n20942__ = ys__n1509 & ys__n20138;
  assign new_new_n20943__ = ~new_new_n20941__ & ~new_new_n20942__;
  assign new_new_n20944__ = ~ys__n1508 & ~new_new_n20943__;
  assign ys__n20082 = new_new_n20873__ | new_new_n20944__;
  assign new_new_n20946__ = ys__n20140 & new_new_n20865__;
  assign new_new_n20947__ = ys__n1511 & ys__n20140;
  assign new_new_n20948__ = ~new_new_n20946__ & ~new_new_n20947__;
  assign new_new_n20949__ = ~ys__n1509 & ~new_new_n20948__;
  assign new_new_n20950__ = ys__n1509 & ys__n20140;
  assign new_new_n20951__ = ~new_new_n20949__ & ~new_new_n20950__;
  assign new_new_n20952__ = ~ys__n1508 & ~new_new_n20951__;
  assign ys__n20084 = new_new_n20882__ | new_new_n20952__;
  assign new_new_n20954__ = ys__n20142 & new_new_n20865__;
  assign new_new_n20955__ = ys__n1511 & ys__n20142;
  assign new_new_n20956__ = ~new_new_n20954__ & ~new_new_n20955__;
  assign new_new_n20957__ = ~ys__n1509 & ~new_new_n20956__;
  assign new_new_n20958__ = ys__n1509 & ys__n20142;
  assign new_new_n20959__ = ~new_new_n20957__ & ~new_new_n20958__;
  assign new_new_n20960__ = ~ys__n1508 & ~new_new_n20959__;
  assign ys__n20086 = new_new_n20891__ | new_new_n20960__;
  assign new_new_n20962__ = ys__n20144 & new_new_n20865__;
  assign new_new_n20963__ = ys__n1511 & ys__n20144;
  assign new_new_n20964__ = ~new_new_n20962__ & ~new_new_n20963__;
  assign new_new_n20965__ = ~ys__n1509 & ~new_new_n20964__;
  assign new_new_n20966__ = ys__n1509 & ys__n20144;
  assign new_new_n20967__ = ~new_new_n20965__ & ~new_new_n20966__;
  assign new_new_n20968__ = ~ys__n1508 & ~new_new_n20967__;
  assign ys__n20088 = new_new_n20900__ | new_new_n20968__;
  assign new_new_n20970__ = ys__n20146 & new_new_n20865__;
  assign new_new_n20971__ = ys__n1511 & ys__n20146;
  assign new_new_n20972__ = ~new_new_n20970__ & ~new_new_n20971__;
  assign new_new_n20973__ = ~ys__n1509 & ~new_new_n20972__;
  assign new_new_n20974__ = ys__n1509 & ys__n20146;
  assign new_new_n20975__ = ~new_new_n20973__ & ~new_new_n20974__;
  assign new_new_n20976__ = ~ys__n1508 & ~new_new_n20975__;
  assign ys__n20090 = new_new_n20909__ | new_new_n20976__;
  assign new_new_n20978__ = ys__n20148 & new_new_n20865__;
  assign new_new_n20979__ = ys__n1511 & ys__n20148;
  assign new_new_n20980__ = ~new_new_n20978__ & ~new_new_n20979__;
  assign new_new_n20981__ = ~ys__n1509 & ~new_new_n20980__;
  assign new_new_n20982__ = ys__n1509 & ys__n20148;
  assign new_new_n20983__ = ~new_new_n20981__ & ~new_new_n20982__;
  assign new_new_n20984__ = ~ys__n1508 & ~new_new_n20983__;
  assign ys__n20092 = new_new_n20918__ | new_new_n20984__;
  assign new_new_n20986__ = ys__n20150 & new_new_n20865__;
  assign new_new_n20987__ = ys__n1511 & ys__n20150;
  assign new_new_n20988__ = ~new_new_n20986__ & ~new_new_n20987__;
  assign new_new_n20989__ = ~ys__n1509 & ~new_new_n20988__;
  assign new_new_n20990__ = ys__n1509 & ys__n20150;
  assign new_new_n20991__ = ~new_new_n20989__ & ~new_new_n20990__;
  assign new_new_n20992__ = ~ys__n1508 & ~new_new_n20991__;
  assign ys__n20094 = new_new_n20927__ | new_new_n20992__;
  assign new_new_n20994__ = ys__n20152 & new_new_n20865__;
  assign new_new_n20995__ = ys__n1511 & ys__n20152;
  assign new_new_n20996__ = ~new_new_n20994__ & ~new_new_n20995__;
  assign new_new_n20997__ = ~ys__n1509 & ~new_new_n20996__;
  assign new_new_n20998__ = ys__n1509 & ys__n20152;
  assign new_new_n20999__ = ~new_new_n20997__ & ~new_new_n20998__;
  assign new_new_n21000__ = ~ys__n1508 & ~new_new_n20999__;
  assign ys__n20096 = new_new_n20936__ | new_new_n21000__;
  assign new_new_n21002__ = ys__n20186 & new_new_n20865__;
  assign new_new_n21003__ = ys__n1511 & ys__n20186;
  assign new_new_n21004__ = ~new_new_n21002__ & ~new_new_n21003__;
  assign new_new_n21005__ = ~ys__n1509 & ~new_new_n21004__;
  assign new_new_n21006__ = ~new_new_n20870__ & ~new_new_n21005__;
  assign new_new_n21007__ = ~ys__n1508 & ~new_new_n21006__;
  assign ys__n20098 = new_new_n20873__ | new_new_n21007__;
  assign new_new_n21009__ = ys__n20188 & new_new_n20865__;
  assign new_new_n21010__ = ys__n1511 & ys__n20188;
  assign new_new_n21011__ = ~new_new_n21009__ & ~new_new_n21010__;
  assign new_new_n21012__ = ~ys__n1509 & ~new_new_n21011__;
  assign new_new_n21013__ = ~new_new_n20879__ & ~new_new_n21012__;
  assign new_new_n21014__ = ~ys__n1508 & ~new_new_n21013__;
  assign ys__n20100 = new_new_n20882__ | new_new_n21014__;
  assign new_new_n21016__ = ys__n20190 & new_new_n20865__;
  assign new_new_n21017__ = ys__n1511 & ys__n20190;
  assign new_new_n21018__ = ~new_new_n21016__ & ~new_new_n21017__;
  assign new_new_n21019__ = ~ys__n1509 & ~new_new_n21018__;
  assign new_new_n21020__ = ~new_new_n20888__ & ~new_new_n21019__;
  assign new_new_n21021__ = ~ys__n1508 & ~new_new_n21020__;
  assign ys__n20102 = new_new_n20891__ | new_new_n21021__;
  assign new_new_n21023__ = ys__n20192 & new_new_n20865__;
  assign new_new_n21024__ = ys__n1511 & ys__n20192;
  assign new_new_n21025__ = ~new_new_n21023__ & ~new_new_n21024__;
  assign new_new_n21026__ = ~ys__n1509 & ~new_new_n21025__;
  assign new_new_n21027__ = ~new_new_n20897__ & ~new_new_n21026__;
  assign new_new_n21028__ = ~ys__n1508 & ~new_new_n21027__;
  assign ys__n20104 = new_new_n20900__ | new_new_n21028__;
  assign new_new_n21030__ = ys__n20194 & new_new_n20865__;
  assign new_new_n21031__ = ys__n1511 & ys__n20194;
  assign new_new_n21032__ = ~new_new_n21030__ & ~new_new_n21031__;
  assign new_new_n21033__ = ~ys__n1509 & ~new_new_n21032__;
  assign new_new_n21034__ = ~new_new_n20906__ & ~new_new_n21033__;
  assign new_new_n21035__ = ~ys__n1508 & ~new_new_n21034__;
  assign ys__n20106 = new_new_n20909__ | new_new_n21035__;
  assign new_new_n21037__ = ys__n20196 & new_new_n20865__;
  assign new_new_n21038__ = ys__n1511 & ys__n20196;
  assign new_new_n21039__ = ~new_new_n21037__ & ~new_new_n21038__;
  assign new_new_n21040__ = ~ys__n1509 & ~new_new_n21039__;
  assign new_new_n21041__ = ~new_new_n20915__ & ~new_new_n21040__;
  assign new_new_n21042__ = ~ys__n1508 & ~new_new_n21041__;
  assign ys__n20108 = new_new_n20918__ | new_new_n21042__;
  assign new_new_n21044__ = ys__n20198 & new_new_n20865__;
  assign new_new_n21045__ = ys__n1511 & ys__n20198;
  assign new_new_n21046__ = ~new_new_n21044__ & ~new_new_n21045__;
  assign new_new_n21047__ = ~ys__n1509 & ~new_new_n21046__;
  assign new_new_n21048__ = ~new_new_n20924__ & ~new_new_n21047__;
  assign new_new_n21049__ = ~ys__n1508 & ~new_new_n21048__;
  assign ys__n20110 = new_new_n20927__ | new_new_n21049__;
  assign new_new_n21051__ = ys__n20200 & new_new_n20865__;
  assign new_new_n21052__ = ys__n1511 & ys__n20200;
  assign new_new_n21053__ = ~new_new_n21051__ & ~new_new_n21052__;
  assign new_new_n21054__ = ~ys__n1509 & ~new_new_n21053__;
  assign new_new_n21055__ = ~new_new_n20933__ & ~new_new_n21054__;
  assign new_new_n21056__ = ~ys__n1508 & ~new_new_n21055__;
  assign ys__n20112 = new_new_n20936__ | new_new_n21056__;
  assign new_new_n21058__ = ys__n20202 & new_new_n20865__;
  assign new_new_n21059__ = ys__n1511 & ys__n20202;
  assign new_new_n21060__ = ~new_new_n21058__ & ~new_new_n21059__;
  assign new_new_n21061__ = ~ys__n1509 & ~new_new_n21060__;
  assign new_new_n21062__ = ~new_new_n20942__ & ~new_new_n21061__;
  assign new_new_n21063__ = ~ys__n1508 & ~new_new_n21062__;
  assign ys__n20114 = new_new_n20873__ | new_new_n21063__;
  assign new_new_n21065__ = ys__n20204 & new_new_n20865__;
  assign new_new_n21066__ = ys__n1511 & ys__n20204;
  assign new_new_n21067__ = ~new_new_n21065__ & ~new_new_n21066__;
  assign new_new_n21068__ = ~ys__n1509 & ~new_new_n21067__;
  assign new_new_n21069__ = ~new_new_n20950__ & ~new_new_n21068__;
  assign new_new_n21070__ = ~ys__n1508 & ~new_new_n21069__;
  assign ys__n20116 = new_new_n20882__ | new_new_n21070__;
  assign new_new_n21072__ = ys__n20206 & new_new_n20865__;
  assign new_new_n21073__ = ys__n1511 & ys__n20206;
  assign new_new_n21074__ = ~new_new_n21072__ & ~new_new_n21073__;
  assign new_new_n21075__ = ~ys__n1509 & ~new_new_n21074__;
  assign new_new_n21076__ = ~new_new_n20958__ & ~new_new_n21075__;
  assign new_new_n21077__ = ~ys__n1508 & ~new_new_n21076__;
  assign ys__n20118 = new_new_n20891__ | new_new_n21077__;
  assign new_new_n21079__ = ys__n20208 & new_new_n20865__;
  assign new_new_n21080__ = ys__n1511 & ys__n20208;
  assign new_new_n21081__ = ~new_new_n21079__ & ~new_new_n21080__;
  assign new_new_n21082__ = ~ys__n1509 & ~new_new_n21081__;
  assign new_new_n21083__ = ~new_new_n20966__ & ~new_new_n21082__;
  assign new_new_n21084__ = ~ys__n1508 & ~new_new_n21083__;
  assign ys__n20120 = new_new_n20900__ | new_new_n21084__;
  assign new_new_n21086__ = ys__n20210 & new_new_n20865__;
  assign new_new_n21087__ = ys__n1511 & ys__n20210;
  assign new_new_n21088__ = ~new_new_n21086__ & ~new_new_n21087__;
  assign new_new_n21089__ = ~ys__n1509 & ~new_new_n21088__;
  assign new_new_n21090__ = ~new_new_n20974__ & ~new_new_n21089__;
  assign new_new_n21091__ = ~ys__n1508 & ~new_new_n21090__;
  assign ys__n20122 = new_new_n20909__ | new_new_n21091__;
  assign new_new_n21093__ = ys__n20212 & new_new_n20865__;
  assign new_new_n21094__ = ys__n1511 & ys__n20212;
  assign new_new_n21095__ = ~new_new_n21093__ & ~new_new_n21094__;
  assign new_new_n21096__ = ~ys__n1509 & ~new_new_n21095__;
  assign new_new_n21097__ = ~new_new_n20982__ & ~new_new_n21096__;
  assign new_new_n21098__ = ~ys__n1508 & ~new_new_n21097__;
  assign ys__n20124 = new_new_n20918__ | new_new_n21098__;
  assign new_new_n21100__ = ys__n20214 & new_new_n20865__;
  assign new_new_n21101__ = ys__n1511 & ys__n20214;
  assign new_new_n21102__ = ~new_new_n21100__ & ~new_new_n21101__;
  assign new_new_n21103__ = ~ys__n1509 & ~new_new_n21102__;
  assign new_new_n21104__ = ~new_new_n20990__ & ~new_new_n21103__;
  assign new_new_n21105__ = ~ys__n1508 & ~new_new_n21104__;
  assign ys__n20126 = new_new_n20927__ | new_new_n21105__;
  assign new_new_n21107__ = ys__n20216 & new_new_n20865__;
  assign new_new_n21108__ = ys__n1511 & ys__n20216;
  assign new_new_n21109__ = ~new_new_n21107__ & ~new_new_n21108__;
  assign new_new_n21110__ = ~ys__n1509 & ~new_new_n21109__;
  assign new_new_n21111__ = ~new_new_n20998__ & ~new_new_n21110__;
  assign new_new_n21112__ = ~ys__n1508 & ~new_new_n21111__;
  assign ys__n20128 = new_new_n20936__ | new_new_n21112__;
  assign new_new_n21114__ = ys__n23077 & ~new_new_n12308__;
  assign new_new_n21115__ = new_new_n12305__ & new_new_n21114__;
  assign new_new_n21116__ = ys__n23014 & new_new_n12308__;
  assign new_new_n21117__ = ~new_new_n21115__ & ~new_new_n21116__;
  assign new_new_n21118__ = ~new_new_n12306__ & ~new_new_n21117__;
  assign new_new_n21119__ = ys__n22918 & new_new_n12306__;
  assign ys__n22919 = new_new_n21118__ | new_new_n21119__;
  assign new_new_n21121__ = ys__n23078 & ~new_new_n12308__;
  assign new_new_n21122__ = new_new_n12305__ & new_new_n21121__;
  assign new_new_n21123__ = ys__n23016 & new_new_n12308__;
  assign new_new_n21124__ = ~new_new_n21122__ & ~new_new_n21123__;
  assign new_new_n21125__ = ~new_new_n12306__ & ~new_new_n21124__;
  assign new_new_n21126__ = ys__n22921 & new_new_n12306__;
  assign ys__n22922 = new_new_n21125__ | new_new_n21126__;
  assign new_new_n21128__ = ys__n23079 & ~new_new_n12308__;
  assign new_new_n21129__ = new_new_n12305__ & new_new_n21128__;
  assign new_new_n21130__ = ys__n23018 & new_new_n12308__;
  assign new_new_n21131__ = ~new_new_n21129__ & ~new_new_n21130__;
  assign new_new_n21132__ = ~new_new_n12306__ & ~new_new_n21131__;
  assign new_new_n21133__ = ys__n22924 & new_new_n12306__;
  assign ys__n22925 = new_new_n21132__ | new_new_n21133__;
  assign new_new_n21135__ = ys__n23080 & ~new_new_n12308__;
  assign new_new_n21136__ = new_new_n12305__ & new_new_n21135__;
  assign new_new_n21137__ = ys__n23020 & new_new_n12308__;
  assign new_new_n21138__ = ~new_new_n21136__ & ~new_new_n21137__;
  assign new_new_n21139__ = ~new_new_n12306__ & ~new_new_n21138__;
  assign new_new_n21140__ = ys__n22927 & new_new_n12306__;
  assign ys__n22928 = new_new_n21139__ | new_new_n21140__;
  assign new_new_n21142__ = ys__n23081 & ~new_new_n12308__;
  assign new_new_n21143__ = new_new_n12305__ & new_new_n21142__;
  assign new_new_n21144__ = ys__n23022 & new_new_n12308__;
  assign new_new_n21145__ = ~new_new_n21143__ & ~new_new_n21144__;
  assign new_new_n21146__ = ~new_new_n12306__ & ~new_new_n21145__;
  assign new_new_n21147__ = ys__n22930 & new_new_n12306__;
  assign ys__n22931 = new_new_n21146__ | new_new_n21147__;
  assign new_new_n21149__ = ys__n23082 & ~new_new_n12308__;
  assign new_new_n21150__ = new_new_n12305__ & new_new_n21149__;
  assign new_new_n21151__ = ys__n23024 & new_new_n12308__;
  assign new_new_n21152__ = ~new_new_n21150__ & ~new_new_n21151__;
  assign new_new_n21153__ = ~new_new_n12306__ & ~new_new_n21152__;
  assign new_new_n21154__ = ys__n22933 & new_new_n12306__;
  assign ys__n22934 = new_new_n21153__ | new_new_n21154__;
  assign new_new_n21156__ = ys__n23083 & ~new_new_n12308__;
  assign new_new_n21157__ = new_new_n12305__ & new_new_n21156__;
  assign new_new_n21158__ = ys__n23026 & new_new_n12308__;
  assign new_new_n21159__ = ~new_new_n21157__ & ~new_new_n21158__;
  assign new_new_n21160__ = ~new_new_n12306__ & ~new_new_n21159__;
  assign new_new_n21161__ = ys__n22936 & new_new_n12306__;
  assign ys__n22937 = new_new_n21160__ | new_new_n21161__;
  assign new_new_n21163__ = ys__n23084 & ~new_new_n12308__;
  assign new_new_n21164__ = new_new_n12305__ & new_new_n21163__;
  assign new_new_n21165__ = ys__n23028 & new_new_n12308__;
  assign new_new_n21166__ = ~new_new_n21164__ & ~new_new_n21165__;
  assign new_new_n21167__ = ~new_new_n12306__ & ~new_new_n21166__;
  assign new_new_n21168__ = ys__n22939 & new_new_n12306__;
  assign ys__n22940 = new_new_n21167__ | new_new_n21168__;
  assign new_new_n21170__ = ys__n23085 & ~new_new_n12308__;
  assign new_new_n21171__ = new_new_n12305__ & new_new_n21170__;
  assign new_new_n21172__ = ys__n23030 & new_new_n12308__;
  assign new_new_n21173__ = ~new_new_n21171__ & ~new_new_n21172__;
  assign new_new_n21174__ = ~new_new_n12306__ & ~new_new_n21173__;
  assign new_new_n21175__ = ys__n22942 & new_new_n12306__;
  assign ys__n22943 = new_new_n21174__ | new_new_n21175__;
  assign new_new_n21177__ = ys__n23086 & ~new_new_n12308__;
  assign new_new_n21178__ = new_new_n12305__ & new_new_n21177__;
  assign new_new_n21179__ = ys__n23032 & new_new_n12308__;
  assign new_new_n21180__ = ~new_new_n21178__ & ~new_new_n21179__;
  assign new_new_n21181__ = ~new_new_n12306__ & ~new_new_n21180__;
  assign new_new_n21182__ = ys__n22945 & new_new_n12306__;
  assign ys__n22946 = new_new_n21181__ | new_new_n21182__;
  assign new_new_n21184__ = ys__n23087 & ~new_new_n12308__;
  assign new_new_n21185__ = new_new_n12305__ & new_new_n21184__;
  assign new_new_n21186__ = ys__n23034 & new_new_n12308__;
  assign new_new_n21187__ = ~new_new_n21185__ & ~new_new_n21186__;
  assign new_new_n21188__ = ~new_new_n12306__ & ~new_new_n21187__;
  assign new_new_n21189__ = ys__n22948 & new_new_n12306__;
  assign ys__n22949 = new_new_n21188__ | new_new_n21189__;
  assign new_new_n21191__ = ys__n23088 & ~new_new_n12308__;
  assign new_new_n21192__ = new_new_n12305__ & new_new_n21191__;
  assign new_new_n21193__ = ys__n23036 & new_new_n12308__;
  assign new_new_n21194__ = ~new_new_n21192__ & ~new_new_n21193__;
  assign new_new_n21195__ = ~new_new_n12306__ & ~new_new_n21194__;
  assign new_new_n21196__ = ys__n22951 & new_new_n12306__;
  assign ys__n22952 = new_new_n21195__ | new_new_n21196__;
  assign new_new_n21198__ = ys__n23089 & ~new_new_n12308__;
  assign new_new_n21199__ = new_new_n12305__ & new_new_n21198__;
  assign new_new_n21200__ = ys__n23038 & new_new_n12308__;
  assign new_new_n21201__ = ~new_new_n21199__ & ~new_new_n21200__;
  assign new_new_n21202__ = ~new_new_n12306__ & ~new_new_n21201__;
  assign new_new_n21203__ = ys__n22954 & new_new_n12306__;
  assign ys__n22955 = new_new_n21202__ | new_new_n21203__;
  assign new_new_n21205__ = ys__n23090 & ~new_new_n12308__;
  assign new_new_n21206__ = new_new_n12305__ & new_new_n21205__;
  assign new_new_n21207__ = ys__n23040 & new_new_n12308__;
  assign new_new_n21208__ = ~new_new_n21206__ & ~new_new_n21207__;
  assign new_new_n21209__ = ~new_new_n12306__ & ~new_new_n21208__;
  assign new_new_n21210__ = ys__n22957 & new_new_n12306__;
  assign ys__n22958 = new_new_n21209__ | new_new_n21210__;
  assign new_new_n21212__ = ys__n23091 & ~new_new_n12308__;
  assign new_new_n21213__ = new_new_n12305__ & new_new_n21212__;
  assign new_new_n21214__ = ys__n23042 & new_new_n12308__;
  assign new_new_n21215__ = ~new_new_n21213__ & ~new_new_n21214__;
  assign new_new_n21216__ = ~new_new_n12306__ & ~new_new_n21215__;
  assign new_new_n21217__ = ys__n22960 & new_new_n12306__;
  assign ys__n22961 = new_new_n21216__ | new_new_n21217__;
  assign new_new_n21219__ = ys__n23092 & ~new_new_n12308__;
  assign new_new_n21220__ = new_new_n12305__ & new_new_n21219__;
  assign new_new_n21221__ = ys__n23044 & new_new_n12308__;
  assign new_new_n21222__ = ~new_new_n21220__ & ~new_new_n21221__;
  assign new_new_n21223__ = ~new_new_n12306__ & ~new_new_n21222__;
  assign new_new_n21224__ = ys__n22963 & new_new_n12306__;
  assign ys__n22964 = new_new_n21223__ | new_new_n21224__;
  assign new_new_n21226__ = ys__n23093 & ~new_new_n12308__;
  assign new_new_n21227__ = new_new_n12305__ & new_new_n21226__;
  assign new_new_n21228__ = ys__n23046 & new_new_n12308__;
  assign new_new_n21229__ = ~new_new_n21227__ & ~new_new_n21228__;
  assign new_new_n21230__ = ~new_new_n12306__ & ~new_new_n21229__;
  assign new_new_n21231__ = ys__n22966 & new_new_n12306__;
  assign ys__n22967 = new_new_n21230__ | new_new_n21231__;
  assign new_new_n21233__ = ys__n23094 & ~new_new_n12308__;
  assign new_new_n21234__ = new_new_n12305__ & new_new_n21233__;
  assign new_new_n21235__ = ys__n23048 & new_new_n12308__;
  assign new_new_n21236__ = ~new_new_n21234__ & ~new_new_n21235__;
  assign new_new_n21237__ = ~new_new_n12306__ & ~new_new_n21236__;
  assign new_new_n21238__ = ys__n22969 & new_new_n12306__;
  assign ys__n22970 = new_new_n21237__ | new_new_n21238__;
  assign new_new_n21240__ = ys__n23095 & ~new_new_n12308__;
  assign new_new_n21241__ = new_new_n12305__ & new_new_n21240__;
  assign new_new_n21242__ = ys__n23050 & new_new_n12308__;
  assign new_new_n21243__ = ~new_new_n21241__ & ~new_new_n21242__;
  assign new_new_n21244__ = ~new_new_n12306__ & ~new_new_n21243__;
  assign new_new_n21245__ = ys__n22972 & new_new_n12306__;
  assign ys__n22973 = new_new_n21244__ | new_new_n21245__;
  assign new_new_n21247__ = ys__n23096 & ~new_new_n12308__;
  assign new_new_n21248__ = new_new_n12305__ & new_new_n21247__;
  assign new_new_n21249__ = ys__n23052 & new_new_n12308__;
  assign new_new_n21250__ = ~new_new_n21248__ & ~new_new_n21249__;
  assign new_new_n21251__ = ~new_new_n12306__ & ~new_new_n21250__;
  assign new_new_n21252__ = ys__n22975 & new_new_n12306__;
  assign ys__n22976 = new_new_n21251__ | new_new_n21252__;
  assign new_new_n21254__ = ys__n23097 & ~new_new_n12308__;
  assign new_new_n21255__ = new_new_n12305__ & new_new_n21254__;
  assign new_new_n21256__ = ys__n23054 & new_new_n12308__;
  assign new_new_n21257__ = ~new_new_n21255__ & ~new_new_n21256__;
  assign new_new_n21258__ = ~new_new_n12306__ & ~new_new_n21257__;
  assign new_new_n21259__ = ys__n22978 & new_new_n12306__;
  assign ys__n22979 = new_new_n21258__ | new_new_n21259__;
  assign new_new_n21261__ = ys__n23098 & ~new_new_n12308__;
  assign new_new_n21262__ = new_new_n12305__ & new_new_n21261__;
  assign new_new_n21263__ = ys__n23056 & new_new_n12308__;
  assign new_new_n21264__ = ~new_new_n21262__ & ~new_new_n21263__;
  assign new_new_n21265__ = ~new_new_n12306__ & ~new_new_n21264__;
  assign new_new_n21266__ = ys__n22981 & new_new_n12306__;
  assign ys__n22982 = new_new_n21265__ | new_new_n21266__;
  assign new_new_n21268__ = ys__n23099 & ~new_new_n12308__;
  assign new_new_n21269__ = new_new_n12305__ & new_new_n21268__;
  assign new_new_n21270__ = ys__n23058 & new_new_n12308__;
  assign new_new_n21271__ = ~new_new_n21269__ & ~new_new_n21270__;
  assign new_new_n21272__ = ~new_new_n12306__ & ~new_new_n21271__;
  assign new_new_n21273__ = ys__n22984 & new_new_n12306__;
  assign ys__n22985 = new_new_n21272__ | new_new_n21273__;
  assign new_new_n21275__ = ys__n23100 & ~new_new_n12308__;
  assign new_new_n21276__ = new_new_n12305__ & new_new_n21275__;
  assign new_new_n21277__ = ys__n23060 & new_new_n12308__;
  assign new_new_n21278__ = ~new_new_n21276__ & ~new_new_n21277__;
  assign new_new_n21279__ = ~new_new_n12306__ & ~new_new_n21278__;
  assign new_new_n21280__ = ys__n22987 & new_new_n12306__;
  assign ys__n22988 = new_new_n21279__ | new_new_n21280__;
  assign new_new_n21282__ = ys__n23101 & ~new_new_n12308__;
  assign new_new_n21283__ = new_new_n12305__ & new_new_n21282__;
  assign new_new_n21284__ = ys__n23062 & new_new_n12308__;
  assign new_new_n21285__ = ~new_new_n21283__ & ~new_new_n21284__;
  assign new_new_n21286__ = ~new_new_n12306__ & ~new_new_n21285__;
  assign new_new_n21287__ = ys__n22990 & new_new_n12306__;
  assign ys__n22991 = new_new_n21286__ | new_new_n21287__;
  assign new_new_n21289__ = ys__n23102 & ~new_new_n12308__;
  assign new_new_n21290__ = new_new_n12305__ & new_new_n21289__;
  assign new_new_n21291__ = ys__n23064 & new_new_n12308__;
  assign new_new_n21292__ = ~new_new_n21290__ & ~new_new_n21291__;
  assign new_new_n21293__ = ~new_new_n12306__ & ~new_new_n21292__;
  assign new_new_n21294__ = ys__n22993 & new_new_n12306__;
  assign ys__n22994 = new_new_n21293__ | new_new_n21294__;
  assign new_new_n21296__ = ys__n23103 & ~new_new_n12308__;
  assign new_new_n21297__ = new_new_n12305__ & new_new_n21296__;
  assign new_new_n21298__ = ys__n23066 & new_new_n12308__;
  assign new_new_n21299__ = ~new_new_n21297__ & ~new_new_n21298__;
  assign new_new_n21300__ = ~new_new_n12306__ & ~new_new_n21299__;
  assign new_new_n21301__ = ys__n22996 & new_new_n12306__;
  assign ys__n22997 = new_new_n21300__ | new_new_n21301__;
  assign new_new_n21303__ = ys__n23104 & ~new_new_n12308__;
  assign new_new_n21304__ = new_new_n12305__ & new_new_n21303__;
  assign new_new_n21305__ = ys__n23068 & new_new_n12308__;
  assign new_new_n21306__ = ~new_new_n21304__ & ~new_new_n21305__;
  assign new_new_n21307__ = ~new_new_n12306__ & ~new_new_n21306__;
  assign new_new_n21308__ = ys__n22999 & new_new_n12306__;
  assign ys__n23000 = new_new_n21307__ | new_new_n21308__;
  assign new_new_n21310__ = ys__n23105 & ~new_new_n12308__;
  assign new_new_n21311__ = new_new_n12305__ & new_new_n21310__;
  assign new_new_n21312__ = ys__n23070 & new_new_n12308__;
  assign new_new_n21313__ = ~new_new_n21311__ & ~new_new_n21312__;
  assign new_new_n21314__ = ~new_new_n12306__ & ~new_new_n21313__;
  assign new_new_n21315__ = ys__n23002 & new_new_n12306__;
  assign ys__n23003 = new_new_n21314__ | new_new_n21315__;
  assign new_new_n21317__ = ys__n23106 & ~new_new_n12308__;
  assign new_new_n21318__ = new_new_n12305__ & new_new_n21317__;
  assign new_new_n21319__ = ys__n23072 & new_new_n12308__;
  assign new_new_n21320__ = ~new_new_n21318__ & ~new_new_n21319__;
  assign new_new_n21321__ = ~new_new_n12306__ & ~new_new_n21320__;
  assign new_new_n21322__ = ys__n23005 & new_new_n12306__;
  assign ys__n23006 = new_new_n21321__ | new_new_n21322__;
  assign new_new_n21324__ = ys__n23107 & ~new_new_n12308__;
  assign new_new_n21325__ = new_new_n12305__ & new_new_n21324__;
  assign new_new_n21326__ = ys__n23074 & new_new_n12308__;
  assign new_new_n21327__ = ~new_new_n21325__ & ~new_new_n21326__;
  assign new_new_n21328__ = ~new_new_n12306__ & ~new_new_n21327__;
  assign new_new_n21329__ = ys__n23008 & new_new_n12306__;
  assign ys__n23009 = new_new_n21328__ | new_new_n21329__;
  assign new_new_n21331__ = ys__n23108 & ~new_new_n12308__;
  assign new_new_n21332__ = new_new_n12305__ & new_new_n21331__;
  assign new_new_n21333__ = ys__n23076 & new_new_n12308__;
  assign new_new_n21334__ = ~new_new_n21332__ & ~new_new_n21333__;
  assign new_new_n21335__ = ~new_new_n12306__ & ~new_new_n21334__;
  assign new_new_n21336__ = ys__n23011 & new_new_n12306__;
  assign ys__n23012 = new_new_n21335__ | new_new_n21336__;
  assign new_new_n21338__ = ys__n18240 & ~ys__n18241;
  assign new_new_n21339__ = ys__n100 & ys__n18241;
  assign new_new_n21340__ = ~new_new_n21338__ & ~new_new_n21339__;
  assign new_new_n21341__ = ys__n874 & ~new_new_n21340__;
  assign new_new_n21342__ = ys__n18243 & ~ys__n18241;
  assign new_new_n21343__ = ys__n96 & ys__n18241;
  assign new_new_n21344__ = ~new_new_n21342__ & ~new_new_n21343__;
  assign new_new_n21345__ = ys__n874 & ~new_new_n21344__;
  assign new_new_n21346__ = new_new_n21341__ & ~new_new_n21345__;
  assign new_new_n21347__ = ys__n18223 & new_new_n21341__;
  assign new_new_n21348__ = new_new_n21345__ & new_new_n21347__;
  assign ys__n23263 = new_new_n21346__ | new_new_n21348__;
  assign new_new_n21350__ = ~ys__n18223 & ~new_new_n21345__;
  assign new_new_n21351__ = ys__n18223 & new_new_n21345__;
  assign ys__n23264 = new_new_n21350__ | new_new_n21351__;
  assign new_new_n21353__ = ~ys__n22464 & ys__n23339;
  assign new_new_n21354__ = ys__n22464 & ~ys__n23339;
  assign ys__n23483 = new_new_n21353__ | new_new_n21354__;
  assign new_new_n21356__ = new_new_n11276__ & new_new_n11277__;
  assign new_new_n21357__ = ~new_new_n11276__ & ~new_new_n11277__;
  assign ys__n23485 = new_new_n21356__ | new_new_n21357__;
  assign new_new_n21359__ = ~new_new_n11276__ & new_new_n11277__;
  assign new_new_n21360__ = ~new_new_n11272__ & ~new_new_n21359__;
  assign new_new_n21361__ = ~ys__n23550 & ~new_new_n21360__;
  assign new_new_n21362__ = ys__n23550 & new_new_n21360__;
  assign ys__n23487 = new_new_n21361__ | new_new_n21362__;
  assign new_new_n21364__ = ~ys__n23552 & ~new_new_n11280__;
  assign new_new_n21365__ = ys__n23552 & new_new_n11280__;
  assign ys__n23489 = new_new_n21364__ | new_new_n21365__;
  assign new_new_n21367__ = ys__n23552 & ~new_new_n11280__;
  assign new_new_n21368__ = ~ys__n23554 & new_new_n21367__;
  assign new_new_n21369__ = ys__n23554 & ~new_new_n21367__;
  assign ys__n23491 = new_new_n21368__ | new_new_n21369__;
  assign new_new_n21371__ = ~new_new_n11280__ & new_new_n11281__;
  assign new_new_n21372__ = ~ys__n23556 & new_new_n21371__;
  assign new_new_n21373__ = ys__n23556 & ~new_new_n21371__;
  assign ys__n23493 = new_new_n21372__ | new_new_n21373__;
  assign new_new_n21375__ = ys__n23556 & new_new_n21371__;
  assign new_new_n21376__ = ~ys__n23558 & new_new_n21375__;
  assign new_new_n21377__ = ys__n23558 & ~new_new_n21375__;
  assign ys__n23495 = new_new_n21376__ | new_new_n21377__;
  assign new_new_n21379__ = ~ys__n23560 & new_new_n11284__;
  assign new_new_n21380__ = ys__n23560 & ~new_new_n11284__;
  assign ys__n23497 = new_new_n21379__ | new_new_n21380__;
  assign new_new_n21382__ = ys__n23560 & new_new_n11284__;
  assign new_new_n21383__ = ~ys__n23562 & new_new_n21382__;
  assign new_new_n21384__ = ys__n23562 & ~new_new_n21382__;
  assign ys__n23499 = new_new_n21383__ | new_new_n21384__;
  assign new_new_n21386__ = new_new_n11284__ & new_new_n11285__;
  assign new_new_n21387__ = ~ys__n23564 & new_new_n21386__;
  assign new_new_n21388__ = ys__n23564 & ~new_new_n21386__;
  assign ys__n23501 = new_new_n21387__ | new_new_n21388__;
  assign new_new_n21390__ = ys__n23564 & new_new_n21386__;
  assign new_new_n21391__ = ~ys__n23566 & new_new_n21390__;
  assign new_new_n21392__ = ys__n23566 & ~new_new_n21390__;
  assign ys__n23503 = new_new_n21391__ | new_new_n21392__;
  assign new_new_n21394__ = new_new_n11284__ & new_new_n11287__;
  assign new_new_n21395__ = ~ys__n23568 & new_new_n21394__;
  assign new_new_n21396__ = ys__n23568 & ~new_new_n21394__;
  assign ys__n23505 = new_new_n21395__ | new_new_n21396__;
  assign new_new_n21398__ = ys__n23568 & new_new_n21394__;
  assign new_new_n21399__ = ~ys__n23570 & new_new_n21398__;
  assign new_new_n21400__ = ys__n23570 & ~new_new_n21398__;
  assign ys__n23507 = new_new_n21399__ | new_new_n21400__;
  assign new_new_n21402__ = new_new_n11288__ & new_new_n21394__;
  assign new_new_n21403__ = ~ys__n23572 & new_new_n21402__;
  assign new_new_n21404__ = ys__n23572 & ~new_new_n21402__;
  assign ys__n23509 = new_new_n21403__ | new_new_n21404__;
  assign new_new_n21406__ = ys__n23572 & new_new_n21402__;
  assign new_new_n21407__ = ~ys__n23574 & new_new_n21406__;
  assign new_new_n21408__ = ys__n23574 & ~new_new_n21406__;
  assign ys__n23511 = new_new_n21407__ | new_new_n21408__;
  assign new_new_n21410__ = ys__n420 & ~new_new_n11292__;
  assign new_new_n21411__ = ~ys__n420 & new_new_n11292__;
  assign ys__n23513 = new_new_n21410__ | new_new_n21411__;
  assign new_new_n21413__ = ys__n442 & ~new_new_n11292__;
  assign new_new_n21414__ = ys__n420 & ~ys__n442;
  assign new_new_n21415__ = ~ys__n420 & ys__n442;
  assign new_new_n21416__ = ~new_new_n21414__ & ~new_new_n21415__;
  assign new_new_n21417__ = new_new_n11292__ & ~new_new_n21416__;
  assign ys__n23515 = new_new_n21413__ | new_new_n21417__;
  assign new_new_n21419__ = ys__n440 & ~new_new_n11292__;
  assign new_new_n21420__ = ~ys__n440 & new_new_n11294__;
  assign new_new_n21421__ = ys__n440 & ~new_new_n11294__;
  assign new_new_n21422__ = ~new_new_n21420__ & ~new_new_n21421__;
  assign new_new_n21423__ = new_new_n11292__ & ~new_new_n21422__;
  assign ys__n23517 = new_new_n21419__ | new_new_n21423__;
  assign new_new_n21425__ = ys__n444 & ~new_new_n11292__;
  assign new_new_n21426__ = ys__n440 & new_new_n11294__;
  assign new_new_n21427__ = ~ys__n444 & new_new_n21426__;
  assign new_new_n21428__ = ys__n444 & ~new_new_n21426__;
  assign new_new_n21429__ = ~new_new_n21427__ & ~new_new_n21428__;
  assign new_new_n21430__ = new_new_n11292__ & ~new_new_n21429__;
  assign ys__n23519 = new_new_n21425__ | new_new_n21430__;
  assign new_new_n21432__ = ys__n438 & ~new_new_n11292__;
  assign new_new_n21433__ = ~ys__n438 & new_new_n11296__;
  assign new_new_n21434__ = ys__n438 & ~new_new_n11296__;
  assign new_new_n21435__ = ~new_new_n21433__ & ~new_new_n21434__;
  assign new_new_n21436__ = new_new_n11292__ & ~new_new_n21435__;
  assign ys__n23521 = new_new_n21432__ | new_new_n21436__;
  assign new_new_n21438__ = ys__n446 & ~new_new_n11292__;
  assign new_new_n21439__ = ys__n438 & new_new_n11296__;
  assign new_new_n21440__ = ~ys__n446 & new_new_n21439__;
  assign new_new_n21441__ = ys__n446 & ~new_new_n21439__;
  assign new_new_n21442__ = ~new_new_n21440__ & ~new_new_n21441__;
  assign new_new_n21443__ = new_new_n11292__ & ~new_new_n21442__;
  assign ys__n23523 = new_new_n21438__ | new_new_n21443__;
  assign new_new_n21445__ = ys__n434 & ~new_new_n11292__;
  assign new_new_n21446__ = new_new_n11296__ & new_new_n11297__;
  assign new_new_n21447__ = ~ys__n434 & new_new_n21446__;
  assign new_new_n21448__ = ys__n434 & ~new_new_n21446__;
  assign new_new_n21449__ = ~new_new_n21447__ & ~new_new_n21448__;
  assign new_new_n21450__ = new_new_n11292__ & ~new_new_n21449__;
  assign ys__n23525 = new_new_n21445__ | new_new_n21450__;
  assign new_new_n21452__ = ys__n436 & ~new_new_n11292__;
  assign new_new_n21453__ = ys__n434 & new_new_n21446__;
  assign new_new_n21454__ = ~ys__n436 & new_new_n21453__;
  assign new_new_n21455__ = ys__n436 & ~new_new_n21453__;
  assign new_new_n21456__ = ~new_new_n21454__ & ~new_new_n21455__;
  assign new_new_n21457__ = new_new_n11292__ & ~new_new_n21456__;
  assign ys__n23527 = new_new_n21452__ | new_new_n21457__;
  assign new_new_n21459__ = ys__n432 & ~new_new_n11292__;
  assign new_new_n21460__ = ~ys__n432 & new_new_n11300__;
  assign new_new_n21461__ = ys__n432 & ~new_new_n11300__;
  assign new_new_n21462__ = ~new_new_n21460__ & ~new_new_n21461__;
  assign new_new_n21463__ = new_new_n11292__ & ~new_new_n21462__;
  assign ys__n23529 = new_new_n21459__ | new_new_n21463__;
  assign new_new_n21465__ = ys__n448 & ~new_new_n11292__;
  assign new_new_n21466__ = ys__n432 & new_new_n11300__;
  assign new_new_n21467__ = ~ys__n448 & new_new_n21466__;
  assign new_new_n21468__ = ys__n448 & ~new_new_n21466__;
  assign new_new_n21469__ = ~new_new_n21467__ & ~new_new_n21468__;
  assign new_new_n21470__ = new_new_n11292__ & ~new_new_n21469__;
  assign ys__n23531 = new_new_n21465__ | new_new_n21470__;
  assign new_new_n21472__ = ys__n428 & ~new_new_n11292__;
  assign new_new_n21473__ = new_new_n11300__ & new_new_n11301__;
  assign new_new_n21474__ = ~ys__n428 & new_new_n21473__;
  assign new_new_n21475__ = ys__n428 & ~new_new_n21473__;
  assign new_new_n21476__ = ~new_new_n21474__ & ~new_new_n21475__;
  assign new_new_n21477__ = new_new_n11292__ & ~new_new_n21476__;
  assign ys__n23533 = new_new_n21472__ | new_new_n21477__;
  assign new_new_n21479__ = ys__n430 & ~new_new_n11292__;
  assign new_new_n21480__ = ys__n428 & new_new_n21473__;
  assign new_new_n21481__ = ~ys__n430 & new_new_n21480__;
  assign new_new_n21482__ = ys__n430 & ~new_new_n21480__;
  assign new_new_n21483__ = ~new_new_n21481__ & ~new_new_n21482__;
  assign new_new_n21484__ = new_new_n11292__ & ~new_new_n21483__;
  assign ys__n23535 = new_new_n21479__ | new_new_n21484__;
  assign new_new_n21486__ = ys__n426 & ~new_new_n11292__;
  assign new_new_n21487__ = ~ys__n426 & new_new_n11304__;
  assign new_new_n21488__ = ys__n426 & ~new_new_n11304__;
  assign new_new_n21489__ = ~new_new_n21487__ & ~new_new_n21488__;
  assign new_new_n21490__ = new_new_n11292__ & ~new_new_n21489__;
  assign ys__n23537 = new_new_n21486__ | new_new_n21490__;
  assign new_new_n21492__ = ~ys__n256 & ~ys__n18101;
  assign new_new_n21493__ = ~ys__n18105 & ~ys__n18106;
  assign new_new_n21494__ = new_new_n21492__ & new_new_n21493__;
  assign new_new_n21495__ = ~ys__n4566 & new_new_n21494__;
  assign new_new_n21496__ = ~new_new_n10820__ & ~new_new_n11628__;
  assign new_new_n21497__ = new_new_n10820__ & ~new_new_n11628__;
  assign new_new_n21498__ = ~new_new_n11628__ & ~new_new_n21496__;
  assign new_new_n21499__ = ~new_new_n21497__ & new_new_n21498__;
  assign new_new_n21500__ = new_new_n21496__ & ~new_new_n21499__;
  assign new_new_n21501__ = ys__n38398 & ~new_new_n21500__;
  assign new_new_n21502__ = ~ys__n18111 & ~ys__n18112;
  assign new_new_n21503__ = ys__n18109 & ~new_new_n21502__;
  assign new_new_n21504__ = ~ys__n262 & ~new_new_n21503__;
  assign new_new_n21505__ = ~new_new_n21501__ & ~new_new_n21504__;
  assign new_new_n21506__ = ~new_new_n21501__ & ~new_new_n21505__;
  assign new_new_n21507__ = new_new_n21495__ & ~new_new_n21506__;
  assign ys__n23635 = ~new_new_n21495__ | new_new_n21507__;
  assign new_new_n21509__ = new_new_n11180__ & new_new_n21504__;
  assign new_new_n21510__ = new_new_n21495__ & new_new_n21509__;
  assign new_new_n21511__ = new_new_n21497__ & new_new_n21510__;
  assign new_new_n21512__ = ~new_new_n21499__ & new_new_n21511__;
  assign new_new_n21513__ = ~new_new_n21501__ & new_new_n21512__;
  assign ys__n23636 = ~new_new_n21495__ | new_new_n21513__;
  assign new_new_n21515__ = ~ys__n23840 & ys__n38490;
  assign new_new_n21516__ = ys__n23840 & ~ys__n38490;
  assign new_new_n21517__ = ~new_new_n21515__ & ~new_new_n21516__;
  assign new_new_n21518__ = ~ys__n23842 & ys__n38491;
  assign new_new_n21519__ = ys__n23842 & ~ys__n38491;
  assign new_new_n21520__ = ~new_new_n21518__ & ~new_new_n21519__;
  assign new_new_n21521__ = new_new_n21517__ & new_new_n21520__;
  assign new_new_n21522__ = ~ys__n23834 & ys__n38487;
  assign new_new_n21523__ = ys__n23834 & ~ys__n38487;
  assign new_new_n21524__ = ~new_new_n21522__ & ~new_new_n21523__;
  assign new_new_n21525__ = ~ys__n23836 & ys__n38488;
  assign new_new_n21526__ = ys__n23836 & ~ys__n38488;
  assign new_new_n21527__ = ~new_new_n21525__ & ~new_new_n21526__;
  assign new_new_n21528__ = ~ys__n23838 & ys__n38489;
  assign new_new_n21529__ = ys__n23838 & ~ys__n38489;
  assign new_new_n21530__ = ~new_new_n21528__ & ~new_new_n21529__;
  assign new_new_n21531__ = new_new_n21527__ & new_new_n21530__;
  assign new_new_n21532__ = new_new_n21524__ & new_new_n21531__;
  assign new_new_n21533__ = new_new_n21521__ & new_new_n21532__;
  assign new_new_n21534__ = ys__n18114 & new_new_n21533__;
  assign new_new_n21535__ = ~ys__n296 & ~ys__n2251;
  assign new_new_n21536__ = ~ys__n2245 & new_new_n21535__;
  assign new_new_n21537__ = ~ys__n294 & ~ys__n2247;
  assign new_new_n21538__ = new_new_n21536__ & new_new_n21537__;
  assign new_new_n21539__ = ys__n23834 & new_new_n21538__;
  assign new_new_n21540__ = ~new_new_n21534__ & new_new_n21539__;
  assign new_new_n21541__ = ys__n294 & ~ys__n2247;
  assign new_new_n21542__ = new_new_n21536__ & new_new_n21541__;
  assign new_new_n21543__ = ys__n296 & ~ys__n2251;
  assign new_new_n21544__ = ~ys__n2245 & new_new_n21541__;
  assign new_new_n21545__ = new_new_n21543__ & new_new_n21544__;
  assign new_new_n21546__ = ~new_new_n21542__ & ~new_new_n21545__;
  assign new_new_n21547__ = ys__n23834 & ~new_new_n21546__;
  assign new_new_n21548__ = ys__n29220 & new_new_n21533__;
  assign new_new_n21549__ = ~ys__n2245 & new_new_n21543__;
  assign new_new_n21550__ = new_new_n21537__ & new_new_n21549__;
  assign new_new_n21551__ = ys__n23834 & new_new_n21550__;
  assign new_new_n21552__ = ~new_new_n21548__ & new_new_n21551__;
  assign new_new_n21553__ = ~new_new_n21547__ & ~new_new_n21552__;
  assign new_new_n21554__ = ~new_new_n21540__ & new_new_n21553__;
  assign new_new_n21555__ = ~new_new_n21538__ & ~new_new_n21550__;
  assign new_new_n21556__ = new_new_n21546__ & new_new_n21555__;
  assign new_new_n21557__ = ys__n648 & ~ys__n2239;
  assign new_new_n21558__ = ~ys__n650 & ~ys__n2233;
  assign new_new_n21559__ = new_new_n21557__ & new_new_n21558__;
  assign new_new_n21560__ = ys__n644 & ~ys__n646;
  assign new_new_n21561__ = new_new_n21559__ & new_new_n21560__;
  assign new_new_n21562__ = ~new_new_n21556__ & new_new_n21561__;
  assign new_new_n21563__ = ~new_new_n21554__ & new_new_n21562__;
  assign new_new_n21564__ = ys__n23822 & ~ys__n38491;
  assign new_new_n21565__ = ys__n23821 & ~ys__n38490;
  assign new_new_n21566__ = ~ys__n23822 & ys__n38491;
  assign new_new_n21567__ = ~new_new_n21565__ & ~new_new_n21566__;
  assign new_new_n21568__ = ~new_new_n21564__ & new_new_n21567__;
  assign new_new_n21569__ = ys__n23819 & ~ys__n38488;
  assign new_new_n21570__ = ~ys__n23820 & ys__n38489;
  assign new_new_n21571__ = ~new_new_n21569__ & ~new_new_n21570__;
  assign new_new_n21572__ = ys__n23820 & ~ys__n38489;
  assign new_new_n21573__ = ~ys__n23821 & ys__n38490;
  assign new_new_n21574__ = ~new_new_n21572__ & ~new_new_n21573__;
  assign new_new_n21575__ = new_new_n21571__ & new_new_n21574__;
  assign new_new_n21576__ = ~ys__n23818 & ys__n38487;
  assign new_new_n21577__ = ys__n18114 & ~new_new_n21576__;
  assign new_new_n21578__ = ys__n23818 & ~ys__n38487;
  assign new_new_n21579__ = ~ys__n23819 & ys__n38488;
  assign new_new_n21580__ = ~new_new_n21578__ & ~new_new_n21579__;
  assign new_new_n21581__ = new_new_n21577__ & new_new_n21580__;
  assign new_new_n21582__ = new_new_n21575__ & new_new_n21581__;
  assign new_new_n21583__ = new_new_n21568__ & new_new_n21582__;
  assign new_new_n21584__ = ys__n644 & ys__n646;
  assign new_new_n21585__ = ys__n650 & ~ys__n2233;
  assign new_new_n21586__ = new_new_n21557__ & new_new_n21585__;
  assign new_new_n21587__ = new_new_n21584__ & new_new_n21586__;
  assign new_new_n21588__ = ys__n23818 & new_new_n21587__;
  assign new_new_n21589__ = ~new_new_n21583__ & new_new_n21588__;
  assign new_new_n21590__ = new_new_n21559__ & new_new_n21584__;
  assign new_new_n21591__ = ys__n23818 & ~new_new_n21587__;
  assign new_new_n21592__ = new_new_n21590__ & new_new_n21591__;
  assign new_new_n21593__ = ~new_new_n21589__ & ~new_new_n21592__;
  assign new_new_n21594__ = ~new_new_n21561__ & ~new_new_n21593__;
  assign ys__n23795 = new_new_n21563__ | new_new_n21594__;
  assign new_new_n21596__ = ys__n23836 & new_new_n21538__;
  assign new_new_n21597__ = ~new_new_n21534__ & new_new_n21596__;
  assign new_new_n21598__ = ys__n23836 & ~new_new_n21546__;
  assign new_new_n21599__ = ys__n23836 & new_new_n21550__;
  assign new_new_n21600__ = ~new_new_n21548__ & new_new_n21599__;
  assign new_new_n21601__ = ~new_new_n21598__ & ~new_new_n21600__;
  assign new_new_n21602__ = ~new_new_n21597__ & new_new_n21601__;
  assign new_new_n21603__ = new_new_n21562__ & ~new_new_n21602__;
  assign new_new_n21604__ = ys__n23819 & new_new_n21587__;
  assign new_new_n21605__ = ~new_new_n21583__ & new_new_n21604__;
  assign new_new_n21606__ = ys__n23819 & ~new_new_n21587__;
  assign new_new_n21607__ = new_new_n21590__ & new_new_n21606__;
  assign new_new_n21608__ = ~new_new_n21605__ & ~new_new_n21607__;
  assign new_new_n21609__ = ~new_new_n21561__ & ~new_new_n21608__;
  assign ys__n23798 = new_new_n21603__ | new_new_n21609__;
  assign new_new_n21611__ = ys__n23838 & new_new_n21538__;
  assign new_new_n21612__ = ~new_new_n21534__ & new_new_n21611__;
  assign new_new_n21613__ = ys__n23838 & ~new_new_n21546__;
  assign new_new_n21614__ = ys__n23838 & new_new_n21550__;
  assign new_new_n21615__ = ~new_new_n21548__ & new_new_n21614__;
  assign new_new_n21616__ = ~new_new_n21613__ & ~new_new_n21615__;
  assign new_new_n21617__ = ~new_new_n21612__ & new_new_n21616__;
  assign new_new_n21618__ = new_new_n21562__ & ~new_new_n21617__;
  assign new_new_n21619__ = ys__n23820 & new_new_n21587__;
  assign new_new_n21620__ = ~new_new_n21583__ & new_new_n21619__;
  assign new_new_n21621__ = ys__n23820 & ~new_new_n21587__;
  assign new_new_n21622__ = new_new_n21590__ & new_new_n21621__;
  assign new_new_n21623__ = ~new_new_n21620__ & ~new_new_n21622__;
  assign new_new_n21624__ = ~new_new_n21561__ & ~new_new_n21623__;
  assign ys__n23801 = new_new_n21618__ | new_new_n21624__;
  assign new_new_n21626__ = ys__n23840 & new_new_n21538__;
  assign new_new_n21627__ = ~new_new_n21534__ & new_new_n21626__;
  assign new_new_n21628__ = ys__n23840 & ~new_new_n21546__;
  assign new_new_n21629__ = ys__n23840 & new_new_n21550__;
  assign new_new_n21630__ = ~new_new_n21548__ & new_new_n21629__;
  assign new_new_n21631__ = ~new_new_n21628__ & ~new_new_n21630__;
  assign new_new_n21632__ = ~new_new_n21627__ & new_new_n21631__;
  assign new_new_n21633__ = new_new_n21562__ & ~new_new_n21632__;
  assign new_new_n21634__ = ys__n23821 & new_new_n21587__;
  assign new_new_n21635__ = ~new_new_n21583__ & new_new_n21634__;
  assign new_new_n21636__ = ys__n23821 & ~new_new_n21587__;
  assign new_new_n21637__ = new_new_n21590__ & new_new_n21636__;
  assign new_new_n21638__ = ~new_new_n21635__ & ~new_new_n21637__;
  assign new_new_n21639__ = ~new_new_n21561__ & ~new_new_n21638__;
  assign ys__n23804 = new_new_n21633__ | new_new_n21639__;
  assign new_new_n21641__ = ys__n23842 & new_new_n21538__;
  assign new_new_n21642__ = ~new_new_n21534__ & new_new_n21641__;
  assign new_new_n21643__ = ys__n23842 & ~new_new_n21546__;
  assign new_new_n21644__ = ys__n23842 & new_new_n21550__;
  assign new_new_n21645__ = ~new_new_n21548__ & new_new_n21644__;
  assign new_new_n21646__ = ~new_new_n21643__ & ~new_new_n21645__;
  assign new_new_n21647__ = ~new_new_n21642__ & new_new_n21646__;
  assign new_new_n21648__ = new_new_n21562__ & ~new_new_n21647__;
  assign new_new_n21649__ = ys__n23822 & new_new_n21587__;
  assign new_new_n21650__ = ~new_new_n21583__ & new_new_n21649__;
  assign new_new_n21651__ = ys__n23822 & ~new_new_n21587__;
  assign new_new_n21652__ = new_new_n21590__ & new_new_n21651__;
  assign new_new_n21653__ = ~new_new_n21650__ & ~new_new_n21652__;
  assign new_new_n21654__ = ~new_new_n21561__ & ~new_new_n21653__;
  assign ys__n23807 = new_new_n21648__ | new_new_n21654__;
  assign new_new_n21656__ = ~ys__n740 & new_new_n12150__;
  assign new_new_n21657__ = ~new_new_n12430__ & ~new_new_n21656__;
  assign new_new_n21658__ = ~new_new_n12157__ & ~new_new_n21657__;
  assign new_new_n21659__ = ~new_new_n12157__ & ~new_new_n21658__;
  assign new_new_n21660__ = ~new_new_n12146__ & ~new_new_n21659__;
  assign ys__n23853 = new_new_n12146__ | new_new_n21660__;
  assign new_new_n21662__ = ~ys__n23910 & ys__n38498;
  assign new_new_n21663__ = ys__n23910 & ~ys__n38498;
  assign new_new_n21664__ = ~new_new_n21662__ & ~new_new_n21663__;
  assign new_new_n21665__ = ~ys__n23912 & ys__n38499;
  assign new_new_n21666__ = ys__n23912 & ~ys__n38499;
  assign new_new_n21667__ = ~new_new_n21665__ & ~new_new_n21666__;
  assign new_new_n21668__ = new_new_n21664__ & new_new_n21667__;
  assign new_new_n21669__ = ~ys__n23904 & ys__n38495;
  assign new_new_n21670__ = ys__n23904 & ~ys__n38495;
  assign new_new_n21671__ = ~new_new_n21669__ & ~new_new_n21670__;
  assign new_new_n21672__ = ~ys__n23906 & ys__n38496;
  assign new_new_n21673__ = ys__n23906 & ~ys__n38496;
  assign new_new_n21674__ = ~new_new_n21672__ & ~new_new_n21673__;
  assign new_new_n21675__ = ~ys__n23908 & ys__n38497;
  assign new_new_n21676__ = ys__n23908 & ~ys__n38497;
  assign new_new_n21677__ = ~new_new_n21675__ & ~new_new_n21676__;
  assign new_new_n21678__ = new_new_n21674__ & new_new_n21677__;
  assign new_new_n21679__ = new_new_n21671__ & new_new_n21678__;
  assign new_new_n21680__ = new_new_n21668__ & new_new_n21679__;
  assign new_new_n21681__ = ys__n18116 & new_new_n21680__;
  assign new_new_n21682__ = ~ys__n586 & ~ys__n2312;
  assign new_new_n21683__ = ~ys__n2306 & new_new_n21682__;
  assign new_new_n21684__ = ~ys__n588 & ~ys__n2308;
  assign new_new_n21685__ = new_new_n21683__ & new_new_n21684__;
  assign new_new_n21686__ = ys__n23904 & new_new_n21685__;
  assign new_new_n21687__ = ~new_new_n21681__ & new_new_n21686__;
  assign new_new_n21688__ = ys__n588 & ~ys__n2308;
  assign new_new_n21689__ = new_new_n21683__ & new_new_n21688__;
  assign new_new_n21690__ = ys__n586 & ~ys__n2312;
  assign new_new_n21691__ = ~ys__n2306 & new_new_n21688__;
  assign new_new_n21692__ = new_new_n21690__ & new_new_n21691__;
  assign new_new_n21693__ = ~new_new_n21689__ & ~new_new_n21692__;
  assign new_new_n21694__ = ys__n23904 & ~new_new_n21693__;
  assign new_new_n21695__ = ys__n29533 & new_new_n21680__;
  assign new_new_n21696__ = ~ys__n2306 & new_new_n21690__;
  assign new_new_n21697__ = new_new_n21684__ & new_new_n21696__;
  assign new_new_n21698__ = ys__n23904 & new_new_n21697__;
  assign new_new_n21699__ = ~new_new_n21695__ & new_new_n21698__;
  assign new_new_n21700__ = ~new_new_n21694__ & ~new_new_n21699__;
  assign new_new_n21701__ = ~new_new_n21687__ & new_new_n21700__;
  assign new_new_n21702__ = ~new_new_n21685__ & ~new_new_n21697__;
  assign new_new_n21703__ = new_new_n21693__ & new_new_n21702__;
  assign new_new_n21704__ = ys__n656 & ~ys__n2282;
  assign new_new_n21705__ = ~ys__n658 & ~ys__n2276;
  assign new_new_n21706__ = new_new_n21704__ & new_new_n21705__;
  assign new_new_n21707__ = ys__n652 & ~ys__n654;
  assign new_new_n21708__ = new_new_n21706__ & new_new_n21707__;
  assign new_new_n21709__ = ~new_new_n21703__ & new_new_n21708__;
  assign new_new_n21710__ = ~new_new_n21701__ & new_new_n21709__;
  assign new_new_n21711__ = ys__n23892 & ~ys__n38499;
  assign new_new_n21712__ = ys__n23891 & ~ys__n38498;
  assign new_new_n21713__ = ~ys__n23892 & ys__n38499;
  assign new_new_n21714__ = ~new_new_n21712__ & ~new_new_n21713__;
  assign new_new_n21715__ = ~new_new_n21711__ & new_new_n21714__;
  assign new_new_n21716__ = ys__n23889 & ~ys__n38496;
  assign new_new_n21717__ = ~ys__n23890 & ys__n38497;
  assign new_new_n21718__ = ~new_new_n21716__ & ~new_new_n21717__;
  assign new_new_n21719__ = ys__n23890 & ~ys__n38497;
  assign new_new_n21720__ = ~ys__n23891 & ys__n38498;
  assign new_new_n21721__ = ~new_new_n21719__ & ~new_new_n21720__;
  assign new_new_n21722__ = new_new_n21718__ & new_new_n21721__;
  assign new_new_n21723__ = ~ys__n23888 & ys__n38495;
  assign new_new_n21724__ = ys__n18116 & ~new_new_n21723__;
  assign new_new_n21725__ = ys__n23888 & ~ys__n38495;
  assign new_new_n21726__ = ~ys__n23889 & ys__n38496;
  assign new_new_n21727__ = ~new_new_n21725__ & ~new_new_n21726__;
  assign new_new_n21728__ = new_new_n21724__ & new_new_n21727__;
  assign new_new_n21729__ = new_new_n21722__ & new_new_n21728__;
  assign new_new_n21730__ = new_new_n21715__ & new_new_n21729__;
  assign new_new_n21731__ = ys__n652 & ys__n654;
  assign new_new_n21732__ = ys__n658 & ~ys__n2276;
  assign new_new_n21733__ = new_new_n21704__ & new_new_n21732__;
  assign new_new_n21734__ = new_new_n21731__ & new_new_n21733__;
  assign new_new_n21735__ = ys__n23888 & new_new_n21734__;
  assign new_new_n21736__ = ~new_new_n21730__ & new_new_n21735__;
  assign new_new_n21737__ = new_new_n21706__ & new_new_n21731__;
  assign new_new_n21738__ = ys__n23888 & ~new_new_n21734__;
  assign new_new_n21739__ = new_new_n21737__ & new_new_n21738__;
  assign new_new_n21740__ = ~new_new_n21736__ & ~new_new_n21739__;
  assign new_new_n21741__ = ~new_new_n21708__ & ~new_new_n21740__;
  assign ys__n23865 = new_new_n21710__ | new_new_n21741__;
  assign new_new_n21743__ = ys__n23906 & new_new_n21685__;
  assign new_new_n21744__ = ~new_new_n21681__ & new_new_n21743__;
  assign new_new_n21745__ = ys__n23906 & ~new_new_n21693__;
  assign new_new_n21746__ = ys__n23906 & new_new_n21697__;
  assign new_new_n21747__ = ~new_new_n21695__ & new_new_n21746__;
  assign new_new_n21748__ = ~new_new_n21745__ & ~new_new_n21747__;
  assign new_new_n21749__ = ~new_new_n21744__ & new_new_n21748__;
  assign new_new_n21750__ = new_new_n21709__ & ~new_new_n21749__;
  assign new_new_n21751__ = ys__n23889 & new_new_n21734__;
  assign new_new_n21752__ = ~new_new_n21730__ & new_new_n21751__;
  assign new_new_n21753__ = ys__n23889 & ~new_new_n21734__;
  assign new_new_n21754__ = new_new_n21737__ & new_new_n21753__;
  assign new_new_n21755__ = ~new_new_n21752__ & ~new_new_n21754__;
  assign new_new_n21756__ = ~new_new_n21708__ & ~new_new_n21755__;
  assign ys__n23868 = new_new_n21750__ | new_new_n21756__;
  assign new_new_n21758__ = ys__n23908 & new_new_n21685__;
  assign new_new_n21759__ = ~new_new_n21681__ & new_new_n21758__;
  assign new_new_n21760__ = ys__n23908 & ~new_new_n21693__;
  assign new_new_n21761__ = ys__n23908 & new_new_n21697__;
  assign new_new_n21762__ = ~new_new_n21695__ & new_new_n21761__;
  assign new_new_n21763__ = ~new_new_n21760__ & ~new_new_n21762__;
  assign new_new_n21764__ = ~new_new_n21759__ & new_new_n21763__;
  assign new_new_n21765__ = new_new_n21709__ & ~new_new_n21764__;
  assign new_new_n21766__ = ys__n23890 & new_new_n21734__;
  assign new_new_n21767__ = ~new_new_n21730__ & new_new_n21766__;
  assign new_new_n21768__ = ys__n23890 & ~new_new_n21734__;
  assign new_new_n21769__ = new_new_n21737__ & new_new_n21768__;
  assign new_new_n21770__ = ~new_new_n21767__ & ~new_new_n21769__;
  assign new_new_n21771__ = ~new_new_n21708__ & ~new_new_n21770__;
  assign ys__n23871 = new_new_n21765__ | new_new_n21771__;
  assign new_new_n21773__ = ys__n23910 & new_new_n21685__;
  assign new_new_n21774__ = ~new_new_n21681__ & new_new_n21773__;
  assign new_new_n21775__ = ys__n23910 & ~new_new_n21693__;
  assign new_new_n21776__ = ys__n23910 & new_new_n21697__;
  assign new_new_n21777__ = ~new_new_n21695__ & new_new_n21776__;
  assign new_new_n21778__ = ~new_new_n21775__ & ~new_new_n21777__;
  assign new_new_n21779__ = ~new_new_n21774__ & new_new_n21778__;
  assign new_new_n21780__ = new_new_n21709__ & ~new_new_n21779__;
  assign new_new_n21781__ = ys__n23891 & new_new_n21734__;
  assign new_new_n21782__ = ~new_new_n21730__ & new_new_n21781__;
  assign new_new_n21783__ = ys__n23891 & ~new_new_n21734__;
  assign new_new_n21784__ = new_new_n21737__ & new_new_n21783__;
  assign new_new_n21785__ = ~new_new_n21782__ & ~new_new_n21784__;
  assign new_new_n21786__ = ~new_new_n21708__ & ~new_new_n21785__;
  assign ys__n23874 = new_new_n21780__ | new_new_n21786__;
  assign new_new_n21788__ = ys__n23912 & new_new_n21685__;
  assign new_new_n21789__ = ~new_new_n21681__ & new_new_n21788__;
  assign new_new_n21790__ = ys__n23912 & ~new_new_n21693__;
  assign new_new_n21791__ = ys__n23912 & new_new_n21697__;
  assign new_new_n21792__ = ~new_new_n21695__ & new_new_n21791__;
  assign new_new_n21793__ = ~new_new_n21790__ & ~new_new_n21792__;
  assign new_new_n21794__ = ~new_new_n21789__ & new_new_n21793__;
  assign new_new_n21795__ = new_new_n21709__ & ~new_new_n21794__;
  assign new_new_n21796__ = ys__n23892 & new_new_n21734__;
  assign new_new_n21797__ = ~new_new_n21730__ & new_new_n21796__;
  assign new_new_n21798__ = ys__n23892 & ~new_new_n21734__;
  assign new_new_n21799__ = new_new_n21737__ & new_new_n21798__;
  assign new_new_n21800__ = ~new_new_n21797__ & ~new_new_n21799__;
  assign new_new_n21801__ = ~new_new_n21708__ & ~new_new_n21800__;
  assign ys__n23877 = new_new_n21795__ | new_new_n21801__;
  assign new_new_n21803__ = ~ys__n740 & new_new_n12161__;
  assign new_new_n21804__ = ~new_new_n12451__ & ~new_new_n21803__;
  assign new_new_n21805__ = ~new_new_n12168__ & ~new_new_n21804__;
  assign new_new_n21806__ = ~new_new_n12168__ & ~new_new_n21805__;
  assign new_new_n21807__ = ~new_new_n12146__ & ~new_new_n21806__;
  assign ys__n23921 = new_new_n12146__ | new_new_n21807__;
  assign new_new_n21809__ = ~ys__n23983 & ys__n38506;
  assign new_new_n21810__ = ys__n23983 & ~ys__n38506;
  assign new_new_n21811__ = ~new_new_n21809__ & ~new_new_n21810__;
  assign new_new_n21812__ = ~ys__n23985 & ys__n38507;
  assign new_new_n21813__ = ys__n23985 & ~ys__n38507;
  assign new_new_n21814__ = ~new_new_n21812__ & ~new_new_n21813__;
  assign new_new_n21815__ = new_new_n21811__ & new_new_n21814__;
  assign new_new_n21816__ = ~ys__n23977 & ys__n38503;
  assign new_new_n21817__ = ys__n23977 & ~ys__n38503;
  assign new_new_n21818__ = ~new_new_n21816__ & ~new_new_n21817__;
  assign new_new_n21819__ = ~ys__n23979 & ys__n38504;
  assign new_new_n21820__ = ys__n23979 & ~ys__n38504;
  assign new_new_n21821__ = ~new_new_n21819__ & ~new_new_n21820__;
  assign new_new_n21822__ = ~ys__n23981 & ys__n38505;
  assign new_new_n21823__ = ys__n23981 & ~ys__n38505;
  assign new_new_n21824__ = ~new_new_n21822__ & ~new_new_n21823__;
  assign new_new_n21825__ = new_new_n21821__ & new_new_n21824__;
  assign new_new_n21826__ = new_new_n21818__ & new_new_n21825__;
  assign new_new_n21827__ = new_new_n21815__ & new_new_n21826__;
  assign new_new_n21828__ = ys__n18118 & new_new_n21827__;
  assign new_new_n21829__ = ~ys__n194 & ~ys__n2433;
  assign new_new_n21830__ = ~ys__n2427 & new_new_n21829__;
  assign new_new_n21831__ = ~ys__n304 & ~ys__n2429;
  assign new_new_n21832__ = new_new_n21830__ & new_new_n21831__;
  assign new_new_n21833__ = ys__n23977 & new_new_n21832__;
  assign new_new_n21834__ = ~new_new_n21828__ & new_new_n21833__;
  assign new_new_n21835__ = ys__n304 & ~ys__n2429;
  assign new_new_n21836__ = new_new_n21830__ & new_new_n21835__;
  assign new_new_n21837__ = ys__n194 & ~ys__n2433;
  assign new_new_n21838__ = ~ys__n2427 & new_new_n21835__;
  assign new_new_n21839__ = new_new_n21837__ & new_new_n21838__;
  assign new_new_n21840__ = ~new_new_n21836__ & ~new_new_n21839__;
  assign new_new_n21841__ = ys__n23977 & ~new_new_n21840__;
  assign new_new_n21842__ = ys__n29808 & new_new_n21827__;
  assign new_new_n21843__ = ~ys__n2427 & new_new_n21837__;
  assign new_new_n21844__ = new_new_n21831__ & new_new_n21843__;
  assign new_new_n21845__ = ys__n23977 & new_new_n21844__;
  assign new_new_n21846__ = ~new_new_n21842__ & new_new_n21845__;
  assign new_new_n21847__ = ~new_new_n21841__ & ~new_new_n21846__;
  assign new_new_n21848__ = ~new_new_n21834__ & new_new_n21847__;
  assign new_new_n21849__ = ~new_new_n21832__ & ~new_new_n21844__;
  assign new_new_n21850__ = new_new_n21840__ & new_new_n21849__;
  assign new_new_n21851__ = ys__n662 & ys__n668;
  assign new_new_n21852__ = ~ys__n660 & ~ys__n666;
  assign new_new_n21853__ = new_new_n21851__ & new_new_n21852__;
  assign new_new_n21854__ = ys__n626 & ~ys__n664;
  assign new_new_n21855__ = new_new_n21853__ & new_new_n21854__;
  assign new_new_n21856__ = ~new_new_n21850__ & new_new_n21855__;
  assign new_new_n21857__ = ~new_new_n21848__ & new_new_n21856__;
  assign new_new_n21858__ = ys__n23960 & ~ys__n38507;
  assign new_new_n21859__ = ys__n23959 & ~ys__n38506;
  assign new_new_n21860__ = ~ys__n23960 & ys__n38507;
  assign new_new_n21861__ = ~new_new_n21859__ & ~new_new_n21860__;
  assign new_new_n21862__ = ~new_new_n21858__ & new_new_n21861__;
  assign new_new_n21863__ = ys__n23957 & ~ys__n38504;
  assign new_new_n21864__ = ~ys__n23958 & ys__n38505;
  assign new_new_n21865__ = ~new_new_n21863__ & ~new_new_n21864__;
  assign new_new_n21866__ = ys__n23958 & ~ys__n38505;
  assign new_new_n21867__ = ~ys__n23959 & ys__n38506;
  assign new_new_n21868__ = ~new_new_n21866__ & ~new_new_n21867__;
  assign new_new_n21869__ = new_new_n21865__ & new_new_n21868__;
  assign new_new_n21870__ = ~ys__n23956 & ys__n38503;
  assign new_new_n21871__ = ys__n18118 & ~new_new_n21870__;
  assign new_new_n21872__ = ys__n23956 & ~ys__n38503;
  assign new_new_n21873__ = ~ys__n23957 & ys__n38504;
  assign new_new_n21874__ = ~new_new_n21872__ & ~new_new_n21873__;
  assign new_new_n21875__ = new_new_n21871__ & new_new_n21874__;
  assign new_new_n21876__ = new_new_n21869__ & new_new_n21875__;
  assign new_new_n21877__ = new_new_n21862__ & new_new_n21876__;
  assign new_new_n21878__ = ys__n626 & ys__n664;
  assign new_new_n21879__ = ~ys__n660 & ys__n666;
  assign new_new_n21880__ = new_new_n21851__ & new_new_n21879__;
  assign new_new_n21881__ = new_new_n21878__ & new_new_n21880__;
  assign new_new_n21882__ = ys__n23956 & new_new_n21881__;
  assign new_new_n21883__ = ~new_new_n21877__ & new_new_n21882__;
  assign new_new_n21884__ = new_new_n21853__ & new_new_n21878__;
  assign new_new_n21885__ = ys__n23956 & ~new_new_n21881__;
  assign new_new_n21886__ = new_new_n21884__ & new_new_n21885__;
  assign new_new_n21887__ = ~new_new_n21883__ & ~new_new_n21886__;
  assign new_new_n21888__ = ~new_new_n21855__ & ~new_new_n21887__;
  assign ys__n23933 = new_new_n21857__ | new_new_n21888__;
  assign new_new_n21890__ = ys__n23979 & new_new_n21832__;
  assign new_new_n21891__ = ~new_new_n21828__ & new_new_n21890__;
  assign new_new_n21892__ = ys__n23979 & ~new_new_n21840__;
  assign new_new_n21893__ = ys__n23979 & new_new_n21844__;
  assign new_new_n21894__ = ~new_new_n21842__ & new_new_n21893__;
  assign new_new_n21895__ = ~new_new_n21892__ & ~new_new_n21894__;
  assign new_new_n21896__ = ~new_new_n21891__ & new_new_n21895__;
  assign new_new_n21897__ = new_new_n21856__ & ~new_new_n21896__;
  assign new_new_n21898__ = ys__n23957 & new_new_n21881__;
  assign new_new_n21899__ = ~new_new_n21877__ & new_new_n21898__;
  assign new_new_n21900__ = ys__n23957 & ~new_new_n21881__;
  assign new_new_n21901__ = new_new_n21884__ & new_new_n21900__;
  assign new_new_n21902__ = ~new_new_n21899__ & ~new_new_n21901__;
  assign new_new_n21903__ = ~new_new_n21855__ & ~new_new_n21902__;
  assign ys__n23936 = new_new_n21897__ | new_new_n21903__;
  assign new_new_n21905__ = ys__n23981 & new_new_n21832__;
  assign new_new_n21906__ = ~new_new_n21828__ & new_new_n21905__;
  assign new_new_n21907__ = ys__n23981 & ~new_new_n21840__;
  assign new_new_n21908__ = ys__n23981 & new_new_n21844__;
  assign new_new_n21909__ = ~new_new_n21842__ & new_new_n21908__;
  assign new_new_n21910__ = ~new_new_n21907__ & ~new_new_n21909__;
  assign new_new_n21911__ = ~new_new_n21906__ & new_new_n21910__;
  assign new_new_n21912__ = new_new_n21856__ & ~new_new_n21911__;
  assign new_new_n21913__ = ys__n23958 & new_new_n21881__;
  assign new_new_n21914__ = ~new_new_n21877__ & new_new_n21913__;
  assign new_new_n21915__ = ys__n23958 & ~new_new_n21881__;
  assign new_new_n21916__ = new_new_n21884__ & new_new_n21915__;
  assign new_new_n21917__ = ~new_new_n21914__ & ~new_new_n21916__;
  assign new_new_n21918__ = ~new_new_n21855__ & ~new_new_n21917__;
  assign ys__n23939 = new_new_n21912__ | new_new_n21918__;
  assign new_new_n21920__ = ys__n23983 & new_new_n21832__;
  assign new_new_n21921__ = ~new_new_n21828__ & new_new_n21920__;
  assign new_new_n21922__ = ys__n23983 & ~new_new_n21840__;
  assign new_new_n21923__ = ys__n23983 & new_new_n21844__;
  assign new_new_n21924__ = ~new_new_n21842__ & new_new_n21923__;
  assign new_new_n21925__ = ~new_new_n21922__ & ~new_new_n21924__;
  assign new_new_n21926__ = ~new_new_n21921__ & new_new_n21925__;
  assign new_new_n21927__ = new_new_n21856__ & ~new_new_n21926__;
  assign new_new_n21928__ = ys__n23959 & new_new_n21881__;
  assign new_new_n21929__ = ~new_new_n21877__ & new_new_n21928__;
  assign new_new_n21930__ = ys__n23959 & ~new_new_n21881__;
  assign new_new_n21931__ = new_new_n21884__ & new_new_n21930__;
  assign new_new_n21932__ = ~new_new_n21929__ & ~new_new_n21931__;
  assign new_new_n21933__ = ~new_new_n21855__ & ~new_new_n21932__;
  assign ys__n23942 = new_new_n21927__ | new_new_n21933__;
  assign new_new_n21935__ = ys__n23985 & new_new_n21832__;
  assign new_new_n21936__ = ~new_new_n21828__ & new_new_n21935__;
  assign new_new_n21937__ = ys__n23985 & ~new_new_n21840__;
  assign new_new_n21938__ = ys__n23985 & new_new_n21844__;
  assign new_new_n21939__ = ~new_new_n21842__ & new_new_n21938__;
  assign new_new_n21940__ = ~new_new_n21937__ & ~new_new_n21939__;
  assign new_new_n21941__ = ~new_new_n21936__ & new_new_n21940__;
  assign new_new_n21942__ = new_new_n21856__ & ~new_new_n21941__;
  assign new_new_n21943__ = ys__n23960 & new_new_n21881__;
  assign new_new_n21944__ = ~new_new_n21877__ & new_new_n21943__;
  assign new_new_n21945__ = ys__n23960 & ~new_new_n21881__;
  assign new_new_n21946__ = new_new_n21884__ & new_new_n21945__;
  assign new_new_n21947__ = ~new_new_n21944__ & ~new_new_n21946__;
  assign new_new_n21948__ = ~new_new_n21855__ & ~new_new_n21947__;
  assign ys__n23945 = new_new_n21942__ | new_new_n21948__;
  assign new_new_n21950__ = ~ys__n740 & new_new_n12194__;
  assign new_new_n21951__ = ~new_new_n12459__ & ~new_new_n21950__;
  assign new_new_n21952__ = ~new_new_n12201__ & ~new_new_n21951__;
  assign new_new_n21953__ = ~new_new_n12201__ & ~new_new_n21952__;
  assign new_new_n21954__ = ~new_new_n12146__ & ~new_new_n21953__;
  assign ys__n24099 = new_new_n12146__ | new_new_n21954__;
  assign ys__n24101 = ys__n24106 & ~ys__n24107;
  assign new_new_n21957__ = ~ys__n416 & ~ys__n38526;
  assign new_new_n21958__ = ys__n416 & ys__n38526;
  assign new_new_n21959__ = ~new_new_n21957__ & ~new_new_n21958__;
  assign new_new_n21960__ = ~ys__n24112 & ~new_new_n21959__;
  assign new_new_n21961__ = ~ys__n418 & ys__n24112;
  assign new_new_n21962__ = ~new_new_n21960__ & ~new_new_n21961__;
  assign new_new_n21963__ = ~ys__n1029 & ys__n1030;
  assign new_new_n21964__ = ~new_new_n21962__ & new_new_n21963__;
  assign new_new_n21965__ = ys__n1029 & ys__n24101;
  assign ys__n24102 = new_new_n21964__ | new_new_n21965__;
  assign ys__n24104 = ~ys__n24107 & ys__n24108;
  assign new_new_n21968__ = ys__n416 & ~ys__n686;
  assign new_new_n21969__ = ~ys__n416 & ys__n686;
  assign ys__n35705 = new_new_n21968__ | new_new_n21969__;
  assign new_new_n21971__ = ~ys__n38527 & ys__n35705;
  assign new_new_n21972__ = ys__n38527 & ~ys__n35705;
  assign new_new_n21973__ = ~new_new_n21971__ & ~new_new_n21972__;
  assign new_new_n21974__ = ~ys__n24112 & ~new_new_n21973__;
  assign new_new_n21975__ = ys__n418 & ~ys__n35704;
  assign new_new_n21976__ = ~ys__n418 & ys__n35704;
  assign new_new_n21977__ = ~new_new_n21975__ & ~new_new_n21976__;
  assign new_new_n21978__ = ys__n24112 & ~new_new_n21977__;
  assign new_new_n21979__ = ~new_new_n21974__ & ~new_new_n21978__;
  assign new_new_n21980__ = new_new_n21963__ & ~new_new_n21979__;
  assign new_new_n21981__ = ys__n1029 & ys__n24104;
  assign ys__n24105 = new_new_n21980__ | new_new_n21981__;
  assign new_new_n21983__ = ys__n47663 & new_new_n11634__;
  assign new_new_n21984__ = ys__n22826 & ~new_new_n11180__;
  assign new_new_n21985__ = new_new_n11175__ & new_new_n21984__;
  assign new_new_n21986__ = ~new_new_n16283__ & ~new_new_n21985__;
  assign new_new_n21987__ = ~new_new_n11186__ & ~new_new_n21986__;
  assign new_new_n21988__ = ys__n23548 & new_new_n11186__;
  assign new_new_n21989__ = ~new_new_n21987__ & ~new_new_n21988__;
  assign new_new_n21990__ = ~new_new_n11270__ & ~new_new_n21989__;
  assign new_new_n21991__ = new_new_n11270__ & ys__n23485;
  assign new_new_n21992__ = ~new_new_n21990__ & ~new_new_n21991__;
  assign new_new_n21993__ = new_new_n11324__ & ~new_new_n21992__;
  assign new_new_n21994__ = ys__n528 & ~new_new_n11324__;
  assign new_new_n21995__ = ~new_new_n21993__ & ~new_new_n21994__;
  assign new_new_n21996__ = ~new_new_n11343__ & ~new_new_n21995__;
  assign new_new_n21997__ = new_new_n11372__ & new_new_n11390__;
  assign new_new_n21998__ = ~new_new_n11372__ & ~new_new_n11390__;
  assign new_new_n21999__ = ~new_new_n21997__ & ~new_new_n21998__;
  assign new_new_n22000__ = new_new_n11343__ & ~new_new_n21999__;
  assign new_new_n22001__ = ~new_new_n21996__ & ~new_new_n22000__;
  assign new_new_n22002__ = new_new_n11629__ & ~new_new_n22001__;
  assign new_new_n22003__ = ~new_new_n21983__ & ~new_new_n22002__;
  assign new_new_n22004__ = new_new_n11640__ & ~new_new_n22003__;
  assign new_new_n22005__ = ys__n47663 & new_new_n11644__;
  assign new_new_n22006__ = new_new_n11642__ & ~new_new_n22001__;
  assign new_new_n22007__ = ~new_new_n22005__ & ~new_new_n22006__;
  assign new_new_n22008__ = new_new_n11650__ & ~new_new_n22007__;
  assign ys__n24116 = new_new_n22004__ | new_new_n22008__;
  assign new_new_n22010__ = ~ys__n18121 & ys__n24106;
  assign new_new_n22011__ = ys__n418 & ys__n18121;
  assign new_new_n22012__ = ~new_new_n22010__ & ~new_new_n22011__;
  assign new_new_n22013__ = new_new_n11041__ & new_new_n15897__;
  assign new_new_n22014__ = new_new_n12227__ & new_new_n22013__;
  assign new_new_n22015__ = ys__n1029 & new_new_n22014__;
  assign new_new_n22016__ = ~new_new_n22012__ & ~new_new_n22015__;
  assign new_new_n22017__ = ys__n24116 & new_new_n22015__;
  assign ys__n24118 = new_new_n22016__ | new_new_n22017__;
  assign new_new_n22019__ = ys__n1036 & ~ys__n1048;
  assign new_new_n22020__ = ~ys__n24123 & ys__n24124;
  assign new_new_n22021__ = new_new_n22019__ & new_new_n22020__;
  assign new_new_n22022__ = ys__n1048 & ~ys__n18007;
  assign new_new_n22023__ = ~new_new_n22021__ & ~new_new_n22022__;
  assign new_new_n22024__ = ~ys__n140 & ~new_new_n22023__;
  assign ys__n24120 = ys__n140 | new_new_n22024__;
  assign new_new_n22026__ = ~ys__n1036 & ~ys__n24123;
  assign new_new_n22027__ = ys__n24124 & new_new_n22026__;
  assign ys__n24126 = ys__n24123 | new_new_n22027__;
  assign new_new_n22029__ = ys__n1029 & ~ys__n1036;
  assign new_new_n22030__ = ys__n24131 & new_new_n22029__;
  assign new_new_n22031__ = ys__n1036 & ~ys__n24123;
  assign ys__n24130 = new_new_n22030__ | new_new_n22031__;
  assign new_new_n22033__ = ~ys__n18121 & ys__n18122;
  assign new_new_n22034__ = ~ys__n18124 & new_new_n22033__;
  assign new_new_n22035__ = new_new_n12439__ & new_new_n22034__;
  assign new_new_n22036__ = ys__n678 & ys__n680;
  assign new_new_n22037__ = ys__n682 & ys__n684;
  assign new_new_n22038__ = new_new_n22036__ & new_new_n22037__;
  assign new_new_n22039__ = ys__n670 & ys__n672;
  assign new_new_n22040__ = ys__n674 & ys__n676;
  assign new_new_n22041__ = new_new_n22039__ & new_new_n22040__;
  assign new_new_n22042__ = new_new_n22038__ & new_new_n22041__;
  assign new_new_n22043__ = ~ys__n38524 & ~new_new_n22042__;
  assign new_new_n22044__ = ~ys__n33423 & new_new_n10600__;
  assign new_new_n22045__ = new_new_n22014__ & new_new_n22044__;
  assign new_new_n22046__ = ~new_new_n22043__ & new_new_n22045__;
  assign new_new_n22047__ = ~ys__n18120 & new_new_n22046__;
  assign new_new_n22048__ = ~new_new_n10597__ & new_new_n22047__;
  assign ys__n24134 = new_new_n22035__ | new_new_n22048__;
  assign new_new_n22050__ = ~ys__n18122 & ys__n24143;
  assign new_new_n22051__ = ~ys__n24158 & new_new_n22050__;
  assign new_new_n22052__ = ~new_new_n10855__ & ~new_new_n22051__;
  assign new_new_n22053__ = ~ys__n18121 & ~new_new_n22052__;
  assign new_new_n22054__ = ys__n416 & ys__n686;
  assign new_new_n22055__ = ys__n18124 & new_new_n22054__;
  assign new_new_n22056__ = ys__n18121 & new_new_n22055__;
  assign ys__n24140 = new_new_n22053__ | new_new_n22056__;
  assign new_new_n22058__ = ~ys__n1029 & ys__n1038;
  assign new_new_n22059__ = ~ys__n18120 & new_new_n22015__;
  assign new_new_n22060__ = ~new_new_n10597__ & new_new_n22059__;
  assign new_new_n22061__ = ~ys__n33423 & new_new_n22060__;
  assign new_new_n22062__ = ~ys__n18120 & ~new_new_n22061__;
  assign new_new_n22063__ = ~ys__n18120 & new_new_n22014__;
  assign new_new_n22064__ = ~new_new_n10597__ & new_new_n22063__;
  assign new_new_n22065__ = ~new_new_n22062__ & new_new_n22064__;
  assign new_new_n22066__ = ~ys__n24158 & new_new_n10600__;
  assign new_new_n22067__ = ~new_new_n22065__ & new_new_n22066__;
  assign new_new_n22068__ = ~new_new_n22058__ & ~new_new_n22067__;
  assign new_new_n22069__ = ~ys__n1036 & ~new_new_n22068__;
  assign new_new_n22070__ = ys__n1036 & ys__n24123;
  assign ys__n24145 = new_new_n22069__ | new_new_n22070__;
  assign new_new_n22072__ = ys__n18121 & new_new_n12439__;
  assign new_new_n22073__ = ~new_new_n22055__ & new_new_n22072__;
  assign new_new_n22074__ = new_new_n22043__ & new_new_n22045__;
  assign new_new_n22075__ = ~ys__n18120 & new_new_n22074__;
  assign new_new_n22076__ = ~new_new_n10597__ & new_new_n22075__;
  assign new_new_n22077__ = new_new_n22060__ & new_new_n22076__;
  assign ys__n24149 = new_new_n22073__ | new_new_n22077__;
  assign ys__n38521 = ys__n24143 & ys__n24158;
  assign new_new_n22080__ = new_new_n12434__ & new_new_n12439__;
  assign new_new_n22081__ = ys__n38521 & new_new_n22080__;
  assign new_new_n22082__ = ys__n24158 & new_new_n10600__;
  assign new_new_n22083__ = ~new_new_n22060__ & new_new_n22082__;
  assign ys__n24154 = new_new_n22081__ | new_new_n22083__;
  assign new_new_n22085__ = ~ys__n30974 & ~ys__n33272;
  assign new_new_n22086__ = ~ys__n33274 & ~ys__n33276;
  assign new_new_n22087__ = new_new_n22085__ & new_new_n22086__;
  assign new_new_n22088__ = ~ys__n33278 & ~new_new_n22087__;
  assign new_new_n22089__ = ~ys__n33274 & new_new_n22085__;
  assign new_new_n22090__ = ~ys__n33276 & ~new_new_n22089__;
  assign new_new_n22091__ = ys__n33278 & new_new_n22087__;
  assign new_new_n22092__ = ~new_new_n22090__ & ~new_new_n22091__;
  assign new_new_n22093__ = ~new_new_n22088__ & new_new_n22092__;
  assign new_new_n22094__ = ys__n30974 & ~ys__n33272;
  assign new_new_n22095__ = ~ys__n30974 & ys__n33272;
  assign new_new_n22096__ = ~ys__n30974 & ~new_new_n22095__;
  assign new_new_n22097__ = ~new_new_n22094__ & new_new_n22096__;
  assign new_new_n22098__ = ys__n33274 & new_new_n22085__;
  assign new_new_n22099__ = ~ys__n33274 & ~new_new_n22085__;
  assign new_new_n22100__ = ~new_new_n22098__ & ~new_new_n22099__;
  assign new_new_n22101__ = new_new_n22097__ & new_new_n22100__;
  assign new_new_n22102__ = ~ys__n33278 & new_new_n22087__;
  assign new_new_n22103__ = ys__n33276 & new_new_n22089__;
  assign new_new_n22104__ = new_new_n22102__ & ~new_new_n22103__;
  assign new_new_n22105__ = new_new_n22101__ & new_new_n22104__;
  assign new_new_n22106__ = new_new_n22093__ & new_new_n22105__;
  assign new_new_n22107__ = ~ys__n38561 & ~new_new_n22106__;
  assign ys__n24160 = ~ys__n1084 & ~new_new_n22107__;
  assign ys__n24162 = ~ys__n24107 & ys__n24167;
  assign new_new_n22110__ = ~ys__n318 & ~ys__n38564;
  assign new_new_n22111__ = ys__n318 & ys__n38564;
  assign new_new_n22112__ = ~new_new_n22110__ & ~new_new_n22111__;
  assign new_new_n22113__ = ~ys__n24112 & ~new_new_n22112__;
  assign new_new_n22114__ = ~ys__n306 & ys__n24112;
  assign new_new_n22115__ = ~new_new_n22113__ & ~new_new_n22114__;
  assign new_new_n22116__ = ~ys__n1072 & ys__n1073;
  assign new_new_n22117__ = ~new_new_n22115__ & new_new_n22116__;
  assign new_new_n22118__ = ys__n1072 & ys__n24162;
  assign ys__n24163 = new_new_n22117__ | new_new_n22118__;
  assign ys__n24165 = ~ys__n24107 & ys__n24168;
  assign new_new_n22121__ = ys__n318 & ~ys__n624;
  assign new_new_n22122__ = ~ys__n318 & ys__n624;
  assign ys__n38566 = new_new_n22121__ | new_new_n22122__;
  assign new_new_n22124__ = ~ys__n38565 & ys__n38566;
  assign new_new_n22125__ = ys__n38565 & ~ys__n38566;
  assign new_new_n22126__ = ~new_new_n22124__ & ~new_new_n22125__;
  assign new_new_n22127__ = ~ys__n24112 & ~new_new_n22126__;
  assign new_new_n22128__ = ys__n306 & ~ys__n38568;
  assign new_new_n22129__ = ~ys__n306 & ys__n38568;
  assign new_new_n22130__ = ~new_new_n22128__ & ~new_new_n22129__;
  assign new_new_n22131__ = ys__n24112 & ~new_new_n22130__;
  assign new_new_n22132__ = ~new_new_n22127__ & ~new_new_n22131__;
  assign new_new_n22133__ = new_new_n22116__ & ~new_new_n22132__;
  assign new_new_n22134__ = ys__n1072 & ys__n24165;
  assign ys__n24166 = new_new_n22133__ | new_new_n22134__;
  assign new_new_n22136__ = ys__n24167 & ~ys__n24177;
  assign new_new_n22137__ = ys__n306 & ys__n24177;
  assign new_new_n22138__ = ~new_new_n22136__ & ~new_new_n22137__;
  assign new_new_n22139__ = ys__n1072 & new_new_n16924__;
  assign new_new_n22140__ = ~new_new_n22138__ & ~new_new_n22139__;
  assign new_new_n22141__ = ys__n24116 & new_new_n22139__;
  assign ys__n24176 = new_new_n22140__ | new_new_n22141__;
  assign new_new_n22143__ = ys__n47665 & new_new_n11634__;
  assign new_new_n22144__ = ys__n22830 & ~new_new_n11180__;
  assign new_new_n22145__ = new_new_n11175__ & new_new_n22144__;
  assign new_new_n22146__ = ~new_new_n16295__ & ~new_new_n22145__;
  assign new_new_n22147__ = ~new_new_n11186__ & ~new_new_n22146__;
  assign new_new_n22148__ = ys__n23552 & new_new_n11186__;
  assign new_new_n22149__ = ~new_new_n22147__ & ~new_new_n22148__;
  assign new_new_n22150__ = ~new_new_n11270__ & ~new_new_n22149__;
  assign new_new_n22151__ = new_new_n11270__ & ys__n23489;
  assign new_new_n22152__ = ~new_new_n22150__ & ~new_new_n22151__;
  assign new_new_n22153__ = new_new_n11324__ & ~new_new_n22152__;
  assign new_new_n22154__ = ys__n524 & ~new_new_n11324__;
  assign new_new_n22155__ = ~new_new_n22153__ & ~new_new_n22154__;
  assign new_new_n22156__ = ~new_new_n11343__ & ~new_new_n22155__;
  assign new_new_n22157__ = ~new_new_n11397__ & new_new_n11442__;
  assign new_new_n22158__ = new_new_n11397__ & ~new_new_n11442__;
  assign new_new_n22159__ = ~new_new_n22157__ & ~new_new_n22158__;
  assign new_new_n22160__ = new_new_n11343__ & ~new_new_n22159__;
  assign new_new_n22161__ = ~new_new_n22156__ & ~new_new_n22160__;
  assign new_new_n22162__ = new_new_n11629__ & ~new_new_n22161__;
  assign new_new_n22163__ = ~new_new_n22143__ & ~new_new_n22162__;
  assign new_new_n22164__ = new_new_n11640__ & ~new_new_n22163__;
  assign new_new_n22165__ = ys__n47665 & new_new_n11644__;
  assign new_new_n22166__ = new_new_n11642__ & ~new_new_n22161__;
  assign new_new_n22167__ = ~new_new_n22165__ & ~new_new_n22166__;
  assign new_new_n22168__ = new_new_n11650__ & ~new_new_n22167__;
  assign ys__n24179 = new_new_n22164__ | new_new_n22168__;
  assign new_new_n22170__ = ~ys__n1084 & ~ys__n24177;
  assign new_new_n22171__ = ys__n24197 & new_new_n22170__;
  assign new_new_n22172__ = ys__n24177 & ys__n24209;
  assign new_new_n22173__ = ~new_new_n22171__ & ~new_new_n22172__;
  assign new_new_n22174__ = ~ys__n1078 & ~new_new_n22173__;
  assign new_new_n22175__ = ys__n1078 & ys__n24197;
  assign new_new_n22176__ = ~new_new_n22174__ & ~new_new_n22175__;
  assign new_new_n22177__ = ~new_new_n22139__ & ~new_new_n22176__;
  assign new_new_n22178__ = new_new_n22139__ & ys__n24179;
  assign ys__n24180 = new_new_n22177__ | new_new_n22178__;
  assign new_new_n22180__ = ys__n47666 & new_new_n11634__;
  assign new_new_n22181__ = ys__n22832 & ~new_new_n11180__;
  assign new_new_n22182__ = new_new_n11175__ & new_new_n22181__;
  assign new_new_n22183__ = ~new_new_n16301__ & ~new_new_n22182__;
  assign new_new_n22184__ = ~new_new_n11186__ & ~new_new_n22183__;
  assign new_new_n22185__ = ys__n23554 & new_new_n11186__;
  assign new_new_n22186__ = ~new_new_n22184__ & ~new_new_n22185__;
  assign new_new_n22187__ = ~new_new_n11270__ & ~new_new_n22186__;
  assign new_new_n22188__ = new_new_n11270__ & ys__n23491;
  assign new_new_n22189__ = ~new_new_n22187__ & ~new_new_n22188__;
  assign new_new_n22190__ = new_new_n11324__ & ~new_new_n22189__;
  assign new_new_n22191__ = ys__n522 & ~new_new_n11324__;
  assign new_new_n22192__ = ~new_new_n22190__ & ~new_new_n22191__;
  assign new_new_n22193__ = ~new_new_n11343__ & ~new_new_n22192__;
  assign new_new_n22194__ = ~new_new_n11397__ & ~new_new_n11442__;
  assign new_new_n22195__ = ~new_new_n11447__ & ~new_new_n22194__;
  assign new_new_n22196__ = new_new_n11431__ & ~new_new_n22195__;
  assign new_new_n22197__ = ~new_new_n11431__ & new_new_n22195__;
  assign new_new_n22198__ = ~new_new_n22196__ & ~new_new_n22197__;
  assign new_new_n22199__ = new_new_n11343__ & ~new_new_n22198__;
  assign new_new_n22200__ = ~new_new_n22193__ & ~new_new_n22199__;
  assign new_new_n22201__ = new_new_n11629__ & ~new_new_n22200__;
  assign new_new_n22202__ = ~new_new_n22180__ & ~new_new_n22201__;
  assign new_new_n22203__ = new_new_n11640__ & ~new_new_n22202__;
  assign new_new_n22204__ = ys__n47666 & new_new_n11644__;
  assign new_new_n22205__ = new_new_n11642__ & ~new_new_n22200__;
  assign new_new_n22206__ = ~new_new_n22204__ & ~new_new_n22205__;
  assign new_new_n22207__ = new_new_n11650__ & ~new_new_n22206__;
  assign ys__n24182 = new_new_n22203__ | new_new_n22207__;
  assign new_new_n22209__ = ys__n24199 & new_new_n22170__;
  assign new_new_n22210__ = ys__n24177 & ys__n24211;
  assign new_new_n22211__ = ~new_new_n22209__ & ~new_new_n22210__;
  assign new_new_n22212__ = ~ys__n1078 & ~new_new_n22211__;
  assign new_new_n22213__ = ys__n1078 & ys__n24199;
  assign new_new_n22214__ = ~new_new_n22212__ & ~new_new_n22213__;
  assign new_new_n22215__ = ~new_new_n22139__ & ~new_new_n22214__;
  assign new_new_n22216__ = new_new_n22139__ & ys__n24182;
  assign ys__n24183 = new_new_n22215__ | new_new_n22216__;
  assign new_new_n22218__ = ys__n47667 & new_new_n11634__;
  assign new_new_n22219__ = ys__n22834 & ~new_new_n11180__;
  assign new_new_n22220__ = new_new_n11175__ & new_new_n22219__;
  assign new_new_n22221__ = ~new_new_n16307__ & ~new_new_n22220__;
  assign new_new_n22222__ = ~new_new_n11186__ & ~new_new_n22221__;
  assign new_new_n22223__ = ys__n23556 & new_new_n11186__;
  assign new_new_n22224__ = ~new_new_n22222__ & ~new_new_n22223__;
  assign new_new_n22225__ = ~new_new_n11270__ & ~new_new_n22224__;
  assign new_new_n22226__ = new_new_n11270__ & ys__n23493;
  assign new_new_n22227__ = ~new_new_n22225__ & ~new_new_n22226__;
  assign new_new_n22228__ = new_new_n11324__ & ~new_new_n22227__;
  assign new_new_n22229__ = ys__n530 & ~new_new_n11324__;
  assign new_new_n22230__ = ~new_new_n22228__ & ~new_new_n22229__;
  assign new_new_n22231__ = ~new_new_n11343__ & ~new_new_n22230__;
  assign new_new_n22232__ = ~new_new_n11397__ & new_new_n11443__;
  assign new_new_n22233__ = new_new_n11449__ & ~new_new_n22232__;
  assign new_new_n22234__ = new_new_n11419__ & ~new_new_n22233__;
  assign new_new_n22235__ = ~new_new_n11419__ & new_new_n22233__;
  assign new_new_n22236__ = ~new_new_n22234__ & ~new_new_n22235__;
  assign new_new_n22237__ = new_new_n11343__ & ~new_new_n22236__;
  assign new_new_n22238__ = ~new_new_n22231__ & ~new_new_n22237__;
  assign new_new_n22239__ = new_new_n11629__ & ~new_new_n22238__;
  assign new_new_n22240__ = ~new_new_n22218__ & ~new_new_n22239__;
  assign new_new_n22241__ = new_new_n11640__ & ~new_new_n22240__;
  assign new_new_n22242__ = ys__n47667 & new_new_n11644__;
  assign new_new_n22243__ = new_new_n11642__ & ~new_new_n22238__;
  assign new_new_n22244__ = ~new_new_n22242__ & ~new_new_n22243__;
  assign new_new_n22245__ = new_new_n11650__ & ~new_new_n22244__;
  assign ys__n24185 = new_new_n22241__ | new_new_n22245__;
  assign new_new_n22247__ = ys__n24201 & new_new_n22170__;
  assign new_new_n22248__ = ys__n24177 & ys__n24213;
  assign new_new_n22249__ = ~new_new_n22247__ & ~new_new_n22248__;
  assign new_new_n22250__ = ~ys__n1078 & ~new_new_n22249__;
  assign new_new_n22251__ = ys__n1078 & ys__n24201;
  assign new_new_n22252__ = ~new_new_n22250__ & ~new_new_n22251__;
  assign new_new_n22253__ = ~new_new_n22139__ & ~new_new_n22252__;
  assign new_new_n22254__ = new_new_n22139__ & ys__n24185;
  assign ys__n24186 = new_new_n22253__ | new_new_n22254__;
  assign new_new_n22256__ = ys__n22836 & ~new_new_n11180__;
  assign new_new_n22257__ = new_new_n11175__ & new_new_n22256__;
  assign new_new_n22258__ = ~new_new_n16313__ & ~new_new_n22257__;
  assign new_new_n22259__ = ~new_new_n11186__ & ~new_new_n22258__;
  assign new_new_n22260__ = ys__n23558 & new_new_n11186__;
  assign new_new_n22261__ = ~new_new_n22259__ & ~new_new_n22260__;
  assign new_new_n22262__ = ~new_new_n11270__ & ~new_new_n22261__;
  assign new_new_n22263__ = new_new_n11270__ & ys__n23495;
  assign new_new_n22264__ = ~new_new_n22262__ & ~new_new_n22263__;
  assign new_new_n22265__ = new_new_n11324__ & ~new_new_n22264__;
  assign new_new_n22266__ = ys__n752 & ~new_new_n11324__;
  assign new_new_n22267__ = ~new_new_n22265__ & ~new_new_n22266__;
  assign new_new_n22268__ = ~new_new_n11343__ & ~new_new_n22267__;
  assign new_new_n22269__ = ~new_new_n11419__ & ~new_new_n22233__;
  assign new_new_n22270__ = ~new_new_n11452__ & ~new_new_n22269__;
  assign new_new_n22271__ = new_new_n11408__ & ~new_new_n22270__;
  assign new_new_n22272__ = ~new_new_n11408__ & new_new_n22270__;
  assign new_new_n22273__ = ~new_new_n22271__ & ~new_new_n22272__;
  assign new_new_n22274__ = new_new_n11343__ & ~new_new_n22273__;
  assign new_new_n22275__ = ~new_new_n22268__ & ~new_new_n22274__;
  assign new_new_n22276__ = new_new_n11629__ & ~new_new_n22275__;
  assign new_new_n22277__ = ~ys__n935 & new_new_n11628__;
  assign new_new_n22278__ = ys__n47668 & new_new_n11634__;
  assign new_new_n22279__ = ~new_new_n22277__ & ~new_new_n22278__;
  assign new_new_n22280__ = ~new_new_n22276__ & new_new_n22279__;
  assign new_new_n22281__ = new_new_n11640__ & ~new_new_n22280__;
  assign new_new_n22282__ = new_new_n11642__ & ~new_new_n22275__;
  assign new_new_n22283__ = ys__n47668 & new_new_n11644__;
  assign new_new_n22284__ = ~new_new_n22277__ & ~new_new_n22283__;
  assign new_new_n22285__ = ~new_new_n22282__ & new_new_n22284__;
  assign new_new_n22286__ = new_new_n11650__ & ~new_new_n22285__;
  assign ys__n24188 = new_new_n22281__ | new_new_n22286__;
  assign new_new_n22288__ = ys__n24203 & new_new_n22170__;
  assign new_new_n22289__ = ys__n24177 & ys__n24215;
  assign new_new_n22290__ = ~new_new_n22288__ & ~new_new_n22289__;
  assign new_new_n22291__ = ~ys__n1078 & ~new_new_n22290__;
  assign new_new_n22292__ = ys__n1078 & ys__n24203;
  assign new_new_n22293__ = ~new_new_n22291__ & ~new_new_n22292__;
  assign new_new_n22294__ = ~new_new_n22139__ & ~new_new_n22293__;
  assign new_new_n22295__ = new_new_n22139__ & ys__n24188;
  assign ys__n24189 = new_new_n22294__ | new_new_n22295__;
  assign new_new_n22297__ = ys__n22838 & ~new_new_n11180__;
  assign new_new_n22298__ = new_new_n11175__ & new_new_n22297__;
  assign new_new_n22299__ = ~new_new_n16319__ & ~new_new_n22298__;
  assign new_new_n22300__ = ~new_new_n11186__ & ~new_new_n22299__;
  assign new_new_n22301__ = ys__n23560 & new_new_n11186__;
  assign new_new_n22302__ = ~new_new_n22300__ & ~new_new_n22301__;
  assign new_new_n22303__ = ~new_new_n11270__ & ~new_new_n22302__;
  assign new_new_n22304__ = new_new_n11270__ & ys__n23497;
  assign new_new_n22305__ = ~new_new_n22303__ & ~new_new_n22304__;
  assign new_new_n22306__ = new_new_n11324__ & ~new_new_n22305__;
  assign new_new_n22307__ = ys__n736 & ~new_new_n11324__;
  assign new_new_n22308__ = ~new_new_n22306__ & ~new_new_n22307__;
  assign new_new_n22309__ = ~new_new_n11343__ & ~new_new_n22308__;
  assign new_new_n22310__ = ~new_new_n11456__ & new_new_n11535__;
  assign new_new_n22311__ = new_new_n11456__ & ~new_new_n11535__;
  assign new_new_n22312__ = ~new_new_n22310__ & ~new_new_n22311__;
  assign new_new_n22313__ = new_new_n11343__ & ~new_new_n22312__;
  assign new_new_n22314__ = ~new_new_n22309__ & ~new_new_n22313__;
  assign new_new_n22315__ = new_new_n11629__ & ~new_new_n22314__;
  assign new_new_n22316__ = new_new_n11628__ & new_new_n11631__;
  assign new_new_n22317__ = ys__n47669 & new_new_n11634__;
  assign new_new_n22318__ = ~new_new_n22316__ & ~new_new_n22317__;
  assign new_new_n22319__ = ~new_new_n22315__ & new_new_n22318__;
  assign new_new_n22320__ = new_new_n11640__ & ~new_new_n22319__;
  assign new_new_n22321__ = new_new_n11642__ & ~new_new_n22314__;
  assign new_new_n22322__ = ys__n47669 & new_new_n11644__;
  assign new_new_n22323__ = ~new_new_n22316__ & ~new_new_n22322__;
  assign new_new_n22324__ = ~new_new_n22321__ & new_new_n22323__;
  assign new_new_n22325__ = new_new_n11650__ & ~new_new_n22324__;
  assign ys__n24191 = new_new_n22320__ | new_new_n22325__;
  assign new_new_n22327__ = ys__n24205 & new_new_n22170__;
  assign new_new_n22328__ = ys__n24177 & ys__n24217;
  assign new_new_n22329__ = ~new_new_n22327__ & ~new_new_n22328__;
  assign new_new_n22330__ = ~ys__n1078 & ~new_new_n22329__;
  assign new_new_n22331__ = ys__n1078 & ys__n24205;
  assign new_new_n22332__ = ~new_new_n22330__ & ~new_new_n22331__;
  assign new_new_n22333__ = ~new_new_n22139__ & ~new_new_n22332__;
  assign new_new_n22334__ = new_new_n22139__ & ys__n24191;
  assign ys__n24192 = new_new_n22333__ | new_new_n22334__;
  assign new_new_n22336__ = ys__n22840 & ~new_new_n11180__;
  assign new_new_n22337__ = new_new_n11175__ & new_new_n22336__;
  assign new_new_n22338__ = ~new_new_n16325__ & ~new_new_n22337__;
  assign new_new_n22339__ = ~new_new_n11186__ & ~new_new_n22338__;
  assign new_new_n22340__ = ys__n23562 & new_new_n11186__;
  assign new_new_n22341__ = ~new_new_n22339__ & ~new_new_n22340__;
  assign new_new_n22342__ = ~new_new_n11270__ & ~new_new_n22341__;
  assign new_new_n22343__ = new_new_n11270__ & ys__n23499;
  assign new_new_n22344__ = ~new_new_n22342__ & ~new_new_n22343__;
  assign new_new_n22345__ = new_new_n11324__ & ~new_new_n22344__;
  assign new_new_n22346__ = ys__n4488 & ~new_new_n11324__;
  assign new_new_n22347__ = ~new_new_n22345__ & ~new_new_n22346__;
  assign new_new_n22348__ = ~new_new_n11343__ & ~new_new_n22347__;
  assign new_new_n22349__ = ~new_new_n11456__ & ~new_new_n11535__;
  assign new_new_n22350__ = ~new_new_n11541__ & ~new_new_n22349__;
  assign new_new_n22351__ = new_new_n11525__ & ~new_new_n22350__;
  assign new_new_n22352__ = ~new_new_n11525__ & new_new_n22350__;
  assign new_new_n22353__ = ~new_new_n22351__ & ~new_new_n22352__;
  assign new_new_n22354__ = new_new_n11343__ & ~new_new_n22353__;
  assign new_new_n22355__ = ~new_new_n22348__ & ~new_new_n22354__;
  assign new_new_n22356__ = new_new_n11629__ & ~new_new_n22355__;
  assign new_new_n22357__ = ys__n935 & new_new_n11628__;
  assign new_new_n22358__ = ys__n47670 & new_new_n11634__;
  assign new_new_n22359__ = ~new_new_n22357__ & ~new_new_n22358__;
  assign new_new_n22360__ = ~new_new_n22356__ & new_new_n22359__;
  assign new_new_n22361__ = new_new_n11640__ & ~new_new_n22360__;
  assign new_new_n22362__ = new_new_n11642__ & ~new_new_n22355__;
  assign new_new_n22363__ = ys__n47670 & new_new_n11644__;
  assign new_new_n22364__ = ~new_new_n22357__ & ~new_new_n22363__;
  assign new_new_n22365__ = ~new_new_n22362__ & new_new_n22364__;
  assign new_new_n22366__ = new_new_n11650__ & ~new_new_n22365__;
  assign ys__n24194 = new_new_n22361__ | new_new_n22366__;
  assign new_new_n22368__ = ~ys__n1084 & ys__n24207;
  assign new_new_n22369__ = ys__n312 & ys__n1084;
  assign new_new_n22370__ = ~new_new_n22368__ & ~new_new_n22369__;
  assign new_new_n22371__ = ~ys__n24177 & ~new_new_n22370__;
  assign new_new_n22372__ = ys__n24177 & ys__n24219;
  assign new_new_n22373__ = ~new_new_n22371__ & ~new_new_n22372__;
  assign new_new_n22374__ = ~ys__n1078 & ~new_new_n22373__;
  assign new_new_n22375__ = ys__n1078 & ys__n24207;
  assign new_new_n22376__ = ~new_new_n22374__ & ~new_new_n22375__;
  assign new_new_n22377__ = ~new_new_n22139__ & ~new_new_n22376__;
  assign new_new_n22378__ = new_new_n22139__ & ys__n24194;
  assign ys__n24195 = new_new_n22377__ | new_new_n22378__;
  assign new_new_n22380__ = ys__n318 & ys__n624;
  assign new_new_n22381__ = ys__n18124 & new_new_n22380__;
  assign new_new_n22382__ = ys__n24177 & ~ys__n1079;
  assign new_new_n22383__ = ~new_new_n22381__ & new_new_n22382__;
  assign new_new_n22384__ = ys__n38561 & new_new_n22106__;
  assign new_new_n22385__ = new_new_n22139__ & ~new_new_n22384__;
  assign new_new_n22386__ = ~ys__n18120 & new_new_n22385__;
  assign new_new_n22387__ = new_new_n10596__ & new_new_n22386__;
  assign new_new_n22388__ = ys__n1072 & ~ys__n24228;
  assign new_new_n22389__ = ~ys__n33442 & new_new_n22388__;
  assign new_new_n22390__ = new_new_n16924__ & new_new_n22389__;
  assign new_new_n22391__ = ~ys__n18120 & new_new_n22390__;
  assign new_new_n22392__ = new_new_n22387__ & new_new_n22391__;
  assign ys__n24222 = new_new_n22383__ | new_new_n22392__;
  assign new_new_n22394__ = ys__n1072 & ~ys__n1076;
  assign new_new_n22395__ = ys__n24228 & new_new_n22394__;
  assign new_new_n22396__ = ys__n1076 & ~ys__n24235;
  assign ys__n24227 = new_new_n22395__ | new_new_n22396__;
  assign new_new_n22398__ = ~ys__n24177 & ys__n24233;
  assign new_new_n22399__ = ~ys__n24243 & new_new_n22398__;
  assign new_new_n22400__ = ys__n24177 & new_new_n22381__;
  assign ys__n24231 = new_new_n22399__ | new_new_n22400__;
  assign new_new_n22402__ = ~ys__n1072 & ys__n1078;
  assign new_new_n22403__ = ~ys__n33442 & new_new_n22387__;
  assign new_new_n22404__ = ~ys__n18120 & ~new_new_n22403__;
  assign new_new_n22405__ = ~ys__n18120 & new_new_n16924__;
  assign new_new_n22406__ = ~new_new_n22404__ & new_new_n22405__;
  assign new_new_n22407__ = ~ys__n24243 & new_new_n22388__;
  assign new_new_n22408__ = ~new_new_n22406__ & new_new_n22407__;
  assign new_new_n22409__ = ~new_new_n22402__ & ~new_new_n22408__;
  assign new_new_n22410__ = ~ys__n1076 & ~new_new_n22409__;
  assign new_new_n22411__ = ys__n1076 & ys__n24235;
  assign ys__n24236 = new_new_n22410__ | new_new_n22411__;
  assign ys__n38556 = ys__n24233 & ys__n24243;
  assign new_new_n22414__ = ~ys__n24177 & ~ys__n1079;
  assign new_new_n22415__ = ys__n38556 & new_new_n22414__;
  assign new_new_n22416__ = ys__n24243 & new_new_n22388__;
  assign new_new_n22417__ = ~new_new_n22387__ & new_new_n22416__;
  assign ys__n24240 = new_new_n22415__ | new_new_n22417__;
  assign new_new_n22419__ = ~ys__n1084 & ys__n24248;
  assign new_new_n22420__ = new_new_n22396__ & new_new_n22419__;
  assign new_new_n22421__ = ys__n1084 & ~ys__n18015;
  assign new_new_n22422__ = ~new_new_n22420__ & ~new_new_n22421__;
  assign new_new_n22423__ = ~ys__n140 & ~new_new_n22422__;
  assign ys__n24245 = ys__n140 | new_new_n22423__;
  assign new_new_n22425__ = ~ys__n1076 & ~ys__n24235;
  assign new_new_n22426__ = ys__n24248 & new_new_n22425__;
  assign ys__n24250 = ys__n24235 | new_new_n22426__;
  assign new_new_n22428__ = ~ys__n24464 & ys__n24483;
  assign new_new_n22429__ = ys__n24464 & new_new_n16582__;
  assign new_new_n22430__ = ~new_new_n22428__ & ~new_new_n22429__;
  assign new_new_n22431__ = ~ys__n24463 & ~new_new_n22430__;
  assign new_new_n22432__ = ~new_new_n13990__ & ~new_new_n22431__;
  assign new_new_n22433__ = ~ys__n1120 & ~ys__n24461;
  assign new_new_n22434__ = ~new_new_n22432__ & new_new_n22433__;
  assign new_new_n22435__ = ~ys__n1120 & ~new_new_n22434__;
  assign new_new_n22436__ = ~ys__n1116 & ~ys__n1117;
  assign new_new_n22437__ = ~ys__n1119 & new_new_n22436__;
  assign new_new_n22438__ = ~new_new_n22435__ & new_new_n22437__;
  assign new_new_n22439__ = ys__n690 & ys__n692;
  assign new_new_n22440__ = ys__n694 & ys__n696;
  assign new_new_n22441__ = new_new_n22439__ & new_new_n22440__;
  assign new_new_n22442__ = ys__n606 & ys__n608;
  assign new_new_n22443__ = ys__n610 & ys__n688;
  assign new_new_n22444__ = new_new_n22442__ & new_new_n22443__;
  assign new_new_n22445__ = new_new_n22441__ & new_new_n22444__;
  assign new_new_n22446__ = ~ys__n38654 & ~new_new_n22445__;
  assign new_new_n22447__ = new_new_n16582__ & new_new_n22446__;
  assign new_new_n22448__ = ys__n140 & ys__n1119;
  assign new_new_n22449__ = new_new_n22447__ & new_new_n22448__;
  assign new_new_n22450__ = ~new_new_n22438__ & ~new_new_n22449__;
  assign new_new_n22451__ = new_new_n12497__ & ~new_new_n22450__;
  assign new_new_n22452__ = ~ys__n1110 & ~new_new_n22451__;
  assign new_new_n22453__ = ~ys__n1099 & ~ys__n1109;
  assign new_new_n22454__ = new_new_n12475__ & new_new_n22453__;
  assign new_new_n22455__ = ~new_new_n22452__ & new_new_n22454__;
  assign new_new_n22456__ = ys__n1099 & ys__n24506;
  assign new_new_n22457__ = ~new_new_n22455__ & ~new_new_n22456__;
  assign new_new_n22458__ = ~ys__n1106 & ~new_new_n22457__;
  assign new_new_n22459__ = ys__n1106 & ys__n33495;
  assign new_new_n22460__ = new_new_n16582__ & new_new_n22459__;
  assign new_new_n22461__ = ~ys__n4696 & new_new_n22460__;
  assign new_new_n22462__ = ys__n33481 & new_new_n22461__;
  assign new_new_n22463__ = ~ys__n33493 & ys__n4696;
  assign new_new_n22464__ = ys__n33495 & ~new_new_n22446__;
  assign new_new_n22465__ = ~ys__n33497 & ~new_new_n12472__;
  assign new_new_n22466__ = ys__n1106 & ys__n33491;
  assign new_new_n22467__ = ~new_new_n22465__ & new_new_n22466__;
  assign new_new_n22468__ = ~ys__n24567 & ~ys__n33495;
  assign new_new_n22469__ = ~ys__n33497 & ~ys__n33499;
  assign new_new_n22470__ = new_new_n22468__ & new_new_n22469__;
  assign new_new_n22471__ = new_new_n16582__ & ~new_new_n22470__;
  assign new_new_n22472__ = ~new_new_n22467__ & new_new_n22471__;
  assign new_new_n22473__ = ~ys__n4566 & new_new_n22472__;
  assign new_new_n22474__ = ~new_new_n22464__ & new_new_n22473__;
  assign new_new_n22475__ = ~new_new_n22463__ & new_new_n22474__;
  assign new_new_n22476__ = ~new_new_n22462__ & new_new_n22475__;
  assign new_new_n22477__ = ys__n1106 & ~new_new_n22476__;
  assign new_new_n22478__ = ~new_new_n22458__ & ~new_new_n22477__;
  assign ys__n24502 = ~ys__n1094 & ~new_new_n22478__;
  assign new_new_n22480__ = ys__n1106 & ~ys__n33493;
  assign new_new_n22481__ = ~new_new_n22446__ & new_new_n22480__;
  assign new_new_n22482__ = ~ys__n33493 & ys__n1088;
  assign new_new_n22483__ = ys__n1106 & ys__n33479;
  assign new_new_n22484__ = ~ys__n1119 & ~new_new_n22483__;
  assign new_new_n22485__ = ~new_new_n22482__ & new_new_n22484__;
  assign new_new_n22486__ = ~new_new_n22481__ & new_new_n22485__;
  assign new_new_n22487__ = ~ys__n33495 & ~ys__n33497;
  assign new_new_n22488__ = new_new_n16582__ & ~new_new_n22487__;
  assign new_new_n22489__ = ~new_new_n22486__ & new_new_n22488__;
  assign ys__n24271 = ~ys__n4696 & new_new_n22489__;
  assign new_new_n22491__ = ys__n1106 & ~new_new_n22467__;
  assign new_new_n22492__ = new_new_n22446__ & new_new_n22491__;
  assign new_new_n22493__ = ~ys__n4566 & new_new_n22492__;
  assign new_new_n22494__ = new_new_n22461__ & new_new_n22493__;
  assign ys__n33457 = ~ys__n24271 & new_new_n22494__;
  assign new_new_n22496__ = ys__n24502 & ys__n33457;
  assign ys__n33455 = ys__n24519 & ~new_new_n12476__;
  assign new_new_n22498__ = ys__n38631 & ~ys__n4696;
  assign ys__n38633 = ys__n33455 | new_new_n22498__;
  assign ys__n24258 = ys__n38624 | ~new_new_n16582__;
  assign new_new_n22501__ = ys__n24256 & ~ys__n24258;
  assign new_new_n22502__ = ys__n33497 & ys__n24258;
  assign new_new_n22503__ = ~ys__n4566 & new_new_n22502__;
  assign ys__n24259 = new_new_n22501__ | new_new_n22503__;
  assign new_new_n22505__ = ~ys__n1511 & ys__n30216;
  assign new_new_n22506__ = ~ys__n24258 & new_new_n22505__;
  assign new_new_n22507__ = ~ys__n4566 & new_new_n22506__;
  assign new_new_n22508__ = ys__n38670 & ys__n24258;
  assign new_new_n22509__ = ~ys__n4566 & new_new_n22508__;
  assign ys__n24265 = new_new_n22507__ | new_new_n22509__;
  assign new_new_n22511__ = ~ys__n24259 & ~ys__n24265;
  assign new_new_n22512__ = ~ys__n1106 & ~ys__n1119;
  assign new_new_n22513__ = ~ys__n1120 & ~ys__n24463;
  assign new_new_n22514__ = ~ys__n24464 & new_new_n22513__;
  assign new_new_n22515__ = new_new_n22512__ & new_new_n22514__;
  assign new_new_n22516__ = ~new_new_n22511__ & ~new_new_n22515__;
  assign new_new_n22517__ = ys__n38633 & new_new_n22516__;
  assign new_new_n22518__ = ~new_new_n22496__ & new_new_n22517__;
  assign new_new_n22519__ = ~ys__n33464 & ys__n33488;
  assign new_new_n22520__ = new_new_n12483__ & new_new_n22519__;
  assign ys__n38628 = ~ys__n33481 & new_new_n22461__;
  assign new_new_n22522__ = ~new_new_n12483__ & ys__n38628;
  assign new_new_n22523__ = ~new_new_n22520__ & ~new_new_n22522__;
  assign new_new_n22524__ = ~ys__n24271 & ~new_new_n22523__;
  assign new_new_n22525__ = ys__n24271 & new_new_n22520__;
  assign ys__n24272 = new_new_n22524__ | new_new_n22525__;
  assign new_new_n22527__ = ys__n33552 & ys__n24272;
  assign new_new_n22528__ = new_new_n22511__ & ~new_new_n22527__;
  assign new_new_n22529__ = ys__n38633 & ~new_new_n22515__;
  assign new_new_n22530__ = new_new_n22496__ & new_new_n22529__;
  assign new_new_n22531__ = ~new_new_n22528__ & new_new_n22530__;
  assign ys__n24255 = new_new_n22518__ | new_new_n22531__;
  assign ys__n24260 = ys__n30216 & ~ys__n4566;
  assign new_new_n22534__ = ~ys__n24258 & ys__n24260;
  assign new_new_n22535__ = ys__n33495 & ys__n24258;
  assign new_new_n22536__ = ~ys__n4566 & new_new_n22535__;
  assign ys__n24262 = new_new_n22534__ | new_new_n22536__;
  assign new_new_n22538__ = ~ys__n1511 & ys__n30219;
  assign new_new_n22539__ = ~ys__n24258 & new_new_n22538__;
  assign new_new_n22540__ = ~ys__n4566 & new_new_n22539__;
  assign new_new_n22541__ = ys__n33493 & ys__n24258;
  assign new_new_n22542__ = ~ys__n4566 & new_new_n22541__;
  assign ys__n24268 = new_new_n22540__ | new_new_n22542__;
  assign ys__n24274 = ~ys__n24107 & ys__n24279;
  assign new_new_n22545__ = ~ys__n454 & ~ys__n38693;
  assign new_new_n22546__ = ys__n454 & ys__n38693;
  assign new_new_n22547__ = ~new_new_n22545__ & ~new_new_n22546__;
  assign new_new_n22548__ = ~ys__n24112 & ~new_new_n22547__;
  assign new_new_n22549__ = ~ys__n452 & ys__n24112;
  assign new_new_n22550__ = ~new_new_n22548__ & ~new_new_n22549__;
  assign new_new_n22551__ = ~ys__n1088 & ys__n1089;
  assign new_new_n22552__ = ~new_new_n22550__ & new_new_n22551__;
  assign new_new_n22553__ = ys__n1088 & ys__n24274;
  assign ys__n24275 = new_new_n22552__ | new_new_n22553__;
  assign ys__n24277 = ~ys__n24107 & ys__n24280;
  assign new_new_n22556__ = ys__n454 & ~ys__n712;
  assign new_new_n22557__ = ~ys__n454 & ys__n712;
  assign ys__n35425 = new_new_n22556__ | new_new_n22557__;
  assign new_new_n22559__ = ~ys__n38694 & ys__n35425;
  assign new_new_n22560__ = ys__n38694 & ~ys__n35425;
  assign new_new_n22561__ = ~new_new_n22559__ & ~new_new_n22560__;
  assign new_new_n22562__ = ~ys__n24112 & ~new_new_n22561__;
  assign new_new_n22563__ = ys__n452 & ~ys__n35426;
  assign new_new_n22564__ = ~ys__n452 & ys__n35426;
  assign new_new_n22565__ = ~new_new_n22563__ & ~new_new_n22564__;
  assign new_new_n22566__ = ys__n24112 & ~new_new_n22565__;
  assign new_new_n22567__ = ~new_new_n22562__ & ~new_new_n22566__;
  assign new_new_n22568__ = new_new_n22551__ & ~new_new_n22567__;
  assign new_new_n22569__ = ys__n1088 & ys__n24277;
  assign ys__n24278 = new_new_n22568__ | new_new_n22569__;
  assign new_new_n22571__ = ~ys__n80 & ~ys__n82;
  assign new_new_n22572__ = ys__n84 & ys__n86;
  assign new_new_n22573__ = new_new_n22571__ & new_new_n22572__;
  assign new_new_n22574__ = ys__n84 & ~ys__n86;
  assign new_new_n22575__ = new_new_n22571__ & new_new_n22574__;
  assign new_new_n22576__ = ~new_new_n22573__ & ~new_new_n22575__;
  assign new_new_n22577__ = ~ys__n84 & ys__n86;
  assign new_new_n22578__ = new_new_n22571__ & new_new_n22577__;
  assign new_new_n22579__ = ~ys__n84 & ~ys__n86;
  assign new_new_n22580__ = new_new_n22571__ & new_new_n22579__;
  assign new_new_n22581__ = ~new_new_n22578__ & ~new_new_n22580__;
  assign new_new_n22582__ = new_new_n22576__ & new_new_n22581__;
  assign new_new_n22583__ = ys__n80 & ~ys__n82;
  assign new_new_n22584__ = new_new_n22574__ & new_new_n22583__;
  assign new_new_n22585__ = new_new_n22579__ & new_new_n22583__;
  assign new_new_n22586__ = ~new_new_n22584__ & ~new_new_n22585__;
  assign new_new_n22587__ = new_new_n22582__ & new_new_n22586__;
  assign new_new_n22588__ = ys__n80 & ys__n82;
  assign new_new_n22589__ = new_new_n22579__ & new_new_n22588__;
  assign new_new_n22590__ = new_new_n22587__ & ~new_new_n22589__;
  assign new_new_n22591__ = ~new_new_n22587__ & ~new_new_n22590__;
  assign new_new_n22592__ = ys__n47194 & ~new_new_n22591__;
  assign new_new_n22593__ = ~new_new_n22575__ & ~new_new_n22584__;
  assign new_new_n22594__ = ys__n47193 & ~new_new_n22593__;
  assign new_new_n22595__ = ~new_new_n22580__ & ~new_new_n22585__;
  assign new_new_n22596__ = ys__n47201 & ~new_new_n22595__;
  assign new_new_n22597__ = ys__n47009 & new_new_n22578__;
  assign new_new_n22598__ = ys__n47001 & new_new_n22573__;
  assign new_new_n22599__ = ~new_new_n22597__ & ~new_new_n22598__;
  assign new_new_n22600__ = ~new_new_n22596__ & new_new_n22599__;
  assign new_new_n22601__ = ~new_new_n22594__ & new_new_n22600__;
  assign new_new_n22602__ = ~new_new_n22573__ & ~new_new_n22578__;
  assign new_new_n22603__ = new_new_n22593__ & new_new_n22595__;
  assign new_new_n22604__ = new_new_n22602__ & new_new_n22603__;
  assign new_new_n22605__ = ys__n38898 & ~new_new_n22604__;
  assign new_new_n22606__ = ~new_new_n22601__ & new_new_n22605__;
  assign new_new_n22607__ = new_new_n22591__ & new_new_n22606__;
  assign new_new_n22608__ = ~new_new_n22592__ & ~new_new_n22607__;
  assign new_new_n22609__ = ys__n18149 & ys__n18137;
  assign new_new_n22610__ = new_new_n16221__ & new_new_n22609__;
  assign new_new_n22611__ = ~ys__n1154 & ~ys__n38805;
  assign new_new_n22612__ = ~new_new_n22610__ & new_new_n22611__;
  assign new_new_n22613__ = new_new_n10609__ & ~new_new_n22612__;
  assign new_new_n22614__ = ~new_new_n22608__ & ~new_new_n22613__;
  assign new_new_n22615__ = ~ys__n1106 & ~ys__n1109;
  assign new_new_n22616__ = ~ys__n1116 & new_new_n22615__;
  assign new_new_n22617__ = new_new_n22614__ & new_new_n22616__;
  assign new_new_n22618__ = ~ys__n4176 & new_new_n10609__;
  assign new_new_n22619__ = ys__n33407 & new_new_n22618__;
  assign new_new_n22620__ = ys__n28932 & new_new_n22619__;
  assign new_new_n22621__ = ys__n33409 & new_new_n22618__;
  assign new_new_n22622__ = ys__n29286 & new_new_n22621__;
  assign new_new_n22623__ = ys__n33411 & new_new_n22618__;
  assign new_new_n22624__ = ys__n29593 & new_new_n22623__;
  assign new_new_n22625__ = ys__n29594 & ~new_new_n22623__;
  assign new_new_n22626__ = ~new_new_n22624__ & ~new_new_n22625__;
  assign new_new_n22627__ = ~new_new_n22621__ & ~new_new_n22626__;
  assign new_new_n22628__ = ~new_new_n22622__ & ~new_new_n22627__;
  assign new_new_n22629__ = ~new_new_n22619__ & ~new_new_n22628__;
  assign new_new_n22630__ = ~new_new_n22620__ & ~new_new_n22629__;
  assign new_new_n22631__ = ~new_new_n22616__ & ~new_new_n22630__;
  assign ys__n24286 = new_new_n22617__ | new_new_n22631__;
  assign new_new_n22633__ = ys__n47195 & ~new_new_n22591__;
  assign new_new_n22634__ = ~new_new_n22607__ & ~new_new_n22633__;
  assign new_new_n22635__ = ~new_new_n22613__ & ~new_new_n22634__;
  assign new_new_n22636__ = new_new_n22616__ & new_new_n22635__;
  assign new_new_n22637__ = ys__n28935 & new_new_n22619__;
  assign new_new_n22638__ = ys__n29288 & new_new_n22621__;
  assign new_new_n22639__ = ys__n29595 & new_new_n22623__;
  assign new_new_n22640__ = ys__n29596 & ~new_new_n22623__;
  assign new_new_n22641__ = ~new_new_n22639__ & ~new_new_n22640__;
  assign new_new_n22642__ = ~new_new_n22621__ & ~new_new_n22641__;
  assign new_new_n22643__ = ~new_new_n22638__ & ~new_new_n22642__;
  assign new_new_n22644__ = ~new_new_n22619__ & ~new_new_n22643__;
  assign new_new_n22645__ = ~new_new_n22637__ & ~new_new_n22644__;
  assign new_new_n22646__ = ~new_new_n22616__ & ~new_new_n22645__;
  assign ys__n24289 = new_new_n22636__ | new_new_n22646__;
  assign new_new_n22648__ = ys__n47196 & ~new_new_n22591__;
  assign new_new_n22649__ = ~new_new_n22607__ & ~new_new_n22648__;
  assign new_new_n22650__ = ~new_new_n22613__ & ~new_new_n22649__;
  assign new_new_n22651__ = new_new_n22616__ & new_new_n22650__;
  assign new_new_n22652__ = ys__n28938 & new_new_n22619__;
  assign new_new_n22653__ = ys__n29290 & new_new_n22621__;
  assign new_new_n22654__ = ys__n29597 & new_new_n22623__;
  assign new_new_n22655__ = ys__n29598 & ~new_new_n22623__;
  assign new_new_n22656__ = ~new_new_n22654__ & ~new_new_n22655__;
  assign new_new_n22657__ = ~new_new_n22621__ & ~new_new_n22656__;
  assign new_new_n22658__ = ~new_new_n22653__ & ~new_new_n22657__;
  assign new_new_n22659__ = ~new_new_n22619__ & ~new_new_n22658__;
  assign new_new_n22660__ = ~new_new_n22652__ & ~new_new_n22659__;
  assign new_new_n22661__ = ~new_new_n22616__ & ~new_new_n22660__;
  assign ys__n24291 = new_new_n22651__ | new_new_n22661__;
  assign new_new_n22663__ = ys__n47197 & ~new_new_n22591__;
  assign new_new_n22664__ = ~new_new_n22607__ & ~new_new_n22663__;
  assign new_new_n22665__ = ~new_new_n22613__ & ~new_new_n22664__;
  assign new_new_n22666__ = new_new_n22616__ & new_new_n22665__;
  assign new_new_n22667__ = ys__n28941 & new_new_n22619__;
  assign new_new_n22668__ = ys__n29292 & new_new_n22621__;
  assign new_new_n22669__ = ys__n29599 & new_new_n22623__;
  assign new_new_n22670__ = ys__n29600 & ~new_new_n22623__;
  assign new_new_n22671__ = ~new_new_n22669__ & ~new_new_n22670__;
  assign new_new_n22672__ = ~new_new_n22621__ & ~new_new_n22671__;
  assign new_new_n22673__ = ~new_new_n22668__ & ~new_new_n22672__;
  assign new_new_n22674__ = ~new_new_n22619__ & ~new_new_n22673__;
  assign new_new_n22675__ = ~new_new_n22667__ & ~new_new_n22674__;
  assign new_new_n22676__ = ~new_new_n22616__ & ~new_new_n22675__;
  assign ys__n24293 = new_new_n22666__ | new_new_n22676__;
  assign new_new_n22678__ = ys__n47198 & ~new_new_n22591__;
  assign new_new_n22679__ = ~new_new_n22607__ & ~new_new_n22678__;
  assign new_new_n22680__ = ~new_new_n22613__ & ~new_new_n22679__;
  assign new_new_n22681__ = new_new_n22616__ & new_new_n22680__;
  assign new_new_n22682__ = ys__n28944 & new_new_n22619__;
  assign new_new_n22683__ = ys__n29294 & new_new_n22621__;
  assign new_new_n22684__ = ys__n29601 & new_new_n22623__;
  assign new_new_n22685__ = ys__n29602 & ~new_new_n22623__;
  assign new_new_n22686__ = ~new_new_n22684__ & ~new_new_n22685__;
  assign new_new_n22687__ = ~new_new_n22621__ & ~new_new_n22686__;
  assign new_new_n22688__ = ~new_new_n22683__ & ~new_new_n22687__;
  assign new_new_n22689__ = ~new_new_n22619__ & ~new_new_n22688__;
  assign new_new_n22690__ = ~new_new_n22682__ & ~new_new_n22689__;
  assign new_new_n22691__ = ~new_new_n22616__ & ~new_new_n22690__;
  assign ys__n24295 = new_new_n22681__ | new_new_n22691__;
  assign new_new_n22693__ = ys__n47199 & ~new_new_n22591__;
  assign new_new_n22694__ = ~new_new_n22607__ & ~new_new_n22693__;
  assign new_new_n22695__ = ~new_new_n22613__ & ~new_new_n22694__;
  assign new_new_n22696__ = new_new_n22616__ & new_new_n22695__;
  assign new_new_n22697__ = ys__n28947 & new_new_n22619__;
  assign new_new_n22698__ = ys__n29296 & new_new_n22621__;
  assign new_new_n22699__ = ys__n29603 & new_new_n22623__;
  assign new_new_n22700__ = ys__n29604 & ~new_new_n22623__;
  assign new_new_n22701__ = ~new_new_n22699__ & ~new_new_n22700__;
  assign new_new_n22702__ = ~new_new_n22621__ & ~new_new_n22701__;
  assign new_new_n22703__ = ~new_new_n22698__ & ~new_new_n22702__;
  assign new_new_n22704__ = ~new_new_n22619__ & ~new_new_n22703__;
  assign new_new_n22705__ = ~new_new_n22697__ & ~new_new_n22704__;
  assign new_new_n22706__ = ~new_new_n22616__ & ~new_new_n22705__;
  assign ys__n24297 = new_new_n22696__ | new_new_n22706__;
  assign new_new_n22708__ = ys__n47200 & ~new_new_n22591__;
  assign new_new_n22709__ = ~new_new_n22607__ & ~new_new_n22708__;
  assign new_new_n22710__ = ~new_new_n22613__ & ~new_new_n22709__;
  assign new_new_n22711__ = new_new_n22616__ & new_new_n22710__;
  assign new_new_n22712__ = ys__n28950 & new_new_n22619__;
  assign new_new_n22713__ = ys__n29298 & new_new_n22621__;
  assign new_new_n22714__ = ys__n29605 & new_new_n22623__;
  assign new_new_n22715__ = ys__n29606 & ~new_new_n22623__;
  assign new_new_n22716__ = ~new_new_n22714__ & ~new_new_n22715__;
  assign new_new_n22717__ = ~new_new_n22621__ & ~new_new_n22716__;
  assign new_new_n22718__ = ~new_new_n22713__ & ~new_new_n22717__;
  assign new_new_n22719__ = ~new_new_n22619__ & ~new_new_n22718__;
  assign new_new_n22720__ = ~new_new_n22712__ & ~new_new_n22719__;
  assign new_new_n22721__ = ~new_new_n22616__ & ~new_new_n22720__;
  assign ys__n24299 = new_new_n22711__ | new_new_n22721__;
  assign new_new_n22723__ = ys__n47201 & ~new_new_n22591__;
  assign new_new_n22724__ = ~new_new_n22607__ & ~new_new_n22723__;
  assign new_new_n22725__ = ~new_new_n22613__ & ~new_new_n22724__;
  assign new_new_n22726__ = new_new_n22616__ & new_new_n22725__;
  assign new_new_n22727__ = ys__n28953 & new_new_n22619__;
  assign new_new_n22728__ = ys__n29300 & new_new_n22621__;
  assign new_new_n22729__ = ys__n29607 & new_new_n22623__;
  assign new_new_n22730__ = ys__n29608 & ~new_new_n22623__;
  assign new_new_n22731__ = ~new_new_n22729__ & ~new_new_n22730__;
  assign new_new_n22732__ = ~new_new_n22621__ & ~new_new_n22731__;
  assign new_new_n22733__ = ~new_new_n22728__ & ~new_new_n22732__;
  assign new_new_n22734__ = ~new_new_n22619__ & ~new_new_n22733__;
  assign new_new_n22735__ = ~new_new_n22727__ & ~new_new_n22734__;
  assign new_new_n22736__ = ~new_new_n22616__ & ~new_new_n22735__;
  assign ys__n24301 = new_new_n22726__ | new_new_n22736__;
  assign new_new_n22738__ = ~ys__n33469 & new_new_n12473__;
  assign new_new_n22739__ = ys__n1107 & ys__n2693;
  assign new_new_n22740__ = new_new_n13987__ & new_new_n22739__;
  assign new_new_n22741__ = ~new_new_n22738__ & ~new_new_n22740__;
  assign new_new_n22742__ = ys__n24286 & new_new_n22741__;
  assign new_new_n22743__ = ys__n24303 & new_new_n22740__;
  assign ys__n24305 = new_new_n22742__ | new_new_n22743__;
  assign new_new_n22745__ = ys__n24289 & new_new_n22741__;
  assign new_new_n22746__ = ys__n24306 & new_new_n22740__;
  assign ys__n24307 = new_new_n22745__ | new_new_n22746__;
  assign new_new_n22748__ = ys__n24291 & new_new_n22741__;
  assign new_new_n22749__ = ys__n24308 & new_new_n22740__;
  assign ys__n24309 = new_new_n22748__ | new_new_n22749__;
  assign new_new_n22751__ = ys__n24293 & new_new_n22741__;
  assign new_new_n22752__ = ys__n24310 & new_new_n22740__;
  assign ys__n24311 = new_new_n22751__ | new_new_n22752__;
  assign new_new_n22754__ = ys__n24295 & new_new_n22741__;
  assign new_new_n22755__ = ys__n24312 & new_new_n22740__;
  assign ys__n24313 = new_new_n22754__ | new_new_n22755__;
  assign new_new_n22757__ = ys__n24297 & new_new_n22741__;
  assign new_new_n22758__ = ys__n24314 & new_new_n22740__;
  assign ys__n24315 = new_new_n22757__ | new_new_n22758__;
  assign new_new_n22760__ = ys__n24299 & new_new_n22741__;
  assign new_new_n22761__ = ys__n24316 & new_new_n22740__;
  assign ys__n24317 = new_new_n22760__ | new_new_n22761__;
  assign new_new_n22763__ = ys__n24301 & new_new_n22741__;
  assign new_new_n22764__ = ys__n24318 & new_new_n22740__;
  assign ys__n24319 = new_new_n22763__ | new_new_n22764__;
  assign new_new_n22766__ = ys__n47002 & ~new_new_n22591__;
  assign new_new_n22767__ = ~new_new_n22607__ & ~new_new_n22766__;
  assign new_new_n22768__ = ~new_new_n22613__ & ~new_new_n22767__;
  assign new_new_n22769__ = new_new_n22616__ & new_new_n22768__;
  assign new_new_n22770__ = ys__n28908 & new_new_n22619__;
  assign new_new_n22771__ = ys__n29270 & new_new_n22621__;
  assign new_new_n22772__ = ys__n29577 & new_new_n22623__;
  assign new_new_n22773__ = ys__n29578 & ~new_new_n22623__;
  assign new_new_n22774__ = ~new_new_n22772__ & ~new_new_n22773__;
  assign new_new_n22775__ = ~new_new_n22621__ & ~new_new_n22774__;
  assign new_new_n22776__ = ~new_new_n22771__ & ~new_new_n22775__;
  assign new_new_n22777__ = ~new_new_n22619__ & ~new_new_n22776__;
  assign new_new_n22778__ = ~new_new_n22770__ & ~new_new_n22777__;
  assign new_new_n22779__ = ~new_new_n22616__ & ~new_new_n22778__;
  assign ys__n24320 = new_new_n22769__ | new_new_n22779__;
  assign new_new_n22781__ = ys__n47003 & ~new_new_n22591__;
  assign new_new_n22782__ = ~new_new_n22607__ & ~new_new_n22781__;
  assign new_new_n22783__ = ~new_new_n22613__ & ~new_new_n22782__;
  assign new_new_n22784__ = new_new_n22616__ & new_new_n22783__;
  assign new_new_n22785__ = ys__n28911 & new_new_n22619__;
  assign new_new_n22786__ = ys__n29272 & new_new_n22621__;
  assign new_new_n22787__ = ys__n29579 & new_new_n22623__;
  assign new_new_n22788__ = ys__n29580 & ~new_new_n22623__;
  assign new_new_n22789__ = ~new_new_n22787__ & ~new_new_n22788__;
  assign new_new_n22790__ = ~new_new_n22621__ & ~new_new_n22789__;
  assign new_new_n22791__ = ~new_new_n22786__ & ~new_new_n22790__;
  assign new_new_n22792__ = ~new_new_n22619__ & ~new_new_n22791__;
  assign new_new_n22793__ = ~new_new_n22785__ & ~new_new_n22792__;
  assign new_new_n22794__ = ~new_new_n22616__ & ~new_new_n22793__;
  assign ys__n24323 = new_new_n22784__ | new_new_n22794__;
  assign new_new_n22796__ = ys__n47004 & ~new_new_n22591__;
  assign new_new_n22797__ = ~new_new_n22607__ & ~new_new_n22796__;
  assign new_new_n22798__ = ~new_new_n22613__ & ~new_new_n22797__;
  assign new_new_n22799__ = new_new_n22616__ & new_new_n22798__;
  assign new_new_n22800__ = ys__n28914 & new_new_n22619__;
  assign new_new_n22801__ = ys__n29274 & new_new_n22621__;
  assign new_new_n22802__ = ys__n29581 & new_new_n22623__;
  assign new_new_n22803__ = ys__n29582 & ~new_new_n22623__;
  assign new_new_n22804__ = ~new_new_n22802__ & ~new_new_n22803__;
  assign new_new_n22805__ = ~new_new_n22621__ & ~new_new_n22804__;
  assign new_new_n22806__ = ~new_new_n22801__ & ~new_new_n22805__;
  assign new_new_n22807__ = ~new_new_n22619__ & ~new_new_n22806__;
  assign new_new_n22808__ = ~new_new_n22800__ & ~new_new_n22807__;
  assign new_new_n22809__ = ~new_new_n22616__ & ~new_new_n22808__;
  assign ys__n24325 = new_new_n22799__ | new_new_n22809__;
  assign new_new_n22811__ = ys__n47005 & ~new_new_n22591__;
  assign new_new_n22812__ = ~new_new_n22607__ & ~new_new_n22811__;
  assign new_new_n22813__ = ~new_new_n22613__ & ~new_new_n22812__;
  assign new_new_n22814__ = new_new_n22616__ & new_new_n22813__;
  assign new_new_n22815__ = ys__n28917 & new_new_n22619__;
  assign new_new_n22816__ = ys__n29276 & new_new_n22621__;
  assign new_new_n22817__ = ys__n29583 & new_new_n22623__;
  assign new_new_n22818__ = ys__n29584 & ~new_new_n22623__;
  assign new_new_n22819__ = ~new_new_n22817__ & ~new_new_n22818__;
  assign new_new_n22820__ = ~new_new_n22621__ & ~new_new_n22819__;
  assign new_new_n22821__ = ~new_new_n22816__ & ~new_new_n22820__;
  assign new_new_n22822__ = ~new_new_n22619__ & ~new_new_n22821__;
  assign new_new_n22823__ = ~new_new_n22815__ & ~new_new_n22822__;
  assign new_new_n22824__ = ~new_new_n22616__ & ~new_new_n22823__;
  assign ys__n24327 = new_new_n22814__ | new_new_n22824__;
  assign new_new_n22826__ = ys__n47006 & ~new_new_n22591__;
  assign new_new_n22827__ = ~new_new_n22607__ & ~new_new_n22826__;
  assign new_new_n22828__ = ~new_new_n22613__ & ~new_new_n22827__;
  assign new_new_n22829__ = new_new_n22616__ & new_new_n22828__;
  assign new_new_n22830__ = ys__n28920 & new_new_n22619__;
  assign new_new_n22831__ = ys__n29278 & new_new_n22621__;
  assign new_new_n22832__ = ys__n29585 & new_new_n22623__;
  assign new_new_n22833__ = ys__n29586 & ~new_new_n22623__;
  assign new_new_n22834__ = ~new_new_n22832__ & ~new_new_n22833__;
  assign new_new_n22835__ = ~new_new_n22621__ & ~new_new_n22834__;
  assign new_new_n22836__ = ~new_new_n22831__ & ~new_new_n22835__;
  assign new_new_n22837__ = ~new_new_n22619__ & ~new_new_n22836__;
  assign new_new_n22838__ = ~new_new_n22830__ & ~new_new_n22837__;
  assign new_new_n22839__ = ~new_new_n22616__ & ~new_new_n22838__;
  assign ys__n24329 = new_new_n22829__ | new_new_n22839__;
  assign new_new_n22841__ = ys__n47007 & ~new_new_n22591__;
  assign new_new_n22842__ = ~new_new_n22607__ & ~new_new_n22841__;
  assign new_new_n22843__ = ~new_new_n22613__ & ~new_new_n22842__;
  assign new_new_n22844__ = new_new_n22616__ & new_new_n22843__;
  assign new_new_n22845__ = ys__n28923 & new_new_n22619__;
  assign new_new_n22846__ = ys__n29280 & new_new_n22621__;
  assign new_new_n22847__ = ys__n29587 & new_new_n22623__;
  assign new_new_n22848__ = ys__n29588 & ~new_new_n22623__;
  assign new_new_n22849__ = ~new_new_n22847__ & ~new_new_n22848__;
  assign new_new_n22850__ = ~new_new_n22621__ & ~new_new_n22849__;
  assign new_new_n22851__ = ~new_new_n22846__ & ~new_new_n22850__;
  assign new_new_n22852__ = ~new_new_n22619__ & ~new_new_n22851__;
  assign new_new_n22853__ = ~new_new_n22845__ & ~new_new_n22852__;
  assign new_new_n22854__ = ~new_new_n22616__ & ~new_new_n22853__;
  assign ys__n24331 = new_new_n22844__ | new_new_n22854__;
  assign new_new_n22856__ = ys__n47008 & ~new_new_n22591__;
  assign new_new_n22857__ = ~new_new_n22607__ & ~new_new_n22856__;
  assign new_new_n22858__ = ~new_new_n22613__ & ~new_new_n22857__;
  assign new_new_n22859__ = new_new_n22616__ & new_new_n22858__;
  assign new_new_n22860__ = ys__n28926 & new_new_n22619__;
  assign new_new_n22861__ = ys__n29282 & new_new_n22621__;
  assign new_new_n22862__ = ys__n29589 & new_new_n22623__;
  assign new_new_n22863__ = ys__n29590 & ~new_new_n22623__;
  assign new_new_n22864__ = ~new_new_n22862__ & ~new_new_n22863__;
  assign new_new_n22865__ = ~new_new_n22621__ & ~new_new_n22864__;
  assign new_new_n22866__ = ~new_new_n22861__ & ~new_new_n22865__;
  assign new_new_n22867__ = ~new_new_n22619__ & ~new_new_n22866__;
  assign new_new_n22868__ = ~new_new_n22860__ & ~new_new_n22867__;
  assign new_new_n22869__ = ~new_new_n22616__ & ~new_new_n22868__;
  assign ys__n24333 = new_new_n22859__ | new_new_n22869__;
  assign new_new_n22871__ = ys__n47009 & ~new_new_n22591__;
  assign new_new_n22872__ = ~new_new_n22607__ & ~new_new_n22871__;
  assign new_new_n22873__ = ~new_new_n22613__ & ~new_new_n22872__;
  assign new_new_n22874__ = new_new_n22616__ & new_new_n22873__;
  assign new_new_n22875__ = ys__n28929 & new_new_n22619__;
  assign new_new_n22876__ = ys__n29284 & new_new_n22621__;
  assign new_new_n22877__ = ys__n29591 & new_new_n22623__;
  assign new_new_n22878__ = ys__n29592 & ~new_new_n22623__;
  assign new_new_n22879__ = ~new_new_n22877__ & ~new_new_n22878__;
  assign new_new_n22880__ = ~new_new_n22621__ & ~new_new_n22879__;
  assign new_new_n22881__ = ~new_new_n22876__ & ~new_new_n22880__;
  assign new_new_n22882__ = ~new_new_n22619__ & ~new_new_n22881__;
  assign new_new_n22883__ = ~new_new_n22875__ & ~new_new_n22882__;
  assign new_new_n22884__ = ~new_new_n22616__ & ~new_new_n22883__;
  assign ys__n24335 = new_new_n22874__ | new_new_n22884__;
  assign new_new_n22886__ = ~ys__n33471 & new_new_n12473__;
  assign new_new_n22887__ = ys__n16 & ys__n1107;
  assign new_new_n22888__ = new_new_n13987__ & new_new_n22887__;
  assign new_new_n22889__ = ~new_new_n22886__ & ~new_new_n22888__;
  assign new_new_n22890__ = ys__n24320 & new_new_n22889__;
  assign new_new_n22891__ = ys__n24337 & new_new_n22888__;
  assign ys__n24339 = new_new_n22890__ | new_new_n22891__;
  assign new_new_n22893__ = ys__n24323 & new_new_n22889__;
  assign new_new_n22894__ = ys__n24340 & new_new_n22888__;
  assign ys__n24341 = new_new_n22893__ | new_new_n22894__;
  assign new_new_n22896__ = ys__n24325 & new_new_n22889__;
  assign new_new_n22897__ = ys__n24342 & new_new_n22888__;
  assign ys__n24343 = new_new_n22896__ | new_new_n22897__;
  assign new_new_n22899__ = ys__n24327 & new_new_n22889__;
  assign new_new_n22900__ = ys__n24344 & new_new_n22888__;
  assign ys__n24345 = new_new_n22899__ | new_new_n22900__;
  assign new_new_n22902__ = ys__n24329 & new_new_n22889__;
  assign new_new_n22903__ = ys__n24346 & new_new_n22888__;
  assign ys__n24347 = new_new_n22902__ | new_new_n22903__;
  assign new_new_n22905__ = ys__n24331 & new_new_n22889__;
  assign new_new_n22906__ = ys__n24348 & new_new_n22888__;
  assign ys__n24349 = new_new_n22905__ | new_new_n22906__;
  assign new_new_n22908__ = ys__n24333 & new_new_n22889__;
  assign new_new_n22909__ = ys__n24350 & new_new_n22888__;
  assign ys__n24351 = new_new_n22908__ | new_new_n22909__;
  assign new_new_n22911__ = ys__n24335 & new_new_n22889__;
  assign new_new_n22912__ = ys__n24352 & new_new_n22888__;
  assign ys__n24353 = new_new_n22911__ | new_new_n22912__;
  assign new_new_n22914__ = new_new_n22581__ & ~new_new_n22585__;
  assign new_new_n22915__ = ~new_new_n22584__ & ~new_new_n22589__;
  assign new_new_n22916__ = new_new_n22576__ & new_new_n22915__;
  assign new_new_n22917__ = new_new_n22914__ & new_new_n22916__;
  assign new_new_n22918__ = ~new_new_n22914__ & ~new_new_n22917__;
  assign new_new_n22919__ = ys__n47186 & ~new_new_n22918__;
  assign new_new_n22920__ = ys__n47194 & new_new_n22918__;
  assign new_new_n22921__ = ~new_new_n22919__ & ~new_new_n22920__;
  assign new_new_n22922__ = new_new_n22586__ & ~new_new_n22589__;
  assign new_new_n22923__ = new_new_n22582__ & new_new_n22922__;
  assign new_new_n22924__ = ~new_new_n22582__ & ~new_new_n22923__;
  assign new_new_n22925__ = ~new_new_n22921__ & ~new_new_n22924__;
  assign new_new_n22926__ = new_new_n22606__ & new_new_n22924__;
  assign new_new_n22927__ = ~new_new_n22925__ & ~new_new_n22926__;
  assign new_new_n22928__ = ~new_new_n22613__ & ~new_new_n22927__;
  assign new_new_n22929__ = new_new_n22616__ & new_new_n22928__;
  assign new_new_n22930__ = ys__n28884 & new_new_n22619__;
  assign new_new_n22931__ = ys__n29254 & new_new_n22621__;
  assign new_new_n22932__ = ys__n29561 & new_new_n22623__;
  assign new_new_n22933__ = ys__n29562 & ~new_new_n22623__;
  assign new_new_n22934__ = ~new_new_n22932__ & ~new_new_n22933__;
  assign new_new_n22935__ = ~new_new_n22621__ & ~new_new_n22934__;
  assign new_new_n22936__ = ~new_new_n22931__ & ~new_new_n22935__;
  assign new_new_n22937__ = ~new_new_n22619__ & ~new_new_n22936__;
  assign new_new_n22938__ = ~new_new_n22930__ & ~new_new_n22937__;
  assign new_new_n22939__ = ~new_new_n22616__ & ~new_new_n22938__;
  assign ys__n24354 = new_new_n22929__ | new_new_n22939__;
  assign new_new_n22941__ = ys__n47187 & ~new_new_n22918__;
  assign new_new_n22942__ = ys__n47195 & new_new_n22918__;
  assign new_new_n22943__ = ~new_new_n22941__ & ~new_new_n22942__;
  assign new_new_n22944__ = ~new_new_n22924__ & ~new_new_n22943__;
  assign new_new_n22945__ = ~new_new_n22926__ & ~new_new_n22944__;
  assign new_new_n22946__ = ~new_new_n22613__ & ~new_new_n22945__;
  assign new_new_n22947__ = new_new_n22616__ & new_new_n22946__;
  assign new_new_n22948__ = ys__n28887 & new_new_n22619__;
  assign new_new_n22949__ = ys__n29256 & new_new_n22621__;
  assign new_new_n22950__ = ys__n29563 & new_new_n22623__;
  assign new_new_n22951__ = ys__n29564 & ~new_new_n22623__;
  assign new_new_n22952__ = ~new_new_n22950__ & ~new_new_n22951__;
  assign new_new_n22953__ = ~new_new_n22621__ & ~new_new_n22952__;
  assign new_new_n22954__ = ~new_new_n22949__ & ~new_new_n22953__;
  assign new_new_n22955__ = ~new_new_n22619__ & ~new_new_n22954__;
  assign new_new_n22956__ = ~new_new_n22948__ & ~new_new_n22955__;
  assign new_new_n22957__ = ~new_new_n22616__ & ~new_new_n22956__;
  assign ys__n24357 = new_new_n22947__ | new_new_n22957__;
  assign new_new_n22959__ = ys__n47188 & ~new_new_n22918__;
  assign new_new_n22960__ = ys__n47196 & new_new_n22918__;
  assign new_new_n22961__ = ~new_new_n22959__ & ~new_new_n22960__;
  assign new_new_n22962__ = ~new_new_n22924__ & ~new_new_n22961__;
  assign new_new_n22963__ = ~new_new_n22926__ & ~new_new_n22962__;
  assign new_new_n22964__ = ~new_new_n22613__ & ~new_new_n22963__;
  assign new_new_n22965__ = new_new_n22616__ & new_new_n22964__;
  assign new_new_n22966__ = ys__n28890 & new_new_n22619__;
  assign new_new_n22967__ = ys__n29258 & new_new_n22621__;
  assign new_new_n22968__ = ys__n29565 & new_new_n22623__;
  assign new_new_n22969__ = ys__n29566 & ~new_new_n22623__;
  assign new_new_n22970__ = ~new_new_n22968__ & ~new_new_n22969__;
  assign new_new_n22971__ = ~new_new_n22621__ & ~new_new_n22970__;
  assign new_new_n22972__ = ~new_new_n22967__ & ~new_new_n22971__;
  assign new_new_n22973__ = ~new_new_n22619__ & ~new_new_n22972__;
  assign new_new_n22974__ = ~new_new_n22966__ & ~new_new_n22973__;
  assign new_new_n22975__ = ~new_new_n22616__ & ~new_new_n22974__;
  assign ys__n24359 = new_new_n22965__ | new_new_n22975__;
  assign new_new_n22977__ = ys__n47189 & ~new_new_n22918__;
  assign new_new_n22978__ = ys__n47197 & new_new_n22918__;
  assign new_new_n22979__ = ~new_new_n22977__ & ~new_new_n22978__;
  assign new_new_n22980__ = ~new_new_n22924__ & ~new_new_n22979__;
  assign new_new_n22981__ = ~new_new_n22926__ & ~new_new_n22980__;
  assign new_new_n22982__ = ~new_new_n22613__ & ~new_new_n22981__;
  assign new_new_n22983__ = new_new_n22616__ & new_new_n22982__;
  assign new_new_n22984__ = ys__n28893 & new_new_n22619__;
  assign new_new_n22985__ = ys__n29260 & new_new_n22621__;
  assign new_new_n22986__ = ys__n29567 & new_new_n22623__;
  assign new_new_n22987__ = ys__n29568 & ~new_new_n22623__;
  assign new_new_n22988__ = ~new_new_n22986__ & ~new_new_n22987__;
  assign new_new_n22989__ = ~new_new_n22621__ & ~new_new_n22988__;
  assign new_new_n22990__ = ~new_new_n22985__ & ~new_new_n22989__;
  assign new_new_n22991__ = ~new_new_n22619__ & ~new_new_n22990__;
  assign new_new_n22992__ = ~new_new_n22984__ & ~new_new_n22991__;
  assign new_new_n22993__ = ~new_new_n22616__ & ~new_new_n22992__;
  assign ys__n24361 = new_new_n22983__ | new_new_n22993__;
  assign new_new_n22995__ = ys__n47190 & ~new_new_n22918__;
  assign new_new_n22996__ = ys__n47198 & new_new_n22918__;
  assign new_new_n22997__ = ~new_new_n22995__ & ~new_new_n22996__;
  assign new_new_n22998__ = ~new_new_n22924__ & ~new_new_n22997__;
  assign new_new_n22999__ = ~new_new_n22926__ & ~new_new_n22998__;
  assign new_new_n23000__ = ~new_new_n22613__ & ~new_new_n22999__;
  assign new_new_n23001__ = new_new_n22616__ & new_new_n23000__;
  assign new_new_n23002__ = ys__n28896 & new_new_n22619__;
  assign new_new_n23003__ = ys__n29262 & new_new_n22621__;
  assign new_new_n23004__ = ys__n29569 & new_new_n22623__;
  assign new_new_n23005__ = ys__n29570 & ~new_new_n22623__;
  assign new_new_n23006__ = ~new_new_n23004__ & ~new_new_n23005__;
  assign new_new_n23007__ = ~new_new_n22621__ & ~new_new_n23006__;
  assign new_new_n23008__ = ~new_new_n23003__ & ~new_new_n23007__;
  assign new_new_n23009__ = ~new_new_n22619__ & ~new_new_n23008__;
  assign new_new_n23010__ = ~new_new_n23002__ & ~new_new_n23009__;
  assign new_new_n23011__ = ~new_new_n22616__ & ~new_new_n23010__;
  assign ys__n24363 = new_new_n23001__ | new_new_n23011__;
  assign new_new_n23013__ = ys__n47191 & ~new_new_n22918__;
  assign new_new_n23014__ = ys__n47199 & new_new_n22918__;
  assign new_new_n23015__ = ~new_new_n23013__ & ~new_new_n23014__;
  assign new_new_n23016__ = ~new_new_n22924__ & ~new_new_n23015__;
  assign new_new_n23017__ = ~new_new_n22926__ & ~new_new_n23016__;
  assign new_new_n23018__ = ~new_new_n22613__ & ~new_new_n23017__;
  assign new_new_n23019__ = new_new_n22616__ & new_new_n23018__;
  assign new_new_n23020__ = ys__n28899 & new_new_n22619__;
  assign new_new_n23021__ = ys__n29264 & new_new_n22621__;
  assign new_new_n23022__ = ys__n29571 & new_new_n22623__;
  assign new_new_n23023__ = ys__n29572 & ~new_new_n22623__;
  assign new_new_n23024__ = ~new_new_n23022__ & ~new_new_n23023__;
  assign new_new_n23025__ = ~new_new_n22621__ & ~new_new_n23024__;
  assign new_new_n23026__ = ~new_new_n23021__ & ~new_new_n23025__;
  assign new_new_n23027__ = ~new_new_n22619__ & ~new_new_n23026__;
  assign new_new_n23028__ = ~new_new_n23020__ & ~new_new_n23027__;
  assign new_new_n23029__ = ~new_new_n22616__ & ~new_new_n23028__;
  assign ys__n24365 = new_new_n23019__ | new_new_n23029__;
  assign new_new_n23031__ = ys__n47192 & ~new_new_n22918__;
  assign new_new_n23032__ = ys__n47200 & new_new_n22918__;
  assign new_new_n23033__ = ~new_new_n23031__ & ~new_new_n23032__;
  assign new_new_n23034__ = ~new_new_n22924__ & ~new_new_n23033__;
  assign new_new_n23035__ = ~new_new_n22926__ & ~new_new_n23034__;
  assign new_new_n23036__ = ~new_new_n22613__ & ~new_new_n23035__;
  assign new_new_n23037__ = new_new_n22616__ & new_new_n23036__;
  assign new_new_n23038__ = ys__n28902 & new_new_n22619__;
  assign new_new_n23039__ = ys__n29266 & new_new_n22621__;
  assign new_new_n23040__ = ys__n29573 & new_new_n22623__;
  assign new_new_n23041__ = ys__n29574 & ~new_new_n22623__;
  assign new_new_n23042__ = ~new_new_n23040__ & ~new_new_n23041__;
  assign new_new_n23043__ = ~new_new_n22621__ & ~new_new_n23042__;
  assign new_new_n23044__ = ~new_new_n23039__ & ~new_new_n23043__;
  assign new_new_n23045__ = ~new_new_n22619__ & ~new_new_n23044__;
  assign new_new_n23046__ = ~new_new_n23038__ & ~new_new_n23045__;
  assign new_new_n23047__ = ~new_new_n22616__ & ~new_new_n23046__;
  assign ys__n24367 = new_new_n23037__ | new_new_n23047__;
  assign new_new_n23049__ = ys__n47193 & ~new_new_n22918__;
  assign new_new_n23050__ = ys__n47201 & new_new_n22918__;
  assign new_new_n23051__ = ~new_new_n23049__ & ~new_new_n23050__;
  assign new_new_n23052__ = ~new_new_n22924__ & ~new_new_n23051__;
  assign new_new_n23053__ = ~new_new_n22926__ & ~new_new_n23052__;
  assign new_new_n23054__ = ~new_new_n22613__ & ~new_new_n23053__;
  assign new_new_n23055__ = new_new_n22616__ & new_new_n23054__;
  assign new_new_n23056__ = ys__n28905 & new_new_n22619__;
  assign new_new_n23057__ = ys__n29268 & new_new_n22621__;
  assign new_new_n23058__ = ys__n29575 & new_new_n22623__;
  assign new_new_n23059__ = ys__n29576 & ~new_new_n22623__;
  assign new_new_n23060__ = ~new_new_n23058__ & ~new_new_n23059__;
  assign new_new_n23061__ = ~new_new_n22621__ & ~new_new_n23060__;
  assign new_new_n23062__ = ~new_new_n23057__ & ~new_new_n23061__;
  assign new_new_n23063__ = ~new_new_n22619__ & ~new_new_n23062__;
  assign new_new_n23064__ = ~new_new_n23056__ & ~new_new_n23063__;
  assign new_new_n23065__ = ~new_new_n22616__ & ~new_new_n23064__;
  assign ys__n24369 = new_new_n23055__ | new_new_n23065__;
  assign new_new_n23067__ = ~ys__n33473 & new_new_n12473__;
  assign new_new_n23068__ = ys__n14 & ys__n1107;
  assign new_new_n23069__ = new_new_n13987__ & new_new_n23068__;
  assign new_new_n23070__ = ~new_new_n23067__ & ~new_new_n23069__;
  assign new_new_n23071__ = ys__n24354 & new_new_n23070__;
  assign new_new_n23072__ = ys__n24371 & new_new_n23069__;
  assign ys__n24373 = new_new_n23071__ | new_new_n23072__;
  assign new_new_n23074__ = ys__n24357 & new_new_n23070__;
  assign new_new_n23075__ = ys__n24374 & new_new_n23069__;
  assign ys__n24375 = new_new_n23074__ | new_new_n23075__;
  assign new_new_n23077__ = ys__n24359 & new_new_n23070__;
  assign new_new_n23078__ = ys__n24376 & new_new_n23069__;
  assign ys__n24377 = new_new_n23077__ | new_new_n23078__;
  assign new_new_n23080__ = ys__n24361 & new_new_n23070__;
  assign new_new_n23081__ = ys__n24378 & new_new_n23069__;
  assign ys__n24379 = new_new_n23080__ | new_new_n23081__;
  assign new_new_n23083__ = ys__n24363 & new_new_n23070__;
  assign new_new_n23084__ = ys__n24380 & new_new_n23069__;
  assign ys__n24381 = new_new_n23083__ | new_new_n23084__;
  assign new_new_n23086__ = ys__n24365 & new_new_n23070__;
  assign new_new_n23087__ = ys__n24382 & new_new_n23069__;
  assign ys__n24383 = new_new_n23086__ | new_new_n23087__;
  assign new_new_n23089__ = ys__n24367 & new_new_n23070__;
  assign new_new_n23090__ = ys__n24384 & new_new_n23069__;
  assign ys__n24385 = new_new_n23089__ | new_new_n23090__;
  assign new_new_n23092__ = ys__n24369 & new_new_n23070__;
  assign new_new_n23093__ = ys__n24386 & new_new_n23069__;
  assign ys__n24387 = new_new_n23092__ | new_new_n23093__;
  assign new_new_n23095__ = ~ys__n1154 & ys__n24575;
  assign new_new_n23096__ = ~ys__n90 & ~ys__n4736;
  assign new_new_n23097__ = ~ys__n88 & ~ys__n4736;
  assign new_new_n23098__ = ys__n1154 & ys__n47448;
  assign new_new_n23099__ = ~new_new_n23097__ & new_new_n23098__;
  assign new_new_n23100__ = ~new_new_n23096__ & new_new_n23099__;
  assign new_new_n23101__ = ~new_new_n23095__ & ~new_new_n23100__;
  assign new_new_n23102__ = new_new_n22613__ & ~new_new_n23101__;
  assign new_new_n23103__ = ys__n46994 & ~new_new_n22918__;
  assign new_new_n23104__ = ys__n47002 & new_new_n22918__;
  assign new_new_n23105__ = ~new_new_n23103__ & ~new_new_n23104__;
  assign new_new_n23106__ = ~new_new_n22575__ & ~new_new_n22580__;
  assign new_new_n23107__ = new_new_n22602__ & new_new_n23106__;
  assign new_new_n23108__ = new_new_n22922__ & new_new_n23107__;
  assign new_new_n23109__ = ~new_new_n23106__ & ~new_new_n23108__;
  assign new_new_n23110__ = ~new_new_n23105__ & ~new_new_n23109__;
  assign new_new_n23111__ = ~new_new_n22921__ & new_new_n23109__;
  assign new_new_n23112__ = ~new_new_n23110__ & ~new_new_n23111__;
  assign new_new_n23113__ = ~new_new_n22613__ & ~new_new_n23112__;
  assign new_new_n23114__ = ~new_new_n23102__ & ~new_new_n23113__;
  assign new_new_n23115__ = new_new_n22616__ & ~new_new_n23114__;
  assign new_new_n23116__ = ys__n28859 & new_new_n22619__;
  assign new_new_n23117__ = ys__n29237 & new_new_n22621__;
  assign new_new_n23118__ = ys__n29550 & new_new_n22623__;
  assign new_new_n23119__ = ys__n28462 & ~new_new_n22623__;
  assign new_new_n23120__ = ~new_new_n23118__ & ~new_new_n23119__;
  assign new_new_n23121__ = ~new_new_n22621__ & ~new_new_n23120__;
  assign new_new_n23122__ = ~new_new_n23117__ & ~new_new_n23121__;
  assign new_new_n23123__ = ~new_new_n22619__ & ~new_new_n23122__;
  assign new_new_n23124__ = ~new_new_n23116__ & ~new_new_n23123__;
  assign new_new_n23125__ = ~new_new_n22616__ & ~new_new_n23124__;
  assign ys__n24388 = new_new_n23115__ | new_new_n23125__;
  assign new_new_n23127__ = ys__n46995 & ~new_new_n22918__;
  assign new_new_n23128__ = ys__n47003 & new_new_n22918__;
  assign new_new_n23129__ = ~new_new_n23127__ & ~new_new_n23128__;
  assign new_new_n23130__ = ~new_new_n23109__ & ~new_new_n23129__;
  assign new_new_n23131__ = ~new_new_n22943__ & new_new_n23109__;
  assign new_new_n23132__ = ~new_new_n23130__ & ~new_new_n23131__;
  assign new_new_n23133__ = ~new_new_n22613__ & ~new_new_n23132__;
  assign new_new_n23134__ = new_new_n22616__ & new_new_n23133__;
  assign new_new_n23135__ = ys__n28863 & new_new_n22619__;
  assign new_new_n23136__ = ys__n29240 & new_new_n22621__;
  assign new_new_n23137__ = ys__n29552 & new_new_n22623__;
  assign new_new_n23138__ = ys__n28464 & ~new_new_n22623__;
  assign new_new_n23139__ = ~new_new_n23137__ & ~new_new_n23138__;
  assign new_new_n23140__ = ~new_new_n22621__ & ~new_new_n23139__;
  assign new_new_n23141__ = ~new_new_n23136__ & ~new_new_n23140__;
  assign new_new_n23142__ = ~new_new_n22619__ & ~new_new_n23141__;
  assign new_new_n23143__ = ~new_new_n23135__ & ~new_new_n23142__;
  assign new_new_n23144__ = ~new_new_n22616__ & ~new_new_n23143__;
  assign ys__n24392 = new_new_n23134__ | new_new_n23144__;
  assign new_new_n23146__ = ys__n46996 & ~new_new_n22918__;
  assign new_new_n23147__ = ys__n47004 & new_new_n22918__;
  assign new_new_n23148__ = ~new_new_n23146__ & ~new_new_n23147__;
  assign new_new_n23149__ = ~new_new_n23109__ & ~new_new_n23148__;
  assign new_new_n23150__ = ~new_new_n22961__ & new_new_n23109__;
  assign new_new_n23151__ = ~new_new_n23149__ & ~new_new_n23150__;
  assign new_new_n23152__ = ~new_new_n22613__ & ~new_new_n23151__;
  assign new_new_n23153__ = new_new_n22616__ & new_new_n23152__;
  assign new_new_n23154__ = ys__n28866 & new_new_n22619__;
  assign new_new_n23155__ = ys__n29242 & new_new_n22621__;
  assign new_new_n23156__ = ys__n29553 & new_new_n22623__;
  assign new_new_n23157__ = ys__n28466 & ~new_new_n22623__;
  assign new_new_n23158__ = ~new_new_n23156__ & ~new_new_n23157__;
  assign new_new_n23159__ = ~new_new_n22621__ & ~new_new_n23158__;
  assign new_new_n23160__ = ~new_new_n23155__ & ~new_new_n23159__;
  assign new_new_n23161__ = ~new_new_n22619__ & ~new_new_n23160__;
  assign new_new_n23162__ = ~new_new_n23154__ & ~new_new_n23161__;
  assign new_new_n23163__ = ~new_new_n22616__ & ~new_new_n23162__;
  assign ys__n24394 = new_new_n23153__ | new_new_n23163__;
  assign new_new_n23165__ = ys__n46997 & ~new_new_n22918__;
  assign new_new_n23166__ = ys__n47005 & new_new_n22918__;
  assign new_new_n23167__ = ~new_new_n23165__ & ~new_new_n23166__;
  assign new_new_n23168__ = ~new_new_n23109__ & ~new_new_n23167__;
  assign new_new_n23169__ = ~new_new_n22979__ & new_new_n23109__;
  assign new_new_n23170__ = ~new_new_n23168__ & ~new_new_n23169__;
  assign new_new_n23171__ = ~new_new_n22613__ & ~new_new_n23170__;
  assign new_new_n23172__ = new_new_n22616__ & new_new_n23171__;
  assign new_new_n23173__ = ys__n28869 & new_new_n22619__;
  assign new_new_n23174__ = ys__n29244 & new_new_n22621__;
  assign new_new_n23175__ = ys__n29554 & new_new_n22623__;
  assign new_new_n23176__ = ys__n28468 & ~new_new_n22623__;
  assign new_new_n23177__ = ~new_new_n23175__ & ~new_new_n23176__;
  assign new_new_n23178__ = ~new_new_n22621__ & ~new_new_n23177__;
  assign new_new_n23179__ = ~new_new_n23174__ & ~new_new_n23178__;
  assign new_new_n23180__ = ~new_new_n22619__ & ~new_new_n23179__;
  assign new_new_n23181__ = ~new_new_n23173__ & ~new_new_n23180__;
  assign new_new_n23182__ = ~new_new_n22616__ & ~new_new_n23181__;
  assign ys__n24396 = new_new_n23172__ | new_new_n23182__;
  assign new_new_n23184__ = ys__n46998 & ~new_new_n22918__;
  assign new_new_n23185__ = ys__n47006 & new_new_n22918__;
  assign new_new_n23186__ = ~new_new_n23184__ & ~new_new_n23185__;
  assign new_new_n23187__ = ~new_new_n23109__ & ~new_new_n23186__;
  assign new_new_n23188__ = ~new_new_n22997__ & new_new_n23109__;
  assign new_new_n23189__ = ~new_new_n23187__ & ~new_new_n23188__;
  assign new_new_n23190__ = ~new_new_n22613__ & ~new_new_n23189__;
  assign new_new_n23191__ = new_new_n22616__ & new_new_n23190__;
  assign new_new_n23192__ = ys__n28872 & new_new_n22619__;
  assign new_new_n23193__ = ys__n29246 & new_new_n22621__;
  assign new_new_n23194__ = ys__n29555 & new_new_n22623__;
  assign new_new_n23195__ = ys__n28470 & ~new_new_n22623__;
  assign new_new_n23196__ = ~new_new_n23194__ & ~new_new_n23195__;
  assign new_new_n23197__ = ~new_new_n22621__ & ~new_new_n23196__;
  assign new_new_n23198__ = ~new_new_n23193__ & ~new_new_n23197__;
  assign new_new_n23199__ = ~new_new_n22619__ & ~new_new_n23198__;
  assign new_new_n23200__ = ~new_new_n23192__ & ~new_new_n23199__;
  assign new_new_n23201__ = ~new_new_n22616__ & ~new_new_n23200__;
  assign ys__n24398 = new_new_n23191__ | new_new_n23201__;
  assign new_new_n23203__ = ys__n46999 & ~new_new_n22918__;
  assign new_new_n23204__ = ys__n47007 & new_new_n22918__;
  assign new_new_n23205__ = ~new_new_n23203__ & ~new_new_n23204__;
  assign new_new_n23206__ = ~new_new_n23109__ & ~new_new_n23205__;
  assign new_new_n23207__ = ~new_new_n23015__ & new_new_n23109__;
  assign new_new_n23208__ = ~new_new_n23206__ & ~new_new_n23207__;
  assign new_new_n23209__ = ~new_new_n22613__ & ~new_new_n23208__;
  assign new_new_n23210__ = new_new_n22616__ & new_new_n23209__;
  assign new_new_n23211__ = ys__n28875 & new_new_n22619__;
  assign new_new_n23212__ = ys__n29248 & new_new_n22621__;
  assign new_new_n23213__ = ys__n29556 & new_new_n22623__;
  assign new_new_n23214__ = ys__n28472 & ~new_new_n22623__;
  assign new_new_n23215__ = ~new_new_n23213__ & ~new_new_n23214__;
  assign new_new_n23216__ = ~new_new_n22621__ & ~new_new_n23215__;
  assign new_new_n23217__ = ~new_new_n23212__ & ~new_new_n23216__;
  assign new_new_n23218__ = ~new_new_n22619__ & ~new_new_n23217__;
  assign new_new_n23219__ = ~new_new_n23211__ & ~new_new_n23218__;
  assign new_new_n23220__ = ~new_new_n22616__ & ~new_new_n23219__;
  assign ys__n24400 = new_new_n23210__ | new_new_n23220__;
  assign new_new_n23222__ = ys__n47000 & ~new_new_n22918__;
  assign new_new_n23223__ = ys__n47008 & new_new_n22918__;
  assign new_new_n23224__ = ~new_new_n23222__ & ~new_new_n23223__;
  assign new_new_n23225__ = ~new_new_n23109__ & ~new_new_n23224__;
  assign new_new_n23226__ = ~new_new_n23033__ & new_new_n23109__;
  assign new_new_n23227__ = ~new_new_n23225__ & ~new_new_n23226__;
  assign new_new_n23228__ = ~new_new_n22613__ & ~new_new_n23227__;
  assign new_new_n23229__ = new_new_n22616__ & new_new_n23228__;
  assign new_new_n23230__ = ys__n28878 & new_new_n22619__;
  assign new_new_n23231__ = ys__n29250 & new_new_n22621__;
  assign new_new_n23232__ = ys__n29557 & new_new_n22623__;
  assign new_new_n23233__ = ys__n29558 & ~new_new_n22623__;
  assign new_new_n23234__ = ~new_new_n23232__ & ~new_new_n23233__;
  assign new_new_n23235__ = ~new_new_n22621__ & ~new_new_n23234__;
  assign new_new_n23236__ = ~new_new_n23231__ & ~new_new_n23235__;
  assign new_new_n23237__ = ~new_new_n22619__ & ~new_new_n23236__;
  assign new_new_n23238__ = ~new_new_n23230__ & ~new_new_n23237__;
  assign new_new_n23239__ = ~new_new_n22616__ & ~new_new_n23238__;
  assign ys__n24402 = new_new_n23229__ | new_new_n23239__;
  assign new_new_n23241__ = ys__n47001 & ~new_new_n22918__;
  assign new_new_n23242__ = ys__n47009 & new_new_n22918__;
  assign new_new_n23243__ = ~new_new_n23241__ & ~new_new_n23242__;
  assign new_new_n23244__ = ~new_new_n23109__ & ~new_new_n23243__;
  assign new_new_n23245__ = ~new_new_n23051__ & new_new_n23109__;
  assign new_new_n23246__ = ~new_new_n23244__ & ~new_new_n23245__;
  assign new_new_n23247__ = ~new_new_n22613__ & ~new_new_n23246__;
  assign new_new_n23248__ = new_new_n22616__ & new_new_n23247__;
  assign new_new_n23249__ = ys__n28881 & new_new_n22619__;
  assign new_new_n23250__ = ys__n29252 & new_new_n22621__;
  assign new_new_n23251__ = ys__n29559 & new_new_n22623__;
  assign new_new_n23252__ = ys__n29560 & ~new_new_n22623__;
  assign new_new_n23253__ = ~new_new_n23251__ & ~new_new_n23252__;
  assign new_new_n23254__ = ~new_new_n22621__ & ~new_new_n23253__;
  assign new_new_n23255__ = ~new_new_n23250__ & ~new_new_n23254__;
  assign new_new_n23256__ = ~new_new_n22619__ & ~new_new_n23255__;
  assign new_new_n23257__ = ~new_new_n23249__ & ~new_new_n23256__;
  assign new_new_n23258__ = ~new_new_n22616__ & ~new_new_n23257__;
  assign ys__n24404 = new_new_n23248__ | new_new_n23258__;
  assign new_new_n23260__ = ~ys__n33475 & new_new_n12473__;
  assign new_new_n23261__ = ys__n24388 & ~new_new_n23260__;
  assign new_new_n23262__ = ys__n24389 & new_new_n23260__;
  assign new_new_n23263__ = ~new_new_n23261__ & ~new_new_n23262__;
  assign new_new_n23264__ = ys__n1107 & ys__n4688;
  assign new_new_n23265__ = new_new_n13987__ & new_new_n23264__;
  assign new_new_n23266__ = ~new_new_n23263__ & ~new_new_n23265__;
  assign new_new_n23267__ = ys__n24406 & new_new_n23265__;
  assign ys__n24408 = new_new_n23266__ | new_new_n23267__;
  assign new_new_n23269__ = ~new_new_n23260__ & ~new_new_n23265__;
  assign new_new_n23270__ = ys__n24392 & new_new_n23269__;
  assign new_new_n23271__ = ys__n24409 & new_new_n23265__;
  assign ys__n24410 = new_new_n23270__ | new_new_n23271__;
  assign new_new_n23273__ = ys__n24394 & new_new_n23269__;
  assign new_new_n23274__ = ys__n24411 & new_new_n23265__;
  assign ys__n24412 = new_new_n23273__ | new_new_n23274__;
  assign new_new_n23276__ = ys__n24396 & new_new_n23269__;
  assign new_new_n23277__ = ys__n24413 & new_new_n23265__;
  assign ys__n24414 = new_new_n23276__ | new_new_n23277__;
  assign new_new_n23279__ = ys__n24398 & new_new_n23269__;
  assign new_new_n23280__ = ys__n24415 & new_new_n23265__;
  assign ys__n24416 = new_new_n23279__ | new_new_n23280__;
  assign new_new_n23282__ = ys__n24400 & new_new_n23269__;
  assign new_new_n23283__ = ys__n24417 & new_new_n23265__;
  assign ys__n24418 = new_new_n23282__ | new_new_n23283__;
  assign new_new_n23285__ = ys__n24402 & new_new_n23269__;
  assign new_new_n23286__ = ys__n24419 & new_new_n23265__;
  assign ys__n24420 = new_new_n23285__ | new_new_n23286__;
  assign new_new_n23288__ = ys__n24404 & new_new_n23269__;
  assign new_new_n23289__ = ys__n24421 & new_new_n23265__;
  assign ys__n24422 = new_new_n23288__ | new_new_n23289__;
  assign new_new_n23291__ = ~ys__n1116 & new_new_n12476__;
  assign new_new_n23292__ = ys__n24279 & new_new_n23291__;
  assign new_new_n23293__ = ys__n452 & ~new_new_n23291__;
  assign new_new_n23294__ = ~new_new_n23292__ & ~new_new_n23293__;
  assign new_new_n23295__ = ~ys__n1109 & ~ys__n1116;
  assign new_new_n23296__ = ~ys__n1117 & new_new_n23295__;
  assign new_new_n23297__ = ~new_new_n23294__ & new_new_n23296__;
  assign new_new_n23298__ = ys__n24427 & ~new_new_n23296__;
  assign new_new_n23299__ = ~new_new_n23297__ & ~new_new_n23298__;
  assign new_new_n23300__ = ys__n33495 & new_new_n22446__;
  assign new_new_n23301__ = ~ys__n24258 & ~new_new_n22515__;
  assign new_new_n23302__ = ~new_new_n23300__ & new_new_n23301__;
  assign new_new_n23303__ = ~new_new_n23299__ & ~new_new_n23302__;
  assign new_new_n23304__ = ys__n20008 & new_new_n23302__;
  assign ys__n24425 = new_new_n23303__ | new_new_n23304__;
  assign new_new_n23306__ = ys__n1094 & ~ys__n1147;
  assign new_new_n23307__ = ~ys__n24433 & ys__n24434;
  assign new_new_n23308__ = new_new_n23306__ & new_new_n23307__;
  assign new_new_n23309__ = ys__n1147 & ~ys__n18019;
  assign new_new_n23310__ = ~new_new_n23308__ & ~new_new_n23309__;
  assign new_new_n23311__ = ~ys__n140 & ~new_new_n23310__;
  assign ys__n24430 = ys__n140 | new_new_n23311__;
  assign new_new_n23313__ = ~ys__n1094 & ~ys__n24433;
  assign new_new_n23314__ = ys__n24434 & new_new_n23313__;
  assign ys__n24436 = ys__n24433 | new_new_n23314__;
  assign new_new_n23316__ = ys__n454 & ys__n712;
  assign ys__n24470 = ys__n24519 & new_new_n23316__;
  assign new_new_n23318__ = ~ys__n1098 & ~ys__n1099;
  assign new_new_n23319__ = ys__n1107 & new_new_n23318__;
  assign new_new_n23320__ = ~ys__n24470 & new_new_n23319__;
  assign new_new_n23321__ = ys__n1099 & ~ys__n24506;
  assign new_new_n23322__ = ys__n33488 & new_new_n23321__;
  assign ys__n24440 = new_new_n23320__ | new_new_n23322__;
  assign new_new_n23324__ = ys__n1098 & ~ys__n1099;
  assign new_new_n23325__ = ~ys__n24470 & new_new_n23324__;
  assign new_new_n23326__ = ~ys__n33488 & new_new_n23321__;
  assign ys__n24445 = new_new_n23325__ | new_new_n23326__;
  assign new_new_n23328__ = ~ys__n1107 & ~ys__n1110;
  assign new_new_n23329__ = new_new_n22615__ & new_new_n23328__;
  assign new_new_n23330__ = new_new_n23318__ & new_new_n23329__;
  assign new_new_n23331__ = ~ys__n1129 & ~ys__n24461;
  assign new_new_n23332__ = ~ys__n24463 & new_new_n23331__;
  assign new_new_n23333__ = new_new_n12500__ & new_new_n22436__;
  assign new_new_n23334__ = new_new_n23332__ & new_new_n23333__;
  assign new_new_n23335__ = new_new_n23330__ & new_new_n23334__;
  assign new_new_n23336__ = new_new_n16590__ & new_new_n23335__;
  assign new_new_n23337__ = ys__n33493 & new_new_n16582__;
  assign new_new_n23338__ = ys__n1106 & ~ys__n33491;
  assign new_new_n23339__ = new_new_n23337__ & new_new_n23338__;
  assign new_new_n23340__ = ~ys__n4566 & new_new_n23339__;
  assign new_new_n23341__ = ys__n4696 & new_new_n23340__;
  assign new_new_n23342__ = ~new_new_n23336__ & ~new_new_n23341__;
  assign ys__n24447 = ~ys__n1094 & ~new_new_n23342__;
  assign new_new_n23344__ = new_new_n12475__ & new_new_n12488__;
  assign new_new_n23345__ = new_new_n23333__ & new_new_n23344__;
  assign new_new_n23346__ = ~ys__n24483 & ys__n24485;
  assign new_new_n23347__ = ~ys__n24567 & new_new_n23346__;
  assign new_new_n23348__ = ~ys__n24463 & ~ys__n24464;
  assign new_new_n23349__ = new_new_n23331__ & new_new_n23348__;
  assign new_new_n23350__ = new_new_n23347__ & new_new_n23349__;
  assign new_new_n23351__ = new_new_n23345__ & new_new_n23350__;
  assign new_new_n23352__ = ys__n1098 & ys__n24470;
  assign new_new_n23353__ = ~new_new_n23351__ & ~new_new_n23352__;
  assign new_new_n23354__ = ~ys__n1099 & new_new_n12483__;
  assign new_new_n23355__ = ~new_new_n23353__ & new_new_n23354__;
  assign new_new_n23356__ = ys__n1094 & ys__n24433;
  assign ys__n24466 = new_new_n23355__ | new_new_n23356__;
  assign new_new_n23358__ = ys__n1119 & ~ys__n1129;
  assign new_new_n23359__ = new_new_n23328__ & new_new_n23358__;
  assign new_new_n23360__ = new_new_n22615__ & new_new_n23318__;
  assign new_new_n23361__ = new_new_n23359__ & new_new_n23360__;
  assign new_new_n23362__ = new_new_n16582__ & new_new_n23361__;
  assign new_new_n23363__ = ~new_new_n22446__ & new_new_n23362__;
  assign new_new_n23364__ = ys__n33481 & ys__n33497;
  assign new_new_n23365__ = new_new_n23338__ & new_new_n23364__;
  assign new_new_n23366__ = new_new_n16582__ & new_new_n23365__;
  assign new_new_n23367__ = ~new_new_n22446__ & new_new_n23366__;
  assign new_new_n23368__ = ~ys__n4566 & new_new_n23367__;
  assign new_new_n23369__ = ~ys__n4696 & new_new_n23368__;
  assign ys__n24488 = new_new_n23363__ | new_new_n23369__;
  assign new_new_n23371__ = ~ys__n1094 & ys__n1106;
  assign new_new_n23372__ = ys__n33499 & new_new_n22487__;
  assign new_new_n23373__ = new_new_n23371__ & new_new_n23372__;
  assign new_new_n23374__ = new_new_n16582__ & new_new_n23373__;
  assign new_new_n23375__ = ~ys__n4566 & new_new_n23374__;
  assign new_new_n23376__ = ys__n1094 & ~ys__n24433;
  assign ys__n24499 = new_new_n23375__ | new_new_n23376__;
  assign new_new_n23378__ = ~ys__n140 & ys__n1119;
  assign new_new_n23379__ = ~ys__n1129 & new_new_n23378__;
  assign new_new_n23380__ = new_new_n22447__ & new_new_n23379__;
  assign new_new_n23381__ = ys__n1129 & ~ys__n24470;
  assign ys__n24522 = new_new_n23380__ | new_new_n23381__;
  assign new_new_n23383__ = ~ys__n24461 & ys__n24463;
  assign new_new_n23384__ = ~ys__n24519 & new_new_n23383__;
  assign ys__n24532 = ys__n24461 | new_new_n23384__;
  assign new_new_n23386__ = ~ys__n1129 & new_new_n23328__;
  assign new_new_n23387__ = new_new_n23360__ & new_new_n23386__;
  assign new_new_n23388__ = new_new_n16583__ & new_new_n23387__;
  assign new_new_n23389__ = ~ys__n4696 & new_new_n23340__;
  assign new_new_n23390__ = ~new_new_n23388__ & ~new_new_n23389__;
  assign ys__n24541 = ~ys__n1094 & ~new_new_n23390__;
  assign ys__n38677 = ys__n24485 & ys__n24567;
  assign new_new_n23393__ = new_new_n23360__ & ys__n38677;
  assign new_new_n23394__ = ~ys__n24483 & new_new_n23348__;
  assign new_new_n23395__ = new_new_n12500__ & new_new_n23331__;
  assign new_new_n23396__ = new_new_n22436__ & new_new_n23328__;
  assign new_new_n23397__ = new_new_n23395__ & new_new_n23396__;
  assign new_new_n23398__ = new_new_n23394__ & new_new_n23397__;
  assign new_new_n23399__ = new_new_n23393__ & new_new_n23398__;
  assign new_new_n23400__ = ys__n1106 & ys__n24567;
  assign new_new_n23401__ = ~ys__n33499 & new_new_n22487__;
  assign new_new_n23402__ = new_new_n23400__ & new_new_n23401__;
  assign new_new_n23403__ = new_new_n16582__ & new_new_n23402__;
  assign new_new_n23404__ = ~new_new_n22467__ & new_new_n23403__;
  assign new_new_n23405__ = ~ys__n4566 & new_new_n23404__;
  assign ys__n24552 = new_new_n23399__ | new_new_n23405__;
  assign new_new_n23407__ = ~ys__n18227 & ys__n24260;
  assign new_new_n23408__ = ys__n18150 & ~ys__n4566;
  assign new_new_n23409__ = ys__n18227 & new_new_n23408__;
  assign ys__n24570 = new_new_n23407__ | new_new_n23409__;
  assign new_new_n23411__ = new_new_n16550__ & ys__n33521;
  assign new_new_n23412__ = ys__n18143 & ~ys__n4566;
  assign new_new_n23413__ = ys__n18227 & new_new_n23412__;
  assign ys__n24573 = new_new_n23411__ | new_new_n23413__;
  assign new_new_n23415__ = ~ys__n14 & ~ys__n4688;
  assign new_new_n23416__ = ys__n30011 & ~new_new_n23415__;
  assign new_new_n23417__ = ys__n30044 & new_new_n23415__;
  assign new_new_n23418__ = ~new_new_n23416__ & ~new_new_n23417__;
  assign new_new_n23419__ = ~ys__n16 & ~ys__n4688;
  assign new_new_n23420__ = ~new_new_n23418__ & ~new_new_n23419__;
  assign new_new_n23421__ = ys__n30028 & ~new_new_n23415__;
  assign new_new_n23422__ = ys__n30060 & new_new_n23415__;
  assign new_new_n23423__ = ~new_new_n23421__ & ~new_new_n23422__;
  assign new_new_n23424__ = new_new_n23419__ & ~new_new_n23423__;
  assign new_new_n23425__ = ~new_new_n23420__ & ~new_new_n23424__;
  assign new_new_n23426__ = ys__n33552 & ys__n38680;
  assign new_new_n23427__ = new_new_n22483__ & new_new_n23426__;
  assign new_new_n23428__ = ~new_new_n23425__ & ~new_new_n23427__;
  assign new_new_n23429__ = ys__n30011 & new_new_n23427__;
  assign new_new_n23430__ = ~new_new_n23428__ & ~new_new_n23429__;
  assign new_new_n23431__ = new_new_n12500__ & ~new_new_n23427__;
  assign new_new_n23432__ = ~new_new_n23430__ & ~new_new_n23431__;
  assign new_new_n23433__ = ys__n24389 & new_new_n23431__;
  assign new_new_n23434__ = ~new_new_n23432__ & ~new_new_n23433__;
  assign new_new_n23435__ = ~ys__n4176 & ~ys__n4696;
  assign new_new_n23436__ = new_new_n10609__ & ~new_new_n23435__;
  assign new_new_n23437__ = ys__n33497 & ys__n1088;
  assign new_new_n23438__ = ~ys__n1117 & ~ys__n1119;
  assign new_new_n23439__ = new_new_n13991__ & new_new_n23438__;
  assign new_new_n23440__ = ~new_new_n23427__ & new_new_n23439__;
  assign new_new_n23441__ = ~new_new_n23437__ & new_new_n23440__;
  assign new_new_n23442__ = ~new_new_n23436__ & ~new_new_n23441__;
  assign new_new_n23443__ = ~new_new_n23434__ & new_new_n23442__;
  assign new_new_n23444__ = ~new_new_n23124__ & ~new_new_n23442__;
  assign new_new_n23445__ = ~new_new_n23443__ & ~new_new_n23444__;
  assign new_new_n23446__ = ys__n1151 & ~ys__n33522;
  assign new_new_n23447__ = new_new_n16563__ & new_new_n23446__;
  assign new_new_n23448__ = ~new_new_n23445__ & ~new_new_n23447__;
  assign new_new_n23449__ = ys__n24575 & new_new_n23447__;
  assign ys__n24577 = new_new_n23448__ | new_new_n23449__;
  assign new_new_n23451__ = ys__n1151 & ys__n18143;
  assign new_new_n23452__ = new_new_n16555__ & new_new_n23451__;
  assign new_new_n23453__ = new_new_n16555__ & new_new_n16558__;
  assign new_new_n23454__ = new_new_n12517__ & ~ys__n18137;
  assign new_new_n23455__ = ~ys__n18227 & ~new_new_n23454__;
  assign new_new_n23456__ = ~new_new_n23453__ & new_new_n23455__;
  assign new_new_n23457__ = ~new_new_n23452__ & new_new_n23456__;
  assign new_new_n23458__ = ys__n24578 & ~new_new_n23457__;
  assign new_new_n23459__ = ys__n20008 & new_new_n23457__;
  assign ys__n24579 = new_new_n23458__ | new_new_n23459__;
  assign new_new_n23461__ = ~ys__n140 & ys__n1151;
  assign ys__n24581 = ~new_new_n16589__ & new_new_n23461__;
  assign new_new_n23463__ = ~ys__n1157 & new_new_n12517__;
  assign ys__n38801 = ys__n24590 & ys__n24591;
  assign new_new_n23465__ = ~ys__n18137 & ys__n38801;
  assign new_new_n23466__ = new_new_n23463__ & new_new_n23465__;
  assign new_new_n23467__ = ys__n1151 & new_new_n16593__;
  assign ys__n24585 = new_new_n23466__ | new_new_n23467__;
  assign new_new_n23469__ = ys__n1154 & ~ys__n18137;
  assign new_new_n23470__ = ~new_new_n16548__ & new_new_n23469__;
  assign new_new_n23471__ = ys__n1151 & ~new_new_n16592__;
  assign new_new_n23472__ = ~new_new_n23470__ & ~new_new_n23471__;
  assign ys__n24604 = ~ys__n140 & ~new_new_n23472__;
  assign ys__n24713 = new_new_n12127__ & ys__n19183;
  assign ys__n24714 = ~new_new_n12127__ & new_new_n16918__;
  assign new_new_n23476__ = ~ys__n44906 & ~ys__n44907;
  assign new_new_n23477__ = ~ys__n44908 & new_new_n23476__;
  assign new_new_n23478__ = ys__n30819 & ys__n31031;
  assign new_new_n23479__ = ~new_new_n23477__ & new_new_n23478__;
  assign new_new_n23480__ = ~ys__n2779 & ~new_new_n23479__;
  assign new_new_n23481__ = ys__n31031 & ys__n47026;
  assign new_new_n23482__ = new_new_n23480__ & new_new_n23481__;
  assign new_new_n23483__ = ys__n34762 & ys__n34764;
  assign new_new_n23484__ = ys__n34766 & new_new_n23483__;
  assign new_new_n23485__ = ~ys__n34762 & ~ys__n34764;
  assign new_new_n23486__ = ys__n34766 & new_new_n23485__;
  assign new_new_n23487__ = ~new_new_n23484__ & ~new_new_n23486__;
  assign new_new_n23488__ = ~ys__n34762 & ys__n34764;
  assign new_new_n23489__ = ~ys__n34766 & new_new_n23488__;
  assign new_new_n23490__ = ys__n34762 & ~ys__n34764;
  assign new_new_n23491__ = ~ys__n34766 & new_new_n23490__;
  assign new_new_n23492__ = ~new_new_n23489__ & ~new_new_n23491__;
  assign new_new_n23493__ = new_new_n23487__ & new_new_n23492__;
  assign new_new_n23494__ = ys__n34770 & ys__n34772;
  assign new_new_n23495__ = ys__n34768 & ys__n34770;
  assign new_new_n23496__ = ys__n34768 & ys__n34772;
  assign new_new_n23497__ = ~new_new_n23495__ & ~new_new_n23496__;
  assign new_new_n23498__ = ~new_new_n23494__ & new_new_n23497__;
  assign new_new_n23499__ = new_new_n23493__ & ~new_new_n23498__;
  assign new_new_n23500__ = ~new_new_n23493__ & new_new_n23498__;
  assign new_new_n23501__ = ~new_new_n23499__ & ~new_new_n23500__;
  assign new_new_n23502__ = ys__n34852 & ys__n34854;
  assign new_new_n23503__ = ys__n34856 & new_new_n23502__;
  assign new_new_n23504__ = ~ys__n34852 & ~ys__n34854;
  assign new_new_n23505__ = ys__n34856 & new_new_n23504__;
  assign new_new_n23506__ = ~new_new_n23503__ & ~new_new_n23505__;
  assign new_new_n23507__ = ~ys__n34852 & ys__n34854;
  assign new_new_n23508__ = ~ys__n34856 & new_new_n23507__;
  assign new_new_n23509__ = ys__n34852 & ~ys__n34854;
  assign new_new_n23510__ = ~ys__n34856 & new_new_n23509__;
  assign new_new_n23511__ = ~new_new_n23508__ & ~new_new_n23510__;
  assign new_new_n23512__ = new_new_n23506__ & new_new_n23511__;
  assign new_new_n23513__ = ys__n34860 & ys__n34862;
  assign new_new_n23514__ = ys__n34858 & ys__n34860;
  assign new_new_n23515__ = ys__n34858 & ys__n34862;
  assign new_new_n23516__ = ~new_new_n23514__ & ~new_new_n23515__;
  assign new_new_n23517__ = ~new_new_n23513__ & new_new_n23516__;
  assign new_new_n23518__ = ~new_new_n23512__ & ~new_new_n23517__;
  assign new_new_n23519__ = new_new_n23512__ & ~new_new_n23517__;
  assign new_new_n23520__ = ~new_new_n23512__ & new_new_n23517__;
  assign new_new_n23521__ = ~new_new_n23519__ & ~new_new_n23520__;
  assign new_new_n23522__ = ys__n34862 & new_new_n23514__;
  assign new_new_n23523__ = ~ys__n34858 & ~ys__n34860;
  assign new_new_n23524__ = ys__n34862 & new_new_n23523__;
  assign new_new_n23525__ = ~new_new_n23522__ & ~new_new_n23524__;
  assign new_new_n23526__ = ~ys__n34858 & ys__n34860;
  assign new_new_n23527__ = ~ys__n34862 & new_new_n23526__;
  assign new_new_n23528__ = ys__n34858 & ~ys__n34860;
  assign new_new_n23529__ = ~ys__n34862 & new_new_n23528__;
  assign new_new_n23530__ = ~new_new_n23527__ & ~new_new_n23529__;
  assign new_new_n23531__ = new_new_n23525__ & new_new_n23530__;
  assign new_new_n23532__ = ys__n34866 & ys__n34868;
  assign new_new_n23533__ = ys__n34864 & ys__n34866;
  assign new_new_n23534__ = ys__n34864 & ys__n34868;
  assign new_new_n23535__ = ~new_new_n23533__ & ~new_new_n23534__;
  assign new_new_n23536__ = ~new_new_n23532__ & new_new_n23535__;
  assign new_new_n23537__ = ~new_new_n23531__ & ~new_new_n23536__;
  assign new_new_n23538__ = ~new_new_n23521__ & new_new_n23537__;
  assign new_new_n23539__ = ~new_new_n23518__ & ~new_new_n23538__;
  assign new_new_n23540__ = ys__n34840 & ys__n34842;
  assign new_new_n23541__ = ys__n34844 & new_new_n23540__;
  assign new_new_n23542__ = ~ys__n34840 & ~ys__n34842;
  assign new_new_n23543__ = ys__n34844 & new_new_n23542__;
  assign new_new_n23544__ = ~new_new_n23541__ & ~new_new_n23543__;
  assign new_new_n23545__ = ~ys__n34840 & ys__n34842;
  assign new_new_n23546__ = ~ys__n34844 & new_new_n23545__;
  assign new_new_n23547__ = ys__n34840 & ~ys__n34842;
  assign new_new_n23548__ = ~ys__n34844 & new_new_n23547__;
  assign new_new_n23549__ = ~new_new_n23546__ & ~new_new_n23548__;
  assign new_new_n23550__ = new_new_n23544__ & new_new_n23549__;
  assign new_new_n23551__ = ys__n34848 & ys__n34850;
  assign new_new_n23552__ = ys__n34846 & ys__n34848;
  assign new_new_n23553__ = ys__n34846 & ys__n34850;
  assign new_new_n23554__ = ~new_new_n23552__ & ~new_new_n23553__;
  assign new_new_n23555__ = ~new_new_n23551__ & new_new_n23554__;
  assign new_new_n23556__ = new_new_n23550__ & ~new_new_n23555__;
  assign new_new_n23557__ = ~new_new_n23550__ & new_new_n23555__;
  assign new_new_n23558__ = ~new_new_n23556__ & ~new_new_n23557__;
  assign new_new_n23559__ = ys__n34850 & new_new_n23552__;
  assign new_new_n23560__ = ~ys__n34846 & ~ys__n34848;
  assign new_new_n23561__ = ys__n34850 & new_new_n23560__;
  assign new_new_n23562__ = ~new_new_n23559__ & ~new_new_n23561__;
  assign new_new_n23563__ = ~ys__n34846 & ys__n34848;
  assign new_new_n23564__ = ~ys__n34850 & new_new_n23563__;
  assign new_new_n23565__ = ys__n34846 & ~ys__n34848;
  assign new_new_n23566__ = ~ys__n34850 & new_new_n23565__;
  assign new_new_n23567__ = ~new_new_n23564__ & ~new_new_n23566__;
  assign new_new_n23568__ = new_new_n23562__ & new_new_n23567__;
  assign new_new_n23569__ = ys__n34854 & ys__n34856;
  assign new_new_n23570__ = ys__n34852 & ys__n34856;
  assign new_new_n23571__ = ~new_new_n23502__ & ~new_new_n23570__;
  assign new_new_n23572__ = ~new_new_n23569__ & new_new_n23571__;
  assign new_new_n23573__ = new_new_n23568__ & ~new_new_n23572__;
  assign new_new_n23574__ = ~new_new_n23568__ & new_new_n23572__;
  assign new_new_n23575__ = ~new_new_n23573__ & ~new_new_n23574__;
  assign new_new_n23576__ = ~new_new_n23558__ & ~new_new_n23575__;
  assign new_new_n23577__ = ~new_new_n23539__ & new_new_n23576__;
  assign new_new_n23578__ = ~new_new_n23550__ & ~new_new_n23555__;
  assign new_new_n23579__ = ~new_new_n23568__ & ~new_new_n23572__;
  assign new_new_n23580__ = ~new_new_n23558__ & new_new_n23579__;
  assign new_new_n23581__ = ~new_new_n23578__ & ~new_new_n23580__;
  assign new_new_n23582__ = ~new_new_n23577__ & new_new_n23581__;
  assign new_new_n23583__ = ys__n34816 & ys__n34818;
  assign new_new_n23584__ = ys__n34820 & new_new_n23583__;
  assign new_new_n23585__ = ~ys__n34816 & ~ys__n34818;
  assign new_new_n23586__ = ys__n34820 & new_new_n23585__;
  assign new_new_n23587__ = ~new_new_n23584__ & ~new_new_n23586__;
  assign new_new_n23588__ = ~ys__n34816 & ys__n34818;
  assign new_new_n23589__ = ~ys__n34820 & new_new_n23588__;
  assign new_new_n23590__ = ys__n34816 & ~ys__n34818;
  assign new_new_n23591__ = ~ys__n34820 & new_new_n23590__;
  assign new_new_n23592__ = ~new_new_n23589__ & ~new_new_n23591__;
  assign new_new_n23593__ = new_new_n23587__ & new_new_n23592__;
  assign new_new_n23594__ = ys__n34824 & ys__n34826;
  assign new_new_n23595__ = ys__n34822 & ys__n34824;
  assign new_new_n23596__ = ys__n34822 & ys__n34826;
  assign new_new_n23597__ = ~new_new_n23595__ & ~new_new_n23596__;
  assign new_new_n23598__ = ~new_new_n23594__ & new_new_n23597__;
  assign new_new_n23599__ = new_new_n23593__ & ~new_new_n23598__;
  assign new_new_n23600__ = ~new_new_n23593__ & new_new_n23598__;
  assign new_new_n23601__ = ~new_new_n23599__ & ~new_new_n23600__;
  assign new_new_n23602__ = ys__n34826 & new_new_n23595__;
  assign new_new_n23603__ = ~ys__n34822 & ~ys__n34824;
  assign new_new_n23604__ = ys__n34826 & new_new_n23603__;
  assign new_new_n23605__ = ~new_new_n23602__ & ~new_new_n23604__;
  assign new_new_n23606__ = ~ys__n34822 & ys__n34824;
  assign new_new_n23607__ = ~ys__n34826 & new_new_n23606__;
  assign new_new_n23608__ = ys__n34822 & ~ys__n34824;
  assign new_new_n23609__ = ~ys__n34826 & new_new_n23608__;
  assign new_new_n23610__ = ~new_new_n23607__ & ~new_new_n23609__;
  assign new_new_n23611__ = new_new_n23605__ & new_new_n23610__;
  assign new_new_n23612__ = ys__n34830 & ys__n34832;
  assign new_new_n23613__ = ys__n34828 & ys__n34830;
  assign new_new_n23614__ = ys__n34828 & ys__n34832;
  assign new_new_n23615__ = ~new_new_n23613__ & ~new_new_n23614__;
  assign new_new_n23616__ = ~new_new_n23612__ & new_new_n23615__;
  assign new_new_n23617__ = new_new_n23611__ & ~new_new_n23616__;
  assign new_new_n23618__ = ~new_new_n23611__ & new_new_n23616__;
  assign new_new_n23619__ = ~new_new_n23617__ & ~new_new_n23618__;
  assign new_new_n23620__ = ~new_new_n23601__ & ~new_new_n23619__;
  assign new_new_n23621__ = ys__n34832 & new_new_n23613__;
  assign new_new_n23622__ = ~ys__n34828 & ~ys__n34830;
  assign new_new_n23623__ = ys__n34832 & new_new_n23622__;
  assign new_new_n23624__ = ~new_new_n23621__ & ~new_new_n23623__;
  assign new_new_n23625__ = ~ys__n34828 & ys__n34830;
  assign new_new_n23626__ = ~ys__n34832 & new_new_n23625__;
  assign new_new_n23627__ = ys__n34828 & ~ys__n34830;
  assign new_new_n23628__ = ~ys__n34832 & new_new_n23627__;
  assign new_new_n23629__ = ~new_new_n23626__ & ~new_new_n23628__;
  assign new_new_n23630__ = new_new_n23624__ & new_new_n23629__;
  assign new_new_n23631__ = ys__n34836 & ys__n34838;
  assign new_new_n23632__ = ys__n34834 & ys__n34836;
  assign new_new_n23633__ = ys__n34834 & ys__n34838;
  assign new_new_n23634__ = ~new_new_n23632__ & ~new_new_n23633__;
  assign new_new_n23635__ = ~new_new_n23631__ & new_new_n23634__;
  assign new_new_n23636__ = new_new_n23630__ & ~new_new_n23635__;
  assign new_new_n23637__ = ~new_new_n23630__ & new_new_n23635__;
  assign new_new_n23638__ = ~new_new_n23636__ & ~new_new_n23637__;
  assign new_new_n23639__ = ys__n34838 & new_new_n23632__;
  assign new_new_n23640__ = ~ys__n34834 & ~ys__n34836;
  assign new_new_n23641__ = ys__n34838 & new_new_n23640__;
  assign new_new_n23642__ = ~new_new_n23639__ & ~new_new_n23641__;
  assign new_new_n23643__ = ~ys__n34834 & ys__n34836;
  assign new_new_n23644__ = ~ys__n34838 & new_new_n23643__;
  assign new_new_n23645__ = ys__n34834 & ~ys__n34836;
  assign new_new_n23646__ = ~ys__n34838 & new_new_n23645__;
  assign new_new_n23647__ = ~new_new_n23644__ & ~new_new_n23646__;
  assign new_new_n23648__ = new_new_n23642__ & new_new_n23647__;
  assign new_new_n23649__ = ys__n34842 & ys__n34844;
  assign new_new_n23650__ = ys__n34840 & ys__n34844;
  assign new_new_n23651__ = ~new_new_n23540__ & ~new_new_n23650__;
  assign new_new_n23652__ = ~new_new_n23649__ & new_new_n23651__;
  assign new_new_n23653__ = new_new_n23648__ & ~new_new_n23652__;
  assign new_new_n23654__ = ~new_new_n23648__ & new_new_n23652__;
  assign new_new_n23655__ = ~new_new_n23653__ & ~new_new_n23654__;
  assign new_new_n23656__ = ~new_new_n23638__ & ~new_new_n23655__;
  assign new_new_n23657__ = new_new_n23620__ & new_new_n23656__;
  assign new_new_n23658__ = ~new_new_n23582__ & new_new_n23657__;
  assign new_new_n23659__ = ~new_new_n23630__ & ~new_new_n23635__;
  assign new_new_n23660__ = ~new_new_n23648__ & ~new_new_n23652__;
  assign new_new_n23661__ = ~new_new_n23638__ & new_new_n23660__;
  assign new_new_n23662__ = ~new_new_n23659__ & ~new_new_n23661__;
  assign new_new_n23663__ = new_new_n23620__ & ~new_new_n23662__;
  assign new_new_n23664__ = ~new_new_n23593__ & ~new_new_n23598__;
  assign new_new_n23665__ = ~new_new_n23611__ & ~new_new_n23616__;
  assign new_new_n23666__ = ~new_new_n23601__ & new_new_n23665__;
  assign new_new_n23667__ = ~new_new_n23664__ & ~new_new_n23666__;
  assign new_new_n23668__ = ~new_new_n23663__ & new_new_n23667__;
  assign new_new_n23669__ = ~new_new_n23658__ & new_new_n23668__;
  assign new_new_n23670__ = ys__n34772 & new_new_n23495__;
  assign new_new_n23671__ = ~ys__n34768 & ~ys__n34770;
  assign new_new_n23672__ = ys__n34772 & new_new_n23671__;
  assign new_new_n23673__ = ~new_new_n23670__ & ~new_new_n23672__;
  assign new_new_n23674__ = ~ys__n34768 & ys__n34770;
  assign new_new_n23675__ = ~ys__n34772 & new_new_n23674__;
  assign new_new_n23676__ = ys__n34768 & ~ys__n34770;
  assign new_new_n23677__ = ~ys__n34772 & new_new_n23676__;
  assign new_new_n23678__ = ~new_new_n23675__ & ~new_new_n23677__;
  assign new_new_n23679__ = new_new_n23673__ & new_new_n23678__;
  assign new_new_n23680__ = ys__n34776 & ys__n34778;
  assign new_new_n23681__ = ys__n34774 & ys__n34776;
  assign new_new_n23682__ = ys__n34774 & ys__n34778;
  assign new_new_n23683__ = ~new_new_n23681__ & ~new_new_n23682__;
  assign new_new_n23684__ = ~new_new_n23680__ & new_new_n23683__;
  assign new_new_n23685__ = new_new_n23679__ & ~new_new_n23684__;
  assign new_new_n23686__ = ~new_new_n23679__ & new_new_n23684__;
  assign new_new_n23687__ = ~new_new_n23685__ & ~new_new_n23686__;
  assign new_new_n23688__ = ys__n34778 & new_new_n23681__;
  assign new_new_n23689__ = ~ys__n34774 & ~ys__n34776;
  assign new_new_n23690__ = ys__n34778 & new_new_n23689__;
  assign new_new_n23691__ = ~new_new_n23688__ & ~new_new_n23690__;
  assign new_new_n23692__ = ~ys__n34774 & ys__n34776;
  assign new_new_n23693__ = ~ys__n34778 & new_new_n23692__;
  assign new_new_n23694__ = ys__n34774 & ~ys__n34776;
  assign new_new_n23695__ = ~ys__n34778 & new_new_n23694__;
  assign new_new_n23696__ = ~new_new_n23693__ & ~new_new_n23695__;
  assign new_new_n23697__ = new_new_n23691__ & new_new_n23696__;
  assign new_new_n23698__ = ys__n34782 & ys__n34784;
  assign new_new_n23699__ = ys__n34780 & ys__n34782;
  assign new_new_n23700__ = ys__n34780 & ys__n34784;
  assign new_new_n23701__ = ~new_new_n23699__ & ~new_new_n23700__;
  assign new_new_n23702__ = ~new_new_n23698__ & new_new_n23701__;
  assign new_new_n23703__ = new_new_n23697__ & ~new_new_n23702__;
  assign new_new_n23704__ = ~new_new_n23697__ & new_new_n23702__;
  assign new_new_n23705__ = ~new_new_n23703__ & ~new_new_n23704__;
  assign new_new_n23706__ = ~new_new_n23687__ & ~new_new_n23705__;
  assign new_new_n23707__ = ys__n34784 & new_new_n23699__;
  assign new_new_n23708__ = ~ys__n34780 & ~ys__n34782;
  assign new_new_n23709__ = ys__n34784 & new_new_n23708__;
  assign new_new_n23710__ = ~new_new_n23707__ & ~new_new_n23709__;
  assign new_new_n23711__ = ~ys__n34780 & ys__n34782;
  assign new_new_n23712__ = ~ys__n34784 & new_new_n23711__;
  assign new_new_n23713__ = ys__n34780 & ~ys__n34782;
  assign new_new_n23714__ = ~ys__n34784 & new_new_n23713__;
  assign new_new_n23715__ = ~new_new_n23712__ & ~new_new_n23714__;
  assign new_new_n23716__ = new_new_n23710__ & new_new_n23715__;
  assign new_new_n23717__ = ys__n34788 & ys__n34790;
  assign new_new_n23718__ = ys__n34786 & ys__n34788;
  assign new_new_n23719__ = ys__n34786 & ys__n34790;
  assign new_new_n23720__ = ~new_new_n23718__ & ~new_new_n23719__;
  assign new_new_n23721__ = ~new_new_n23717__ & new_new_n23720__;
  assign new_new_n23722__ = new_new_n23716__ & ~new_new_n23721__;
  assign new_new_n23723__ = ~new_new_n23716__ & new_new_n23721__;
  assign new_new_n23724__ = ~new_new_n23722__ & ~new_new_n23723__;
  assign new_new_n23725__ = ys__n34790 & new_new_n23718__;
  assign new_new_n23726__ = ~ys__n34786 & ~ys__n34788;
  assign new_new_n23727__ = ys__n34790 & new_new_n23726__;
  assign new_new_n23728__ = ~new_new_n23725__ & ~new_new_n23727__;
  assign new_new_n23729__ = ~ys__n34786 & ys__n34788;
  assign new_new_n23730__ = ~ys__n34790 & new_new_n23729__;
  assign new_new_n23731__ = ys__n34786 & ~ys__n34788;
  assign new_new_n23732__ = ~ys__n34790 & new_new_n23731__;
  assign new_new_n23733__ = ~new_new_n23730__ & ~new_new_n23732__;
  assign new_new_n23734__ = new_new_n23728__ & new_new_n23733__;
  assign new_new_n23735__ = ys__n34794 & ys__n34796;
  assign new_new_n23736__ = ys__n34792 & ys__n34794;
  assign new_new_n23737__ = ys__n34792 & ys__n34796;
  assign new_new_n23738__ = ~new_new_n23736__ & ~new_new_n23737__;
  assign new_new_n23739__ = ~new_new_n23735__ & new_new_n23738__;
  assign new_new_n23740__ = new_new_n23734__ & ~new_new_n23739__;
  assign new_new_n23741__ = ~new_new_n23734__ & new_new_n23739__;
  assign new_new_n23742__ = ~new_new_n23740__ & ~new_new_n23741__;
  assign new_new_n23743__ = ~new_new_n23724__ & ~new_new_n23742__;
  assign new_new_n23744__ = new_new_n23706__ & new_new_n23743__;
  assign new_new_n23745__ = ys__n34796 & new_new_n23736__;
  assign new_new_n23746__ = ~ys__n34792 & ~ys__n34794;
  assign new_new_n23747__ = ys__n34796 & new_new_n23746__;
  assign new_new_n23748__ = ~new_new_n23745__ & ~new_new_n23747__;
  assign new_new_n23749__ = ~ys__n34792 & ys__n34794;
  assign new_new_n23750__ = ~ys__n34796 & new_new_n23749__;
  assign new_new_n23751__ = ys__n34792 & ~ys__n34794;
  assign new_new_n23752__ = ~ys__n34796 & new_new_n23751__;
  assign new_new_n23753__ = ~new_new_n23750__ & ~new_new_n23752__;
  assign new_new_n23754__ = new_new_n23748__ & new_new_n23753__;
  assign new_new_n23755__ = ys__n34800 & ys__n34802;
  assign new_new_n23756__ = ys__n34798 & ys__n34800;
  assign new_new_n23757__ = ys__n34798 & ys__n34802;
  assign new_new_n23758__ = ~new_new_n23756__ & ~new_new_n23757__;
  assign new_new_n23759__ = ~new_new_n23755__ & new_new_n23758__;
  assign new_new_n23760__ = new_new_n23754__ & ~new_new_n23759__;
  assign new_new_n23761__ = ~new_new_n23754__ & new_new_n23759__;
  assign new_new_n23762__ = ~new_new_n23760__ & ~new_new_n23761__;
  assign new_new_n23763__ = ys__n34802 & new_new_n23756__;
  assign new_new_n23764__ = ~ys__n34798 & ~ys__n34800;
  assign new_new_n23765__ = ys__n34802 & new_new_n23764__;
  assign new_new_n23766__ = ~new_new_n23763__ & ~new_new_n23765__;
  assign new_new_n23767__ = ~ys__n34798 & ys__n34800;
  assign new_new_n23768__ = ~ys__n34802 & new_new_n23767__;
  assign new_new_n23769__ = ys__n34798 & ~ys__n34800;
  assign new_new_n23770__ = ~ys__n34802 & new_new_n23769__;
  assign new_new_n23771__ = ~new_new_n23768__ & ~new_new_n23770__;
  assign new_new_n23772__ = new_new_n23766__ & new_new_n23771__;
  assign new_new_n23773__ = ys__n34806 & ys__n34808;
  assign new_new_n23774__ = ys__n34804 & ys__n34806;
  assign new_new_n23775__ = ys__n34804 & ys__n34808;
  assign new_new_n23776__ = ~new_new_n23774__ & ~new_new_n23775__;
  assign new_new_n23777__ = ~new_new_n23773__ & new_new_n23776__;
  assign new_new_n23778__ = new_new_n23772__ & ~new_new_n23777__;
  assign new_new_n23779__ = ~new_new_n23772__ & new_new_n23777__;
  assign new_new_n23780__ = ~new_new_n23778__ & ~new_new_n23779__;
  assign new_new_n23781__ = ~new_new_n23762__ & ~new_new_n23780__;
  assign new_new_n23782__ = ys__n34808 & new_new_n23774__;
  assign new_new_n23783__ = ~ys__n34804 & ~ys__n34806;
  assign new_new_n23784__ = ys__n34808 & new_new_n23783__;
  assign new_new_n23785__ = ~new_new_n23782__ & ~new_new_n23784__;
  assign new_new_n23786__ = ~ys__n34804 & ys__n34806;
  assign new_new_n23787__ = ~ys__n34808 & new_new_n23786__;
  assign new_new_n23788__ = ys__n34804 & ~ys__n34806;
  assign new_new_n23789__ = ~ys__n34808 & new_new_n23788__;
  assign new_new_n23790__ = ~new_new_n23787__ & ~new_new_n23789__;
  assign new_new_n23791__ = new_new_n23785__ & new_new_n23790__;
  assign new_new_n23792__ = ys__n34812 & ys__n34814;
  assign new_new_n23793__ = ys__n34810 & ys__n34812;
  assign new_new_n23794__ = ys__n34810 & ys__n34814;
  assign new_new_n23795__ = ~new_new_n23793__ & ~new_new_n23794__;
  assign new_new_n23796__ = ~new_new_n23792__ & new_new_n23795__;
  assign new_new_n23797__ = new_new_n23791__ & ~new_new_n23796__;
  assign new_new_n23798__ = ~new_new_n23791__ & new_new_n23796__;
  assign new_new_n23799__ = ~new_new_n23797__ & ~new_new_n23798__;
  assign new_new_n23800__ = ys__n34814 & new_new_n23793__;
  assign new_new_n23801__ = ~ys__n34810 & ~ys__n34812;
  assign new_new_n23802__ = ys__n34814 & new_new_n23801__;
  assign new_new_n23803__ = ~new_new_n23800__ & ~new_new_n23802__;
  assign new_new_n23804__ = ~ys__n34810 & ys__n34812;
  assign new_new_n23805__ = ~ys__n34814 & new_new_n23804__;
  assign new_new_n23806__ = ys__n34810 & ~ys__n34812;
  assign new_new_n23807__ = ~ys__n34814 & new_new_n23806__;
  assign new_new_n23808__ = ~new_new_n23805__ & ~new_new_n23807__;
  assign new_new_n23809__ = new_new_n23803__ & new_new_n23808__;
  assign new_new_n23810__ = ys__n34818 & ys__n34820;
  assign new_new_n23811__ = ys__n34816 & ys__n34820;
  assign new_new_n23812__ = ~new_new_n23583__ & ~new_new_n23811__;
  assign new_new_n23813__ = ~new_new_n23810__ & new_new_n23812__;
  assign new_new_n23814__ = new_new_n23809__ & ~new_new_n23813__;
  assign new_new_n23815__ = ~new_new_n23809__ & new_new_n23813__;
  assign new_new_n23816__ = ~new_new_n23814__ & ~new_new_n23815__;
  assign new_new_n23817__ = ~new_new_n23799__ & ~new_new_n23816__;
  assign new_new_n23818__ = new_new_n23781__ & new_new_n23817__;
  assign new_new_n23819__ = new_new_n23744__ & new_new_n23818__;
  assign new_new_n23820__ = ~new_new_n23669__ & new_new_n23819__;
  assign new_new_n23821__ = ~new_new_n23791__ & ~new_new_n23796__;
  assign new_new_n23822__ = ~new_new_n23809__ & ~new_new_n23813__;
  assign new_new_n23823__ = ~new_new_n23799__ & new_new_n23822__;
  assign new_new_n23824__ = ~new_new_n23821__ & ~new_new_n23823__;
  assign new_new_n23825__ = new_new_n23781__ & ~new_new_n23824__;
  assign new_new_n23826__ = ~new_new_n23754__ & ~new_new_n23759__;
  assign new_new_n23827__ = ~new_new_n23772__ & ~new_new_n23777__;
  assign new_new_n23828__ = ~new_new_n23762__ & new_new_n23827__;
  assign new_new_n23829__ = ~new_new_n23826__ & ~new_new_n23828__;
  assign new_new_n23830__ = ~new_new_n23825__ & new_new_n23829__;
  assign new_new_n23831__ = new_new_n23744__ & ~new_new_n23830__;
  assign new_new_n23832__ = ~new_new_n23716__ & ~new_new_n23721__;
  assign new_new_n23833__ = ~new_new_n23734__ & ~new_new_n23739__;
  assign new_new_n23834__ = ~new_new_n23724__ & new_new_n23833__;
  assign new_new_n23835__ = ~new_new_n23832__ & ~new_new_n23834__;
  assign new_new_n23836__ = new_new_n23706__ & ~new_new_n23835__;
  assign new_new_n23837__ = ~new_new_n23679__ & ~new_new_n23684__;
  assign new_new_n23838__ = ~new_new_n23697__ & ~new_new_n23702__;
  assign new_new_n23839__ = ~new_new_n23687__ & new_new_n23838__;
  assign new_new_n23840__ = ~new_new_n23837__ & ~new_new_n23839__;
  assign new_new_n23841__ = ~new_new_n23836__ & new_new_n23840__;
  assign new_new_n23842__ = ~new_new_n23831__ & new_new_n23841__;
  assign new_new_n23843__ = ~new_new_n23820__ & new_new_n23842__;
  assign new_new_n23844__ = ys__n34938 & ys__n34940;
  assign new_new_n23845__ = ys__n34942 & new_new_n23844__;
  assign new_new_n23846__ = ~ys__n34938 & ~ys__n34940;
  assign new_new_n23847__ = ys__n34942 & new_new_n23846__;
  assign new_new_n23848__ = ~new_new_n23845__ & ~new_new_n23847__;
  assign new_new_n23849__ = ~ys__n34938 & ys__n34940;
  assign new_new_n23850__ = ~ys__n34942 & new_new_n23849__;
  assign new_new_n23851__ = ys__n34938 & ~ys__n34940;
  assign new_new_n23852__ = ~ys__n34942 & new_new_n23851__;
  assign new_new_n23853__ = ~new_new_n23850__ & ~new_new_n23852__;
  assign new_new_n23854__ = new_new_n23848__ & new_new_n23853__;
  assign new_new_n23855__ = ys__n34944 & ys__n34946;
  assign new_new_n23856__ = new_new_n23854__ & new_new_n23855__;
  assign new_new_n23857__ = ~new_new_n23854__ & ~new_new_n23855__;
  assign new_new_n23858__ = ~new_new_n23856__ & ~new_new_n23857__;
  assign new_new_n23859__ = ~ys__n34934 & ys__n34936;
  assign new_new_n23860__ = ys__n34934 & ~ys__n34936;
  assign new_new_n23861__ = ~new_new_n23859__ & ~new_new_n23860__;
  assign new_new_n23862__ = ys__n34940 & ys__n34942;
  assign new_new_n23863__ = ys__n34938 & ys__n34942;
  assign new_new_n23864__ = ~new_new_n23844__ & ~new_new_n23863__;
  assign new_new_n23865__ = ~new_new_n23862__ & new_new_n23864__;
  assign new_new_n23866__ = new_new_n23861__ & ~new_new_n23865__;
  assign new_new_n23867__ = ~new_new_n23861__ & new_new_n23865__;
  assign new_new_n23868__ = ~new_new_n23866__ & ~new_new_n23867__;
  assign new_new_n23869__ = ~ys__n34944 & ys__n34946;
  assign new_new_n23870__ = ys__n34944 & ~ys__n34946;
  assign new_new_n23871__ = ~new_new_n23869__ & ~new_new_n23870__;
  assign new_new_n23872__ = ys__n34948 & ys__n34950;
  assign new_new_n23873__ = ~new_new_n23871__ & new_new_n23872__;
  assign new_new_n23874__ = ~new_new_n23868__ & new_new_n23873__;
  assign new_new_n23875__ = ~new_new_n23858__ & new_new_n23874__;
  assign new_new_n23876__ = ~new_new_n23861__ & ~new_new_n23865__;
  assign new_new_n23877__ = ~new_new_n23854__ & new_new_n23855__;
  assign new_new_n23878__ = ~new_new_n23868__ & new_new_n23877__;
  assign new_new_n23879__ = ~new_new_n23876__ & ~new_new_n23878__;
  assign new_new_n23880__ = ~new_new_n23875__ & new_new_n23879__;
  assign new_new_n23881__ = ys__n34912 & ys__n34914;
  assign new_new_n23882__ = ys__n34916 & new_new_n23881__;
  assign new_new_n23883__ = ~ys__n34912 & ~ys__n34914;
  assign new_new_n23884__ = ys__n34916 & new_new_n23883__;
  assign new_new_n23885__ = ~new_new_n23882__ & ~new_new_n23884__;
  assign new_new_n23886__ = ~ys__n34912 & ys__n34914;
  assign new_new_n23887__ = ~ys__n34916 & new_new_n23886__;
  assign new_new_n23888__ = ys__n34912 & ~ys__n34914;
  assign new_new_n23889__ = ~ys__n34916 & new_new_n23888__;
  assign new_new_n23890__ = ~new_new_n23887__ & ~new_new_n23889__;
  assign new_new_n23891__ = new_new_n23885__ & new_new_n23890__;
  assign new_new_n23892__ = ys__n34920 & ys__n34922;
  assign new_new_n23893__ = ys__n34918 & ys__n34920;
  assign new_new_n23894__ = ys__n34918 & ys__n34922;
  assign new_new_n23895__ = ~new_new_n23893__ & ~new_new_n23894__;
  assign new_new_n23896__ = ~new_new_n23892__ & new_new_n23895__;
  assign new_new_n23897__ = new_new_n23891__ & ~new_new_n23896__;
  assign new_new_n23898__ = ~new_new_n23891__ & new_new_n23896__;
  assign new_new_n23899__ = ~new_new_n23897__ & ~new_new_n23898__;
  assign new_new_n23900__ = ys__n34922 & new_new_n23893__;
  assign new_new_n23901__ = ~ys__n34918 & ~ys__n34920;
  assign new_new_n23902__ = ys__n34922 & new_new_n23901__;
  assign new_new_n23903__ = ~new_new_n23900__ & ~new_new_n23902__;
  assign new_new_n23904__ = ~ys__n34918 & ys__n34920;
  assign new_new_n23905__ = ~ys__n34922 & new_new_n23904__;
  assign new_new_n23906__ = ys__n34918 & ~ys__n34920;
  assign new_new_n23907__ = ~ys__n34922 & new_new_n23906__;
  assign new_new_n23908__ = ~new_new_n23905__ & ~new_new_n23907__;
  assign new_new_n23909__ = new_new_n23903__ & new_new_n23908__;
  assign new_new_n23910__ = ys__n34926 & ys__n34928;
  assign new_new_n23911__ = ys__n34924 & ys__n34926;
  assign new_new_n23912__ = ys__n34924 & ys__n34928;
  assign new_new_n23913__ = ~new_new_n23911__ & ~new_new_n23912__;
  assign new_new_n23914__ = ~new_new_n23910__ & new_new_n23913__;
  assign new_new_n23915__ = new_new_n23909__ & ~new_new_n23914__;
  assign new_new_n23916__ = ~new_new_n23909__ & new_new_n23914__;
  assign new_new_n23917__ = ~new_new_n23915__ & ~new_new_n23916__;
  assign new_new_n23918__ = ~new_new_n23899__ & ~new_new_n23917__;
  assign new_new_n23919__ = ys__n34928 & new_new_n23911__;
  assign new_new_n23920__ = ~ys__n34924 & ~ys__n34926;
  assign new_new_n23921__ = ys__n34928 & new_new_n23920__;
  assign new_new_n23922__ = ~new_new_n23919__ & ~new_new_n23921__;
  assign new_new_n23923__ = ~ys__n34924 & ys__n34926;
  assign new_new_n23924__ = ~ys__n34928 & new_new_n23923__;
  assign new_new_n23925__ = ys__n34924 & ~ys__n34926;
  assign new_new_n23926__ = ~ys__n34928 & new_new_n23925__;
  assign new_new_n23927__ = ~new_new_n23924__ & ~new_new_n23926__;
  assign new_new_n23928__ = new_new_n23922__ & new_new_n23927__;
  assign new_new_n23929__ = ys__n34930 & ys__n34932;
  assign new_new_n23930__ = new_new_n23928__ & new_new_n23929__;
  assign new_new_n23931__ = ~new_new_n23928__ & ~new_new_n23929__;
  assign new_new_n23932__ = ~new_new_n23930__ & ~new_new_n23931__;
  assign new_new_n23933__ = ~ys__n34930 & ys__n34932;
  assign new_new_n23934__ = ys__n34930 & ~ys__n34932;
  assign new_new_n23935__ = ~new_new_n23933__ & ~new_new_n23934__;
  assign new_new_n23936__ = ys__n34934 & ys__n34936;
  assign new_new_n23937__ = new_new_n23935__ & new_new_n23936__;
  assign new_new_n23938__ = ~new_new_n23935__ & ~new_new_n23936__;
  assign new_new_n23939__ = ~new_new_n23937__ & ~new_new_n23938__;
  assign new_new_n23940__ = ~new_new_n23932__ & ~new_new_n23939__;
  assign new_new_n23941__ = new_new_n23918__ & new_new_n23940__;
  assign new_new_n23942__ = ~new_new_n23880__ & new_new_n23941__;
  assign new_new_n23943__ = ~new_new_n23928__ & new_new_n23929__;
  assign new_new_n23944__ = ~new_new_n23935__ & new_new_n23936__;
  assign new_new_n23945__ = ~new_new_n23932__ & new_new_n23944__;
  assign new_new_n23946__ = ~new_new_n23943__ & ~new_new_n23945__;
  assign new_new_n23947__ = new_new_n23918__ & ~new_new_n23946__;
  assign new_new_n23948__ = ~new_new_n23891__ & ~new_new_n23896__;
  assign new_new_n23949__ = ~new_new_n23909__ & ~new_new_n23914__;
  assign new_new_n23950__ = ~new_new_n23899__ & new_new_n23949__;
  assign new_new_n23951__ = ~new_new_n23948__ & ~new_new_n23950__;
  assign new_new_n23952__ = ~new_new_n23947__ & new_new_n23951__;
  assign new_new_n23953__ = ~new_new_n23942__ & new_new_n23952__;
  assign new_new_n23954__ = ys__n34868 & new_new_n23533__;
  assign new_new_n23955__ = ~ys__n34864 & ~ys__n34866;
  assign new_new_n23956__ = ys__n34868 & new_new_n23955__;
  assign new_new_n23957__ = ~new_new_n23954__ & ~new_new_n23956__;
  assign new_new_n23958__ = ~ys__n34864 & ys__n34866;
  assign new_new_n23959__ = ~ys__n34868 & new_new_n23958__;
  assign new_new_n23960__ = ys__n34864 & ~ys__n34866;
  assign new_new_n23961__ = ~ys__n34868 & new_new_n23960__;
  assign new_new_n23962__ = ~new_new_n23959__ & ~new_new_n23961__;
  assign new_new_n23963__ = new_new_n23957__ & new_new_n23962__;
  assign new_new_n23964__ = ys__n34872 & ys__n34874;
  assign new_new_n23965__ = ys__n34870 & ys__n34872;
  assign new_new_n23966__ = ys__n34870 & ys__n34874;
  assign new_new_n23967__ = ~new_new_n23965__ & ~new_new_n23966__;
  assign new_new_n23968__ = ~new_new_n23964__ & new_new_n23967__;
  assign new_new_n23969__ = new_new_n23963__ & ~new_new_n23968__;
  assign new_new_n23970__ = ~new_new_n23963__ & new_new_n23968__;
  assign new_new_n23971__ = ~new_new_n23969__ & ~new_new_n23970__;
  assign new_new_n23972__ = ys__n34874 & new_new_n23965__;
  assign new_new_n23973__ = ~ys__n34870 & ~ys__n34872;
  assign new_new_n23974__ = ys__n34874 & new_new_n23973__;
  assign new_new_n23975__ = ~new_new_n23972__ & ~new_new_n23974__;
  assign new_new_n23976__ = ~ys__n34870 & ys__n34872;
  assign new_new_n23977__ = ~ys__n34874 & new_new_n23976__;
  assign new_new_n23978__ = ys__n34870 & ~ys__n34872;
  assign new_new_n23979__ = ~ys__n34874 & new_new_n23978__;
  assign new_new_n23980__ = ~new_new_n23977__ & ~new_new_n23979__;
  assign new_new_n23981__ = new_new_n23975__ & new_new_n23980__;
  assign new_new_n23982__ = ys__n34878 & ys__n34880;
  assign new_new_n23983__ = ys__n34876 & ys__n34878;
  assign new_new_n23984__ = ys__n34876 & ys__n34880;
  assign new_new_n23985__ = ~new_new_n23983__ & ~new_new_n23984__;
  assign new_new_n23986__ = ~new_new_n23982__ & new_new_n23985__;
  assign new_new_n23987__ = new_new_n23981__ & ~new_new_n23986__;
  assign new_new_n23988__ = ~new_new_n23981__ & new_new_n23986__;
  assign new_new_n23989__ = ~new_new_n23987__ & ~new_new_n23988__;
  assign new_new_n23990__ = ~new_new_n23971__ & ~new_new_n23989__;
  assign new_new_n23991__ = ys__n34880 & new_new_n23983__;
  assign new_new_n23992__ = ~ys__n34876 & ~ys__n34878;
  assign new_new_n23993__ = ys__n34880 & new_new_n23992__;
  assign new_new_n23994__ = ~new_new_n23991__ & ~new_new_n23993__;
  assign new_new_n23995__ = ~ys__n34876 & ys__n34878;
  assign new_new_n23996__ = ~ys__n34880 & new_new_n23995__;
  assign new_new_n23997__ = ys__n34876 & ~ys__n34878;
  assign new_new_n23998__ = ~ys__n34880 & new_new_n23997__;
  assign new_new_n23999__ = ~new_new_n23996__ & ~new_new_n23998__;
  assign new_new_n24000__ = new_new_n23994__ & new_new_n23999__;
  assign new_new_n24001__ = ys__n34884 & ys__n34886;
  assign new_new_n24002__ = ys__n34882 & ys__n34884;
  assign new_new_n24003__ = ys__n34882 & ys__n34886;
  assign new_new_n24004__ = ~new_new_n24002__ & ~new_new_n24003__;
  assign new_new_n24005__ = ~new_new_n24001__ & new_new_n24004__;
  assign new_new_n24006__ = new_new_n24000__ & ~new_new_n24005__;
  assign new_new_n24007__ = ~new_new_n24000__ & new_new_n24005__;
  assign new_new_n24008__ = ~new_new_n24006__ & ~new_new_n24007__;
  assign new_new_n24009__ = ys__n34886 & new_new_n24002__;
  assign new_new_n24010__ = ~ys__n34882 & ~ys__n34884;
  assign new_new_n24011__ = ys__n34886 & new_new_n24010__;
  assign new_new_n24012__ = ~new_new_n24009__ & ~new_new_n24011__;
  assign new_new_n24013__ = ~ys__n34882 & ys__n34884;
  assign new_new_n24014__ = ~ys__n34886 & new_new_n24013__;
  assign new_new_n24015__ = ys__n34882 & ~ys__n34884;
  assign new_new_n24016__ = ~ys__n34886 & new_new_n24015__;
  assign new_new_n24017__ = ~new_new_n24014__ & ~new_new_n24016__;
  assign new_new_n24018__ = new_new_n24012__ & new_new_n24017__;
  assign new_new_n24019__ = ys__n34890 & ys__n34892;
  assign new_new_n24020__ = ys__n34888 & ys__n34890;
  assign new_new_n24021__ = ys__n34888 & ys__n34892;
  assign new_new_n24022__ = ~new_new_n24020__ & ~new_new_n24021__;
  assign new_new_n24023__ = ~new_new_n24019__ & new_new_n24022__;
  assign new_new_n24024__ = new_new_n24018__ & ~new_new_n24023__;
  assign new_new_n24025__ = ~new_new_n24018__ & new_new_n24023__;
  assign new_new_n24026__ = ~new_new_n24024__ & ~new_new_n24025__;
  assign new_new_n24027__ = ~new_new_n24008__ & ~new_new_n24026__;
  assign new_new_n24028__ = new_new_n23990__ & new_new_n24027__;
  assign new_new_n24029__ = ys__n34892 & new_new_n24020__;
  assign new_new_n24030__ = ~ys__n34888 & ~ys__n34890;
  assign new_new_n24031__ = ys__n34892 & new_new_n24030__;
  assign new_new_n24032__ = ~new_new_n24029__ & ~new_new_n24031__;
  assign new_new_n24033__ = ~ys__n34888 & ys__n34890;
  assign new_new_n24034__ = ~ys__n34892 & new_new_n24033__;
  assign new_new_n24035__ = ys__n34888 & ~ys__n34890;
  assign new_new_n24036__ = ~ys__n34892 & new_new_n24035__;
  assign new_new_n24037__ = ~new_new_n24034__ & ~new_new_n24036__;
  assign new_new_n24038__ = new_new_n24032__ & new_new_n24037__;
  assign new_new_n24039__ = ys__n34896 & ys__n34898;
  assign new_new_n24040__ = ys__n34894 & ys__n34896;
  assign new_new_n24041__ = ys__n34894 & ys__n34898;
  assign new_new_n24042__ = ~new_new_n24040__ & ~new_new_n24041__;
  assign new_new_n24043__ = ~new_new_n24039__ & new_new_n24042__;
  assign new_new_n24044__ = new_new_n24038__ & ~new_new_n24043__;
  assign new_new_n24045__ = ~new_new_n24038__ & new_new_n24043__;
  assign new_new_n24046__ = ~new_new_n24044__ & ~new_new_n24045__;
  assign new_new_n24047__ = ys__n34898 & new_new_n24040__;
  assign new_new_n24048__ = ~ys__n34894 & ~ys__n34896;
  assign new_new_n24049__ = ys__n34898 & new_new_n24048__;
  assign new_new_n24050__ = ~new_new_n24047__ & ~new_new_n24049__;
  assign new_new_n24051__ = ~ys__n34894 & ys__n34896;
  assign new_new_n24052__ = ~ys__n34898 & new_new_n24051__;
  assign new_new_n24053__ = ys__n34894 & ~ys__n34896;
  assign new_new_n24054__ = ~ys__n34898 & new_new_n24053__;
  assign new_new_n24055__ = ~new_new_n24052__ & ~new_new_n24054__;
  assign new_new_n24056__ = new_new_n24050__ & new_new_n24055__;
  assign new_new_n24057__ = ys__n34902 & ys__n34904;
  assign new_new_n24058__ = ys__n34900 & ys__n34902;
  assign new_new_n24059__ = ys__n34900 & ys__n34904;
  assign new_new_n24060__ = ~new_new_n24058__ & ~new_new_n24059__;
  assign new_new_n24061__ = ~new_new_n24057__ & new_new_n24060__;
  assign new_new_n24062__ = new_new_n24056__ & ~new_new_n24061__;
  assign new_new_n24063__ = ~new_new_n24056__ & new_new_n24061__;
  assign new_new_n24064__ = ~new_new_n24062__ & ~new_new_n24063__;
  assign new_new_n24065__ = ~new_new_n24046__ & ~new_new_n24064__;
  assign new_new_n24066__ = ys__n34904 & new_new_n24058__;
  assign new_new_n24067__ = ~ys__n34900 & ~ys__n34902;
  assign new_new_n24068__ = ys__n34904 & new_new_n24067__;
  assign new_new_n24069__ = ~new_new_n24066__ & ~new_new_n24068__;
  assign new_new_n24070__ = ~ys__n34900 & ys__n34902;
  assign new_new_n24071__ = ~ys__n34904 & new_new_n24070__;
  assign new_new_n24072__ = ys__n34900 & ~ys__n34902;
  assign new_new_n24073__ = ~ys__n34904 & new_new_n24072__;
  assign new_new_n24074__ = ~new_new_n24071__ & ~new_new_n24073__;
  assign new_new_n24075__ = new_new_n24069__ & new_new_n24074__;
  assign new_new_n24076__ = ys__n34908 & ys__n34910;
  assign new_new_n24077__ = ys__n34906 & ys__n34908;
  assign new_new_n24078__ = ys__n34906 & ys__n34910;
  assign new_new_n24079__ = ~new_new_n24077__ & ~new_new_n24078__;
  assign new_new_n24080__ = ~new_new_n24076__ & new_new_n24079__;
  assign new_new_n24081__ = new_new_n24075__ & ~new_new_n24080__;
  assign new_new_n24082__ = ~new_new_n24075__ & new_new_n24080__;
  assign new_new_n24083__ = ~new_new_n24081__ & ~new_new_n24082__;
  assign new_new_n24084__ = ys__n34910 & new_new_n24077__;
  assign new_new_n24085__ = ~ys__n34906 & ~ys__n34908;
  assign new_new_n24086__ = ys__n34910 & new_new_n24085__;
  assign new_new_n24087__ = ~new_new_n24084__ & ~new_new_n24086__;
  assign new_new_n24088__ = ~ys__n34906 & ys__n34908;
  assign new_new_n24089__ = ~ys__n34910 & new_new_n24088__;
  assign new_new_n24090__ = ys__n34906 & ~ys__n34908;
  assign new_new_n24091__ = ~ys__n34910 & new_new_n24090__;
  assign new_new_n24092__ = ~new_new_n24089__ & ~new_new_n24091__;
  assign new_new_n24093__ = new_new_n24087__ & new_new_n24092__;
  assign new_new_n24094__ = ys__n34914 & ys__n34916;
  assign new_new_n24095__ = ys__n34912 & ys__n34916;
  assign new_new_n24096__ = ~new_new_n23881__ & ~new_new_n24095__;
  assign new_new_n24097__ = ~new_new_n24094__ & new_new_n24096__;
  assign new_new_n24098__ = new_new_n24093__ & ~new_new_n24097__;
  assign new_new_n24099__ = ~new_new_n24093__ & new_new_n24097__;
  assign new_new_n24100__ = ~new_new_n24098__ & ~new_new_n24099__;
  assign new_new_n24101__ = ~new_new_n24083__ & ~new_new_n24100__;
  assign new_new_n24102__ = new_new_n24065__ & new_new_n24101__;
  assign new_new_n24103__ = new_new_n24028__ & new_new_n24102__;
  assign new_new_n24104__ = ~new_new_n23953__ & new_new_n24103__;
  assign new_new_n24105__ = ~new_new_n24075__ & ~new_new_n24080__;
  assign new_new_n24106__ = ~new_new_n24093__ & ~new_new_n24097__;
  assign new_new_n24107__ = ~new_new_n24083__ & new_new_n24106__;
  assign new_new_n24108__ = ~new_new_n24105__ & ~new_new_n24107__;
  assign new_new_n24109__ = new_new_n24065__ & ~new_new_n24108__;
  assign new_new_n24110__ = ~new_new_n24038__ & ~new_new_n24043__;
  assign new_new_n24111__ = ~new_new_n24056__ & ~new_new_n24061__;
  assign new_new_n24112__ = ~new_new_n24046__ & new_new_n24111__;
  assign new_new_n24113__ = ~new_new_n24110__ & ~new_new_n24112__;
  assign new_new_n24114__ = ~new_new_n24109__ & new_new_n24113__;
  assign new_new_n24115__ = new_new_n24028__ & ~new_new_n24114__;
  assign new_new_n24116__ = ~new_new_n24000__ & ~new_new_n24005__;
  assign new_new_n24117__ = ~new_new_n24018__ & ~new_new_n24023__;
  assign new_new_n24118__ = ~new_new_n24008__ & new_new_n24117__;
  assign new_new_n24119__ = ~new_new_n24116__ & ~new_new_n24118__;
  assign new_new_n24120__ = new_new_n23990__ & ~new_new_n24119__;
  assign new_new_n24121__ = ~new_new_n23963__ & ~new_new_n23968__;
  assign new_new_n24122__ = ~new_new_n23981__ & ~new_new_n23986__;
  assign new_new_n24123__ = ~new_new_n23971__ & new_new_n24122__;
  assign new_new_n24124__ = ~new_new_n24121__ & ~new_new_n24123__;
  assign new_new_n24125__ = ~new_new_n24120__ & new_new_n24124__;
  assign new_new_n24126__ = ~new_new_n24115__ & new_new_n24125__;
  assign new_new_n24127__ = ~new_new_n24104__ & new_new_n24126__;
  assign new_new_n24128__ = ~new_new_n23843__ & new_new_n24127__;
  assign new_new_n24129__ = ~new_new_n23669__ & new_new_n23818__;
  assign new_new_n24130__ = new_new_n23830__ & ~new_new_n24129__;
  assign new_new_n24131__ = new_new_n23743__ & ~new_new_n24130__;
  assign new_new_n24132__ = new_new_n23835__ & ~new_new_n24131__;
  assign new_new_n24133__ = ~new_new_n23705__ & ~new_new_n24132__;
  assign new_new_n24134__ = ~new_new_n23838__ & ~new_new_n24133__;
  assign new_new_n24135__ = new_new_n23687__ & ~new_new_n24134__;
  assign new_new_n24136__ = ~new_new_n23687__ & new_new_n24134__;
  assign new_new_n24137__ = ~new_new_n24135__ & ~new_new_n24136__;
  assign new_new_n24138__ = ~new_new_n23669__ & new_new_n23817__;
  assign new_new_n24139__ = new_new_n23824__ & ~new_new_n24138__;
  assign new_new_n24140__ = ~new_new_n23780__ & ~new_new_n24139__;
  assign new_new_n24141__ = ~new_new_n23827__ & ~new_new_n24140__;
  assign new_new_n24142__ = new_new_n23762__ & ~new_new_n24141__;
  assign new_new_n24143__ = ~new_new_n23762__ & new_new_n24141__;
  assign new_new_n24144__ = ~new_new_n24142__ & ~new_new_n24143__;
  assign new_new_n24145__ = new_new_n23780__ & ~new_new_n24139__;
  assign new_new_n24146__ = ~new_new_n23780__ & new_new_n24139__;
  assign new_new_n24147__ = ~new_new_n24145__ & ~new_new_n24146__;
  assign new_new_n24148__ = ~new_new_n23669__ & ~new_new_n23816__;
  assign new_new_n24149__ = ~new_new_n23822__ & ~new_new_n24148__;
  assign new_new_n24150__ = new_new_n23799__ & ~new_new_n24149__;
  assign new_new_n24151__ = ~new_new_n23799__ & new_new_n24149__;
  assign new_new_n24152__ = ~new_new_n24150__ & ~new_new_n24151__;
  assign new_new_n24153__ = ~new_new_n23669__ & new_new_n23816__;
  assign new_new_n24154__ = new_new_n23669__ & ~new_new_n23816__;
  assign new_new_n24155__ = ~new_new_n24153__ & ~new_new_n24154__;
  assign new_new_n24156__ = ~new_new_n24152__ & ~new_new_n24155__;
  assign new_new_n24157__ = ~new_new_n24147__ & new_new_n24156__;
  assign new_new_n24158__ = ~new_new_n24144__ & new_new_n24157__;
  assign new_new_n24159__ = ~new_new_n23742__ & ~new_new_n24130__;
  assign new_new_n24160__ = ~new_new_n23833__ & ~new_new_n24159__;
  assign new_new_n24161__ = new_new_n23724__ & ~new_new_n24160__;
  assign new_new_n24162__ = ~new_new_n23724__ & new_new_n24160__;
  assign new_new_n24163__ = ~new_new_n24161__ & ~new_new_n24162__;
  assign new_new_n24164__ = new_new_n23742__ & ~new_new_n24130__;
  assign new_new_n24165__ = ~new_new_n23742__ & new_new_n24130__;
  assign new_new_n24166__ = ~new_new_n24164__ & ~new_new_n24165__;
  assign new_new_n24167__ = ~new_new_n24163__ & ~new_new_n24166__;
  assign new_new_n24168__ = new_new_n23705__ & ~new_new_n24132__;
  assign new_new_n24169__ = ~new_new_n23705__ & new_new_n24132__;
  assign new_new_n24170__ = ~new_new_n24168__ & ~new_new_n24169__;
  assign new_new_n24171__ = ~new_new_n23582__ & new_new_n23656__;
  assign new_new_n24172__ = new_new_n23662__ & ~new_new_n24171__;
  assign new_new_n24173__ = ~new_new_n23619__ & ~new_new_n24172__;
  assign new_new_n24174__ = ~new_new_n23665__ & ~new_new_n24173__;
  assign new_new_n24175__ = new_new_n23601__ & ~new_new_n24174__;
  assign new_new_n24176__ = ~new_new_n23601__ & new_new_n24174__;
  assign new_new_n24177__ = ~new_new_n24175__ & ~new_new_n24176__;
  assign new_new_n24178__ = ~new_new_n23582__ & ~new_new_n23655__;
  assign new_new_n24179__ = ~new_new_n23660__ & ~new_new_n24178__;
  assign new_new_n24180__ = new_new_n23638__ & ~new_new_n24179__;
  assign new_new_n24181__ = ~new_new_n23638__ & new_new_n24179__;
  assign new_new_n24182__ = ~new_new_n24180__ & ~new_new_n24181__;
  assign new_new_n24183__ = ~new_new_n23582__ & new_new_n23655__;
  assign new_new_n24184__ = new_new_n23582__ & ~new_new_n23655__;
  assign new_new_n24185__ = ~new_new_n24183__ & ~new_new_n24184__;
  assign new_new_n24186__ = ~new_new_n24182__ & ~new_new_n24185__;
  assign new_new_n24187__ = new_new_n23619__ & ~new_new_n24172__;
  assign new_new_n24188__ = ~new_new_n23619__ & new_new_n24172__;
  assign new_new_n24189__ = ~new_new_n24187__ & ~new_new_n24188__;
  assign new_new_n24190__ = ~new_new_n23539__ & ~new_new_n23575__;
  assign new_new_n24191__ = ~new_new_n23579__ & ~new_new_n24190__;
  assign new_new_n24192__ = new_new_n23558__ & ~new_new_n24191__;
  assign new_new_n24193__ = ~new_new_n23558__ & new_new_n24191__;
  assign new_new_n24194__ = ~new_new_n24192__ & ~new_new_n24193__;
  assign new_new_n24195__ = ~new_new_n23539__ & new_new_n23575__;
  assign new_new_n24196__ = new_new_n23539__ & ~new_new_n23575__;
  assign new_new_n24197__ = ~new_new_n24195__ & ~new_new_n24196__;
  assign new_new_n24198__ = new_new_n23521__ & new_new_n23537__;
  assign new_new_n24199__ = ~new_new_n23521__ & ~new_new_n23537__;
  assign new_new_n24200__ = ~new_new_n24198__ & ~new_new_n24199__;
  assign new_new_n24201__ = new_new_n23531__ & ~new_new_n23536__;
  assign new_new_n24202__ = ~new_new_n23531__ & new_new_n23536__;
  assign new_new_n24203__ = ~new_new_n24201__ & ~new_new_n24202__;
  assign new_new_n24204__ = ~new_new_n24200__ & ~new_new_n24203__;
  assign new_new_n24205__ = ~new_new_n24197__ & new_new_n24204__;
  assign new_new_n24206__ = ~new_new_n24194__ & new_new_n24205__;
  assign new_new_n24207__ = ~new_new_n24189__ & new_new_n24206__;
  assign new_new_n24208__ = new_new_n24186__ & new_new_n24207__;
  assign new_new_n24209__ = ~new_new_n24177__ & new_new_n24208__;
  assign new_new_n24210__ = ~new_new_n24170__ & new_new_n24209__;
  assign new_new_n24211__ = new_new_n24167__ & new_new_n24210__;
  assign new_new_n24212__ = new_new_n24158__ & new_new_n24211__;
  assign new_new_n24213__ = ~new_new_n24137__ & new_new_n24212__;
  assign new_new_n24214__ = new_new_n23843__ & new_new_n24213__;
  assign new_new_n24215__ = ~new_new_n23843__ & ~new_new_n24213__;
  assign new_new_n24216__ = ~new_new_n24214__ & ~new_new_n24215__;
  assign new_new_n24217__ = ~new_new_n24127__ & ~new_new_n24216__;
  assign new_new_n24218__ = ~new_new_n24128__ & ~new_new_n24217__;
  assign new_new_n24219__ = ~ys__n33749 & ~new_new_n24218__;
  assign new_new_n24220__ = ~ys__n33749 & ~new_new_n24219__;
  assign new_new_n24221__ = ~new_new_n23501__ & new_new_n24220__;
  assign new_new_n24222__ = new_new_n23501__ & ~new_new_n24220__;
  assign new_new_n24223__ = ~new_new_n24221__ & ~new_new_n24222__;
  assign new_new_n24224__ = ys__n33749 & ~new_new_n24218__;
  assign new_new_n24225__ = ~new_new_n24223__ & ~new_new_n24224__;
  assign new_new_n24226__ = ~new_new_n23501__ & new_new_n24224__;
  assign new_new_n24227__ = ~new_new_n24225__ & ~new_new_n24226__;
  assign new_new_n24228__ = ~new_new_n23480__ & ~new_new_n24227__;
  assign new_new_n24229__ = ~new_new_n23482__ & ~new_new_n24228__;
  assign new_new_n24230__ = ys__n31031 & new_new_n12216__;
  assign new_new_n24231__ = ~new_new_n24229__ & ~new_new_n24230__;
  assign new_new_n24232__ = ~ys__n34948 & ys__n34950;
  assign new_new_n24233__ = ys__n34948 & ~ys__n34950;
  assign new_new_n24234__ = ~new_new_n24232__ & ~new_new_n24233__;
  assign new_new_n24235__ = new_new_n24230__ & ~new_new_n24234__;
  assign new_new_n24236__ = ~new_new_n24231__ & ~new_new_n24235__;
  assign new_new_n24237__ = ys__n2779 & ~ys__n2535;
  assign new_new_n24238__ = ~new_new_n24236__ & new_new_n24237__;
  assign new_new_n24239__ = ys__n2535 & ~new_new_n24236__;
  assign new_new_n24240__ = ~new_new_n24238__ & ~new_new_n24239__;
  assign new_new_n24241__ = ~new_new_n12574__ & ~new_new_n24240__;
  assign new_new_n24242__ = ys__n166 & ys__n30819;
  assign new_new_n24243__ = ~new_new_n23477__ & new_new_n24242__;
  assign new_new_n24244__ = ys__n168 & ys__n30816;
  assign new_new_n24245__ = ys__n30818 & new_new_n24244__;
  assign new_new_n24246__ = ys__n168 & ys__n30820;
  assign new_new_n24247__ = ~new_new_n23477__ & new_new_n24246__;
  assign new_new_n24248__ = ~new_new_n24245__ & ~new_new_n24247__;
  assign new_new_n24249__ = ~new_new_n24243__ & new_new_n24248__;
  assign new_new_n24250__ = ~ys__n166 & ys__n168;
  assign new_new_n24251__ = ys__n47074 & new_new_n24250__;
  assign new_new_n24252__ = ys__n166 & ~ys__n168;
  assign new_new_n24253__ = ys__n47010 & new_new_n24252__;
  assign new_new_n24254__ = ~new_new_n24251__ & ~new_new_n24253__;
  assign new_new_n24255__ = ~new_new_n24250__ & ~new_new_n24252__;
  assign new_new_n24256__ = ~new_new_n24254__ & ~new_new_n24255__;
  assign new_new_n24257__ = new_new_n24249__ & new_new_n24256__;
  assign new_new_n24258__ = new_new_n24127__ & ~new_new_n24203__;
  assign new_new_n24259__ = ~new_new_n24127__ & new_new_n24203__;
  assign new_new_n24260__ = ~new_new_n24258__ & ~new_new_n24259__;
  assign new_new_n24261__ = ~new_new_n24249__ & ~new_new_n24260__;
  assign new_new_n24262__ = ~new_new_n24257__ & ~new_new_n24261__;
  assign new_new_n24263__ = ys__n166 & ys__n30815;
  assign new_new_n24264__ = ys__n30816 & new_new_n24263__;
  assign new_new_n24265__ = ~ys__n2779 & ~new_new_n24264__;
  assign new_new_n24266__ = ~new_new_n24262__ & new_new_n24265__;
  assign new_new_n24267__ = ys__n314 & ~new_new_n24265__;
  assign new_new_n24268__ = ~new_new_n24266__ & ~new_new_n24267__;
  assign new_new_n24269__ = new_new_n12574__ & ~new_new_n24268__;
  assign new_new_n24270__ = ~new_new_n24241__ & ~new_new_n24269__;
  assign new_new_n24271__ = ~ys__n1598 & ~new_new_n24270__;
  assign new_new_n24272__ = ys__n24741 & ys__n1598;
  assign ys__n24742 = new_new_n24271__ | new_new_n24272__;
  assign new_new_n24274__ = ys__n31031 & ys__n47027;
  assign new_new_n24275__ = new_new_n23480__ & new_new_n24274__;
  assign new_new_n24276__ = ys__n34756 & ys__n34758;
  assign new_new_n24277__ = ys__n34760 & new_new_n24276__;
  assign new_new_n24278__ = ~ys__n34756 & ~ys__n34758;
  assign new_new_n24279__ = ys__n34760 & new_new_n24278__;
  assign new_new_n24280__ = ~new_new_n24277__ & ~new_new_n24279__;
  assign new_new_n24281__ = ~ys__n34756 & ys__n34758;
  assign new_new_n24282__ = ~ys__n34760 & new_new_n24281__;
  assign new_new_n24283__ = ys__n34756 & ~ys__n34758;
  assign new_new_n24284__ = ~ys__n34760 & new_new_n24283__;
  assign new_new_n24285__ = ~new_new_n24282__ & ~new_new_n24284__;
  assign new_new_n24286__ = new_new_n24280__ & new_new_n24285__;
  assign new_new_n24287__ = ys__n34764 & ys__n34766;
  assign new_new_n24288__ = ys__n34762 & ys__n34766;
  assign new_new_n24289__ = ~new_new_n23483__ & ~new_new_n24288__;
  assign new_new_n24290__ = ~new_new_n24287__ & new_new_n24289__;
  assign new_new_n24291__ = new_new_n24286__ & ~new_new_n24290__;
  assign new_new_n24292__ = ~new_new_n24286__ & new_new_n24290__;
  assign new_new_n24293__ = ~new_new_n24291__ & ~new_new_n24292__;
  assign new_new_n24294__ = ~new_new_n23493__ & ~new_new_n23498__;
  assign new_new_n24295__ = new_new_n24293__ & new_new_n24294__;
  assign new_new_n24296__ = ~new_new_n24293__ & ~new_new_n24294__;
  assign new_new_n24297__ = ~new_new_n24295__ & ~new_new_n24296__;
  assign new_new_n24298__ = new_new_n24220__ & ~new_new_n24297__;
  assign new_new_n24299__ = ~new_new_n23501__ & new_new_n24297__;
  assign new_new_n24300__ = new_new_n23501__ & ~new_new_n24297__;
  assign new_new_n24301__ = ~new_new_n24299__ & ~new_new_n24300__;
  assign new_new_n24302__ = ~new_new_n24220__ & ~new_new_n24301__;
  assign new_new_n24303__ = ~new_new_n24298__ & ~new_new_n24302__;
  assign new_new_n24304__ = ~new_new_n24224__ & ~new_new_n24303__;
  assign new_new_n24305__ = new_new_n24224__ & new_new_n24297__;
  assign new_new_n24306__ = ~new_new_n24304__ & ~new_new_n24305__;
  assign new_new_n24307__ = ~new_new_n23480__ & ~new_new_n24306__;
  assign new_new_n24308__ = ~new_new_n24275__ & ~new_new_n24307__;
  assign new_new_n24309__ = ~new_new_n24230__ & ~new_new_n24308__;
  assign new_new_n24310__ = new_new_n23871__ & new_new_n23872__;
  assign new_new_n24311__ = ~new_new_n23871__ & ~new_new_n23872__;
  assign new_new_n24312__ = ~new_new_n24310__ & ~new_new_n24311__;
  assign new_new_n24313__ = new_new_n24230__ & ~new_new_n24312__;
  assign new_new_n24314__ = ~new_new_n24309__ & ~new_new_n24313__;
  assign new_new_n24315__ = new_new_n24237__ & ~new_new_n24314__;
  assign new_new_n24316__ = ys__n2535 & ~new_new_n24314__;
  assign new_new_n24317__ = ~new_new_n24315__ & ~new_new_n24316__;
  assign new_new_n24318__ = ~new_new_n12574__ & ~new_new_n24317__;
  assign new_new_n24319__ = ys__n47075 & new_new_n24250__;
  assign new_new_n24320__ = ys__n47011 & new_new_n24252__;
  assign new_new_n24321__ = ~new_new_n24319__ & ~new_new_n24320__;
  assign new_new_n24322__ = ~new_new_n24255__ & ~new_new_n24321__;
  assign new_new_n24323__ = new_new_n24249__ & new_new_n24322__;
  assign new_new_n24324__ = new_new_n24127__ & ~new_new_n24200__;
  assign new_new_n24325__ = new_new_n24200__ & ~new_new_n24203__;
  assign new_new_n24326__ = ~new_new_n24200__ & new_new_n24203__;
  assign new_new_n24327__ = ~new_new_n24325__ & ~new_new_n24326__;
  assign new_new_n24328__ = ~new_new_n24127__ & ~new_new_n24327__;
  assign new_new_n24329__ = ~new_new_n24324__ & ~new_new_n24328__;
  assign new_new_n24330__ = ~new_new_n24249__ & ~new_new_n24329__;
  assign new_new_n24331__ = ~new_new_n24323__ & ~new_new_n24330__;
  assign new_new_n24332__ = new_new_n24265__ & ~new_new_n24331__;
  assign new_new_n24333__ = ys__n170 & ~new_new_n24265__;
  assign new_new_n24334__ = ~new_new_n24332__ & ~new_new_n24333__;
  assign new_new_n24335__ = new_new_n12574__ & ~new_new_n24334__;
  assign new_new_n24336__ = ~new_new_n24318__ & ~new_new_n24335__;
  assign new_new_n24337__ = ~ys__n1598 & ~new_new_n24336__;
  assign new_new_n24338__ = ys__n24744 & ys__n1598;
  assign ys__n24745 = new_new_n24337__ | new_new_n24338__;
  assign new_new_n24340__ = ys__n31031 & ys__n47028;
  assign new_new_n24341__ = new_new_n23480__ & new_new_n24340__;
  assign new_new_n24342__ = ys__n34750 & ys__n34752;
  assign new_new_n24343__ = ys__n34754 & new_new_n24342__;
  assign new_new_n24344__ = ~ys__n34750 & ~ys__n34752;
  assign new_new_n24345__ = ys__n34754 & new_new_n24344__;
  assign new_new_n24346__ = ~new_new_n24343__ & ~new_new_n24345__;
  assign new_new_n24347__ = ~ys__n34750 & ys__n34752;
  assign new_new_n24348__ = ~ys__n34754 & new_new_n24347__;
  assign new_new_n24349__ = ys__n34750 & ~ys__n34752;
  assign new_new_n24350__ = ~ys__n34754 & new_new_n24349__;
  assign new_new_n24351__ = ~new_new_n24348__ & ~new_new_n24350__;
  assign new_new_n24352__ = new_new_n24346__ & new_new_n24351__;
  assign new_new_n24353__ = ys__n34758 & ys__n34760;
  assign new_new_n24354__ = ys__n34756 & ys__n34760;
  assign new_new_n24355__ = ~new_new_n24276__ & ~new_new_n24354__;
  assign new_new_n24356__ = ~new_new_n24353__ & new_new_n24355__;
  assign new_new_n24357__ = new_new_n24352__ & ~new_new_n24356__;
  assign new_new_n24358__ = ~new_new_n24352__ & new_new_n24356__;
  assign new_new_n24359__ = ~new_new_n24357__ & ~new_new_n24358__;
  assign new_new_n24360__ = ~new_new_n24286__ & ~new_new_n24290__;
  assign new_new_n24361__ = ~new_new_n24293__ & new_new_n24294__;
  assign new_new_n24362__ = ~new_new_n24360__ & ~new_new_n24361__;
  assign new_new_n24363__ = new_new_n24359__ & ~new_new_n24362__;
  assign new_new_n24364__ = ~new_new_n24359__ & new_new_n24362__;
  assign new_new_n24365__ = ~new_new_n24363__ & ~new_new_n24364__;
  assign new_new_n24366__ = new_new_n24220__ & ~new_new_n24365__;
  assign new_new_n24367__ = ~new_new_n23501__ & ~new_new_n24297__;
  assign new_new_n24368__ = new_new_n24365__ & new_new_n24367__;
  assign new_new_n24369__ = ~new_new_n24365__ & ~new_new_n24367__;
  assign new_new_n24370__ = ~new_new_n24368__ & ~new_new_n24369__;
  assign new_new_n24371__ = ~new_new_n24220__ & ~new_new_n24370__;
  assign new_new_n24372__ = ~new_new_n24366__ & ~new_new_n24371__;
  assign new_new_n24373__ = ~new_new_n24224__ & ~new_new_n24372__;
  assign new_new_n24374__ = ~new_new_n24297__ & new_new_n24365__;
  assign new_new_n24375__ = new_new_n24297__ & ~new_new_n24365__;
  assign new_new_n24376__ = ~new_new_n24374__ & ~new_new_n24375__;
  assign new_new_n24377__ = new_new_n24224__ & ~new_new_n24376__;
  assign new_new_n24378__ = ~new_new_n24373__ & ~new_new_n24377__;
  assign new_new_n24379__ = ~new_new_n23480__ & ~new_new_n24378__;
  assign new_new_n24380__ = ~new_new_n24341__ & ~new_new_n24379__;
  assign new_new_n24381__ = ~new_new_n24230__ & ~new_new_n24380__;
  assign new_new_n24382__ = new_new_n23858__ & new_new_n23873__;
  assign new_new_n24383__ = ~new_new_n23858__ & ~new_new_n23873__;
  assign new_new_n24384__ = ~new_new_n24382__ & ~new_new_n24383__;
  assign new_new_n24385__ = new_new_n24230__ & ~new_new_n24384__;
  assign new_new_n24386__ = ~new_new_n24381__ & ~new_new_n24385__;
  assign new_new_n24387__ = new_new_n24237__ & ~new_new_n24386__;
  assign new_new_n24388__ = ys__n2535 & ~new_new_n24386__;
  assign new_new_n24389__ = ~new_new_n24387__ & ~new_new_n24388__;
  assign new_new_n24390__ = ~new_new_n12574__ & ~new_new_n24389__;
  assign new_new_n24391__ = ys__n47076 & new_new_n24250__;
  assign new_new_n24392__ = ys__n47012 & new_new_n24252__;
  assign new_new_n24393__ = ~new_new_n24391__ & ~new_new_n24392__;
  assign new_new_n24394__ = ~new_new_n24255__ & ~new_new_n24393__;
  assign new_new_n24395__ = new_new_n24249__ & new_new_n24394__;
  assign new_new_n24396__ = new_new_n24127__ & ~new_new_n24197__;
  assign new_new_n24397__ = new_new_n24197__ & new_new_n24204__;
  assign new_new_n24398__ = ~new_new_n24197__ & ~new_new_n24204__;
  assign new_new_n24399__ = ~new_new_n24397__ & ~new_new_n24398__;
  assign new_new_n24400__ = ~new_new_n24127__ & ~new_new_n24399__;
  assign new_new_n24401__ = ~new_new_n24396__ & ~new_new_n24400__;
  assign new_new_n24402__ = ~new_new_n24249__ & ~new_new_n24401__;
  assign new_new_n24403__ = ~new_new_n24395__ & ~new_new_n24402__;
  assign new_new_n24404__ = new_new_n24265__ & ~new_new_n24403__;
  assign new_new_n24405__ = ys__n380 & ~new_new_n24265__;
  assign new_new_n24406__ = ~new_new_n24404__ & ~new_new_n24405__;
  assign new_new_n24407__ = new_new_n12574__ & ~new_new_n24406__;
  assign new_new_n24408__ = ~new_new_n24390__ & ~new_new_n24407__;
  assign new_new_n24409__ = ~ys__n1598 & ~new_new_n24408__;
  assign new_new_n24410__ = ys__n24747 & ys__n1598;
  assign ys__n24748 = new_new_n24409__ | new_new_n24410__;
  assign new_new_n24412__ = ys__n31031 & ys__n47029;
  assign new_new_n24413__ = new_new_n23480__ & new_new_n24412__;
  assign new_new_n24414__ = ys__n34744 & ys__n34746;
  assign new_new_n24415__ = ys__n34748 & new_new_n24414__;
  assign new_new_n24416__ = ~ys__n34744 & ~ys__n34746;
  assign new_new_n24417__ = ys__n34748 & new_new_n24416__;
  assign new_new_n24418__ = ~new_new_n24415__ & ~new_new_n24417__;
  assign new_new_n24419__ = ~ys__n34744 & ys__n34746;
  assign new_new_n24420__ = ~ys__n34748 & new_new_n24419__;
  assign new_new_n24421__ = ys__n34744 & ~ys__n34746;
  assign new_new_n24422__ = ~ys__n34748 & new_new_n24421__;
  assign new_new_n24423__ = ~new_new_n24420__ & ~new_new_n24422__;
  assign new_new_n24424__ = new_new_n24418__ & new_new_n24423__;
  assign new_new_n24425__ = ys__n34752 & ys__n34754;
  assign new_new_n24426__ = ys__n34750 & ys__n34754;
  assign new_new_n24427__ = ~new_new_n24342__ & ~new_new_n24426__;
  assign new_new_n24428__ = ~new_new_n24425__ & new_new_n24427__;
  assign new_new_n24429__ = new_new_n24424__ & ~new_new_n24428__;
  assign new_new_n24430__ = ~new_new_n24424__ & new_new_n24428__;
  assign new_new_n24431__ = ~new_new_n24429__ & ~new_new_n24430__;
  assign new_new_n24432__ = ~new_new_n24352__ & ~new_new_n24356__;
  assign new_new_n24433__ = ~new_new_n24359__ & ~new_new_n24362__;
  assign new_new_n24434__ = ~new_new_n24432__ & ~new_new_n24433__;
  assign new_new_n24435__ = new_new_n24431__ & ~new_new_n24434__;
  assign new_new_n24436__ = ~new_new_n24431__ & new_new_n24434__;
  assign new_new_n24437__ = ~new_new_n24435__ & ~new_new_n24436__;
  assign new_new_n24438__ = new_new_n24220__ & ~new_new_n24437__;
  assign new_new_n24439__ = ~new_new_n24365__ & new_new_n24367__;
  assign new_new_n24440__ = new_new_n24437__ & new_new_n24439__;
  assign new_new_n24441__ = ~new_new_n24437__ & ~new_new_n24439__;
  assign new_new_n24442__ = ~new_new_n24440__ & ~new_new_n24441__;
  assign new_new_n24443__ = ~new_new_n24220__ & ~new_new_n24442__;
  assign new_new_n24444__ = ~new_new_n24438__ & ~new_new_n24443__;
  assign new_new_n24445__ = ~new_new_n24224__ & ~new_new_n24444__;
  assign new_new_n24446__ = ~new_new_n24297__ & ~new_new_n24365__;
  assign new_new_n24447__ = new_new_n24437__ & new_new_n24446__;
  assign new_new_n24448__ = ~new_new_n24437__ & ~new_new_n24446__;
  assign new_new_n24449__ = ~new_new_n24447__ & ~new_new_n24448__;
  assign new_new_n24450__ = new_new_n24224__ & ~new_new_n24449__;
  assign new_new_n24451__ = ~new_new_n24445__ & ~new_new_n24450__;
  assign new_new_n24452__ = ~new_new_n23480__ & ~new_new_n24451__;
  assign new_new_n24453__ = ~new_new_n24413__ & ~new_new_n24452__;
  assign new_new_n24454__ = ~new_new_n24230__ & ~new_new_n24453__;
  assign new_new_n24455__ = ~new_new_n23858__ & new_new_n23873__;
  assign new_new_n24456__ = ~new_new_n23877__ & ~new_new_n24455__;
  assign new_new_n24457__ = new_new_n23868__ & ~new_new_n24456__;
  assign new_new_n24458__ = ~new_new_n23868__ & new_new_n24456__;
  assign new_new_n24459__ = ~new_new_n24457__ & ~new_new_n24458__;
  assign new_new_n24460__ = new_new_n24230__ & ~new_new_n24459__;
  assign new_new_n24461__ = ~new_new_n24454__ & ~new_new_n24460__;
  assign new_new_n24462__ = new_new_n24237__ & ~new_new_n24461__;
  assign new_new_n24463__ = ys__n2535 & ~new_new_n24461__;
  assign new_new_n24464__ = ~new_new_n24462__ & ~new_new_n24463__;
  assign new_new_n24465__ = ~new_new_n12574__ & ~new_new_n24464__;
  assign new_new_n24466__ = ys__n47077 & new_new_n24250__;
  assign new_new_n24467__ = ys__n47013 & new_new_n24252__;
  assign new_new_n24468__ = ~new_new_n24466__ & ~new_new_n24467__;
  assign new_new_n24469__ = ~new_new_n24255__ & ~new_new_n24468__;
  assign new_new_n24470__ = new_new_n24249__ & new_new_n24469__;
  assign new_new_n24471__ = new_new_n24127__ & ~new_new_n24194__;
  assign new_new_n24472__ = new_new_n24194__ & new_new_n24205__;
  assign new_new_n24473__ = ~new_new_n24194__ & ~new_new_n24205__;
  assign new_new_n24474__ = ~new_new_n24472__ & ~new_new_n24473__;
  assign new_new_n24475__ = ~new_new_n24127__ & ~new_new_n24474__;
  assign new_new_n24476__ = ~new_new_n24471__ & ~new_new_n24475__;
  assign new_new_n24477__ = ~new_new_n24249__ & ~new_new_n24476__;
  assign new_new_n24478__ = ~new_new_n24470__ & ~new_new_n24477__;
  assign new_new_n24479__ = new_new_n24265__ & ~new_new_n24478__;
  assign new_new_n24480__ = ys__n378 & ~new_new_n24265__;
  assign new_new_n24481__ = ~new_new_n24479__ & ~new_new_n24480__;
  assign new_new_n24482__ = new_new_n12574__ & ~new_new_n24481__;
  assign new_new_n24483__ = ~new_new_n24465__ & ~new_new_n24482__;
  assign new_new_n24484__ = ~ys__n1598 & ~new_new_n24483__;
  assign new_new_n24485__ = ys__n24750 & ys__n1598;
  assign ys__n24751 = new_new_n24484__ | new_new_n24485__;
  assign new_new_n24487__ = ys__n31031 & ys__n47030;
  assign new_new_n24488__ = new_new_n23480__ & new_new_n24487__;
  assign new_new_n24489__ = ys__n34738 & ys__n34740;
  assign new_new_n24490__ = ys__n34742 & new_new_n24489__;
  assign new_new_n24491__ = ~ys__n34738 & ~ys__n34740;
  assign new_new_n24492__ = ys__n34742 & new_new_n24491__;
  assign new_new_n24493__ = ~new_new_n24490__ & ~new_new_n24492__;
  assign new_new_n24494__ = ~ys__n34738 & ys__n34740;
  assign new_new_n24495__ = ~ys__n34742 & new_new_n24494__;
  assign new_new_n24496__ = ys__n34738 & ~ys__n34740;
  assign new_new_n24497__ = ~ys__n34742 & new_new_n24496__;
  assign new_new_n24498__ = ~new_new_n24495__ & ~new_new_n24497__;
  assign new_new_n24499__ = new_new_n24493__ & new_new_n24498__;
  assign new_new_n24500__ = ys__n34746 & ys__n34748;
  assign new_new_n24501__ = ys__n34744 & ys__n34748;
  assign new_new_n24502__ = ~new_new_n24414__ & ~new_new_n24501__;
  assign new_new_n24503__ = ~new_new_n24500__ & new_new_n24502__;
  assign new_new_n24504__ = new_new_n24499__ & ~new_new_n24503__;
  assign new_new_n24505__ = ~new_new_n24499__ & new_new_n24503__;
  assign new_new_n24506__ = ~new_new_n24504__ & ~new_new_n24505__;
  assign new_new_n24507__ = ~new_new_n24359__ & ~new_new_n24431__;
  assign new_new_n24508__ = ~new_new_n24362__ & new_new_n24507__;
  assign new_new_n24509__ = ~new_new_n24424__ & ~new_new_n24428__;
  assign new_new_n24510__ = ~new_new_n24431__ & new_new_n24432__;
  assign new_new_n24511__ = ~new_new_n24509__ & ~new_new_n24510__;
  assign new_new_n24512__ = ~new_new_n24508__ & new_new_n24511__;
  assign new_new_n24513__ = new_new_n24506__ & ~new_new_n24512__;
  assign new_new_n24514__ = ~new_new_n24506__ & new_new_n24512__;
  assign new_new_n24515__ = ~new_new_n24513__ & ~new_new_n24514__;
  assign new_new_n24516__ = new_new_n24220__ & ~new_new_n24515__;
  assign new_new_n24517__ = ~new_new_n24365__ & ~new_new_n24437__;
  assign new_new_n24518__ = new_new_n24367__ & new_new_n24517__;
  assign new_new_n24519__ = new_new_n24515__ & new_new_n24518__;
  assign new_new_n24520__ = ~new_new_n24515__ & ~new_new_n24518__;
  assign new_new_n24521__ = ~new_new_n24519__ & ~new_new_n24520__;
  assign new_new_n24522__ = ~new_new_n24220__ & ~new_new_n24521__;
  assign new_new_n24523__ = ~new_new_n24516__ & ~new_new_n24522__;
  assign new_new_n24524__ = ~new_new_n24224__ & ~new_new_n24523__;
  assign new_new_n24525__ = ~new_new_n24297__ & new_new_n24517__;
  assign new_new_n24526__ = new_new_n24515__ & new_new_n24525__;
  assign new_new_n24527__ = ~new_new_n24515__ & ~new_new_n24525__;
  assign new_new_n24528__ = ~new_new_n24526__ & ~new_new_n24527__;
  assign new_new_n24529__ = new_new_n24224__ & ~new_new_n24528__;
  assign new_new_n24530__ = ~new_new_n24524__ & ~new_new_n24529__;
  assign new_new_n24531__ = ~new_new_n23480__ & ~new_new_n24530__;
  assign new_new_n24532__ = ~new_new_n24488__ & ~new_new_n24531__;
  assign new_new_n24533__ = ~new_new_n24230__ & ~new_new_n24532__;
  assign new_new_n24534__ = ~new_new_n23880__ & new_new_n23939__;
  assign new_new_n24535__ = new_new_n23880__ & ~new_new_n23939__;
  assign new_new_n24536__ = ~new_new_n24534__ & ~new_new_n24535__;
  assign new_new_n24537__ = new_new_n24230__ & ~new_new_n24536__;
  assign new_new_n24538__ = ~new_new_n24533__ & ~new_new_n24537__;
  assign new_new_n24539__ = new_new_n24237__ & ~new_new_n24538__;
  assign new_new_n24540__ = ys__n2535 & ~new_new_n24538__;
  assign new_new_n24541__ = ~new_new_n24539__ & ~new_new_n24540__;
  assign new_new_n24542__ = ~new_new_n12574__ & ~new_new_n24541__;
  assign new_new_n24543__ = ys__n47078 & new_new_n24250__;
  assign new_new_n24544__ = ys__n47014 & new_new_n24252__;
  assign new_new_n24545__ = ~new_new_n24543__ & ~new_new_n24544__;
  assign new_new_n24546__ = ~new_new_n24255__ & ~new_new_n24545__;
  assign new_new_n24547__ = new_new_n24249__ & new_new_n24546__;
  assign new_new_n24548__ = new_new_n24127__ & ~new_new_n24185__;
  assign new_new_n24549__ = new_new_n24185__ & new_new_n24206__;
  assign new_new_n24550__ = ~new_new_n24185__ & ~new_new_n24206__;
  assign new_new_n24551__ = ~new_new_n24549__ & ~new_new_n24550__;
  assign new_new_n24552__ = ~new_new_n24127__ & ~new_new_n24551__;
  assign new_new_n24553__ = ~new_new_n24548__ & ~new_new_n24552__;
  assign new_new_n24554__ = ~new_new_n24249__ & ~new_new_n24553__;
  assign new_new_n24555__ = ~new_new_n24547__ & ~new_new_n24554__;
  assign new_new_n24556__ = new_new_n24265__ & ~new_new_n24555__;
  assign new_new_n24557__ = ys__n382 & ~new_new_n24265__;
  assign new_new_n24558__ = ~new_new_n24556__ & ~new_new_n24557__;
  assign new_new_n24559__ = new_new_n12574__ & ~new_new_n24558__;
  assign new_new_n24560__ = ~new_new_n24542__ & ~new_new_n24559__;
  assign new_new_n24561__ = ~ys__n1598 & ~new_new_n24560__;
  assign new_new_n24562__ = ys__n24753 & ys__n1598;
  assign ys__n24754 = new_new_n24561__ | new_new_n24562__;
  assign new_new_n24564__ = ys__n31031 & ys__n47031;
  assign new_new_n24565__ = new_new_n23480__ & new_new_n24564__;
  assign new_new_n24566__ = ys__n34732 & ys__n34734;
  assign new_new_n24567__ = ys__n34736 & new_new_n24566__;
  assign new_new_n24568__ = ~ys__n34732 & ~ys__n34734;
  assign new_new_n24569__ = ys__n34736 & new_new_n24568__;
  assign new_new_n24570__ = ~new_new_n24567__ & ~new_new_n24569__;
  assign new_new_n24571__ = ~ys__n34732 & ys__n34734;
  assign new_new_n24572__ = ~ys__n34736 & new_new_n24571__;
  assign new_new_n24573__ = ys__n34732 & ~ys__n34734;
  assign new_new_n24574__ = ~ys__n34736 & new_new_n24573__;
  assign new_new_n24575__ = ~new_new_n24572__ & ~new_new_n24574__;
  assign new_new_n24576__ = new_new_n24570__ & new_new_n24575__;
  assign new_new_n24577__ = ys__n34740 & ys__n34742;
  assign new_new_n24578__ = ys__n34738 & ys__n34742;
  assign new_new_n24579__ = ~new_new_n24489__ & ~new_new_n24578__;
  assign new_new_n24580__ = ~new_new_n24577__ & new_new_n24579__;
  assign new_new_n24581__ = new_new_n24576__ & ~new_new_n24580__;
  assign new_new_n24582__ = ~new_new_n24576__ & new_new_n24580__;
  assign new_new_n24583__ = ~new_new_n24581__ & ~new_new_n24582__;
  assign new_new_n24584__ = ~new_new_n24499__ & ~new_new_n24503__;
  assign new_new_n24585__ = ~new_new_n24506__ & ~new_new_n24512__;
  assign new_new_n24586__ = ~new_new_n24584__ & ~new_new_n24585__;
  assign new_new_n24587__ = new_new_n24583__ & ~new_new_n24586__;
  assign new_new_n24588__ = ~new_new_n24583__ & new_new_n24586__;
  assign new_new_n24589__ = ~new_new_n24587__ & ~new_new_n24588__;
  assign new_new_n24590__ = new_new_n24220__ & ~new_new_n24589__;
  assign new_new_n24591__ = ~new_new_n24515__ & new_new_n24518__;
  assign new_new_n24592__ = new_new_n24589__ & new_new_n24591__;
  assign new_new_n24593__ = ~new_new_n24589__ & ~new_new_n24591__;
  assign new_new_n24594__ = ~new_new_n24592__ & ~new_new_n24593__;
  assign new_new_n24595__ = ~new_new_n24220__ & ~new_new_n24594__;
  assign new_new_n24596__ = ~new_new_n24590__ & ~new_new_n24595__;
  assign new_new_n24597__ = ~new_new_n24224__ & ~new_new_n24596__;
  assign new_new_n24598__ = ~new_new_n24515__ & new_new_n24525__;
  assign new_new_n24599__ = new_new_n24589__ & new_new_n24598__;
  assign new_new_n24600__ = ~new_new_n24589__ & ~new_new_n24598__;
  assign new_new_n24601__ = ~new_new_n24599__ & ~new_new_n24600__;
  assign new_new_n24602__ = new_new_n24224__ & ~new_new_n24601__;
  assign new_new_n24603__ = ~new_new_n24597__ & ~new_new_n24602__;
  assign new_new_n24604__ = ~new_new_n23480__ & ~new_new_n24603__;
  assign new_new_n24605__ = ~new_new_n24565__ & ~new_new_n24604__;
  assign new_new_n24606__ = ~new_new_n24230__ & ~new_new_n24605__;
  assign new_new_n24607__ = ~new_new_n23880__ & ~new_new_n23939__;
  assign new_new_n24608__ = ~new_new_n23944__ & ~new_new_n24607__;
  assign new_new_n24609__ = new_new_n23932__ & ~new_new_n24608__;
  assign new_new_n24610__ = ~new_new_n23932__ & new_new_n24608__;
  assign new_new_n24611__ = ~new_new_n24609__ & ~new_new_n24610__;
  assign new_new_n24612__ = new_new_n24230__ & ~new_new_n24611__;
  assign new_new_n24613__ = ~new_new_n24606__ & ~new_new_n24612__;
  assign new_new_n24614__ = new_new_n24237__ & ~new_new_n24613__;
  assign new_new_n24615__ = ys__n2535 & ~new_new_n24613__;
  assign new_new_n24616__ = ~new_new_n24614__ & ~new_new_n24615__;
  assign new_new_n24617__ = ~new_new_n12574__ & ~new_new_n24616__;
  assign new_new_n24618__ = ys__n47079 & new_new_n24250__;
  assign new_new_n24619__ = ys__n47015 & new_new_n24252__;
  assign new_new_n24620__ = ~new_new_n24618__ & ~new_new_n24619__;
  assign new_new_n24621__ = ~new_new_n24255__ & ~new_new_n24620__;
  assign new_new_n24622__ = new_new_n24249__ & new_new_n24621__;
  assign new_new_n24623__ = new_new_n24127__ & ~new_new_n24182__;
  assign new_new_n24624__ = ~new_new_n24185__ & new_new_n24206__;
  assign new_new_n24625__ = new_new_n24182__ & new_new_n24624__;
  assign new_new_n24626__ = ~new_new_n24182__ & ~new_new_n24624__;
  assign new_new_n24627__ = ~new_new_n24625__ & ~new_new_n24626__;
  assign new_new_n24628__ = ~new_new_n24127__ & ~new_new_n24627__;
  assign new_new_n24629__ = ~new_new_n24623__ & ~new_new_n24628__;
  assign new_new_n24630__ = ~new_new_n24249__ & ~new_new_n24629__;
  assign new_new_n24631__ = ~new_new_n24622__ & ~new_new_n24630__;
  assign new_new_n24632__ = new_new_n24265__ & ~new_new_n24631__;
  assign new_new_n24633__ = ys__n374 & ~new_new_n24265__;
  assign new_new_n24634__ = ~new_new_n24632__ & ~new_new_n24633__;
  assign new_new_n24635__ = new_new_n12574__ & ~new_new_n24634__;
  assign new_new_n24636__ = ~new_new_n24617__ & ~new_new_n24635__;
  assign new_new_n24637__ = ~ys__n1598 & ~new_new_n24636__;
  assign new_new_n24638__ = ys__n24756 & ys__n1598;
  assign ys__n24757 = new_new_n24637__ | new_new_n24638__;
  assign new_new_n24640__ = ys__n31031 & ys__n47032;
  assign new_new_n24641__ = new_new_n23480__ & new_new_n24640__;
  assign new_new_n24642__ = ys__n34726 & ys__n34728;
  assign new_new_n24643__ = ys__n34730 & new_new_n24642__;
  assign new_new_n24644__ = ~ys__n34726 & ~ys__n34728;
  assign new_new_n24645__ = ys__n34730 & new_new_n24644__;
  assign new_new_n24646__ = ~new_new_n24643__ & ~new_new_n24645__;
  assign new_new_n24647__ = ~ys__n34726 & ys__n34728;
  assign new_new_n24648__ = ~ys__n34730 & new_new_n24647__;
  assign new_new_n24649__ = ys__n34726 & ~ys__n34728;
  assign new_new_n24650__ = ~ys__n34730 & new_new_n24649__;
  assign new_new_n24651__ = ~new_new_n24648__ & ~new_new_n24650__;
  assign new_new_n24652__ = new_new_n24646__ & new_new_n24651__;
  assign new_new_n24653__ = ys__n34734 & ys__n34736;
  assign new_new_n24654__ = ys__n34732 & ys__n34736;
  assign new_new_n24655__ = ~new_new_n24566__ & ~new_new_n24654__;
  assign new_new_n24656__ = ~new_new_n24653__ & new_new_n24655__;
  assign new_new_n24657__ = new_new_n24652__ & ~new_new_n24656__;
  assign new_new_n24658__ = ~new_new_n24652__ & new_new_n24656__;
  assign new_new_n24659__ = ~new_new_n24657__ & ~new_new_n24658__;
  assign new_new_n24660__ = ~new_new_n24576__ & ~new_new_n24580__;
  assign new_new_n24661__ = ~new_new_n24583__ & new_new_n24584__;
  assign new_new_n24662__ = ~new_new_n24660__ & ~new_new_n24661__;
  assign new_new_n24663__ = ~new_new_n24506__ & ~new_new_n24583__;
  assign new_new_n24664__ = ~new_new_n24512__ & new_new_n24663__;
  assign new_new_n24665__ = new_new_n24662__ & ~new_new_n24664__;
  assign new_new_n24666__ = new_new_n24659__ & ~new_new_n24665__;
  assign new_new_n24667__ = ~new_new_n24659__ & new_new_n24665__;
  assign new_new_n24668__ = ~new_new_n24666__ & ~new_new_n24667__;
  assign new_new_n24669__ = new_new_n24220__ & ~new_new_n24668__;
  assign new_new_n24670__ = ~new_new_n24515__ & ~new_new_n24589__;
  assign new_new_n24671__ = new_new_n24518__ & new_new_n24670__;
  assign new_new_n24672__ = new_new_n24668__ & new_new_n24671__;
  assign new_new_n24673__ = ~new_new_n24668__ & ~new_new_n24671__;
  assign new_new_n24674__ = ~new_new_n24672__ & ~new_new_n24673__;
  assign new_new_n24675__ = ~new_new_n24220__ & ~new_new_n24674__;
  assign new_new_n24676__ = ~new_new_n24669__ & ~new_new_n24675__;
  assign new_new_n24677__ = ~new_new_n24224__ & ~new_new_n24676__;
  assign new_new_n24678__ = new_new_n24525__ & new_new_n24670__;
  assign new_new_n24679__ = new_new_n24668__ & new_new_n24678__;
  assign new_new_n24680__ = ~new_new_n24668__ & ~new_new_n24678__;
  assign new_new_n24681__ = ~new_new_n24679__ & ~new_new_n24680__;
  assign new_new_n24682__ = new_new_n24224__ & ~new_new_n24681__;
  assign new_new_n24683__ = ~new_new_n24677__ & ~new_new_n24682__;
  assign new_new_n24684__ = ~new_new_n23480__ & ~new_new_n24683__;
  assign new_new_n24685__ = ~new_new_n24641__ & ~new_new_n24684__;
  assign new_new_n24686__ = ~new_new_n24230__ & ~new_new_n24685__;
  assign new_new_n24687__ = ~new_new_n23880__ & new_new_n23940__;
  assign new_new_n24688__ = new_new_n23946__ & ~new_new_n24687__;
  assign new_new_n24689__ = new_new_n23917__ & ~new_new_n24688__;
  assign new_new_n24690__ = ~new_new_n23917__ & new_new_n24688__;
  assign new_new_n24691__ = ~new_new_n24689__ & ~new_new_n24690__;
  assign new_new_n24692__ = new_new_n24230__ & ~new_new_n24691__;
  assign new_new_n24693__ = ~new_new_n24686__ & ~new_new_n24692__;
  assign new_new_n24694__ = new_new_n24237__ & ~new_new_n24693__;
  assign new_new_n24695__ = ys__n2535 & ~new_new_n24693__;
  assign new_new_n24696__ = ~new_new_n24694__ & ~new_new_n24695__;
  assign new_new_n24697__ = ~new_new_n12574__ & ~new_new_n24696__;
  assign new_new_n24698__ = ys__n47080 & new_new_n24250__;
  assign new_new_n24699__ = ys__n47016 & new_new_n24252__;
  assign new_new_n24700__ = ~new_new_n24698__ & ~new_new_n24699__;
  assign new_new_n24701__ = ~new_new_n24255__ & ~new_new_n24700__;
  assign new_new_n24702__ = new_new_n24249__ & new_new_n24701__;
  assign new_new_n24703__ = new_new_n24127__ & ~new_new_n24189__;
  assign new_new_n24704__ = new_new_n24186__ & new_new_n24206__;
  assign new_new_n24705__ = new_new_n24189__ & new_new_n24704__;
  assign new_new_n24706__ = ~new_new_n24189__ & ~new_new_n24704__;
  assign new_new_n24707__ = ~new_new_n24705__ & ~new_new_n24706__;
  assign new_new_n24708__ = ~new_new_n24127__ & ~new_new_n24707__;
  assign new_new_n24709__ = ~new_new_n24703__ & ~new_new_n24708__;
  assign new_new_n24710__ = ~new_new_n24249__ & ~new_new_n24709__;
  assign new_new_n24711__ = ~new_new_n24702__ & ~new_new_n24710__;
  assign new_new_n24712__ = new_new_n24265__ & ~new_new_n24711__;
  assign new_new_n24713__ = ys__n376 & ~new_new_n24265__;
  assign new_new_n24714__ = ~new_new_n24712__ & ~new_new_n24713__;
  assign new_new_n24715__ = new_new_n12574__ & ~new_new_n24714__;
  assign new_new_n24716__ = ~new_new_n24697__ & ~new_new_n24715__;
  assign new_new_n24717__ = ~ys__n1598 & ~new_new_n24716__;
  assign new_new_n24718__ = ys__n24759 & ys__n1598;
  assign ys__n24760 = new_new_n24717__ | new_new_n24718__;
  assign new_new_n24720__ = ys__n31031 & ys__n47033;
  assign new_new_n24721__ = new_new_n23480__ & new_new_n24720__;
  assign new_new_n24722__ = ys__n34720 & ys__n34722;
  assign new_new_n24723__ = ys__n34724 & new_new_n24722__;
  assign new_new_n24724__ = ~ys__n34720 & ~ys__n34722;
  assign new_new_n24725__ = ys__n34724 & new_new_n24724__;
  assign new_new_n24726__ = ~new_new_n24723__ & ~new_new_n24725__;
  assign new_new_n24727__ = ~ys__n34720 & ys__n34722;
  assign new_new_n24728__ = ~ys__n34724 & new_new_n24727__;
  assign new_new_n24729__ = ys__n34720 & ~ys__n34722;
  assign new_new_n24730__ = ~ys__n34724 & new_new_n24729__;
  assign new_new_n24731__ = ~new_new_n24728__ & ~new_new_n24730__;
  assign new_new_n24732__ = new_new_n24726__ & new_new_n24731__;
  assign new_new_n24733__ = ys__n34728 & ys__n34730;
  assign new_new_n24734__ = ys__n34726 & ys__n34730;
  assign new_new_n24735__ = ~new_new_n24642__ & ~new_new_n24734__;
  assign new_new_n24736__ = ~new_new_n24733__ & new_new_n24735__;
  assign new_new_n24737__ = new_new_n24732__ & ~new_new_n24736__;
  assign new_new_n24738__ = ~new_new_n24732__ & new_new_n24736__;
  assign new_new_n24739__ = ~new_new_n24737__ & ~new_new_n24738__;
  assign new_new_n24740__ = ~new_new_n24652__ & ~new_new_n24656__;
  assign new_new_n24741__ = ~new_new_n24659__ & ~new_new_n24665__;
  assign new_new_n24742__ = ~new_new_n24740__ & ~new_new_n24741__;
  assign new_new_n24743__ = new_new_n24739__ & ~new_new_n24742__;
  assign new_new_n24744__ = ~new_new_n24739__ & new_new_n24742__;
  assign new_new_n24745__ = ~new_new_n24743__ & ~new_new_n24744__;
  assign new_new_n24746__ = new_new_n24220__ & ~new_new_n24745__;
  assign new_new_n24747__ = ~new_new_n24668__ & new_new_n24671__;
  assign new_new_n24748__ = new_new_n24745__ & new_new_n24747__;
  assign new_new_n24749__ = ~new_new_n24745__ & ~new_new_n24747__;
  assign new_new_n24750__ = ~new_new_n24748__ & ~new_new_n24749__;
  assign new_new_n24751__ = ~new_new_n24220__ & ~new_new_n24750__;
  assign new_new_n24752__ = ~new_new_n24746__ & ~new_new_n24751__;
  assign new_new_n24753__ = ~new_new_n24224__ & ~new_new_n24752__;
  assign new_new_n24754__ = ~new_new_n24668__ & new_new_n24678__;
  assign new_new_n24755__ = new_new_n24745__ & new_new_n24754__;
  assign new_new_n24756__ = ~new_new_n24745__ & ~new_new_n24754__;
  assign new_new_n24757__ = ~new_new_n24755__ & ~new_new_n24756__;
  assign new_new_n24758__ = new_new_n24224__ & ~new_new_n24757__;
  assign new_new_n24759__ = ~new_new_n24753__ & ~new_new_n24758__;
  assign new_new_n24760__ = ~new_new_n23480__ & ~new_new_n24759__;
  assign new_new_n24761__ = ~new_new_n24721__ & ~new_new_n24760__;
  assign new_new_n24762__ = ~new_new_n24230__ & ~new_new_n24761__;
  assign new_new_n24763__ = ~new_new_n23917__ & ~new_new_n24688__;
  assign new_new_n24764__ = ~new_new_n23949__ & ~new_new_n24763__;
  assign new_new_n24765__ = new_new_n23899__ & ~new_new_n24764__;
  assign new_new_n24766__ = ~new_new_n23899__ & new_new_n24764__;
  assign new_new_n24767__ = ~new_new_n24765__ & ~new_new_n24766__;
  assign new_new_n24768__ = new_new_n24230__ & ~new_new_n24767__;
  assign new_new_n24769__ = ~new_new_n24762__ & ~new_new_n24768__;
  assign new_new_n24770__ = new_new_n24237__ & ~new_new_n24769__;
  assign new_new_n24771__ = ys__n2535 & ~new_new_n24769__;
  assign new_new_n24772__ = ~new_new_n24770__ & ~new_new_n24771__;
  assign new_new_n24773__ = ~new_new_n12574__ & ~new_new_n24772__;
  assign new_new_n24774__ = ys__n47081 & new_new_n24250__;
  assign new_new_n24775__ = ys__n47017 & new_new_n24252__;
  assign new_new_n24776__ = ~new_new_n24774__ & ~new_new_n24775__;
  assign new_new_n24777__ = ~new_new_n24255__ & ~new_new_n24776__;
  assign new_new_n24778__ = new_new_n24249__ & new_new_n24777__;
  assign new_new_n24779__ = new_new_n24127__ & ~new_new_n24177__;
  assign new_new_n24780__ = ~new_new_n24189__ & new_new_n24704__;
  assign new_new_n24781__ = new_new_n24177__ & new_new_n24780__;
  assign new_new_n24782__ = ~new_new_n24177__ & ~new_new_n24780__;
  assign new_new_n24783__ = ~new_new_n24781__ & ~new_new_n24782__;
  assign new_new_n24784__ = ~new_new_n24127__ & ~new_new_n24783__;
  assign new_new_n24785__ = ~new_new_n24779__ & ~new_new_n24784__;
  assign new_new_n24786__ = ~new_new_n24249__ & ~new_new_n24785__;
  assign new_new_n24787__ = ~new_new_n24778__ & ~new_new_n24786__;
  assign new_new_n24788__ = new_new_n24265__ & ~new_new_n24787__;
  assign new_new_n24789__ = ys__n372 & ~new_new_n24265__;
  assign new_new_n24790__ = ~new_new_n24788__ & ~new_new_n24789__;
  assign new_new_n24791__ = new_new_n12574__ & ~new_new_n24790__;
  assign new_new_n24792__ = ~new_new_n24773__ & ~new_new_n24791__;
  assign new_new_n24793__ = ~ys__n1598 & ~new_new_n24792__;
  assign new_new_n24794__ = ys__n24762 & ys__n1598;
  assign ys__n24763 = new_new_n24793__ | new_new_n24794__;
  assign new_new_n24796__ = ys__n31031 & ys__n47034;
  assign new_new_n24797__ = new_new_n23480__ & new_new_n24796__;
  assign new_new_n24798__ = ys__n34714 & ys__n34716;
  assign new_new_n24799__ = ys__n34718 & new_new_n24798__;
  assign new_new_n24800__ = ~ys__n34714 & ~ys__n34716;
  assign new_new_n24801__ = ys__n34718 & new_new_n24800__;
  assign new_new_n24802__ = ~new_new_n24799__ & ~new_new_n24801__;
  assign new_new_n24803__ = ~ys__n34714 & ys__n34716;
  assign new_new_n24804__ = ~ys__n34718 & new_new_n24803__;
  assign new_new_n24805__ = ys__n34714 & ~ys__n34716;
  assign new_new_n24806__ = ~ys__n34718 & new_new_n24805__;
  assign new_new_n24807__ = ~new_new_n24804__ & ~new_new_n24806__;
  assign new_new_n24808__ = new_new_n24802__ & new_new_n24807__;
  assign new_new_n24809__ = ys__n34722 & ys__n34724;
  assign new_new_n24810__ = ys__n34720 & ys__n34724;
  assign new_new_n24811__ = ~new_new_n24722__ & ~new_new_n24810__;
  assign new_new_n24812__ = ~new_new_n24809__ & new_new_n24811__;
  assign new_new_n24813__ = new_new_n24808__ & ~new_new_n24812__;
  assign new_new_n24814__ = ~new_new_n24808__ & new_new_n24812__;
  assign new_new_n24815__ = ~new_new_n24813__ & ~new_new_n24814__;
  assign new_new_n24816__ = ~new_new_n24659__ & ~new_new_n24739__;
  assign new_new_n24817__ = new_new_n24663__ & new_new_n24816__;
  assign new_new_n24818__ = ~new_new_n24512__ & new_new_n24817__;
  assign new_new_n24819__ = ~new_new_n24662__ & new_new_n24816__;
  assign new_new_n24820__ = ~new_new_n24732__ & ~new_new_n24736__;
  assign new_new_n24821__ = ~new_new_n24739__ & new_new_n24740__;
  assign new_new_n24822__ = ~new_new_n24820__ & ~new_new_n24821__;
  assign new_new_n24823__ = ~new_new_n24819__ & new_new_n24822__;
  assign new_new_n24824__ = ~new_new_n24818__ & new_new_n24823__;
  assign new_new_n24825__ = new_new_n24815__ & ~new_new_n24824__;
  assign new_new_n24826__ = ~new_new_n24815__ & new_new_n24824__;
  assign new_new_n24827__ = ~new_new_n24825__ & ~new_new_n24826__;
  assign new_new_n24828__ = new_new_n24220__ & ~new_new_n24827__;
  assign new_new_n24829__ = ~new_new_n24668__ & new_new_n24670__;
  assign new_new_n24830__ = ~new_new_n24745__ & new_new_n24829__;
  assign new_new_n24831__ = new_new_n24518__ & new_new_n24830__;
  assign new_new_n24832__ = new_new_n24827__ & new_new_n24831__;
  assign new_new_n24833__ = ~new_new_n24827__ & ~new_new_n24831__;
  assign new_new_n24834__ = ~new_new_n24832__ & ~new_new_n24833__;
  assign new_new_n24835__ = ~new_new_n24220__ & ~new_new_n24834__;
  assign new_new_n24836__ = ~new_new_n24828__ & ~new_new_n24835__;
  assign new_new_n24837__ = ~new_new_n24224__ & ~new_new_n24836__;
  assign new_new_n24838__ = new_new_n24525__ & new_new_n24830__;
  assign new_new_n24839__ = new_new_n24827__ & new_new_n24838__;
  assign new_new_n24840__ = ~new_new_n24827__ & ~new_new_n24838__;
  assign new_new_n24841__ = ~new_new_n24839__ & ~new_new_n24840__;
  assign new_new_n24842__ = new_new_n24224__ & ~new_new_n24841__;
  assign new_new_n24843__ = ~new_new_n24837__ & ~new_new_n24842__;
  assign new_new_n24844__ = ~new_new_n23480__ & ~new_new_n24843__;
  assign new_new_n24845__ = ~new_new_n24797__ & ~new_new_n24844__;
  assign new_new_n24846__ = ~new_new_n24230__ & ~new_new_n24845__;
  assign new_new_n24847__ = ~new_new_n23953__ & new_new_n24100__;
  assign new_new_n24848__ = new_new_n23953__ & ~new_new_n24100__;
  assign new_new_n24849__ = ~new_new_n24847__ & ~new_new_n24848__;
  assign new_new_n24850__ = new_new_n24230__ & ~new_new_n24849__;
  assign new_new_n24851__ = ~new_new_n24846__ & ~new_new_n24850__;
  assign new_new_n24852__ = new_new_n24237__ & ~new_new_n24851__;
  assign new_new_n24853__ = ys__n2535 & ~new_new_n24851__;
  assign new_new_n24854__ = ~new_new_n24852__ & ~new_new_n24853__;
  assign new_new_n24855__ = ~new_new_n12574__ & ~new_new_n24854__;
  assign new_new_n24856__ = ys__n47082 & new_new_n24250__;
  assign new_new_n24857__ = ys__n47018 & new_new_n24252__;
  assign new_new_n24858__ = ~new_new_n24856__ & ~new_new_n24857__;
  assign new_new_n24859__ = ~new_new_n24255__ & ~new_new_n24858__;
  assign new_new_n24860__ = new_new_n24249__ & new_new_n24859__;
  assign new_new_n24861__ = new_new_n24127__ & ~new_new_n24155__;
  assign new_new_n24862__ = new_new_n24155__ & new_new_n24209__;
  assign new_new_n24863__ = ~new_new_n24155__ & ~new_new_n24209__;
  assign new_new_n24864__ = ~new_new_n24862__ & ~new_new_n24863__;
  assign new_new_n24865__ = ~new_new_n24127__ & ~new_new_n24864__;
  assign new_new_n24866__ = ~new_new_n24861__ & ~new_new_n24865__;
  assign new_new_n24867__ = ~new_new_n24249__ & ~new_new_n24866__;
  assign new_new_n24868__ = ~new_new_n24860__ & ~new_new_n24867__;
  assign new_new_n24869__ = new_new_n24265__ & ~new_new_n24868__;
  assign new_new_n24870__ = ys__n384 & ~new_new_n24265__;
  assign new_new_n24871__ = ~new_new_n24869__ & ~new_new_n24870__;
  assign new_new_n24872__ = new_new_n12574__ & ~new_new_n24871__;
  assign new_new_n24873__ = ~new_new_n24855__ & ~new_new_n24872__;
  assign new_new_n24874__ = ~ys__n1598 & ~new_new_n24873__;
  assign new_new_n24875__ = ys__n24765 & ys__n1598;
  assign ys__n24766 = new_new_n24874__ | new_new_n24875__;
  assign new_new_n24877__ = ys__n31031 & ys__n47035;
  assign new_new_n24878__ = new_new_n23480__ & new_new_n24877__;
  assign new_new_n24879__ = ys__n34708 & ys__n34710;
  assign new_new_n24880__ = ys__n34712 & new_new_n24879__;
  assign new_new_n24881__ = ~ys__n34708 & ~ys__n34710;
  assign new_new_n24882__ = ys__n34712 & new_new_n24881__;
  assign new_new_n24883__ = ~new_new_n24880__ & ~new_new_n24882__;
  assign new_new_n24884__ = ~ys__n34708 & ys__n34710;
  assign new_new_n24885__ = ~ys__n34712 & new_new_n24884__;
  assign new_new_n24886__ = ys__n34708 & ~ys__n34710;
  assign new_new_n24887__ = ~ys__n34712 & new_new_n24886__;
  assign new_new_n24888__ = ~new_new_n24885__ & ~new_new_n24887__;
  assign new_new_n24889__ = new_new_n24883__ & new_new_n24888__;
  assign new_new_n24890__ = ys__n34716 & ys__n34718;
  assign new_new_n24891__ = ys__n34714 & ys__n34718;
  assign new_new_n24892__ = ~new_new_n24798__ & ~new_new_n24891__;
  assign new_new_n24893__ = ~new_new_n24890__ & new_new_n24892__;
  assign new_new_n24894__ = new_new_n24889__ & ~new_new_n24893__;
  assign new_new_n24895__ = ~new_new_n24889__ & new_new_n24893__;
  assign new_new_n24896__ = ~new_new_n24894__ & ~new_new_n24895__;
  assign new_new_n24897__ = ~new_new_n24808__ & ~new_new_n24812__;
  assign new_new_n24898__ = ~new_new_n24815__ & ~new_new_n24824__;
  assign new_new_n24899__ = ~new_new_n24897__ & ~new_new_n24898__;
  assign new_new_n24900__ = new_new_n24896__ & ~new_new_n24899__;
  assign new_new_n24901__ = ~new_new_n24896__ & new_new_n24899__;
  assign new_new_n24902__ = ~new_new_n24900__ & ~new_new_n24901__;
  assign new_new_n24903__ = new_new_n24220__ & ~new_new_n24902__;
  assign new_new_n24904__ = ~new_new_n24827__ & new_new_n24831__;
  assign new_new_n24905__ = new_new_n24902__ & new_new_n24904__;
  assign new_new_n24906__ = ~new_new_n24902__ & ~new_new_n24904__;
  assign new_new_n24907__ = ~new_new_n24905__ & ~new_new_n24906__;
  assign new_new_n24908__ = ~new_new_n24220__ & ~new_new_n24907__;
  assign new_new_n24909__ = ~new_new_n24903__ & ~new_new_n24908__;
  assign new_new_n24910__ = ~new_new_n24224__ & ~new_new_n24909__;
  assign new_new_n24911__ = ~new_new_n24827__ & new_new_n24838__;
  assign new_new_n24912__ = new_new_n24902__ & new_new_n24911__;
  assign new_new_n24913__ = ~new_new_n24902__ & ~new_new_n24911__;
  assign new_new_n24914__ = ~new_new_n24912__ & ~new_new_n24913__;
  assign new_new_n24915__ = new_new_n24224__ & ~new_new_n24914__;
  assign new_new_n24916__ = ~new_new_n24910__ & ~new_new_n24915__;
  assign new_new_n24917__ = ~new_new_n23480__ & ~new_new_n24916__;
  assign new_new_n24918__ = ~new_new_n24878__ & ~new_new_n24917__;
  assign new_new_n24919__ = ~new_new_n24230__ & ~new_new_n24918__;
  assign new_new_n24920__ = ~new_new_n23953__ & ~new_new_n24100__;
  assign new_new_n24921__ = ~new_new_n24106__ & ~new_new_n24920__;
  assign new_new_n24922__ = new_new_n24083__ & ~new_new_n24921__;
  assign new_new_n24923__ = ~new_new_n24083__ & new_new_n24921__;
  assign new_new_n24924__ = ~new_new_n24922__ & ~new_new_n24923__;
  assign new_new_n24925__ = new_new_n24230__ & ~new_new_n24924__;
  assign new_new_n24926__ = ~new_new_n24919__ & ~new_new_n24925__;
  assign new_new_n24927__ = new_new_n24237__ & ~new_new_n24926__;
  assign new_new_n24928__ = ys__n2535 & ~new_new_n24926__;
  assign new_new_n24929__ = ~new_new_n24927__ & ~new_new_n24928__;
  assign new_new_n24930__ = ~new_new_n12574__ & ~new_new_n24929__;
  assign new_new_n24931__ = ys__n47083 & new_new_n24250__;
  assign new_new_n24932__ = ys__n47019 & new_new_n24252__;
  assign new_new_n24933__ = ~new_new_n24931__ & ~new_new_n24932__;
  assign new_new_n24934__ = ~new_new_n24255__ & ~new_new_n24933__;
  assign new_new_n24935__ = new_new_n24249__ & new_new_n24934__;
  assign new_new_n24936__ = new_new_n24127__ & ~new_new_n24152__;
  assign new_new_n24937__ = ~new_new_n24155__ & new_new_n24209__;
  assign new_new_n24938__ = new_new_n24152__ & new_new_n24937__;
  assign new_new_n24939__ = ~new_new_n24152__ & ~new_new_n24937__;
  assign new_new_n24940__ = ~new_new_n24938__ & ~new_new_n24939__;
  assign new_new_n24941__ = ~new_new_n24127__ & ~new_new_n24940__;
  assign new_new_n24942__ = ~new_new_n24936__ & ~new_new_n24941__;
  assign new_new_n24943__ = ~new_new_n24249__ & ~new_new_n24942__;
  assign new_new_n24944__ = ~new_new_n24935__ & ~new_new_n24943__;
  assign new_new_n24945__ = new_new_n24265__ & ~new_new_n24944__;
  assign new_new_n24946__ = ys__n366 & ~new_new_n24265__;
  assign new_new_n24947__ = ~new_new_n24945__ & ~new_new_n24946__;
  assign new_new_n24948__ = new_new_n12574__ & ~new_new_n24947__;
  assign new_new_n24949__ = ~new_new_n24930__ & ~new_new_n24948__;
  assign new_new_n24950__ = ~ys__n1598 & ~new_new_n24949__;
  assign new_new_n24951__ = ys__n24768 & ys__n1598;
  assign ys__n24769 = new_new_n24950__ | new_new_n24951__;
  assign new_new_n24953__ = ys__n31031 & ys__n47036;
  assign new_new_n24954__ = new_new_n23480__ & new_new_n24953__;
  assign new_new_n24955__ = ys__n34702 & ys__n34704;
  assign new_new_n24956__ = ys__n34706 & new_new_n24955__;
  assign new_new_n24957__ = ~ys__n34702 & ~ys__n34704;
  assign new_new_n24958__ = ys__n34706 & new_new_n24957__;
  assign new_new_n24959__ = ~new_new_n24956__ & ~new_new_n24958__;
  assign new_new_n24960__ = ~ys__n34702 & ys__n34704;
  assign new_new_n24961__ = ~ys__n34706 & new_new_n24960__;
  assign new_new_n24962__ = ys__n34702 & ~ys__n34704;
  assign new_new_n24963__ = ~ys__n34706 & new_new_n24962__;
  assign new_new_n24964__ = ~new_new_n24961__ & ~new_new_n24963__;
  assign new_new_n24965__ = new_new_n24959__ & new_new_n24964__;
  assign new_new_n24966__ = ys__n34710 & ys__n34712;
  assign new_new_n24967__ = ys__n34708 & ys__n34712;
  assign new_new_n24968__ = ~new_new_n24879__ & ~new_new_n24967__;
  assign new_new_n24969__ = ~new_new_n24966__ & new_new_n24968__;
  assign new_new_n24970__ = new_new_n24965__ & ~new_new_n24969__;
  assign new_new_n24971__ = ~new_new_n24965__ & new_new_n24969__;
  assign new_new_n24972__ = ~new_new_n24970__ & ~new_new_n24971__;
  assign new_new_n24973__ = ~new_new_n24889__ & ~new_new_n24893__;
  assign new_new_n24974__ = ~new_new_n24896__ & new_new_n24897__;
  assign new_new_n24975__ = ~new_new_n24973__ & ~new_new_n24974__;
  assign new_new_n24976__ = ~new_new_n24815__ & ~new_new_n24896__;
  assign new_new_n24977__ = ~new_new_n24824__ & new_new_n24976__;
  assign new_new_n24978__ = new_new_n24975__ & ~new_new_n24977__;
  assign new_new_n24979__ = new_new_n24972__ & ~new_new_n24978__;
  assign new_new_n24980__ = ~new_new_n24972__ & new_new_n24978__;
  assign new_new_n24981__ = ~new_new_n24979__ & ~new_new_n24980__;
  assign new_new_n24982__ = new_new_n24220__ & ~new_new_n24981__;
  assign new_new_n24983__ = ~new_new_n24827__ & ~new_new_n24902__;
  assign new_new_n24984__ = new_new_n24831__ & new_new_n24983__;
  assign new_new_n24985__ = new_new_n24981__ & new_new_n24984__;
  assign new_new_n24986__ = ~new_new_n24981__ & ~new_new_n24984__;
  assign new_new_n24987__ = ~new_new_n24985__ & ~new_new_n24986__;
  assign new_new_n24988__ = ~new_new_n24220__ & ~new_new_n24987__;
  assign new_new_n24989__ = ~new_new_n24982__ & ~new_new_n24988__;
  assign new_new_n24990__ = ~new_new_n24224__ & ~new_new_n24989__;
  assign new_new_n24991__ = new_new_n24838__ & new_new_n24983__;
  assign new_new_n24992__ = new_new_n24981__ & new_new_n24991__;
  assign new_new_n24993__ = ~new_new_n24981__ & ~new_new_n24991__;
  assign new_new_n24994__ = ~new_new_n24992__ & ~new_new_n24993__;
  assign new_new_n24995__ = new_new_n24224__ & ~new_new_n24994__;
  assign new_new_n24996__ = ~new_new_n24990__ & ~new_new_n24995__;
  assign new_new_n24997__ = ~new_new_n23480__ & ~new_new_n24996__;
  assign new_new_n24998__ = ~new_new_n24954__ & ~new_new_n24997__;
  assign new_new_n24999__ = ~new_new_n24230__ & ~new_new_n24998__;
  assign new_new_n25000__ = ~new_new_n23953__ & new_new_n24101__;
  assign new_new_n25001__ = new_new_n24108__ & ~new_new_n25000__;
  assign new_new_n25002__ = new_new_n24064__ & ~new_new_n25001__;
  assign new_new_n25003__ = ~new_new_n24064__ & new_new_n25001__;
  assign new_new_n25004__ = ~new_new_n25002__ & ~new_new_n25003__;
  assign new_new_n25005__ = new_new_n24230__ & ~new_new_n25004__;
  assign new_new_n25006__ = ~new_new_n24999__ & ~new_new_n25005__;
  assign new_new_n25007__ = new_new_n24237__ & ~new_new_n25006__;
  assign new_new_n25008__ = ys__n2535 & ~new_new_n25006__;
  assign new_new_n25009__ = ~new_new_n25007__ & ~new_new_n25008__;
  assign new_new_n25010__ = ~new_new_n12574__ & ~new_new_n25009__;
  assign new_new_n25011__ = ys__n47084 & new_new_n24250__;
  assign new_new_n25012__ = ys__n47020 & new_new_n24252__;
  assign new_new_n25013__ = ~new_new_n25011__ & ~new_new_n25012__;
  assign new_new_n25014__ = ~new_new_n24255__ & ~new_new_n25013__;
  assign new_new_n25015__ = new_new_n24249__ & new_new_n25014__;
  assign new_new_n25016__ = new_new_n24127__ & ~new_new_n24147__;
  assign new_new_n25017__ = new_new_n24156__ & new_new_n24209__;
  assign new_new_n25018__ = new_new_n24147__ & new_new_n25017__;
  assign new_new_n25019__ = ~new_new_n24147__ & ~new_new_n25017__;
  assign new_new_n25020__ = ~new_new_n25018__ & ~new_new_n25019__;
  assign new_new_n25021__ = ~new_new_n24127__ & ~new_new_n25020__;
  assign new_new_n25022__ = ~new_new_n25016__ & ~new_new_n25021__;
  assign new_new_n25023__ = ~new_new_n24249__ & ~new_new_n25022__;
  assign new_new_n25024__ = ~new_new_n25015__ & ~new_new_n25023__;
  assign new_new_n25025__ = new_new_n24265__ & ~new_new_n25024__;
  assign new_new_n25026__ = ys__n368 & ~new_new_n24265__;
  assign new_new_n25027__ = ~new_new_n25025__ & ~new_new_n25026__;
  assign new_new_n25028__ = new_new_n12574__ & ~new_new_n25027__;
  assign new_new_n25029__ = ~new_new_n25010__ & ~new_new_n25028__;
  assign new_new_n25030__ = ~ys__n1598 & ~new_new_n25029__;
  assign new_new_n25031__ = ys__n24771 & ys__n1598;
  assign ys__n24772 = new_new_n25030__ | new_new_n25031__;
  assign new_new_n25033__ = ys__n31031 & ys__n47037;
  assign new_new_n25034__ = new_new_n23480__ & new_new_n25033__;
  assign new_new_n25035__ = ys__n34696 & ys__n34698;
  assign new_new_n25036__ = ys__n34700 & new_new_n25035__;
  assign new_new_n25037__ = ~ys__n34696 & ~ys__n34698;
  assign new_new_n25038__ = ys__n34700 & new_new_n25037__;
  assign new_new_n25039__ = ~new_new_n25036__ & ~new_new_n25038__;
  assign new_new_n25040__ = ~ys__n34696 & ys__n34698;
  assign new_new_n25041__ = ~ys__n34700 & new_new_n25040__;
  assign new_new_n25042__ = ys__n34696 & ~ys__n34698;
  assign new_new_n25043__ = ~ys__n34700 & new_new_n25042__;
  assign new_new_n25044__ = ~new_new_n25041__ & ~new_new_n25043__;
  assign new_new_n25045__ = new_new_n25039__ & new_new_n25044__;
  assign new_new_n25046__ = ys__n34704 & ys__n34706;
  assign new_new_n25047__ = ys__n34702 & ys__n34706;
  assign new_new_n25048__ = ~new_new_n24955__ & ~new_new_n25047__;
  assign new_new_n25049__ = ~new_new_n25046__ & new_new_n25048__;
  assign new_new_n25050__ = new_new_n25045__ & ~new_new_n25049__;
  assign new_new_n25051__ = ~new_new_n25045__ & new_new_n25049__;
  assign new_new_n25052__ = ~new_new_n25050__ & ~new_new_n25051__;
  assign new_new_n25053__ = ~new_new_n24965__ & ~new_new_n24969__;
  assign new_new_n25054__ = ~new_new_n24972__ & ~new_new_n24978__;
  assign new_new_n25055__ = ~new_new_n25053__ & ~new_new_n25054__;
  assign new_new_n25056__ = new_new_n25052__ & ~new_new_n25055__;
  assign new_new_n25057__ = ~new_new_n25052__ & new_new_n25055__;
  assign new_new_n25058__ = ~new_new_n25056__ & ~new_new_n25057__;
  assign new_new_n25059__ = new_new_n24220__ & ~new_new_n25058__;
  assign new_new_n25060__ = ~new_new_n24981__ & new_new_n24984__;
  assign new_new_n25061__ = new_new_n25058__ & new_new_n25060__;
  assign new_new_n25062__ = ~new_new_n25058__ & ~new_new_n25060__;
  assign new_new_n25063__ = ~new_new_n25061__ & ~new_new_n25062__;
  assign new_new_n25064__ = ~new_new_n24220__ & ~new_new_n25063__;
  assign new_new_n25065__ = ~new_new_n25059__ & ~new_new_n25064__;
  assign new_new_n25066__ = ~new_new_n24224__ & ~new_new_n25065__;
  assign new_new_n25067__ = ~new_new_n24981__ & new_new_n24991__;
  assign new_new_n25068__ = new_new_n25058__ & new_new_n25067__;
  assign new_new_n25069__ = ~new_new_n25058__ & ~new_new_n25067__;
  assign new_new_n25070__ = ~new_new_n25068__ & ~new_new_n25069__;
  assign new_new_n25071__ = new_new_n24224__ & ~new_new_n25070__;
  assign new_new_n25072__ = ~new_new_n25066__ & ~new_new_n25071__;
  assign new_new_n25073__ = ~new_new_n23480__ & ~new_new_n25072__;
  assign new_new_n25074__ = ~new_new_n25034__ & ~new_new_n25073__;
  assign new_new_n25075__ = ~new_new_n24230__ & ~new_new_n25074__;
  assign new_new_n25076__ = ~new_new_n24064__ & ~new_new_n25001__;
  assign new_new_n25077__ = ~new_new_n24111__ & ~new_new_n25076__;
  assign new_new_n25078__ = new_new_n24046__ & ~new_new_n25077__;
  assign new_new_n25079__ = ~new_new_n24046__ & new_new_n25077__;
  assign new_new_n25080__ = ~new_new_n25078__ & ~new_new_n25079__;
  assign new_new_n25081__ = new_new_n24230__ & ~new_new_n25080__;
  assign new_new_n25082__ = ~new_new_n25075__ & ~new_new_n25081__;
  assign new_new_n25083__ = new_new_n24237__ & ~new_new_n25082__;
  assign new_new_n25084__ = ys__n2535 & ~new_new_n25082__;
  assign new_new_n25085__ = ~new_new_n25083__ & ~new_new_n25084__;
  assign new_new_n25086__ = ~new_new_n12574__ & ~new_new_n25085__;
  assign new_new_n25087__ = ys__n47085 & new_new_n24250__;
  assign new_new_n25088__ = ys__n47021 & new_new_n24252__;
  assign new_new_n25089__ = ~new_new_n25087__ & ~new_new_n25088__;
  assign new_new_n25090__ = ~new_new_n24255__ & ~new_new_n25089__;
  assign new_new_n25091__ = new_new_n24249__ & new_new_n25090__;
  assign new_new_n25092__ = new_new_n24127__ & ~new_new_n24144__;
  assign new_new_n25093__ = ~new_new_n24147__ & new_new_n25017__;
  assign new_new_n25094__ = new_new_n24144__ & new_new_n25093__;
  assign new_new_n25095__ = ~new_new_n24144__ & ~new_new_n25093__;
  assign new_new_n25096__ = ~new_new_n25094__ & ~new_new_n25095__;
  assign new_new_n25097__ = ~new_new_n24127__ & ~new_new_n25096__;
  assign new_new_n25098__ = ~new_new_n25092__ & ~new_new_n25097__;
  assign new_new_n25099__ = ~new_new_n24249__ & ~new_new_n25098__;
  assign new_new_n25100__ = ~new_new_n25091__ & ~new_new_n25099__;
  assign new_new_n25101__ = new_new_n24265__ & ~new_new_n25100__;
  assign new_new_n25102__ = ys__n364 & ~new_new_n24265__;
  assign new_new_n25103__ = ~new_new_n25101__ & ~new_new_n25102__;
  assign new_new_n25104__ = new_new_n12574__ & ~new_new_n25103__;
  assign new_new_n25105__ = ~new_new_n25086__ & ~new_new_n25104__;
  assign new_new_n25106__ = ~ys__n1598 & ~new_new_n25105__;
  assign new_new_n25107__ = ys__n24774 & ys__n1598;
  assign ys__n24775 = new_new_n25106__ | new_new_n25107__;
  assign new_new_n25109__ = ys__n31031 & ys__n47038;
  assign new_new_n25110__ = new_new_n23480__ & new_new_n25109__;
  assign new_new_n25111__ = ys__n34690 & ys__n34692;
  assign new_new_n25112__ = ys__n34694 & new_new_n25111__;
  assign new_new_n25113__ = ~ys__n34690 & ~ys__n34692;
  assign new_new_n25114__ = ys__n34694 & new_new_n25113__;
  assign new_new_n25115__ = ~new_new_n25112__ & ~new_new_n25114__;
  assign new_new_n25116__ = ~ys__n34690 & ys__n34692;
  assign new_new_n25117__ = ~ys__n34694 & new_new_n25116__;
  assign new_new_n25118__ = ys__n34690 & ~ys__n34692;
  assign new_new_n25119__ = ~ys__n34694 & new_new_n25118__;
  assign new_new_n25120__ = ~new_new_n25117__ & ~new_new_n25119__;
  assign new_new_n25121__ = new_new_n25115__ & new_new_n25120__;
  assign new_new_n25122__ = ys__n34698 & ys__n34700;
  assign new_new_n25123__ = ys__n34696 & ys__n34700;
  assign new_new_n25124__ = ~new_new_n25035__ & ~new_new_n25123__;
  assign new_new_n25125__ = ~new_new_n25122__ & new_new_n25124__;
  assign new_new_n25126__ = new_new_n25121__ & ~new_new_n25125__;
  assign new_new_n25127__ = ~new_new_n25121__ & new_new_n25125__;
  assign new_new_n25128__ = ~new_new_n25126__ & ~new_new_n25127__;
  assign new_new_n25129__ = ~new_new_n24972__ & ~new_new_n25052__;
  assign new_new_n25130__ = new_new_n24976__ & new_new_n25129__;
  assign new_new_n25131__ = ~new_new_n24824__ & new_new_n25130__;
  assign new_new_n25132__ = ~new_new_n24975__ & new_new_n25129__;
  assign new_new_n25133__ = ~new_new_n25045__ & ~new_new_n25049__;
  assign new_new_n25134__ = ~new_new_n25052__ & new_new_n25053__;
  assign new_new_n25135__ = ~new_new_n25133__ & ~new_new_n25134__;
  assign new_new_n25136__ = ~new_new_n25132__ & new_new_n25135__;
  assign new_new_n25137__ = ~new_new_n25131__ & new_new_n25136__;
  assign new_new_n25138__ = new_new_n25128__ & ~new_new_n25137__;
  assign new_new_n25139__ = ~new_new_n25128__ & new_new_n25137__;
  assign new_new_n25140__ = ~new_new_n25138__ & ~new_new_n25139__;
  assign new_new_n25141__ = new_new_n24220__ & ~new_new_n25140__;
  assign new_new_n25142__ = ~new_new_n24981__ & new_new_n24983__;
  assign new_new_n25143__ = ~new_new_n25058__ & new_new_n25142__;
  assign new_new_n25144__ = new_new_n24831__ & new_new_n25143__;
  assign new_new_n25145__ = new_new_n25140__ & new_new_n25144__;
  assign new_new_n25146__ = ~new_new_n25140__ & ~new_new_n25144__;
  assign new_new_n25147__ = ~new_new_n25145__ & ~new_new_n25146__;
  assign new_new_n25148__ = ~new_new_n24220__ & ~new_new_n25147__;
  assign new_new_n25149__ = ~new_new_n25141__ & ~new_new_n25148__;
  assign new_new_n25150__ = ~new_new_n24224__ & ~new_new_n25149__;
  assign new_new_n25151__ = new_new_n24838__ & new_new_n25143__;
  assign new_new_n25152__ = new_new_n25140__ & new_new_n25151__;
  assign new_new_n25153__ = ~new_new_n25140__ & ~new_new_n25151__;
  assign new_new_n25154__ = ~new_new_n25152__ & ~new_new_n25153__;
  assign new_new_n25155__ = new_new_n24224__ & ~new_new_n25154__;
  assign new_new_n25156__ = ~new_new_n25150__ & ~new_new_n25155__;
  assign new_new_n25157__ = ~new_new_n23480__ & ~new_new_n25156__;
  assign new_new_n25158__ = ~new_new_n25110__ & ~new_new_n25157__;
  assign new_new_n25159__ = ~new_new_n24230__ & ~new_new_n25158__;
  assign new_new_n25160__ = ~new_new_n23953__ & new_new_n24102__;
  assign new_new_n25161__ = new_new_n24114__ & ~new_new_n25160__;
  assign new_new_n25162__ = new_new_n24026__ & ~new_new_n25161__;
  assign new_new_n25163__ = ~new_new_n24026__ & new_new_n25161__;
  assign new_new_n25164__ = ~new_new_n25162__ & ~new_new_n25163__;
  assign new_new_n25165__ = new_new_n24230__ & ~new_new_n25164__;
  assign new_new_n25166__ = ~new_new_n25159__ & ~new_new_n25165__;
  assign new_new_n25167__ = new_new_n24237__ & ~new_new_n25166__;
  assign new_new_n25168__ = ys__n2535 & ~new_new_n25166__;
  assign new_new_n25169__ = ~new_new_n25167__ & ~new_new_n25168__;
  assign new_new_n25170__ = ~new_new_n12574__ & ~new_new_n25169__;
  assign new_new_n25171__ = ys__n47086 & new_new_n24250__;
  assign new_new_n25172__ = ys__n47022 & new_new_n24252__;
  assign new_new_n25173__ = ~new_new_n25171__ & ~new_new_n25172__;
  assign new_new_n25174__ = ~new_new_n24255__ & ~new_new_n25173__;
  assign new_new_n25175__ = new_new_n24249__ & new_new_n25174__;
  assign new_new_n25176__ = new_new_n24127__ & ~new_new_n24166__;
  assign new_new_n25177__ = new_new_n24158__ & new_new_n24209__;
  assign new_new_n25178__ = new_new_n24166__ & new_new_n25177__;
  assign new_new_n25179__ = ~new_new_n24166__ & ~new_new_n25177__;
  assign new_new_n25180__ = ~new_new_n25178__ & ~new_new_n25179__;
  assign new_new_n25181__ = ~new_new_n24127__ & ~new_new_n25180__;
  assign new_new_n25182__ = ~new_new_n25176__ & ~new_new_n25181__;
  assign new_new_n25183__ = ~new_new_n24249__ & ~new_new_n25182__;
  assign new_new_n25184__ = ~new_new_n25175__ & ~new_new_n25183__;
  assign new_new_n25185__ = new_new_n24265__ & ~new_new_n25184__;
  assign new_new_n25186__ = ys__n370 & ~new_new_n24265__;
  assign new_new_n25187__ = ~new_new_n25185__ & ~new_new_n25186__;
  assign new_new_n25188__ = new_new_n12574__ & ~new_new_n25187__;
  assign new_new_n25189__ = ~new_new_n25170__ & ~new_new_n25188__;
  assign new_new_n25190__ = ~ys__n1598 & ~new_new_n25189__;
  assign new_new_n25191__ = ys__n24777 & ys__n1598;
  assign ys__n24778 = new_new_n25190__ | new_new_n25191__;
  assign new_new_n25193__ = ys__n31031 & ys__n47039;
  assign new_new_n25194__ = new_new_n23480__ & new_new_n25193__;
  assign new_new_n25195__ = ys__n34684 & ys__n34686;
  assign new_new_n25196__ = ys__n34688 & new_new_n25195__;
  assign new_new_n25197__ = ~ys__n34684 & ~ys__n34686;
  assign new_new_n25198__ = ys__n34688 & new_new_n25197__;
  assign new_new_n25199__ = ~new_new_n25196__ & ~new_new_n25198__;
  assign new_new_n25200__ = ~ys__n34684 & ys__n34686;
  assign new_new_n25201__ = ~ys__n34688 & new_new_n25200__;
  assign new_new_n25202__ = ys__n34684 & ~ys__n34686;
  assign new_new_n25203__ = ~ys__n34688 & new_new_n25202__;
  assign new_new_n25204__ = ~new_new_n25201__ & ~new_new_n25203__;
  assign new_new_n25205__ = new_new_n25199__ & new_new_n25204__;
  assign new_new_n25206__ = ys__n34692 & ys__n34694;
  assign new_new_n25207__ = ys__n34690 & ys__n34694;
  assign new_new_n25208__ = ~new_new_n25111__ & ~new_new_n25207__;
  assign new_new_n25209__ = ~new_new_n25206__ & new_new_n25208__;
  assign new_new_n25210__ = new_new_n25205__ & ~new_new_n25209__;
  assign new_new_n25211__ = ~new_new_n25205__ & new_new_n25209__;
  assign new_new_n25212__ = ~new_new_n25210__ & ~new_new_n25211__;
  assign new_new_n25213__ = ~new_new_n25121__ & ~new_new_n25125__;
  assign new_new_n25214__ = ~new_new_n25128__ & ~new_new_n25137__;
  assign new_new_n25215__ = ~new_new_n25213__ & ~new_new_n25214__;
  assign new_new_n25216__ = new_new_n25212__ & ~new_new_n25215__;
  assign new_new_n25217__ = ~new_new_n25212__ & new_new_n25215__;
  assign new_new_n25218__ = ~new_new_n25216__ & ~new_new_n25217__;
  assign new_new_n25219__ = new_new_n24220__ & ~new_new_n25218__;
  assign new_new_n25220__ = ~new_new_n25140__ & new_new_n25144__;
  assign new_new_n25221__ = new_new_n25218__ & new_new_n25220__;
  assign new_new_n25222__ = ~new_new_n25218__ & ~new_new_n25220__;
  assign new_new_n25223__ = ~new_new_n25221__ & ~new_new_n25222__;
  assign new_new_n25224__ = ~new_new_n24220__ & ~new_new_n25223__;
  assign new_new_n25225__ = ~new_new_n25219__ & ~new_new_n25224__;
  assign new_new_n25226__ = ~new_new_n24224__ & ~new_new_n25225__;
  assign new_new_n25227__ = ~new_new_n25140__ & new_new_n25151__;
  assign new_new_n25228__ = new_new_n25218__ & new_new_n25227__;
  assign new_new_n25229__ = ~new_new_n25218__ & ~new_new_n25227__;
  assign new_new_n25230__ = ~new_new_n25228__ & ~new_new_n25229__;
  assign new_new_n25231__ = new_new_n24224__ & ~new_new_n25230__;
  assign new_new_n25232__ = ~new_new_n25226__ & ~new_new_n25231__;
  assign new_new_n25233__ = ~new_new_n23480__ & ~new_new_n25232__;
  assign new_new_n25234__ = ~new_new_n25194__ & ~new_new_n25233__;
  assign new_new_n25235__ = ~new_new_n24230__ & ~new_new_n25234__;
  assign new_new_n25236__ = ~new_new_n24026__ & ~new_new_n25161__;
  assign new_new_n25237__ = ~new_new_n24117__ & ~new_new_n25236__;
  assign new_new_n25238__ = new_new_n24008__ & ~new_new_n25237__;
  assign new_new_n25239__ = ~new_new_n24008__ & new_new_n25237__;
  assign new_new_n25240__ = ~new_new_n25238__ & ~new_new_n25239__;
  assign new_new_n25241__ = new_new_n24230__ & ~new_new_n25240__;
  assign new_new_n25242__ = ~new_new_n25235__ & ~new_new_n25241__;
  assign new_new_n25243__ = new_new_n24237__ & ~new_new_n25242__;
  assign new_new_n25244__ = ys__n2535 & ~new_new_n25242__;
  assign new_new_n25245__ = ~new_new_n25243__ & ~new_new_n25244__;
  assign new_new_n25246__ = ~new_new_n12574__ & ~new_new_n25245__;
  assign new_new_n25247__ = ys__n47087 & new_new_n24250__;
  assign new_new_n25248__ = ys__n47023 & new_new_n24252__;
  assign new_new_n25249__ = ~new_new_n25247__ & ~new_new_n25248__;
  assign new_new_n25250__ = ~new_new_n24255__ & ~new_new_n25249__;
  assign new_new_n25251__ = new_new_n24249__ & new_new_n25250__;
  assign new_new_n25252__ = new_new_n24127__ & ~new_new_n24163__;
  assign new_new_n25253__ = ~new_new_n24166__ & new_new_n25177__;
  assign new_new_n25254__ = new_new_n24163__ & new_new_n25253__;
  assign new_new_n25255__ = ~new_new_n24163__ & ~new_new_n25253__;
  assign new_new_n25256__ = ~new_new_n25254__ & ~new_new_n25255__;
  assign new_new_n25257__ = ~new_new_n24127__ & ~new_new_n25256__;
  assign new_new_n25258__ = ~new_new_n25252__ & ~new_new_n25257__;
  assign new_new_n25259__ = ~new_new_n24249__ & ~new_new_n25258__;
  assign new_new_n25260__ = ~new_new_n25251__ & ~new_new_n25259__;
  assign new_new_n25261__ = new_new_n24265__ & ~new_new_n25260__;
  assign new_new_n25262__ = ys__n360 & ~new_new_n24265__;
  assign new_new_n25263__ = ~new_new_n25261__ & ~new_new_n25262__;
  assign new_new_n25264__ = new_new_n12574__ & ~new_new_n25263__;
  assign new_new_n25265__ = ~new_new_n25246__ & ~new_new_n25264__;
  assign new_new_n25266__ = ~ys__n1598 & ~new_new_n25265__;
  assign new_new_n25267__ = ys__n24780 & ys__n1598;
  assign ys__n24781 = new_new_n25266__ | new_new_n25267__;
  assign new_new_n25269__ = ys__n31031 & ys__n47040;
  assign new_new_n25270__ = new_new_n23480__ & new_new_n25269__;
  assign new_new_n25271__ = ys__n34678 & ys__n34680;
  assign new_new_n25272__ = ys__n34682 & new_new_n25271__;
  assign new_new_n25273__ = ~ys__n34678 & ~ys__n34680;
  assign new_new_n25274__ = ys__n34682 & new_new_n25273__;
  assign new_new_n25275__ = ~new_new_n25272__ & ~new_new_n25274__;
  assign new_new_n25276__ = ~ys__n34678 & ys__n34680;
  assign new_new_n25277__ = ~ys__n34682 & new_new_n25276__;
  assign new_new_n25278__ = ys__n34678 & ~ys__n34680;
  assign new_new_n25279__ = ~ys__n34682 & new_new_n25278__;
  assign new_new_n25280__ = ~new_new_n25277__ & ~new_new_n25279__;
  assign new_new_n25281__ = new_new_n25275__ & new_new_n25280__;
  assign new_new_n25282__ = ys__n34686 & ys__n34688;
  assign new_new_n25283__ = ys__n34684 & ys__n34688;
  assign new_new_n25284__ = ~new_new_n25195__ & ~new_new_n25283__;
  assign new_new_n25285__ = ~new_new_n25282__ & new_new_n25284__;
  assign new_new_n25286__ = new_new_n25281__ & ~new_new_n25285__;
  assign new_new_n25287__ = ~new_new_n25281__ & new_new_n25285__;
  assign new_new_n25288__ = ~new_new_n25286__ & ~new_new_n25287__;
  assign new_new_n25289__ = ~new_new_n25128__ & ~new_new_n25212__;
  assign new_new_n25290__ = ~new_new_n25137__ & new_new_n25289__;
  assign new_new_n25291__ = ~new_new_n25205__ & ~new_new_n25209__;
  assign new_new_n25292__ = ~new_new_n25212__ & new_new_n25213__;
  assign new_new_n25293__ = ~new_new_n25291__ & ~new_new_n25292__;
  assign new_new_n25294__ = ~new_new_n25290__ & new_new_n25293__;
  assign new_new_n25295__ = new_new_n25288__ & ~new_new_n25294__;
  assign new_new_n25296__ = ~new_new_n25288__ & new_new_n25294__;
  assign new_new_n25297__ = ~new_new_n25295__ & ~new_new_n25296__;
  assign new_new_n25298__ = new_new_n24220__ & ~new_new_n25297__;
  assign new_new_n25299__ = ~new_new_n25140__ & ~new_new_n25218__;
  assign new_new_n25300__ = new_new_n25144__ & new_new_n25299__;
  assign new_new_n25301__ = new_new_n25297__ & new_new_n25300__;
  assign new_new_n25302__ = ~new_new_n25297__ & ~new_new_n25300__;
  assign new_new_n25303__ = ~new_new_n25301__ & ~new_new_n25302__;
  assign new_new_n25304__ = ~new_new_n24220__ & ~new_new_n25303__;
  assign new_new_n25305__ = ~new_new_n25298__ & ~new_new_n25304__;
  assign new_new_n25306__ = ~new_new_n24224__ & ~new_new_n25305__;
  assign new_new_n25307__ = new_new_n25151__ & new_new_n25299__;
  assign new_new_n25308__ = new_new_n25297__ & new_new_n25307__;
  assign new_new_n25309__ = ~new_new_n25297__ & ~new_new_n25307__;
  assign new_new_n25310__ = ~new_new_n25308__ & ~new_new_n25309__;
  assign new_new_n25311__ = new_new_n24224__ & ~new_new_n25310__;
  assign new_new_n25312__ = ~new_new_n25306__ & ~new_new_n25311__;
  assign new_new_n25313__ = ~new_new_n23480__ & ~new_new_n25312__;
  assign new_new_n25314__ = ~new_new_n25270__ & ~new_new_n25313__;
  assign new_new_n25315__ = ~new_new_n24230__ & ~new_new_n25314__;
  assign new_new_n25316__ = new_new_n24027__ & ~new_new_n25161__;
  assign new_new_n25317__ = new_new_n24119__ & ~new_new_n25316__;
  assign new_new_n25318__ = new_new_n23989__ & ~new_new_n25317__;
  assign new_new_n25319__ = ~new_new_n23989__ & new_new_n25317__;
  assign new_new_n25320__ = ~new_new_n25318__ & ~new_new_n25319__;
  assign new_new_n25321__ = new_new_n24230__ & ~new_new_n25320__;
  assign new_new_n25322__ = ~new_new_n25315__ & ~new_new_n25321__;
  assign new_new_n25323__ = new_new_n24237__ & ~new_new_n25322__;
  assign new_new_n25324__ = ys__n2535 & ~new_new_n25322__;
  assign new_new_n25325__ = ~new_new_n25323__ & ~new_new_n25324__;
  assign new_new_n25326__ = ~new_new_n12574__ & ~new_new_n25325__;
  assign new_new_n25327__ = ys__n47088 & new_new_n24250__;
  assign new_new_n25328__ = ys__n47024 & new_new_n24252__;
  assign new_new_n25329__ = ~new_new_n25327__ & ~new_new_n25328__;
  assign new_new_n25330__ = ~new_new_n24255__ & ~new_new_n25329__;
  assign new_new_n25331__ = new_new_n24249__ & new_new_n25330__;
  assign new_new_n25332__ = new_new_n24127__ & ~new_new_n24170__;
  assign new_new_n25333__ = new_new_n24167__ & new_new_n25177__;
  assign new_new_n25334__ = new_new_n24170__ & new_new_n25333__;
  assign new_new_n25335__ = ~new_new_n24170__ & ~new_new_n25333__;
  assign new_new_n25336__ = ~new_new_n25334__ & ~new_new_n25335__;
  assign new_new_n25337__ = ~new_new_n24127__ & ~new_new_n25336__;
  assign new_new_n25338__ = ~new_new_n25332__ & ~new_new_n25337__;
  assign new_new_n25339__ = ~new_new_n24249__ & ~new_new_n25338__;
  assign new_new_n25340__ = ~new_new_n25331__ & ~new_new_n25339__;
  assign new_new_n25341__ = new_new_n24265__ & ~new_new_n25340__;
  assign new_new_n25342__ = ys__n362 & ~new_new_n24265__;
  assign new_new_n25343__ = ~new_new_n25341__ & ~new_new_n25342__;
  assign new_new_n25344__ = new_new_n12574__ & ~new_new_n25343__;
  assign new_new_n25345__ = ~new_new_n25326__ & ~new_new_n25344__;
  assign new_new_n25346__ = ~ys__n1598 & ~new_new_n25345__;
  assign new_new_n25347__ = ys__n24783 & ys__n1598;
  assign ys__n24784 = new_new_n25346__ | new_new_n25347__;
  assign new_new_n25349__ = ys__n31031 & ys__n47041;
  assign new_new_n25350__ = new_new_n23480__ & new_new_n25349__;
  assign new_new_n25351__ = ~ys__n34674 & ys__n34676;
  assign new_new_n25352__ = ys__n34674 & ~ys__n34676;
  assign new_new_n25353__ = ~new_new_n25351__ & ~new_new_n25352__;
  assign new_new_n25354__ = ys__n34680 & ys__n34682;
  assign new_new_n25355__ = ys__n34678 & ys__n34682;
  assign new_new_n25356__ = ~new_new_n25271__ & ~new_new_n25355__;
  assign new_new_n25357__ = ~new_new_n25354__ & new_new_n25356__;
  assign new_new_n25358__ = new_new_n25353__ & ~new_new_n25357__;
  assign new_new_n25359__ = ~new_new_n25353__ & new_new_n25357__;
  assign new_new_n25360__ = ~new_new_n25358__ & ~new_new_n25359__;
  assign new_new_n25361__ = ~ys__n48324 & ~new_new_n25360__;
  assign new_new_n25362__ = ys__n48324 & new_new_n25360__;
  assign new_new_n25363__ = ~new_new_n25361__ & ~new_new_n25362__;
  assign new_new_n25364__ = ~new_new_n25281__ & ~new_new_n25285__;
  assign new_new_n25365__ = ~new_new_n25288__ & ~new_new_n25294__;
  assign new_new_n25366__ = ~new_new_n25364__ & ~new_new_n25365__;
  assign new_new_n25367__ = new_new_n24220__ & ~new_new_n25366__;
  assign new_new_n25368__ = ~new_new_n25297__ & new_new_n25300__;
  assign new_new_n25369__ = new_new_n25366__ & new_new_n25368__;
  assign new_new_n25370__ = ~new_new_n25366__ & ~new_new_n25368__;
  assign new_new_n25371__ = ~new_new_n25369__ & ~new_new_n25370__;
  assign new_new_n25372__ = ~new_new_n24220__ & ~new_new_n25371__;
  assign new_new_n25373__ = ~new_new_n25367__ & ~new_new_n25372__;
  assign new_new_n25374__ = ~new_new_n24224__ & ~new_new_n25373__;
  assign new_new_n25375__ = ~new_new_n25297__ & new_new_n25307__;
  assign new_new_n25376__ = new_new_n25366__ & new_new_n25375__;
  assign new_new_n25377__ = ~new_new_n25366__ & ~new_new_n25375__;
  assign new_new_n25378__ = ~new_new_n25376__ & ~new_new_n25377__;
  assign new_new_n25379__ = new_new_n24224__ & ~new_new_n25378__;
  assign new_new_n25380__ = ~new_new_n25374__ & ~new_new_n25379__;
  assign new_new_n25381__ = ~new_new_n25363__ & new_new_n25380__;
  assign new_new_n25382__ = ~ys__n48324 & new_new_n25360__;
  assign new_new_n25383__ = ys__n48324 & ~new_new_n25360__;
  assign new_new_n25384__ = ~new_new_n25382__ & ~new_new_n25383__;
  assign new_new_n25385__ = ~new_new_n25380__ & ~new_new_n25384__;
  assign new_new_n25386__ = ~new_new_n25381__ & ~new_new_n25385__;
  assign new_new_n25387__ = ~new_new_n23480__ & ~new_new_n25386__;
  assign new_new_n25388__ = ~new_new_n25350__ & ~new_new_n25387__;
  assign new_new_n25389__ = ~new_new_n24230__ & ~new_new_n25388__;
  assign new_new_n25390__ = ~new_new_n23989__ & ~new_new_n25317__;
  assign new_new_n25391__ = ~new_new_n24122__ & ~new_new_n25390__;
  assign new_new_n25392__ = new_new_n23971__ & ~new_new_n25391__;
  assign new_new_n25393__ = ~new_new_n23971__ & new_new_n25391__;
  assign new_new_n25394__ = ~new_new_n25392__ & ~new_new_n25393__;
  assign new_new_n25395__ = new_new_n24230__ & ~new_new_n25394__;
  assign new_new_n25396__ = ~new_new_n25389__ & ~new_new_n25395__;
  assign new_new_n25397__ = new_new_n24237__ & ~new_new_n25396__;
  assign new_new_n25398__ = ys__n2535 & ~new_new_n25396__;
  assign new_new_n25399__ = ~new_new_n25397__ & ~new_new_n25398__;
  assign new_new_n25400__ = ~new_new_n12574__ & ~new_new_n25399__;
  assign new_new_n25401__ = ys__n47089 & new_new_n24250__;
  assign new_new_n25402__ = ys__n47025 & new_new_n24252__;
  assign new_new_n25403__ = ~new_new_n25401__ & ~new_new_n25402__;
  assign new_new_n25404__ = ~new_new_n24255__ & ~new_new_n25403__;
  assign new_new_n25405__ = new_new_n24249__ & new_new_n25404__;
  assign new_new_n25406__ = new_new_n24127__ & ~new_new_n24137__;
  assign new_new_n25407__ = ~new_new_n24170__ & new_new_n25333__;
  assign new_new_n25408__ = new_new_n24137__ & new_new_n25407__;
  assign new_new_n25409__ = ~new_new_n24137__ & ~new_new_n25407__;
  assign new_new_n25410__ = ~new_new_n25408__ & ~new_new_n25409__;
  assign new_new_n25411__ = ~new_new_n24127__ & ~new_new_n25410__;
  assign new_new_n25412__ = ~new_new_n25406__ & ~new_new_n25411__;
  assign new_new_n25413__ = ~new_new_n24249__ & ~new_new_n25412__;
  assign new_new_n25414__ = ~new_new_n25405__ & ~new_new_n25413__;
  assign new_new_n25415__ = new_new_n24265__ & ~new_new_n25414__;
  assign new_new_n25416__ = ys__n358 & ~new_new_n24265__;
  assign new_new_n25417__ = ~new_new_n25415__ & ~new_new_n25416__;
  assign new_new_n25418__ = new_new_n12574__ & ~new_new_n25417__;
  assign new_new_n25419__ = ~new_new_n25400__ & ~new_new_n25418__;
  assign new_new_n25420__ = ~ys__n1598 & ~new_new_n25419__;
  assign new_new_n25421__ = ys__n24786 & ys__n1598;
  assign ys__n24787 = new_new_n25420__ | new_new_n25421__;
  assign new_new_n25423__ = ~ys__n34670 & ys__n34672;
  assign new_new_n25424__ = ys__n34670 & ~ys__n34672;
  assign new_new_n25425__ = ~new_new_n25423__ & ~new_new_n25424__;
  assign new_new_n25426__ = ys__n34674 & ys__n34676;
  assign new_new_n25427__ = new_new_n25425__ & new_new_n25426__;
  assign new_new_n25428__ = ~new_new_n25425__ & ~new_new_n25426__;
  assign new_new_n25429__ = ~new_new_n25427__ & ~new_new_n25428__;
  assign new_new_n25430__ = ~new_new_n25353__ & ~new_new_n25357__;
  assign new_new_n25431__ = new_new_n25429__ & new_new_n25430__;
  assign new_new_n25432__ = ~new_new_n25429__ & ~new_new_n25430__;
  assign new_new_n25433__ = ~new_new_n25431__ & ~new_new_n25432__;
  assign new_new_n25434__ = ~ys__n48325 & ~new_new_n25433__;
  assign new_new_n25435__ = ys__n48325 & new_new_n25433__;
  assign new_new_n25436__ = ~new_new_n25434__ & ~new_new_n25435__;
  assign new_new_n25437__ = new_new_n25383__ & new_new_n25436__;
  assign new_new_n25438__ = ~new_new_n25383__ & ~new_new_n25436__;
  assign new_new_n25439__ = ~new_new_n25437__ & ~new_new_n25438__;
  assign new_new_n25440__ = new_new_n25380__ & ~new_new_n25439__;
  assign new_new_n25441__ = ~new_new_n25360__ & new_new_n25433__;
  assign new_new_n25442__ = new_new_n25360__ & ~new_new_n25433__;
  assign new_new_n25443__ = ~new_new_n25441__ & ~new_new_n25442__;
  assign new_new_n25444__ = ~ys__n48325 & ~new_new_n25443__;
  assign new_new_n25445__ = ys__n48325 & new_new_n25443__;
  assign new_new_n25446__ = ~new_new_n25444__ & ~new_new_n25445__;
  assign new_new_n25447__ = new_new_n25362__ & new_new_n25446__;
  assign new_new_n25448__ = ~new_new_n25362__ & ~new_new_n25446__;
  assign new_new_n25449__ = ~new_new_n25447__ & ~new_new_n25448__;
  assign new_new_n25450__ = ~new_new_n25380__ & ~new_new_n25449__;
  assign new_new_n25451__ = ~new_new_n25440__ & ~new_new_n25450__;
  assign new_new_n25452__ = ys__n2779 & ~new_new_n25451__;
  assign new_new_n25453__ = ~ys__n34666 & ys__n34668;
  assign new_new_n25454__ = ys__n34666 & ~ys__n34668;
  assign new_new_n25455__ = ~new_new_n25453__ & ~new_new_n25454__;
  assign new_new_n25456__ = ys__n34670 & ys__n34672;
  assign new_new_n25457__ = new_new_n25455__ & new_new_n25456__;
  assign new_new_n25458__ = ~new_new_n25455__ & ~new_new_n25456__;
  assign new_new_n25459__ = ~new_new_n25457__ & ~new_new_n25458__;
  assign new_new_n25460__ = ~new_new_n25425__ & new_new_n25426__;
  assign new_new_n25461__ = ~new_new_n25429__ & new_new_n25430__;
  assign new_new_n25462__ = ~new_new_n25460__ & ~new_new_n25461__;
  assign new_new_n25463__ = new_new_n25459__ & ~new_new_n25462__;
  assign new_new_n25464__ = ~new_new_n25459__ & new_new_n25462__;
  assign new_new_n25465__ = ~new_new_n25463__ & ~new_new_n25464__;
  assign new_new_n25466__ = ~ys__n48327 & ~new_new_n25465__;
  assign new_new_n25467__ = ys__n48327 & new_new_n25465__;
  assign new_new_n25468__ = ~new_new_n25466__ & ~new_new_n25467__;
  assign new_new_n25469__ = ys__n48325 & ~new_new_n25433__;
  assign new_new_n25470__ = new_new_n25383__ & ~new_new_n25436__;
  assign new_new_n25471__ = ~new_new_n25469__ & ~new_new_n25470__;
  assign new_new_n25472__ = new_new_n25468__ & ~new_new_n25471__;
  assign new_new_n25473__ = ~new_new_n25468__ & new_new_n25471__;
  assign new_new_n25474__ = ~new_new_n25472__ & ~new_new_n25473__;
  assign new_new_n25475__ = new_new_n25380__ & ~new_new_n25474__;
  assign new_new_n25476__ = ~new_new_n25360__ & ~new_new_n25433__;
  assign new_new_n25477__ = new_new_n25465__ & new_new_n25476__;
  assign new_new_n25478__ = ~new_new_n25465__ & ~new_new_n25476__;
  assign new_new_n25479__ = ~new_new_n25477__ & ~new_new_n25478__;
  assign new_new_n25480__ = ~ys__n48327 & ~new_new_n25479__;
  assign new_new_n25481__ = ys__n48327 & new_new_n25479__;
  assign new_new_n25482__ = ~new_new_n25480__ & ~new_new_n25481__;
  assign new_new_n25483__ = ys__n48325 & ~new_new_n25443__;
  assign new_new_n25484__ = new_new_n25362__ & ~new_new_n25446__;
  assign new_new_n25485__ = ~new_new_n25483__ & ~new_new_n25484__;
  assign new_new_n25486__ = new_new_n25482__ & ~new_new_n25485__;
  assign new_new_n25487__ = ~new_new_n25482__ & new_new_n25485__;
  assign new_new_n25488__ = ~new_new_n25486__ & ~new_new_n25487__;
  assign new_new_n25489__ = ~new_new_n25380__ & ~new_new_n25488__;
  assign new_new_n25490__ = ~new_new_n25475__ & ~new_new_n25489__;
  assign new_new_n25491__ = new_new_n25452__ & ~new_new_n25490__;
  assign new_new_n25492__ = ys__n314 & ~new_new_n25491__;
  assign new_new_n25493__ = ~ys__n314 & new_new_n25491__;
  assign new_new_n25494__ = ~new_new_n25492__ & ~new_new_n25493__;
  assign new_new_n25495__ = new_new_n24237__ & ~new_new_n25494__;
  assign new_new_n25496__ = ys__n2535 & ~new_new_n24268__;
  assign new_new_n25497__ = ~new_new_n25495__ & ~new_new_n25496__;
  assign new_new_n25498__ = ~new_new_n12574__ & ~new_new_n25497__;
  assign new_new_n25499__ = ys__n47090 & new_new_n24250__;
  assign new_new_n25500__ = ys__n47026 & new_new_n24252__;
  assign new_new_n25501__ = ~new_new_n25499__ & ~new_new_n25500__;
  assign new_new_n25502__ = ~new_new_n24255__ & ~new_new_n25501__;
  assign new_new_n25503__ = new_new_n24249__ & new_new_n25502__;
  assign new_new_n25504__ = ~new_new_n24227__ & ~new_new_n24249__;
  assign new_new_n25505__ = ~new_new_n25503__ & ~new_new_n25504__;
  assign new_new_n25506__ = new_new_n24265__ & ~new_new_n25505__;
  assign new_new_n25507__ = ~new_new_n24234__ & ~new_new_n24265__;
  assign new_new_n25508__ = ~new_new_n25506__ & ~new_new_n25507__;
  assign new_new_n25509__ = new_new_n12574__ & ~new_new_n25508__;
  assign new_new_n25510__ = ~new_new_n25498__ & ~new_new_n25509__;
  assign new_new_n25511__ = ~ys__n1598 & ~new_new_n25510__;
  assign new_new_n25512__ = ys__n24789 & ys__n1598;
  assign ys__n24790 = new_new_n25511__ | new_new_n25512__;
  assign new_new_n25514__ = ys__n170 & ~new_new_n25491__;
  assign new_new_n25515__ = ys__n170 & ys__n314;
  assign new_new_n25516__ = ~ys__n170 & ~ys__n314;
  assign new_new_n25517__ = ~new_new_n25515__ & ~new_new_n25516__;
  assign new_new_n25518__ = new_new_n25491__ & ~new_new_n25517__;
  assign new_new_n25519__ = ~new_new_n25514__ & ~new_new_n25518__;
  assign new_new_n25520__ = new_new_n24237__ & ~new_new_n25519__;
  assign new_new_n25521__ = ys__n2535 & ~new_new_n24334__;
  assign new_new_n25522__ = ~new_new_n25520__ & ~new_new_n25521__;
  assign new_new_n25523__ = ~new_new_n12574__ & ~new_new_n25522__;
  assign new_new_n25524__ = ys__n47091 & new_new_n24250__;
  assign new_new_n25525__ = ys__n47027 & new_new_n24252__;
  assign new_new_n25526__ = ~new_new_n25524__ & ~new_new_n25525__;
  assign new_new_n25527__ = ~new_new_n24255__ & ~new_new_n25526__;
  assign new_new_n25528__ = new_new_n24249__ & new_new_n25527__;
  assign new_new_n25529__ = ~new_new_n24249__ & ~new_new_n24306__;
  assign new_new_n25530__ = ~new_new_n25528__ & ~new_new_n25529__;
  assign new_new_n25531__ = new_new_n24265__ & ~new_new_n25530__;
  assign new_new_n25532__ = ~new_new_n24265__ & ~new_new_n24312__;
  assign new_new_n25533__ = ~new_new_n25531__ & ~new_new_n25532__;
  assign new_new_n25534__ = new_new_n12574__ & ~new_new_n25533__;
  assign new_new_n25535__ = ~new_new_n25523__ & ~new_new_n25534__;
  assign new_new_n25536__ = ~ys__n1598 & ~new_new_n25535__;
  assign new_new_n25537__ = ys__n24792 & ys__n1598;
  assign ys__n24793 = new_new_n25536__ | new_new_n25537__;
  assign new_new_n25539__ = ys__n380 & ~new_new_n25491__;
  assign new_new_n25540__ = ~ys__n170 & ys__n314;
  assign new_new_n25541__ = ~ys__n170 & ~new_new_n25540__;
  assign new_new_n25542__ = ys__n380 & ~new_new_n25541__;
  assign new_new_n25543__ = ~ys__n380 & new_new_n25541__;
  assign new_new_n25544__ = ~new_new_n25542__ & ~new_new_n25543__;
  assign new_new_n25545__ = new_new_n25491__ & ~new_new_n25544__;
  assign new_new_n25546__ = ~new_new_n25539__ & ~new_new_n25545__;
  assign new_new_n25547__ = new_new_n24237__ & ~new_new_n25546__;
  assign new_new_n25548__ = ys__n2535 & ~new_new_n24406__;
  assign new_new_n25549__ = ~new_new_n25547__ & ~new_new_n25548__;
  assign new_new_n25550__ = ~new_new_n12574__ & ~new_new_n25549__;
  assign new_new_n25551__ = ys__n47092 & new_new_n24250__;
  assign new_new_n25552__ = ys__n47028 & new_new_n24252__;
  assign new_new_n25553__ = ~new_new_n25551__ & ~new_new_n25552__;
  assign new_new_n25554__ = ~new_new_n24255__ & ~new_new_n25553__;
  assign new_new_n25555__ = new_new_n24249__ & new_new_n25554__;
  assign new_new_n25556__ = ~new_new_n24249__ & ~new_new_n24378__;
  assign new_new_n25557__ = ~new_new_n25555__ & ~new_new_n25556__;
  assign new_new_n25558__ = new_new_n24265__ & ~new_new_n25557__;
  assign new_new_n25559__ = ~new_new_n24265__ & ~new_new_n24384__;
  assign new_new_n25560__ = ~new_new_n25558__ & ~new_new_n25559__;
  assign new_new_n25561__ = new_new_n12574__ & ~new_new_n25560__;
  assign new_new_n25562__ = ~new_new_n25550__ & ~new_new_n25561__;
  assign new_new_n25563__ = ~ys__n1598 & ~new_new_n25562__;
  assign new_new_n25564__ = ys__n24795 & ys__n1598;
  assign ys__n24796 = new_new_n25563__ | new_new_n25564__;
  assign new_new_n25566__ = ys__n378 & ~new_new_n25491__;
  assign new_new_n25567__ = ~ys__n380 & ~new_new_n25541__;
  assign new_new_n25568__ = ~ys__n380 & ~new_new_n25567__;
  assign new_new_n25569__ = ys__n378 & ~new_new_n25568__;
  assign new_new_n25570__ = ~ys__n378 & new_new_n25568__;
  assign new_new_n25571__ = ~new_new_n25569__ & ~new_new_n25570__;
  assign new_new_n25572__ = new_new_n25491__ & ~new_new_n25571__;
  assign new_new_n25573__ = ~new_new_n25566__ & ~new_new_n25572__;
  assign new_new_n25574__ = new_new_n24237__ & ~new_new_n25573__;
  assign new_new_n25575__ = ys__n2535 & ~new_new_n24481__;
  assign new_new_n25576__ = ~new_new_n25574__ & ~new_new_n25575__;
  assign new_new_n25577__ = ~new_new_n12574__ & ~new_new_n25576__;
  assign new_new_n25578__ = ys__n47093 & new_new_n24250__;
  assign new_new_n25579__ = ys__n47029 & new_new_n24252__;
  assign new_new_n25580__ = ~new_new_n25578__ & ~new_new_n25579__;
  assign new_new_n25581__ = ~new_new_n24255__ & ~new_new_n25580__;
  assign new_new_n25582__ = new_new_n24249__ & new_new_n25581__;
  assign new_new_n25583__ = ~new_new_n24249__ & ~new_new_n24451__;
  assign new_new_n25584__ = ~new_new_n25582__ & ~new_new_n25583__;
  assign new_new_n25585__ = new_new_n24265__ & ~new_new_n25584__;
  assign new_new_n25586__ = ~new_new_n24265__ & ~new_new_n24459__;
  assign new_new_n25587__ = ~new_new_n25585__ & ~new_new_n25586__;
  assign new_new_n25588__ = new_new_n12574__ & ~new_new_n25587__;
  assign new_new_n25589__ = ~new_new_n25577__ & ~new_new_n25588__;
  assign new_new_n25590__ = ~ys__n1598 & ~new_new_n25589__;
  assign new_new_n25591__ = ys__n24798 & ys__n1598;
  assign ys__n24799 = new_new_n25590__ | new_new_n25591__;
  assign new_new_n25593__ = ys__n382 & ~new_new_n25491__;
  assign new_new_n25594__ = ~ys__n378 & ~ys__n380;
  assign new_new_n25595__ = ~new_new_n25541__ & new_new_n25594__;
  assign new_new_n25596__ = ~ys__n378 & ys__n380;
  assign new_new_n25597__ = ~ys__n378 & ~new_new_n25596__;
  assign new_new_n25598__ = ~new_new_n25595__ & new_new_n25597__;
  assign new_new_n25599__ = ys__n382 & ~new_new_n25598__;
  assign new_new_n25600__ = ~ys__n382 & new_new_n25598__;
  assign new_new_n25601__ = ~new_new_n25599__ & ~new_new_n25600__;
  assign new_new_n25602__ = new_new_n25491__ & ~new_new_n25601__;
  assign new_new_n25603__ = ~new_new_n25593__ & ~new_new_n25602__;
  assign new_new_n25604__ = new_new_n24237__ & ~new_new_n25603__;
  assign new_new_n25605__ = ys__n2535 & ~new_new_n24558__;
  assign new_new_n25606__ = ~new_new_n25604__ & ~new_new_n25605__;
  assign new_new_n25607__ = ~new_new_n12574__ & ~new_new_n25606__;
  assign new_new_n25608__ = ys__n47094 & new_new_n24250__;
  assign new_new_n25609__ = ys__n47030 & new_new_n24252__;
  assign new_new_n25610__ = ~new_new_n25608__ & ~new_new_n25609__;
  assign new_new_n25611__ = ~new_new_n24255__ & ~new_new_n25610__;
  assign new_new_n25612__ = new_new_n24249__ & new_new_n25611__;
  assign new_new_n25613__ = ~new_new_n24249__ & ~new_new_n24530__;
  assign new_new_n25614__ = ~new_new_n25612__ & ~new_new_n25613__;
  assign new_new_n25615__ = new_new_n24265__ & ~new_new_n25614__;
  assign new_new_n25616__ = ~new_new_n24265__ & ~new_new_n24536__;
  assign new_new_n25617__ = ~new_new_n25615__ & ~new_new_n25616__;
  assign new_new_n25618__ = new_new_n12574__ & ~new_new_n25617__;
  assign new_new_n25619__ = ~new_new_n25607__ & ~new_new_n25618__;
  assign new_new_n25620__ = ~ys__n1598 & ~new_new_n25619__;
  assign new_new_n25621__ = ys__n24801 & ys__n1598;
  assign ys__n24802 = new_new_n25620__ | new_new_n25621__;
  assign new_new_n25623__ = ys__n374 & ~new_new_n25491__;
  assign new_new_n25624__ = ~ys__n382 & ~new_new_n25598__;
  assign new_new_n25625__ = ~ys__n382 & ~new_new_n25624__;
  assign new_new_n25626__ = ys__n374 & ~new_new_n25625__;
  assign new_new_n25627__ = ~ys__n374 & new_new_n25625__;
  assign new_new_n25628__ = ~new_new_n25626__ & ~new_new_n25627__;
  assign new_new_n25629__ = new_new_n25491__ & ~new_new_n25628__;
  assign new_new_n25630__ = ~new_new_n25623__ & ~new_new_n25629__;
  assign new_new_n25631__ = new_new_n24237__ & ~new_new_n25630__;
  assign new_new_n25632__ = ys__n2535 & ~new_new_n24634__;
  assign new_new_n25633__ = ~new_new_n25631__ & ~new_new_n25632__;
  assign new_new_n25634__ = ~new_new_n12574__ & ~new_new_n25633__;
  assign new_new_n25635__ = ys__n47095 & new_new_n24250__;
  assign new_new_n25636__ = ys__n47031 & new_new_n24252__;
  assign new_new_n25637__ = ~new_new_n25635__ & ~new_new_n25636__;
  assign new_new_n25638__ = ~new_new_n24255__ & ~new_new_n25637__;
  assign new_new_n25639__ = new_new_n24249__ & new_new_n25638__;
  assign new_new_n25640__ = ~new_new_n24249__ & ~new_new_n24603__;
  assign new_new_n25641__ = ~new_new_n25639__ & ~new_new_n25640__;
  assign new_new_n25642__ = new_new_n24265__ & ~new_new_n25641__;
  assign new_new_n25643__ = ~new_new_n24265__ & ~new_new_n24611__;
  assign new_new_n25644__ = ~new_new_n25642__ & ~new_new_n25643__;
  assign new_new_n25645__ = new_new_n12574__ & ~new_new_n25644__;
  assign new_new_n25646__ = ~new_new_n25634__ & ~new_new_n25645__;
  assign new_new_n25647__ = ~ys__n1598 & ~new_new_n25646__;
  assign new_new_n25648__ = ys__n24804 & ys__n1598;
  assign ys__n24805 = new_new_n25647__ | new_new_n25648__;
  assign new_new_n25650__ = ys__n376 & ~new_new_n25491__;
  assign new_new_n25651__ = ~ys__n374 & ys__n382;
  assign new_new_n25652__ = ~ys__n374 & ~new_new_n25651__;
  assign new_new_n25653__ = ~ys__n374 & ~ys__n382;
  assign new_new_n25654__ = ~new_new_n25598__ & new_new_n25653__;
  assign new_new_n25655__ = new_new_n25652__ & ~new_new_n25654__;
  assign new_new_n25656__ = ys__n376 & ~new_new_n25655__;
  assign new_new_n25657__ = ~ys__n376 & new_new_n25655__;
  assign new_new_n25658__ = ~new_new_n25656__ & ~new_new_n25657__;
  assign new_new_n25659__ = new_new_n25491__ & ~new_new_n25658__;
  assign new_new_n25660__ = ~new_new_n25650__ & ~new_new_n25659__;
  assign new_new_n25661__ = new_new_n24237__ & ~new_new_n25660__;
  assign new_new_n25662__ = ys__n2535 & ~new_new_n24714__;
  assign new_new_n25663__ = ~new_new_n25661__ & ~new_new_n25662__;
  assign new_new_n25664__ = ~new_new_n12574__ & ~new_new_n25663__;
  assign new_new_n25665__ = ys__n47096 & new_new_n24250__;
  assign new_new_n25666__ = ys__n47032 & new_new_n24252__;
  assign new_new_n25667__ = ~new_new_n25665__ & ~new_new_n25666__;
  assign new_new_n25668__ = ~new_new_n24255__ & ~new_new_n25667__;
  assign new_new_n25669__ = new_new_n24249__ & new_new_n25668__;
  assign new_new_n25670__ = ~new_new_n24249__ & ~new_new_n24683__;
  assign new_new_n25671__ = ~new_new_n25669__ & ~new_new_n25670__;
  assign new_new_n25672__ = new_new_n24265__ & ~new_new_n25671__;
  assign new_new_n25673__ = ~new_new_n24265__ & ~new_new_n24691__;
  assign new_new_n25674__ = ~new_new_n25672__ & ~new_new_n25673__;
  assign new_new_n25675__ = new_new_n12574__ & ~new_new_n25674__;
  assign new_new_n25676__ = ~new_new_n25664__ & ~new_new_n25675__;
  assign new_new_n25677__ = ~ys__n1598 & ~new_new_n25676__;
  assign new_new_n25678__ = ys__n24807 & ys__n1598;
  assign ys__n24808 = new_new_n25677__ | new_new_n25678__;
  assign new_new_n25680__ = ys__n372 & ~new_new_n25491__;
  assign new_new_n25681__ = ~ys__n376 & ~new_new_n25655__;
  assign new_new_n25682__ = ~ys__n376 & ~new_new_n25681__;
  assign new_new_n25683__ = ys__n372 & ~new_new_n25682__;
  assign new_new_n25684__ = ~ys__n372 & new_new_n25682__;
  assign new_new_n25685__ = ~new_new_n25683__ & ~new_new_n25684__;
  assign new_new_n25686__ = new_new_n25491__ & ~new_new_n25685__;
  assign new_new_n25687__ = ~new_new_n25680__ & ~new_new_n25686__;
  assign new_new_n25688__ = new_new_n24237__ & ~new_new_n25687__;
  assign new_new_n25689__ = ys__n2535 & ~new_new_n24790__;
  assign new_new_n25690__ = ~new_new_n25688__ & ~new_new_n25689__;
  assign new_new_n25691__ = ~new_new_n12574__ & ~new_new_n25690__;
  assign new_new_n25692__ = ys__n47097 & new_new_n24250__;
  assign new_new_n25693__ = ys__n47033 & new_new_n24252__;
  assign new_new_n25694__ = ~new_new_n25692__ & ~new_new_n25693__;
  assign new_new_n25695__ = ~new_new_n24255__ & ~new_new_n25694__;
  assign new_new_n25696__ = new_new_n24249__ & new_new_n25695__;
  assign new_new_n25697__ = ~new_new_n24249__ & ~new_new_n24759__;
  assign new_new_n25698__ = ~new_new_n25696__ & ~new_new_n25697__;
  assign new_new_n25699__ = new_new_n24265__ & ~new_new_n25698__;
  assign new_new_n25700__ = ~new_new_n24265__ & ~new_new_n24767__;
  assign new_new_n25701__ = ~new_new_n25699__ & ~new_new_n25700__;
  assign new_new_n25702__ = new_new_n12574__ & ~new_new_n25701__;
  assign new_new_n25703__ = ~new_new_n25691__ & ~new_new_n25702__;
  assign new_new_n25704__ = ~ys__n1598 & ~new_new_n25703__;
  assign new_new_n25705__ = ys__n24810 & ys__n1598;
  assign ys__n24811 = new_new_n25704__ | new_new_n25705__;
  assign new_new_n25707__ = ys__n384 & ~new_new_n25491__;
  assign new_new_n25708__ = ~ys__n372 & ~ys__n376;
  assign new_new_n25709__ = new_new_n25653__ & new_new_n25708__;
  assign new_new_n25710__ = ~new_new_n25598__ & new_new_n25709__;
  assign new_new_n25711__ = ~new_new_n25652__ & new_new_n25708__;
  assign new_new_n25712__ = ~ys__n372 & ys__n376;
  assign new_new_n25713__ = ~ys__n372 & ~new_new_n25712__;
  assign new_new_n25714__ = ~new_new_n25711__ & new_new_n25713__;
  assign new_new_n25715__ = ~new_new_n25710__ & new_new_n25714__;
  assign new_new_n25716__ = ys__n384 & ~new_new_n25715__;
  assign new_new_n25717__ = ~ys__n384 & new_new_n25715__;
  assign new_new_n25718__ = ~new_new_n25716__ & ~new_new_n25717__;
  assign new_new_n25719__ = new_new_n25491__ & ~new_new_n25718__;
  assign new_new_n25720__ = ~new_new_n25707__ & ~new_new_n25719__;
  assign new_new_n25721__ = new_new_n24237__ & ~new_new_n25720__;
  assign new_new_n25722__ = ys__n2535 & ~new_new_n24871__;
  assign new_new_n25723__ = ~new_new_n25721__ & ~new_new_n25722__;
  assign new_new_n25724__ = ~new_new_n12574__ & ~new_new_n25723__;
  assign new_new_n25725__ = ys__n47098 & new_new_n24250__;
  assign new_new_n25726__ = ys__n47034 & new_new_n24252__;
  assign new_new_n25727__ = ~new_new_n25725__ & ~new_new_n25726__;
  assign new_new_n25728__ = ~new_new_n24255__ & ~new_new_n25727__;
  assign new_new_n25729__ = new_new_n24249__ & new_new_n25728__;
  assign new_new_n25730__ = ~new_new_n24249__ & ~new_new_n24843__;
  assign new_new_n25731__ = ~new_new_n25729__ & ~new_new_n25730__;
  assign new_new_n25732__ = new_new_n24265__ & ~new_new_n25731__;
  assign new_new_n25733__ = ~new_new_n24265__ & ~new_new_n24849__;
  assign new_new_n25734__ = ~new_new_n25732__ & ~new_new_n25733__;
  assign new_new_n25735__ = new_new_n12574__ & ~new_new_n25734__;
  assign new_new_n25736__ = ~new_new_n25724__ & ~new_new_n25735__;
  assign new_new_n25737__ = ~ys__n1598 & ~new_new_n25736__;
  assign new_new_n25738__ = ys__n24813 & ys__n1598;
  assign ys__n24814 = new_new_n25737__ | new_new_n25738__;
  assign new_new_n25740__ = ys__n366 & ~new_new_n25491__;
  assign new_new_n25741__ = ~ys__n384 & ~new_new_n25715__;
  assign new_new_n25742__ = ~ys__n384 & ~new_new_n25741__;
  assign new_new_n25743__ = ys__n366 & ~new_new_n25742__;
  assign new_new_n25744__ = ~ys__n366 & new_new_n25742__;
  assign new_new_n25745__ = ~new_new_n25743__ & ~new_new_n25744__;
  assign new_new_n25746__ = new_new_n25491__ & ~new_new_n25745__;
  assign new_new_n25747__ = ~new_new_n25740__ & ~new_new_n25746__;
  assign new_new_n25748__ = new_new_n24237__ & ~new_new_n25747__;
  assign new_new_n25749__ = ys__n2535 & ~new_new_n24947__;
  assign new_new_n25750__ = ~new_new_n25748__ & ~new_new_n25749__;
  assign new_new_n25751__ = ~new_new_n12574__ & ~new_new_n25750__;
  assign new_new_n25752__ = ys__n47099 & new_new_n24250__;
  assign new_new_n25753__ = ys__n47035 & new_new_n24252__;
  assign new_new_n25754__ = ~new_new_n25752__ & ~new_new_n25753__;
  assign new_new_n25755__ = ~new_new_n24255__ & ~new_new_n25754__;
  assign new_new_n25756__ = new_new_n24249__ & new_new_n25755__;
  assign new_new_n25757__ = ~new_new_n24249__ & ~new_new_n24916__;
  assign new_new_n25758__ = ~new_new_n25756__ & ~new_new_n25757__;
  assign new_new_n25759__ = new_new_n24265__ & ~new_new_n25758__;
  assign new_new_n25760__ = ~new_new_n24265__ & ~new_new_n24924__;
  assign new_new_n25761__ = ~new_new_n25759__ & ~new_new_n25760__;
  assign new_new_n25762__ = new_new_n12574__ & ~new_new_n25761__;
  assign new_new_n25763__ = ~new_new_n25751__ & ~new_new_n25762__;
  assign new_new_n25764__ = ~ys__n1598 & ~new_new_n25763__;
  assign new_new_n25765__ = ys__n24816 & ys__n1598;
  assign ys__n24817 = new_new_n25764__ | new_new_n25765__;
  assign new_new_n25767__ = ys__n368 & ~new_new_n25491__;
  assign new_new_n25768__ = ~ys__n366 & ys__n384;
  assign new_new_n25769__ = ~ys__n366 & ~new_new_n25768__;
  assign new_new_n25770__ = ~ys__n366 & ~ys__n384;
  assign new_new_n25771__ = ~new_new_n25715__ & new_new_n25770__;
  assign new_new_n25772__ = new_new_n25769__ & ~new_new_n25771__;
  assign new_new_n25773__ = ys__n368 & ~new_new_n25772__;
  assign new_new_n25774__ = ~ys__n368 & new_new_n25772__;
  assign new_new_n25775__ = ~new_new_n25773__ & ~new_new_n25774__;
  assign new_new_n25776__ = new_new_n25491__ & ~new_new_n25775__;
  assign new_new_n25777__ = ~new_new_n25767__ & ~new_new_n25776__;
  assign new_new_n25778__ = new_new_n24237__ & ~new_new_n25777__;
  assign new_new_n25779__ = ys__n2535 & ~new_new_n25027__;
  assign new_new_n25780__ = ~new_new_n25778__ & ~new_new_n25779__;
  assign new_new_n25781__ = ~new_new_n12574__ & ~new_new_n25780__;
  assign new_new_n25782__ = ys__n47100 & new_new_n24250__;
  assign new_new_n25783__ = ys__n47036 & new_new_n24252__;
  assign new_new_n25784__ = ~new_new_n25782__ & ~new_new_n25783__;
  assign new_new_n25785__ = ~new_new_n24255__ & ~new_new_n25784__;
  assign new_new_n25786__ = new_new_n24249__ & new_new_n25785__;
  assign new_new_n25787__ = ~new_new_n24249__ & ~new_new_n24996__;
  assign new_new_n25788__ = ~new_new_n25786__ & ~new_new_n25787__;
  assign new_new_n25789__ = new_new_n24265__ & ~new_new_n25788__;
  assign new_new_n25790__ = ~new_new_n24265__ & ~new_new_n25004__;
  assign new_new_n25791__ = ~new_new_n25789__ & ~new_new_n25790__;
  assign new_new_n25792__ = new_new_n12574__ & ~new_new_n25791__;
  assign new_new_n25793__ = ~new_new_n25781__ & ~new_new_n25792__;
  assign new_new_n25794__ = ~ys__n1598 & ~new_new_n25793__;
  assign new_new_n25795__ = ys__n24819 & ys__n1598;
  assign ys__n24820 = new_new_n25794__ | new_new_n25795__;
  assign new_new_n25797__ = ys__n364 & ~new_new_n25491__;
  assign new_new_n25798__ = ~ys__n368 & ~new_new_n25772__;
  assign new_new_n25799__ = ~ys__n368 & ~new_new_n25798__;
  assign new_new_n25800__ = ys__n364 & ~new_new_n25799__;
  assign new_new_n25801__ = ~ys__n364 & new_new_n25799__;
  assign new_new_n25802__ = ~new_new_n25800__ & ~new_new_n25801__;
  assign new_new_n25803__ = new_new_n25491__ & ~new_new_n25802__;
  assign new_new_n25804__ = ~new_new_n25797__ & ~new_new_n25803__;
  assign new_new_n25805__ = new_new_n24237__ & ~new_new_n25804__;
  assign new_new_n25806__ = ys__n2535 & ~new_new_n25103__;
  assign new_new_n25807__ = ~new_new_n25805__ & ~new_new_n25806__;
  assign new_new_n25808__ = ~new_new_n12574__ & ~new_new_n25807__;
  assign new_new_n25809__ = ys__n47101 & new_new_n24250__;
  assign new_new_n25810__ = ys__n47037 & new_new_n24252__;
  assign new_new_n25811__ = ~new_new_n25809__ & ~new_new_n25810__;
  assign new_new_n25812__ = ~new_new_n24255__ & ~new_new_n25811__;
  assign new_new_n25813__ = new_new_n24249__ & new_new_n25812__;
  assign new_new_n25814__ = ~new_new_n24249__ & ~new_new_n25072__;
  assign new_new_n25815__ = ~new_new_n25813__ & ~new_new_n25814__;
  assign new_new_n25816__ = new_new_n24265__ & ~new_new_n25815__;
  assign new_new_n25817__ = ~new_new_n24265__ & ~new_new_n25080__;
  assign new_new_n25818__ = ~new_new_n25816__ & ~new_new_n25817__;
  assign new_new_n25819__ = new_new_n12574__ & ~new_new_n25818__;
  assign new_new_n25820__ = ~new_new_n25808__ & ~new_new_n25819__;
  assign new_new_n25821__ = ~ys__n1598 & ~new_new_n25820__;
  assign new_new_n25822__ = ys__n24822 & ys__n1598;
  assign ys__n24823 = new_new_n25821__ | new_new_n25822__;
  assign new_new_n25824__ = ys__n370 & ~new_new_n25491__;
  assign new_new_n25825__ = ~ys__n364 & ~ys__n368;
  assign new_new_n25826__ = ~new_new_n25769__ & new_new_n25825__;
  assign new_new_n25827__ = ~ys__n364 & ys__n368;
  assign new_new_n25828__ = ~ys__n364 & ~new_new_n25827__;
  assign new_new_n25829__ = ~new_new_n25826__ & new_new_n25828__;
  assign new_new_n25830__ = new_new_n25770__ & new_new_n25825__;
  assign new_new_n25831__ = ~new_new_n25715__ & new_new_n25830__;
  assign new_new_n25832__ = new_new_n25829__ & ~new_new_n25831__;
  assign new_new_n25833__ = ys__n370 & ~new_new_n25832__;
  assign new_new_n25834__ = ~ys__n370 & new_new_n25832__;
  assign new_new_n25835__ = ~new_new_n25833__ & ~new_new_n25834__;
  assign new_new_n25836__ = new_new_n25491__ & ~new_new_n25835__;
  assign new_new_n25837__ = ~new_new_n25824__ & ~new_new_n25836__;
  assign new_new_n25838__ = new_new_n24237__ & ~new_new_n25837__;
  assign new_new_n25839__ = ys__n2535 & ~new_new_n25187__;
  assign new_new_n25840__ = ~new_new_n25838__ & ~new_new_n25839__;
  assign new_new_n25841__ = ~new_new_n12574__ & ~new_new_n25840__;
  assign new_new_n25842__ = ys__n47102 & new_new_n24250__;
  assign new_new_n25843__ = ys__n47038 & new_new_n24252__;
  assign new_new_n25844__ = ~new_new_n25842__ & ~new_new_n25843__;
  assign new_new_n25845__ = ~new_new_n24255__ & ~new_new_n25844__;
  assign new_new_n25846__ = new_new_n24249__ & new_new_n25845__;
  assign new_new_n25847__ = ~new_new_n24249__ & ~new_new_n25156__;
  assign new_new_n25848__ = ~new_new_n25846__ & ~new_new_n25847__;
  assign new_new_n25849__ = new_new_n24265__ & ~new_new_n25848__;
  assign new_new_n25850__ = ~new_new_n24265__ & ~new_new_n25164__;
  assign new_new_n25851__ = ~new_new_n25849__ & ~new_new_n25850__;
  assign new_new_n25852__ = new_new_n12574__ & ~new_new_n25851__;
  assign new_new_n25853__ = ~new_new_n25841__ & ~new_new_n25852__;
  assign new_new_n25854__ = ~ys__n1598 & ~new_new_n25853__;
  assign new_new_n25855__ = ys__n24825 & ys__n1598;
  assign ys__n24826 = new_new_n25854__ | new_new_n25855__;
  assign new_new_n25857__ = ys__n360 & ~new_new_n25491__;
  assign new_new_n25858__ = ~ys__n370 & ~new_new_n25832__;
  assign new_new_n25859__ = ~ys__n370 & ~new_new_n25858__;
  assign new_new_n25860__ = ys__n360 & ~new_new_n25859__;
  assign new_new_n25861__ = ~ys__n360 & new_new_n25859__;
  assign new_new_n25862__ = ~new_new_n25860__ & ~new_new_n25861__;
  assign new_new_n25863__ = new_new_n25491__ & ~new_new_n25862__;
  assign new_new_n25864__ = ~new_new_n25857__ & ~new_new_n25863__;
  assign new_new_n25865__ = new_new_n24237__ & ~new_new_n25864__;
  assign new_new_n25866__ = ys__n2535 & ~new_new_n25263__;
  assign new_new_n25867__ = ~new_new_n25865__ & ~new_new_n25866__;
  assign new_new_n25868__ = ~new_new_n12574__ & ~new_new_n25867__;
  assign new_new_n25869__ = ys__n47103 & new_new_n24250__;
  assign new_new_n25870__ = ys__n47039 & new_new_n24252__;
  assign new_new_n25871__ = ~new_new_n25869__ & ~new_new_n25870__;
  assign new_new_n25872__ = ~new_new_n24255__ & ~new_new_n25871__;
  assign new_new_n25873__ = new_new_n24249__ & new_new_n25872__;
  assign new_new_n25874__ = ~new_new_n24249__ & ~new_new_n25232__;
  assign new_new_n25875__ = ~new_new_n25873__ & ~new_new_n25874__;
  assign new_new_n25876__ = new_new_n24265__ & ~new_new_n25875__;
  assign new_new_n25877__ = ~new_new_n24265__ & ~new_new_n25240__;
  assign new_new_n25878__ = ~new_new_n25876__ & ~new_new_n25877__;
  assign new_new_n25879__ = new_new_n12574__ & ~new_new_n25878__;
  assign new_new_n25880__ = ~new_new_n25868__ & ~new_new_n25879__;
  assign new_new_n25881__ = ~ys__n1598 & ~new_new_n25880__;
  assign new_new_n25882__ = ys__n24828 & ys__n1598;
  assign ys__n24829 = new_new_n25881__ | new_new_n25882__;
  assign new_new_n25884__ = ys__n362 & ~new_new_n25491__;
  assign new_new_n25885__ = ~ys__n360 & ys__n370;
  assign new_new_n25886__ = ~ys__n360 & ~new_new_n25885__;
  assign new_new_n25887__ = ~ys__n360 & ~ys__n370;
  assign new_new_n25888__ = ~new_new_n25832__ & new_new_n25887__;
  assign new_new_n25889__ = new_new_n25886__ & ~new_new_n25888__;
  assign new_new_n25890__ = ys__n362 & ~new_new_n25889__;
  assign new_new_n25891__ = ~ys__n362 & new_new_n25889__;
  assign new_new_n25892__ = ~new_new_n25890__ & ~new_new_n25891__;
  assign new_new_n25893__ = new_new_n25491__ & ~new_new_n25892__;
  assign new_new_n25894__ = ~new_new_n25884__ & ~new_new_n25893__;
  assign new_new_n25895__ = new_new_n24237__ & ~new_new_n25894__;
  assign new_new_n25896__ = ys__n2535 & ~new_new_n25343__;
  assign new_new_n25897__ = ~new_new_n25895__ & ~new_new_n25896__;
  assign new_new_n25898__ = ~new_new_n12574__ & ~new_new_n25897__;
  assign new_new_n25899__ = ys__n47104 & new_new_n24250__;
  assign new_new_n25900__ = ys__n47040 & new_new_n24252__;
  assign new_new_n25901__ = ~new_new_n25899__ & ~new_new_n25900__;
  assign new_new_n25902__ = ~new_new_n24255__ & ~new_new_n25901__;
  assign new_new_n25903__ = new_new_n24249__ & new_new_n25902__;
  assign new_new_n25904__ = ~new_new_n24249__ & ~new_new_n25312__;
  assign new_new_n25905__ = ~new_new_n25903__ & ~new_new_n25904__;
  assign new_new_n25906__ = new_new_n24265__ & ~new_new_n25905__;
  assign new_new_n25907__ = ~new_new_n24265__ & ~new_new_n25320__;
  assign new_new_n25908__ = ~new_new_n25906__ & ~new_new_n25907__;
  assign new_new_n25909__ = new_new_n12574__ & ~new_new_n25908__;
  assign new_new_n25910__ = ~new_new_n25898__ & ~new_new_n25909__;
  assign new_new_n25911__ = ~ys__n1598 & ~new_new_n25910__;
  assign new_new_n25912__ = ys__n24831 & ys__n1598;
  assign ys__n24832 = new_new_n25911__ | new_new_n25912__;
  assign new_new_n25914__ = ys__n358 & ~new_new_n25491__;
  assign new_new_n25915__ = ~ys__n362 & ~new_new_n25889__;
  assign new_new_n25916__ = ~ys__n362 & ~new_new_n25915__;
  assign new_new_n25917__ = ys__n358 & ~new_new_n25916__;
  assign new_new_n25918__ = ~ys__n358 & new_new_n25916__;
  assign new_new_n25919__ = ~new_new_n25917__ & ~new_new_n25918__;
  assign new_new_n25920__ = new_new_n25491__ & ~new_new_n25919__;
  assign new_new_n25921__ = ~new_new_n25914__ & ~new_new_n25920__;
  assign new_new_n25922__ = new_new_n24237__ & ~new_new_n25921__;
  assign new_new_n25923__ = ys__n2535 & ~new_new_n25417__;
  assign new_new_n25924__ = ~new_new_n25922__ & ~new_new_n25923__;
  assign new_new_n25925__ = ~new_new_n12574__ & ~new_new_n25924__;
  assign new_new_n25926__ = ys__n47105 & new_new_n24250__;
  assign new_new_n25927__ = ys__n47041 & new_new_n24252__;
  assign new_new_n25928__ = ~new_new_n25926__ & ~new_new_n25927__;
  assign new_new_n25929__ = ~new_new_n24255__ & ~new_new_n25928__;
  assign new_new_n25930__ = new_new_n24249__ & new_new_n25929__;
  assign new_new_n25931__ = ~new_new_n24249__ & ~new_new_n25386__;
  assign new_new_n25932__ = ~new_new_n25930__ & ~new_new_n25931__;
  assign new_new_n25933__ = new_new_n24265__ & ~new_new_n25932__;
  assign new_new_n25934__ = ~new_new_n24265__ & ~new_new_n25394__;
  assign new_new_n25935__ = ~new_new_n25933__ & ~new_new_n25934__;
  assign new_new_n25936__ = new_new_n12574__ & ~new_new_n25935__;
  assign new_new_n25937__ = ~new_new_n25925__ & ~new_new_n25936__;
  assign new_new_n25938__ = ~ys__n1598 & ~new_new_n25937__;
  assign new_new_n25939__ = ys__n24834 & ys__n1598;
  assign ys__n24835 = new_new_n25938__ | new_new_n25939__;
  assign new_new_n25941__ = ys__n386 & ~new_new_n25491__;
  assign new_new_n25942__ = ~ys__n358 & ~ys__n362;
  assign new_new_n25943__ = new_new_n25887__ & new_new_n25942__;
  assign new_new_n25944__ = new_new_n25830__ & new_new_n25943__;
  assign new_new_n25945__ = ~new_new_n25715__ & new_new_n25944__;
  assign new_new_n25946__ = ~new_new_n25829__ & new_new_n25943__;
  assign new_new_n25947__ = ~new_new_n25886__ & new_new_n25942__;
  assign new_new_n25948__ = ~ys__n358 & ys__n362;
  assign new_new_n25949__ = ~ys__n358 & ~new_new_n25948__;
  assign new_new_n25950__ = ~new_new_n25947__ & new_new_n25949__;
  assign new_new_n25951__ = ~new_new_n25946__ & new_new_n25950__;
  assign new_new_n25952__ = ~new_new_n25945__ & new_new_n25951__;
  assign new_new_n25953__ = ys__n386 & ~new_new_n25952__;
  assign new_new_n25954__ = ~ys__n386 & new_new_n25952__;
  assign new_new_n25955__ = ~new_new_n25953__ & ~new_new_n25954__;
  assign new_new_n25956__ = new_new_n25491__ & ~new_new_n25955__;
  assign new_new_n25957__ = ~new_new_n25941__ & ~new_new_n25956__;
  assign new_new_n25958__ = ~new_new_n12574__ & new_new_n24237__;
  assign new_new_n25959__ = ~new_new_n25957__ & new_new_n25958__;
  assign new_new_n25960__ = ~new_new_n24249__ & new_new_n24265__;
  assign new_new_n25961__ = ~new_new_n25451__ & new_new_n25960__;
  assign new_new_n25962__ = new_new_n12574__ & new_new_n25961__;
  assign new_new_n25963__ = ~new_new_n25959__ & ~new_new_n25962__;
  assign new_new_n25964__ = ~ys__n1598 & ~new_new_n25963__;
  assign ys__n24837 = new_new_n25939__ | new_new_n25964__;
  assign new_new_n25966__ = ys__n356 & ~new_new_n25491__;
  assign new_new_n25967__ = ~ys__n386 & ~new_new_n25952__;
  assign new_new_n25968__ = ~ys__n386 & ~new_new_n25967__;
  assign new_new_n25969__ = ys__n356 & ~new_new_n25968__;
  assign new_new_n25970__ = ~ys__n356 & new_new_n25968__;
  assign new_new_n25971__ = ~new_new_n25969__ & ~new_new_n25970__;
  assign new_new_n25972__ = new_new_n25491__ & ~new_new_n25971__;
  assign new_new_n25973__ = ~new_new_n25966__ & ~new_new_n25972__;
  assign new_new_n25974__ = new_new_n25958__ & ~new_new_n25973__;
  assign ys__n24907 = ~new_new_n25490__ & new_new_n25960__;
  assign new_new_n25976__ = new_new_n12574__ & ys__n24907;
  assign new_new_n25977__ = ~new_new_n25974__ & ~new_new_n25976__;
  assign new_new_n25978__ = ~ys__n1598 & ~new_new_n25977__;
  assign ys__n24839 = new_new_n25939__ | new_new_n25978__;
  assign new_new_n25980__ = ys__n31031 & ys__n47010;
  assign new_new_n25981__ = new_new_n23480__ & new_new_n25980__;
  assign new_new_n25982__ = ~new_new_n23480__ & ~new_new_n24260__;
  assign new_new_n25983__ = ~new_new_n25981__ & ~new_new_n25982__;
  assign new_new_n25984__ = ~new_new_n24230__ & ~new_new_n25983__;
  assign new_new_n25985__ = ys__n314 & new_new_n24230__;
  assign new_new_n25986__ = ~new_new_n25984__ & ~new_new_n25985__;
  assign new_new_n25987__ = new_new_n24237__ & ~new_new_n25986__;
  assign new_new_n25988__ = ys__n2535 & ~new_new_n25986__;
  assign ys__n24910 = new_new_n25987__ | new_new_n25988__;
  assign new_new_n25990__ = ys__n31031 & ys__n47011;
  assign new_new_n25991__ = new_new_n23480__ & new_new_n25990__;
  assign new_new_n25992__ = ~new_new_n23480__ & ~new_new_n24329__;
  assign new_new_n25993__ = ~new_new_n25991__ & ~new_new_n25992__;
  assign new_new_n25994__ = ~new_new_n24230__ & ~new_new_n25993__;
  assign new_new_n25995__ = ys__n170 & new_new_n24230__;
  assign new_new_n25996__ = ~new_new_n25994__ & ~new_new_n25995__;
  assign new_new_n25997__ = new_new_n24237__ & ~new_new_n25996__;
  assign new_new_n25998__ = ys__n2535 & ~new_new_n25996__;
  assign ys__n24913 = new_new_n25997__ | new_new_n25998__;
  assign new_new_n26000__ = ys__n31031 & ys__n47012;
  assign new_new_n26001__ = new_new_n23480__ & new_new_n26000__;
  assign new_new_n26002__ = ~new_new_n23480__ & ~new_new_n24401__;
  assign new_new_n26003__ = ~new_new_n26001__ & ~new_new_n26002__;
  assign new_new_n26004__ = ~new_new_n24230__ & ~new_new_n26003__;
  assign new_new_n26005__ = ys__n380 & new_new_n24230__;
  assign new_new_n26006__ = ~new_new_n26004__ & ~new_new_n26005__;
  assign new_new_n26007__ = new_new_n24237__ & ~new_new_n26006__;
  assign new_new_n26008__ = ys__n2535 & ~new_new_n26006__;
  assign ys__n24916 = new_new_n26007__ | new_new_n26008__;
  assign new_new_n26010__ = ys__n31031 & ys__n47013;
  assign new_new_n26011__ = new_new_n23480__ & new_new_n26010__;
  assign new_new_n26012__ = ~new_new_n23480__ & ~new_new_n24476__;
  assign new_new_n26013__ = ~new_new_n26011__ & ~new_new_n26012__;
  assign new_new_n26014__ = ~new_new_n24230__ & ~new_new_n26013__;
  assign new_new_n26015__ = ys__n378 & new_new_n24230__;
  assign new_new_n26016__ = ~new_new_n26014__ & ~new_new_n26015__;
  assign new_new_n26017__ = new_new_n24237__ & ~new_new_n26016__;
  assign new_new_n26018__ = ys__n2535 & ~new_new_n26016__;
  assign ys__n24919 = new_new_n26017__ | new_new_n26018__;
  assign new_new_n26020__ = ys__n31031 & ys__n47014;
  assign new_new_n26021__ = new_new_n23480__ & new_new_n26020__;
  assign new_new_n26022__ = ~new_new_n23480__ & ~new_new_n24553__;
  assign new_new_n26023__ = ~new_new_n26021__ & ~new_new_n26022__;
  assign new_new_n26024__ = ~new_new_n24230__ & ~new_new_n26023__;
  assign new_new_n26025__ = ys__n382 & new_new_n24230__;
  assign new_new_n26026__ = ~new_new_n26024__ & ~new_new_n26025__;
  assign new_new_n26027__ = new_new_n24237__ & ~new_new_n26026__;
  assign new_new_n26028__ = ys__n2535 & ~new_new_n26026__;
  assign ys__n24922 = new_new_n26027__ | new_new_n26028__;
  assign new_new_n26030__ = ys__n31031 & ys__n47015;
  assign new_new_n26031__ = new_new_n23480__ & new_new_n26030__;
  assign new_new_n26032__ = ~new_new_n23480__ & ~new_new_n24629__;
  assign new_new_n26033__ = ~new_new_n26031__ & ~new_new_n26032__;
  assign new_new_n26034__ = ~new_new_n24230__ & ~new_new_n26033__;
  assign new_new_n26035__ = ys__n374 & new_new_n24230__;
  assign new_new_n26036__ = ~new_new_n26034__ & ~new_new_n26035__;
  assign new_new_n26037__ = new_new_n24237__ & ~new_new_n26036__;
  assign new_new_n26038__ = ys__n2535 & ~new_new_n26036__;
  assign ys__n24925 = new_new_n26037__ | new_new_n26038__;
  assign new_new_n26040__ = ys__n31031 & ys__n47016;
  assign new_new_n26041__ = new_new_n23480__ & new_new_n26040__;
  assign new_new_n26042__ = ~new_new_n23480__ & ~new_new_n24709__;
  assign new_new_n26043__ = ~new_new_n26041__ & ~new_new_n26042__;
  assign new_new_n26044__ = ~new_new_n24230__ & ~new_new_n26043__;
  assign new_new_n26045__ = ys__n376 & new_new_n24230__;
  assign new_new_n26046__ = ~new_new_n26044__ & ~new_new_n26045__;
  assign new_new_n26047__ = new_new_n24237__ & ~new_new_n26046__;
  assign new_new_n26048__ = ys__n2535 & ~new_new_n26046__;
  assign ys__n24928 = new_new_n26047__ | new_new_n26048__;
  assign new_new_n26050__ = ys__n31031 & ys__n47017;
  assign new_new_n26051__ = new_new_n23480__ & new_new_n26050__;
  assign new_new_n26052__ = ~new_new_n23480__ & ~new_new_n24785__;
  assign new_new_n26053__ = ~new_new_n26051__ & ~new_new_n26052__;
  assign new_new_n26054__ = ~new_new_n24230__ & ~new_new_n26053__;
  assign new_new_n26055__ = ys__n372 & new_new_n24230__;
  assign new_new_n26056__ = ~new_new_n26054__ & ~new_new_n26055__;
  assign new_new_n26057__ = new_new_n24237__ & ~new_new_n26056__;
  assign new_new_n26058__ = ys__n2535 & ~new_new_n26056__;
  assign ys__n24931 = new_new_n26057__ | new_new_n26058__;
  assign new_new_n26060__ = ys__n31031 & ys__n47018;
  assign new_new_n26061__ = new_new_n23480__ & new_new_n26060__;
  assign new_new_n26062__ = ~new_new_n23480__ & ~new_new_n24866__;
  assign new_new_n26063__ = ~new_new_n26061__ & ~new_new_n26062__;
  assign new_new_n26064__ = ~new_new_n24230__ & ~new_new_n26063__;
  assign new_new_n26065__ = ys__n384 & new_new_n24230__;
  assign new_new_n26066__ = ~new_new_n26064__ & ~new_new_n26065__;
  assign new_new_n26067__ = new_new_n24237__ & ~new_new_n26066__;
  assign new_new_n26068__ = ys__n2535 & ~new_new_n26066__;
  assign ys__n24934 = new_new_n26067__ | new_new_n26068__;
  assign new_new_n26070__ = ys__n31031 & ys__n47019;
  assign new_new_n26071__ = new_new_n23480__ & new_new_n26070__;
  assign new_new_n26072__ = ~new_new_n23480__ & ~new_new_n24942__;
  assign new_new_n26073__ = ~new_new_n26071__ & ~new_new_n26072__;
  assign new_new_n26074__ = ~new_new_n24230__ & ~new_new_n26073__;
  assign new_new_n26075__ = ys__n366 & new_new_n24230__;
  assign new_new_n26076__ = ~new_new_n26074__ & ~new_new_n26075__;
  assign new_new_n26077__ = new_new_n24237__ & ~new_new_n26076__;
  assign new_new_n26078__ = ys__n2535 & ~new_new_n26076__;
  assign ys__n24937 = new_new_n26077__ | new_new_n26078__;
  assign new_new_n26080__ = ys__n31031 & ys__n47020;
  assign new_new_n26081__ = new_new_n23480__ & new_new_n26080__;
  assign new_new_n26082__ = ~new_new_n23480__ & ~new_new_n25022__;
  assign new_new_n26083__ = ~new_new_n26081__ & ~new_new_n26082__;
  assign new_new_n26084__ = ~new_new_n24230__ & ~new_new_n26083__;
  assign new_new_n26085__ = ys__n368 & new_new_n24230__;
  assign new_new_n26086__ = ~new_new_n26084__ & ~new_new_n26085__;
  assign new_new_n26087__ = new_new_n24237__ & ~new_new_n26086__;
  assign new_new_n26088__ = ys__n2535 & ~new_new_n26086__;
  assign ys__n24940 = new_new_n26087__ | new_new_n26088__;
  assign new_new_n26090__ = ys__n31031 & ys__n47021;
  assign new_new_n26091__ = new_new_n23480__ & new_new_n26090__;
  assign new_new_n26092__ = ~new_new_n23480__ & ~new_new_n25098__;
  assign new_new_n26093__ = ~new_new_n26091__ & ~new_new_n26092__;
  assign new_new_n26094__ = ~new_new_n24230__ & ~new_new_n26093__;
  assign new_new_n26095__ = ys__n364 & new_new_n24230__;
  assign new_new_n26096__ = ~new_new_n26094__ & ~new_new_n26095__;
  assign new_new_n26097__ = new_new_n24237__ & ~new_new_n26096__;
  assign new_new_n26098__ = ys__n2535 & ~new_new_n26096__;
  assign ys__n24943 = new_new_n26097__ | new_new_n26098__;
  assign new_new_n26100__ = ys__n31031 & ys__n47022;
  assign new_new_n26101__ = new_new_n23480__ & new_new_n26100__;
  assign new_new_n26102__ = ~new_new_n23480__ & ~new_new_n25182__;
  assign new_new_n26103__ = ~new_new_n26101__ & ~new_new_n26102__;
  assign new_new_n26104__ = ~new_new_n24230__ & ~new_new_n26103__;
  assign new_new_n26105__ = ys__n370 & new_new_n24230__;
  assign new_new_n26106__ = ~new_new_n26104__ & ~new_new_n26105__;
  assign new_new_n26107__ = new_new_n24237__ & ~new_new_n26106__;
  assign new_new_n26108__ = ys__n2535 & ~new_new_n26106__;
  assign ys__n24946 = new_new_n26107__ | new_new_n26108__;
  assign new_new_n26110__ = ys__n31031 & ys__n47023;
  assign new_new_n26111__ = new_new_n23480__ & new_new_n26110__;
  assign new_new_n26112__ = ~new_new_n23480__ & ~new_new_n25258__;
  assign new_new_n26113__ = ~new_new_n26111__ & ~new_new_n26112__;
  assign new_new_n26114__ = ~new_new_n24230__ & ~new_new_n26113__;
  assign new_new_n26115__ = ys__n360 & new_new_n24230__;
  assign new_new_n26116__ = ~new_new_n26114__ & ~new_new_n26115__;
  assign new_new_n26117__ = new_new_n24237__ & ~new_new_n26116__;
  assign new_new_n26118__ = ys__n2535 & ~new_new_n26116__;
  assign ys__n24949 = new_new_n26117__ | new_new_n26118__;
  assign new_new_n26120__ = ys__n31031 & ys__n47024;
  assign new_new_n26121__ = new_new_n23480__ & new_new_n26120__;
  assign new_new_n26122__ = ~new_new_n23480__ & ~new_new_n25338__;
  assign new_new_n26123__ = ~new_new_n26121__ & ~new_new_n26122__;
  assign new_new_n26124__ = ~new_new_n24230__ & ~new_new_n26123__;
  assign new_new_n26125__ = ys__n362 & new_new_n24230__;
  assign new_new_n26126__ = ~new_new_n26124__ & ~new_new_n26125__;
  assign new_new_n26127__ = new_new_n24237__ & ~new_new_n26126__;
  assign new_new_n26128__ = ys__n2535 & ~new_new_n26126__;
  assign ys__n24952 = new_new_n26127__ | new_new_n26128__;
  assign new_new_n26130__ = ys__n31031 & ys__n47025;
  assign new_new_n26131__ = new_new_n23480__ & new_new_n26130__;
  assign new_new_n26132__ = ~new_new_n23480__ & ~new_new_n25412__;
  assign new_new_n26133__ = ~new_new_n26131__ & ~new_new_n26132__;
  assign new_new_n26134__ = ~new_new_n24230__ & ~new_new_n26133__;
  assign new_new_n26135__ = ys__n358 & new_new_n24230__;
  assign new_new_n26136__ = ~new_new_n26134__ & ~new_new_n26135__;
  assign new_new_n26137__ = new_new_n24237__ & ~new_new_n26136__;
  assign new_new_n26138__ = ys__n2535 & ~new_new_n26136__;
  assign ys__n24955 = new_new_n26137__ | new_new_n26138__;
  assign new_new_n26140__ = ys__n698 & ys__n25300;
  assign new_new_n26141__ = new_new_n15900__ & new_new_n26140__;
  assign new_new_n26142__ = new_new_n13930__ & new_new_n15901__;
  assign ys__n25294 = new_new_n26141__ & new_new_n26142__;
  assign new_new_n26144__ = new_new_n13934__ & new_new_n15903__;
  assign new_new_n26145__ = new_new_n13933__ & new_new_n26144__;
  assign new_new_n26146__ = ~ys__n780 & ys__n2644;
  assign new_new_n26147__ = ys__n25292 & new_new_n26146__;
  assign new_new_n26148__ = ~ys__n772 & ~ys__n782;
  assign new_new_n26149__ = new_new_n15900__ & new_new_n26148__;
  assign new_new_n26150__ = new_new_n26142__ & new_new_n26149__;
  assign new_new_n26151__ = new_new_n26147__ & new_new_n26150__;
  assign new_new_n26152__ = new_new_n26145__ & new_new_n26151__;
  assign ys__n25302 = ys__n4168 | new_new_n26152__;
  assign new_new_n26154__ = ys__n25381 & new_new_n26146__;
  assign new_new_n26155__ = new_new_n26150__ & new_new_n26154__;
  assign ys__n25304 = new_new_n26145__ & new_new_n26155__;
  assign new_new_n26157__ = ys__n25382 & new_new_n26146__;
  assign new_new_n26158__ = new_new_n26150__ & new_new_n26157__;
  assign ys__n25306 = new_new_n26145__ & new_new_n26158__;
  assign new_new_n26160__ = ys__n25383 & new_new_n26146__;
  assign new_new_n26161__ = new_new_n26150__ & new_new_n26160__;
  assign ys__n25308 = new_new_n26145__ & new_new_n26161__;
  assign new_new_n26163__ = ys__n25384 & new_new_n26146__;
  assign new_new_n26164__ = new_new_n26150__ & new_new_n26163__;
  assign ys__n25310 = new_new_n26145__ & new_new_n26164__;
  assign new_new_n26166__ = ys__n29883 & ~new_new_n10603__;
  assign new_new_n26167__ = ~new_new_n10601__ & new_new_n26166__;
  assign new_new_n26168__ = ~ys__n23764 & new_new_n26167__;
  assign new_new_n26169__ = ys__n29899 & ~new_new_n10603__;
  assign new_new_n26170__ = ~new_new_n10601__ & new_new_n26169__;
  assign new_new_n26171__ = ~ys__n22466 & new_new_n26170__;
  assign new_new_n26172__ = ys__n22466 & new_new_n26167__;
  assign new_new_n26173__ = ~new_new_n26171__ & ~new_new_n26172__;
  assign new_new_n26174__ = ys__n23764 & ~new_new_n26173__;
  assign new_new_n26175__ = ~new_new_n26168__ & ~new_new_n26174__;
  assign ys__n25385 = new_new_n10866__ & ~new_new_n26175__;
  assign new_new_n26177__ = ys__n29884 & ~new_new_n10603__;
  assign new_new_n26178__ = ~new_new_n10601__ & new_new_n26177__;
  assign new_new_n26179__ = ~ys__n23764 & new_new_n26178__;
  assign new_new_n26180__ = ys__n29900 & ~new_new_n10603__;
  assign new_new_n26181__ = ~new_new_n10601__ & new_new_n26180__;
  assign new_new_n26182__ = ~ys__n22466 & new_new_n26181__;
  assign new_new_n26183__ = ys__n22466 & new_new_n26178__;
  assign new_new_n26184__ = ~new_new_n26182__ & ~new_new_n26183__;
  assign new_new_n26185__ = ys__n23764 & ~new_new_n26184__;
  assign new_new_n26186__ = ~new_new_n26179__ & ~new_new_n26185__;
  assign ys__n25386 = new_new_n10866__ & ~new_new_n26186__;
  assign new_new_n26188__ = ys__n29885 & ~new_new_n10603__;
  assign new_new_n26189__ = ~new_new_n10601__ & new_new_n26188__;
  assign new_new_n26190__ = ~ys__n23764 & new_new_n26189__;
  assign new_new_n26191__ = ys__n29901 & ~new_new_n10603__;
  assign new_new_n26192__ = ~new_new_n10601__ & new_new_n26191__;
  assign new_new_n26193__ = ~ys__n22466 & new_new_n26192__;
  assign new_new_n26194__ = ys__n22466 & new_new_n26189__;
  assign new_new_n26195__ = ~new_new_n26193__ & ~new_new_n26194__;
  assign new_new_n26196__ = ys__n23764 & ~new_new_n26195__;
  assign new_new_n26197__ = ~new_new_n26190__ & ~new_new_n26196__;
  assign ys__n25387 = new_new_n10866__ & ~new_new_n26197__;
  assign new_new_n26199__ = ~ys__n782 & ys__n2644;
  assign new_new_n26200__ = ys__n25300 & new_new_n26199__;
  assign new_new_n26201__ = new_new_n15906__ & new_new_n15916__;
  assign new_new_n26202__ = new_new_n26200__ & new_new_n26201__;
  assign new_new_n26203__ = ys__n598 & ys__n25300;
  assign new_new_n26204__ = ~new_new_n26202__ & ~new_new_n26203__;
  assign new_new_n26205__ = ~ys__n778 & new_new_n13927__;
  assign new_new_n26206__ = new_new_n13932__ & new_new_n26205__;
  assign new_new_n26207__ = ~new_new_n26204__ & new_new_n26206__;
  assign new_new_n26208__ = ys__n776 & ys__n25300;
  assign new_new_n26209__ = ~new_new_n26207__ & ~new_new_n26208__;
  assign ys__n25390 = ~ys__n4168 & ~new_new_n26209__;
  assign new_new_n26211__ = new_new_n13930__ & new_new_n13933__;
  assign new_new_n26212__ = new_new_n26144__ & new_new_n26211__;
  assign new_new_n26213__ = ys__n25300 & new_new_n15920__;
  assign new_new_n26214__ = new_new_n15902__ & new_new_n26213__;
  assign ys__n25406 = new_new_n26212__ & new_new_n26214__;
  assign new_new_n26216__ = ys__n25300 & new_new_n15900__;
  assign new_new_n26217__ = new_new_n15903__ & new_new_n15909__;
  assign new_new_n26218__ = new_new_n26142__ & new_new_n26217__;
  assign new_new_n26219__ = new_new_n26216__ & new_new_n26218__;
  assign new_new_n26220__ = ys__n4168 & ys__n25300;
  assign ys__n25421 = new_new_n26219__ | new_new_n26220__;
  assign new_new_n26222__ = new_new_n12143__ & ~ys__n18360;
  assign new_new_n26223__ = new_new_n12070__ & new_new_n26222__;
  assign ys__n25430 = new_new_n12127__ & new_new_n26223__;
  assign new_new_n26225__ = ~ys__n19256 & ys__n25386;
  assign new_new_n26226__ = ys__n524 & ys__n19256;
  assign new_new_n26227__ = ~new_new_n26225__ & ~new_new_n26226__;
  assign new_new_n26228__ = ys__n874 & ~new_new_n26227__;
  assign new_new_n26229__ = ~ys__n19256 & ys__n25385;
  assign new_new_n26230__ = ys__n526 & ys__n19256;
  assign new_new_n26231__ = ~new_new_n26229__ & ~new_new_n26230__;
  assign new_new_n26232__ = ys__n874 & ~new_new_n26231__;
  assign new_new_n26233__ = ~ys__n19256 & ys__n25387;
  assign new_new_n26234__ = ys__n522 & ys__n19256;
  assign new_new_n26235__ = ~new_new_n26233__ & ~new_new_n26234__;
  assign new_new_n26236__ = ys__n874 & ~new_new_n26235__;
  assign new_new_n26237__ = ~new_new_n26232__ & new_new_n26236__;
  assign ys__n25431 = ~new_new_n26228__ & new_new_n26237__;
  assign new_new_n26239__ = ys__n604 & ~ys__n776;
  assign new_new_n26240__ = ~ys__n4168 & ~ys__n25300;
  assign ys__n25438 = new_new_n26239__ & new_new_n26240__;
  assign new_new_n26242__ = ~ys__n25300 & new_new_n15937__;
  assign new_new_n26243__ = new_new_n13930__ & new_new_n26242__;
  assign new_new_n26244__ = ys__n602 & ~ys__n25300;
  assign new_new_n26245__ = ~new_new_n26243__ & ~new_new_n26244__;
  assign new_new_n26246__ = ~ys__n778 & ~new_new_n26245__;
  assign new_new_n26247__ = ys__n778 & ~ys__n25300;
  assign new_new_n26248__ = ~new_new_n26246__ & ~new_new_n26247__;
  assign new_new_n26249__ = ~ys__n604 & ~ys__n776;
  assign new_new_n26250__ = ~ys__n4168 & new_new_n26249__;
  assign ys__n25441 = ~new_new_n26248__ & new_new_n26250__;
  assign new_new_n26252__ = ~ys__n600 & ys__n698;
  assign new_new_n26253__ = ~ys__n25300 & new_new_n26252__;
  assign new_new_n26254__ = ys__n600 & ~ys__n25300;
  assign new_new_n26255__ = ~new_new_n26253__ & ~new_new_n26254__;
  assign new_new_n26256__ = ~ys__n602 & ~ys__n604;
  assign new_new_n26257__ = ~ys__n778 & new_new_n15900__;
  assign new_new_n26258__ = new_new_n26256__ & new_new_n26257__;
  assign ys__n25449 = ~new_new_n26255__ & new_new_n26258__;
  assign new_new_n26260__ = ys__n602 & ~ys__n778;
  assign new_new_n26261__ = ys__n25300 & new_new_n26260__;
  assign new_new_n26262__ = ys__n778 & ys__n25300;
  assign new_new_n26263__ = ~new_new_n26261__ & ~new_new_n26262__;
  assign ys__n25456 = new_new_n26250__ & ~new_new_n26263__;
  assign new_new_n26265__ = ys__n25381 & new_new_n15911__;
  assign ys__n25461 = ys__n784 | new_new_n26265__;
  assign ys__n25463 = ys__n25382 & new_new_n15911__;
  assign ys__n25465 = ys__n25383 & new_new_n15911__;
  assign ys__n25467 = ys__n25384 & new_new_n15911__;
  assign ys__n25469 = ys__n25470 & new_new_n15911__;
  assign new_new_n26271__ = ~ys__n25300 & new_new_n15920__;
  assign new_new_n26272__ = ys__n772 & ~ys__n25300;
  assign new_new_n26273__ = ~new_new_n26271__ & ~new_new_n26272__;
  assign new_new_n26274__ = ~ys__n600 & ~ys__n778;
  assign new_new_n26275__ = new_new_n15900__ & new_new_n26274__;
  assign new_new_n26276__ = new_new_n13933__ & new_new_n26256__;
  assign new_new_n26277__ = new_new_n26144__ & new_new_n26276__;
  assign new_new_n26278__ = new_new_n26275__ & new_new_n26277__;
  assign ys__n25472 = ~new_new_n26273__ & new_new_n26278__;
  assign new_new_n26280__ = ~ys__n25300 & new_new_n15900__;
  assign new_new_n26281__ = new_new_n15903__ & new_new_n26274__;
  assign new_new_n26282__ = new_new_n15909__ & new_new_n26256__;
  assign new_new_n26283__ = new_new_n26281__ & new_new_n26282__;
  assign ys__n25486 = new_new_n26280__ & new_new_n26283__;
  assign new_new_n26285__ = ~ys__n600 & ~ys__n698;
  assign new_new_n26286__ = ys__n768 & ys__n25300;
  assign new_new_n26287__ = new_new_n26285__ & new_new_n26286__;
  assign new_new_n26288__ = ys__n600 & ys__n25300;
  assign new_new_n26289__ = ~new_new_n26287__ & ~new_new_n26288__;
  assign ys__n25496 = new_new_n26258__ & ~new_new_n26289__;
  assign new_new_n26291__ = ~ys__n770 & ~ys__n772;
  assign new_new_n26292__ = ~ys__n780 & ys__n782;
  assign new_new_n26293__ = ~ys__n25300 & new_new_n26292__;
  assign new_new_n26294__ = new_new_n26291__ & new_new_n26293__;
  assign new_new_n26295__ = ys__n770 & ~ys__n25300;
  assign new_new_n26296__ = ~new_new_n26294__ & ~new_new_n26295__;
  assign new_new_n26297__ = ~ys__n784 & ~new_new_n26296__;
  assign new_new_n26298__ = ys__n784 & ~ys__n25300;
  assign new_new_n26299__ = ~new_new_n26297__ & ~new_new_n26298__;
  assign new_new_n26300__ = new_new_n15903__ & new_new_n26256__;
  assign new_new_n26301__ = new_new_n13933__ & new_new_n26300__;
  assign new_new_n26302__ = new_new_n26275__ & new_new_n26301__;
  assign ys__n25504 = ~new_new_n26299__ & new_new_n26302__;
  assign new_new_n26304__ = ~ys__n4168 & ys__n25300;
  assign ys__n25519 = new_new_n26239__ & new_new_n26304__;
  assign new_new_n26306__ = ys__n25300 & new_new_n15911__;
  assign new_new_n26307__ = ys__n784 & ys__n25300;
  assign new_new_n26308__ = ~new_new_n26306__ & ~new_new_n26307__;
  assign ys__n25522 = new_new_n26302__ & ~new_new_n26308__;
  assign new_new_n26310__ = ~ys__n782 & ~ys__n784;
  assign new_new_n26311__ = ~ys__n25300 & new_new_n26310__;
  assign new_new_n26312__ = new_new_n26146__ & new_new_n26291__;
  assign new_new_n26313__ = new_new_n13933__ & new_new_n26312__;
  assign new_new_n26314__ = new_new_n26311__ & new_new_n26313__;
  assign new_new_n26315__ = ys__n598 & ~ys__n25300;
  assign new_new_n26316__ = ~new_new_n26314__ & ~new_new_n26315__;
  assign new_new_n26317__ = new_new_n26206__ & ~new_new_n26316__;
  assign new_new_n26318__ = ys__n776 & ~ys__n25300;
  assign new_new_n26319__ = ~new_new_n26317__ & ~new_new_n26318__;
  assign new_new_n26320__ = ~ys__n4168 & ~new_new_n26319__;
  assign new_new_n26321__ = ys__n4168 & ~ys__n25300;
  assign ys__n25534 = new_new_n26320__ | new_new_n26321__;
  assign new_new_n26323__ = ys__n782 & ys__n25300;
  assign new_new_n26324__ = new_new_n15916__ & new_new_n26323__;
  assign new_new_n26325__ = ys__n772 & ys__n25300;
  assign new_new_n26326__ = ~new_new_n26324__ & ~new_new_n26325__;
  assign ys__n25550 = new_new_n26278__ & ~new_new_n26326__;
  assign new_new_n26328__ = ~ys__n778 & ys__n25564;
  assign new_new_n26329__ = ~ys__n326 & ~ys__n332;
  assign new_new_n26330__ = ~ys__n336 & new_new_n12316__;
  assign new_new_n26331__ = new_new_n26329__ & new_new_n26330__;
  assign new_new_n26332__ = ys__n25564 & ~new_new_n26331__;
  assign new_new_n26333__ = ~new_new_n26331__ & ~new_new_n26332__;
  assign new_new_n26334__ = ys__n778 & ~new_new_n26333__;
  assign new_new_n26335__ = ~new_new_n26328__ & ~new_new_n26334__;
  assign new_new_n26336__ = ~ys__n602 & ~new_new_n26335__;
  assign new_new_n26337__ = ys__n25567 & new_new_n26331__;
  assign new_new_n26338__ = ~new_new_n26331__ & ~new_new_n26335__;
  assign new_new_n26339__ = ~new_new_n26337__ & ~new_new_n26338__;
  assign new_new_n26340__ = ys__n602 & ~new_new_n26339__;
  assign ys__n25661 = new_new_n26336__ | new_new_n26340__;
  assign new_new_n26342__ = ~ys__n778 & ys__n25567;
  assign new_new_n26343__ = ys__n778 & ys__n25567;
  assign new_new_n26344__ = ~new_new_n26331__ & new_new_n26343__;
  assign new_new_n26345__ = ~new_new_n26342__ & ~new_new_n26344__;
  assign new_new_n26346__ = ~ys__n602 & ~new_new_n26345__;
  assign new_new_n26347__ = ys__n25570 & new_new_n26331__;
  assign new_new_n26348__ = ~new_new_n26331__ & ~new_new_n26345__;
  assign new_new_n26349__ = ~new_new_n26347__ & ~new_new_n26348__;
  assign new_new_n26350__ = ys__n602 & ~new_new_n26349__;
  assign ys__n25663 = new_new_n26346__ | new_new_n26350__;
  assign new_new_n26352__ = ~ys__n778 & ys__n25570;
  assign new_new_n26353__ = ys__n25570 & ~new_new_n26331__;
  assign new_new_n26354__ = ~new_new_n26331__ & ~new_new_n26353__;
  assign new_new_n26355__ = ys__n778 & ~new_new_n26354__;
  assign new_new_n26356__ = ~new_new_n26352__ & ~new_new_n26355__;
  assign new_new_n26357__ = ~ys__n602 & ~new_new_n26356__;
  assign new_new_n26358__ = ys__n25573 & new_new_n26331__;
  assign new_new_n26359__ = ~new_new_n26331__ & ~new_new_n26356__;
  assign new_new_n26360__ = ~new_new_n26358__ & ~new_new_n26359__;
  assign new_new_n26361__ = ys__n602 & ~new_new_n26360__;
  assign ys__n25665 = new_new_n26357__ | new_new_n26361__;
  assign new_new_n26363__ = ~ys__n778 & ys__n25573;
  assign new_new_n26364__ = ys__n25573 & ~new_new_n26331__;
  assign new_new_n26365__ = ~new_new_n26331__ & ~new_new_n26364__;
  assign new_new_n26366__ = ys__n778 & ~new_new_n26365__;
  assign new_new_n26367__ = ~new_new_n26363__ & ~new_new_n26366__;
  assign new_new_n26368__ = ~ys__n602 & ~new_new_n26367__;
  assign new_new_n26369__ = ys__n25576 & new_new_n26331__;
  assign new_new_n26370__ = ~new_new_n26331__ & ~new_new_n26367__;
  assign new_new_n26371__ = ~new_new_n26369__ & ~new_new_n26370__;
  assign new_new_n26372__ = ys__n602 & ~new_new_n26371__;
  assign ys__n25667 = new_new_n26368__ | new_new_n26372__;
  assign new_new_n26374__ = ~ys__n778 & ys__n25576;
  assign new_new_n26375__ = ys__n778 & ys__n25576;
  assign new_new_n26376__ = ~new_new_n26331__ & new_new_n26375__;
  assign new_new_n26377__ = ~new_new_n26374__ & ~new_new_n26376__;
  assign new_new_n26378__ = ~ys__n602 & ~new_new_n26377__;
  assign new_new_n26379__ = ys__n25579 & new_new_n26331__;
  assign new_new_n26380__ = ~new_new_n26331__ & ~new_new_n26377__;
  assign new_new_n26381__ = ~new_new_n26379__ & ~new_new_n26380__;
  assign new_new_n26382__ = ys__n602 & ~new_new_n26381__;
  assign ys__n25669 = new_new_n26378__ | new_new_n26382__;
  assign new_new_n26384__ = ~ys__n778 & ys__n25579;
  assign new_new_n26385__ = ys__n778 & ys__n25579;
  assign new_new_n26386__ = ~new_new_n26331__ & new_new_n26385__;
  assign new_new_n26387__ = ~new_new_n26384__ & ~new_new_n26386__;
  assign new_new_n26388__ = ~ys__n602 & ~new_new_n26387__;
  assign new_new_n26389__ = ys__n25582 & new_new_n26331__;
  assign new_new_n26390__ = ~new_new_n26331__ & ~new_new_n26387__;
  assign new_new_n26391__ = ~new_new_n26389__ & ~new_new_n26390__;
  assign new_new_n26392__ = ys__n602 & ~new_new_n26391__;
  assign ys__n25671 = new_new_n26388__ | new_new_n26392__;
  assign new_new_n26394__ = ~ys__n778 & ys__n25582;
  assign new_new_n26395__ = ys__n778 & ys__n25582;
  assign new_new_n26396__ = ~new_new_n26331__ & new_new_n26395__;
  assign new_new_n26397__ = ~new_new_n26394__ & ~new_new_n26396__;
  assign new_new_n26398__ = ~ys__n602 & ~new_new_n26397__;
  assign new_new_n26399__ = ys__n25585 & new_new_n26331__;
  assign new_new_n26400__ = ~new_new_n26331__ & ~new_new_n26397__;
  assign new_new_n26401__ = ~new_new_n26399__ & ~new_new_n26400__;
  assign new_new_n26402__ = ys__n602 & ~new_new_n26401__;
  assign ys__n25673 = new_new_n26398__ | new_new_n26402__;
  assign new_new_n26404__ = ~ys__n778 & ys__n25585;
  assign new_new_n26405__ = ys__n778 & ys__n25585;
  assign new_new_n26406__ = ~new_new_n26331__ & new_new_n26405__;
  assign new_new_n26407__ = ~new_new_n26404__ & ~new_new_n26406__;
  assign new_new_n26408__ = ~ys__n602 & ~new_new_n26407__;
  assign new_new_n26409__ = ys__n25588 & new_new_n26331__;
  assign new_new_n26410__ = ~new_new_n26331__ & ~new_new_n26407__;
  assign new_new_n26411__ = ~new_new_n26409__ & ~new_new_n26410__;
  assign new_new_n26412__ = ys__n602 & ~new_new_n26411__;
  assign ys__n25675 = new_new_n26408__ | new_new_n26412__;
  assign new_new_n26414__ = ~ys__n778 & ys__n25588;
  assign new_new_n26415__ = ys__n778 & ys__n25588;
  assign new_new_n26416__ = ~new_new_n26331__ & new_new_n26415__;
  assign new_new_n26417__ = ~new_new_n26414__ & ~new_new_n26416__;
  assign new_new_n26418__ = ~ys__n602 & ~new_new_n26417__;
  assign new_new_n26419__ = ys__n25591 & new_new_n26331__;
  assign new_new_n26420__ = ~new_new_n26331__ & ~new_new_n26417__;
  assign new_new_n26421__ = ~new_new_n26419__ & ~new_new_n26420__;
  assign new_new_n26422__ = ys__n602 & ~new_new_n26421__;
  assign ys__n25677 = new_new_n26418__ | new_new_n26422__;
  assign new_new_n26424__ = ~ys__n778 & ys__n25591;
  assign new_new_n26425__ = ys__n778 & ys__n25591;
  assign new_new_n26426__ = ~new_new_n26331__ & new_new_n26425__;
  assign new_new_n26427__ = ~new_new_n26424__ & ~new_new_n26426__;
  assign new_new_n26428__ = ~ys__n602 & ~new_new_n26427__;
  assign new_new_n26429__ = ys__n25594 & new_new_n26331__;
  assign new_new_n26430__ = ~new_new_n26331__ & ~new_new_n26427__;
  assign new_new_n26431__ = ~new_new_n26429__ & ~new_new_n26430__;
  assign new_new_n26432__ = ys__n602 & ~new_new_n26431__;
  assign ys__n25679 = new_new_n26428__ | new_new_n26432__;
  assign new_new_n26434__ = ~ys__n778 & ys__n25594;
  assign new_new_n26435__ = ys__n778 & ys__n25594;
  assign new_new_n26436__ = ~new_new_n26331__ & new_new_n26435__;
  assign new_new_n26437__ = ~new_new_n26434__ & ~new_new_n26436__;
  assign new_new_n26438__ = ~ys__n602 & ~new_new_n26437__;
  assign new_new_n26439__ = ys__n25597 & new_new_n26331__;
  assign new_new_n26440__ = ~new_new_n26331__ & ~new_new_n26437__;
  assign new_new_n26441__ = ~new_new_n26439__ & ~new_new_n26440__;
  assign new_new_n26442__ = ys__n602 & ~new_new_n26441__;
  assign ys__n25681 = new_new_n26438__ | new_new_n26442__;
  assign new_new_n26444__ = ~ys__n778 & ys__n25597;
  assign new_new_n26445__ = ys__n778 & ys__n25597;
  assign new_new_n26446__ = ~new_new_n26331__ & new_new_n26445__;
  assign new_new_n26447__ = ~new_new_n26444__ & ~new_new_n26446__;
  assign new_new_n26448__ = ~ys__n602 & ~new_new_n26447__;
  assign new_new_n26449__ = ys__n25600 & new_new_n26331__;
  assign new_new_n26450__ = ~new_new_n26331__ & ~new_new_n26447__;
  assign new_new_n26451__ = ~new_new_n26449__ & ~new_new_n26450__;
  assign new_new_n26452__ = ys__n602 & ~new_new_n26451__;
  assign ys__n25683 = new_new_n26448__ | new_new_n26452__;
  assign new_new_n26454__ = ~ys__n778 & ys__n25600;
  assign new_new_n26455__ = ys__n778 & ys__n25600;
  assign new_new_n26456__ = ~new_new_n26331__ & new_new_n26455__;
  assign new_new_n26457__ = ~new_new_n26454__ & ~new_new_n26456__;
  assign new_new_n26458__ = ~ys__n602 & ~new_new_n26457__;
  assign new_new_n26459__ = ys__n25603 & new_new_n26331__;
  assign new_new_n26460__ = ~new_new_n26331__ & ~new_new_n26457__;
  assign new_new_n26461__ = ~new_new_n26459__ & ~new_new_n26460__;
  assign new_new_n26462__ = ys__n602 & ~new_new_n26461__;
  assign ys__n25685 = new_new_n26458__ | new_new_n26462__;
  assign new_new_n26464__ = ~ys__n778 & ys__n25603;
  assign new_new_n26465__ = ys__n778 & ys__n25603;
  assign new_new_n26466__ = ~new_new_n26331__ & new_new_n26465__;
  assign new_new_n26467__ = ~new_new_n26464__ & ~new_new_n26466__;
  assign new_new_n26468__ = ~ys__n602 & ~new_new_n26467__;
  assign new_new_n26469__ = ys__n25606 & new_new_n26331__;
  assign new_new_n26470__ = ~new_new_n26331__ & ~new_new_n26467__;
  assign new_new_n26471__ = ~new_new_n26469__ & ~new_new_n26470__;
  assign new_new_n26472__ = ys__n602 & ~new_new_n26471__;
  assign ys__n25687 = new_new_n26468__ | new_new_n26472__;
  assign new_new_n26474__ = ~ys__n778 & ys__n25606;
  assign new_new_n26475__ = ys__n778 & ys__n25606;
  assign new_new_n26476__ = ~new_new_n26331__ & new_new_n26475__;
  assign new_new_n26477__ = ~new_new_n26474__ & ~new_new_n26476__;
  assign new_new_n26478__ = ~ys__n602 & ~new_new_n26477__;
  assign new_new_n26479__ = ys__n25609 & new_new_n26331__;
  assign new_new_n26480__ = ~new_new_n26331__ & ~new_new_n26477__;
  assign new_new_n26481__ = ~new_new_n26479__ & ~new_new_n26480__;
  assign new_new_n26482__ = ys__n602 & ~new_new_n26481__;
  assign ys__n25689 = new_new_n26478__ | new_new_n26482__;
  assign new_new_n26484__ = ~ys__n778 & ys__n25609;
  assign new_new_n26485__ = ys__n778 & ys__n25609;
  assign new_new_n26486__ = ~new_new_n26331__ & new_new_n26485__;
  assign new_new_n26487__ = ~new_new_n26484__ & ~new_new_n26486__;
  assign new_new_n26488__ = ~ys__n602 & ~new_new_n26487__;
  assign new_new_n26489__ = ys__n25612 & new_new_n26331__;
  assign new_new_n26490__ = ~new_new_n26331__ & ~new_new_n26487__;
  assign new_new_n26491__ = ~new_new_n26489__ & ~new_new_n26490__;
  assign new_new_n26492__ = ys__n602 & ~new_new_n26491__;
  assign ys__n25691 = new_new_n26488__ | new_new_n26492__;
  assign new_new_n26494__ = ~ys__n778 & ys__n25612;
  assign new_new_n26495__ = ys__n778 & ys__n25612;
  assign new_new_n26496__ = ~new_new_n26331__ & new_new_n26495__;
  assign new_new_n26497__ = ~new_new_n26494__ & ~new_new_n26496__;
  assign new_new_n26498__ = ~ys__n602 & ~new_new_n26497__;
  assign new_new_n26499__ = ys__n25615 & new_new_n26331__;
  assign new_new_n26500__ = ~new_new_n26331__ & ~new_new_n26497__;
  assign new_new_n26501__ = ~new_new_n26499__ & ~new_new_n26500__;
  assign new_new_n26502__ = ys__n602 & ~new_new_n26501__;
  assign ys__n25693 = new_new_n26498__ | new_new_n26502__;
  assign new_new_n26504__ = ~ys__n778 & ys__n25615;
  assign new_new_n26505__ = ys__n778 & ys__n25615;
  assign new_new_n26506__ = ~new_new_n26331__ & new_new_n26505__;
  assign new_new_n26507__ = ~new_new_n26504__ & ~new_new_n26506__;
  assign new_new_n26508__ = ~ys__n602 & ~new_new_n26507__;
  assign new_new_n26509__ = ys__n25618 & new_new_n26331__;
  assign new_new_n26510__ = ~new_new_n26331__ & ~new_new_n26507__;
  assign new_new_n26511__ = ~new_new_n26509__ & ~new_new_n26510__;
  assign new_new_n26512__ = ys__n602 & ~new_new_n26511__;
  assign ys__n25695 = new_new_n26508__ | new_new_n26512__;
  assign new_new_n26514__ = ~ys__n778 & ys__n25618;
  assign new_new_n26515__ = ys__n778 & ys__n25618;
  assign new_new_n26516__ = ~new_new_n26331__ & new_new_n26515__;
  assign new_new_n26517__ = ~new_new_n26514__ & ~new_new_n26516__;
  assign new_new_n26518__ = ~ys__n602 & ~new_new_n26517__;
  assign new_new_n26519__ = ys__n25621 & new_new_n26331__;
  assign new_new_n26520__ = ~new_new_n26331__ & ~new_new_n26517__;
  assign new_new_n26521__ = ~new_new_n26519__ & ~new_new_n26520__;
  assign new_new_n26522__ = ys__n602 & ~new_new_n26521__;
  assign ys__n25697 = new_new_n26518__ | new_new_n26522__;
  assign new_new_n26524__ = ~ys__n778 & ys__n25621;
  assign new_new_n26525__ = ys__n25621 & ~new_new_n26331__;
  assign new_new_n26526__ = ~new_new_n26331__ & ~new_new_n26525__;
  assign new_new_n26527__ = ys__n778 & ~new_new_n26526__;
  assign new_new_n26528__ = ~new_new_n26524__ & ~new_new_n26527__;
  assign new_new_n26529__ = ~ys__n602 & ~new_new_n26528__;
  assign new_new_n26530__ = ys__n25624 & new_new_n26331__;
  assign new_new_n26531__ = ~new_new_n26331__ & ~new_new_n26528__;
  assign new_new_n26532__ = ~new_new_n26530__ & ~new_new_n26531__;
  assign new_new_n26533__ = ys__n602 & ~new_new_n26532__;
  assign ys__n25699 = new_new_n26529__ | new_new_n26533__;
  assign new_new_n26535__ = ~ys__n778 & ys__n25624;
  assign new_new_n26536__ = ys__n25624 & ~new_new_n26331__;
  assign new_new_n26537__ = ~new_new_n26331__ & ~new_new_n26536__;
  assign new_new_n26538__ = ys__n778 & ~new_new_n26537__;
  assign new_new_n26539__ = ~new_new_n26535__ & ~new_new_n26538__;
  assign new_new_n26540__ = ~ys__n602 & ~new_new_n26539__;
  assign new_new_n26541__ = ys__n25627 & new_new_n26331__;
  assign new_new_n26542__ = ~new_new_n26331__ & ~new_new_n26539__;
  assign new_new_n26543__ = ~new_new_n26541__ & ~new_new_n26542__;
  assign new_new_n26544__ = ys__n602 & ~new_new_n26543__;
  assign ys__n25701 = new_new_n26540__ | new_new_n26544__;
  assign new_new_n26546__ = ~ys__n778 & ys__n25627;
  assign new_new_n26547__ = ys__n778 & ys__n25627;
  assign new_new_n26548__ = ~new_new_n26331__ & new_new_n26547__;
  assign new_new_n26549__ = ~new_new_n26546__ & ~new_new_n26548__;
  assign new_new_n26550__ = ~ys__n602 & ~new_new_n26549__;
  assign new_new_n26551__ = ys__n25630 & new_new_n26331__;
  assign new_new_n26552__ = ~new_new_n26331__ & ~new_new_n26549__;
  assign new_new_n26553__ = ~new_new_n26551__ & ~new_new_n26552__;
  assign new_new_n26554__ = ys__n602 & ~new_new_n26553__;
  assign ys__n25703 = new_new_n26550__ | new_new_n26554__;
  assign new_new_n26556__ = ~ys__n778 & ys__n25630;
  assign new_new_n26557__ = ys__n778 & ys__n25630;
  assign new_new_n26558__ = ~new_new_n26331__ & new_new_n26557__;
  assign new_new_n26559__ = ~new_new_n26556__ & ~new_new_n26558__;
  assign new_new_n26560__ = ~ys__n602 & ~new_new_n26559__;
  assign new_new_n26561__ = ys__n25633 & new_new_n26331__;
  assign new_new_n26562__ = ~new_new_n26331__ & ~new_new_n26559__;
  assign new_new_n26563__ = ~new_new_n26561__ & ~new_new_n26562__;
  assign new_new_n26564__ = ys__n602 & ~new_new_n26563__;
  assign ys__n25705 = new_new_n26560__ | new_new_n26564__;
  assign new_new_n26566__ = ~ys__n778 & ys__n25633;
  assign new_new_n26567__ = ys__n778 & ys__n25633;
  assign new_new_n26568__ = ~new_new_n26331__ & new_new_n26567__;
  assign new_new_n26569__ = ~new_new_n26566__ & ~new_new_n26568__;
  assign new_new_n26570__ = ~ys__n602 & ~new_new_n26569__;
  assign new_new_n26571__ = ys__n25636 & new_new_n26331__;
  assign new_new_n26572__ = ~new_new_n26331__ & ~new_new_n26569__;
  assign new_new_n26573__ = ~new_new_n26571__ & ~new_new_n26572__;
  assign new_new_n26574__ = ys__n602 & ~new_new_n26573__;
  assign ys__n25707 = new_new_n26570__ | new_new_n26574__;
  assign new_new_n26576__ = ~ys__n778 & ys__n25636;
  assign new_new_n26577__ = ys__n778 & ys__n25636;
  assign new_new_n26578__ = ~new_new_n26331__ & new_new_n26577__;
  assign new_new_n26579__ = ~new_new_n26576__ & ~new_new_n26578__;
  assign new_new_n26580__ = ~ys__n602 & ~new_new_n26579__;
  assign new_new_n26581__ = ys__n25639 & new_new_n26331__;
  assign new_new_n26582__ = ~new_new_n26331__ & ~new_new_n26579__;
  assign new_new_n26583__ = ~new_new_n26581__ & ~new_new_n26582__;
  assign new_new_n26584__ = ys__n602 & ~new_new_n26583__;
  assign ys__n25709 = new_new_n26580__ | new_new_n26584__;
  assign new_new_n26586__ = ~ys__n778 & ys__n25639;
  assign new_new_n26587__ = ys__n778 & ys__n25639;
  assign new_new_n26588__ = ~new_new_n26331__ & new_new_n26587__;
  assign new_new_n26589__ = ~new_new_n26586__ & ~new_new_n26588__;
  assign new_new_n26590__ = ~ys__n602 & ~new_new_n26589__;
  assign new_new_n26591__ = ys__n25642 & new_new_n26331__;
  assign new_new_n26592__ = ~new_new_n26331__ & ~new_new_n26589__;
  assign new_new_n26593__ = ~new_new_n26591__ & ~new_new_n26592__;
  assign new_new_n26594__ = ys__n602 & ~new_new_n26593__;
  assign ys__n25711 = new_new_n26590__ | new_new_n26594__;
  assign new_new_n26596__ = ~ys__n778 & ys__n25642;
  assign new_new_n26597__ = ys__n25642 & ~new_new_n26331__;
  assign new_new_n26598__ = ~new_new_n26331__ & ~new_new_n26597__;
  assign new_new_n26599__ = ys__n778 & ~new_new_n26598__;
  assign new_new_n26600__ = ~new_new_n26596__ & ~new_new_n26599__;
  assign new_new_n26601__ = ~ys__n602 & ~new_new_n26600__;
  assign new_new_n26602__ = ys__n25645 & new_new_n26331__;
  assign new_new_n26603__ = ~new_new_n26331__ & ~new_new_n26600__;
  assign new_new_n26604__ = ~new_new_n26602__ & ~new_new_n26603__;
  assign new_new_n26605__ = ys__n602 & ~new_new_n26604__;
  assign ys__n25713 = new_new_n26601__ | new_new_n26605__;
  assign new_new_n26607__ = ~ys__n778 & ys__n25645;
  assign new_new_n26608__ = ys__n778 & ys__n25645;
  assign new_new_n26609__ = ~new_new_n26331__ & new_new_n26608__;
  assign new_new_n26610__ = ~new_new_n26607__ & ~new_new_n26609__;
  assign new_new_n26611__ = ~ys__n602 & ~new_new_n26610__;
  assign new_new_n26612__ = ys__n25648 & new_new_n26331__;
  assign new_new_n26613__ = ~new_new_n26331__ & ~new_new_n26610__;
  assign new_new_n26614__ = ~new_new_n26612__ & ~new_new_n26613__;
  assign new_new_n26615__ = ys__n602 & ~new_new_n26614__;
  assign ys__n25715 = new_new_n26611__ | new_new_n26615__;
  assign new_new_n26617__ = ~ys__n778 & ys__n25648;
  assign new_new_n26618__ = ys__n778 & ys__n25648;
  assign new_new_n26619__ = ~new_new_n26331__ & new_new_n26618__;
  assign new_new_n26620__ = ~new_new_n26617__ & ~new_new_n26619__;
  assign new_new_n26621__ = ~ys__n602 & ~new_new_n26620__;
  assign new_new_n26622__ = ys__n25651 & new_new_n26331__;
  assign new_new_n26623__ = ~new_new_n26331__ & ~new_new_n26620__;
  assign new_new_n26624__ = ~new_new_n26622__ & ~new_new_n26623__;
  assign new_new_n26625__ = ys__n602 & ~new_new_n26624__;
  assign ys__n25717 = new_new_n26621__ | new_new_n26625__;
  assign new_new_n26627__ = ~ys__n778 & ys__n25651;
  assign new_new_n26628__ = ys__n25651 & ~new_new_n26331__;
  assign new_new_n26629__ = ~new_new_n26331__ & ~new_new_n26628__;
  assign new_new_n26630__ = ys__n778 & ~new_new_n26629__;
  assign new_new_n26631__ = ~new_new_n26627__ & ~new_new_n26630__;
  assign new_new_n26632__ = ~ys__n602 & ~new_new_n26631__;
  assign new_new_n26633__ = ys__n25654 & new_new_n26331__;
  assign new_new_n26634__ = ~new_new_n26331__ & ~new_new_n26631__;
  assign new_new_n26635__ = ~new_new_n26633__ & ~new_new_n26634__;
  assign new_new_n26636__ = ys__n602 & ~new_new_n26635__;
  assign ys__n25719 = new_new_n26632__ | new_new_n26636__;
  assign new_new_n26638__ = ~ys__n778 & ys__n25654;
  assign new_new_n26639__ = ys__n778 & ys__n25654;
  assign new_new_n26640__ = ~new_new_n26331__ & new_new_n26639__;
  assign new_new_n26641__ = ~new_new_n26638__ & ~new_new_n26640__;
  assign new_new_n26642__ = ~ys__n602 & ~new_new_n26641__;
  assign new_new_n26643__ = ys__n25657 & new_new_n26331__;
  assign new_new_n26644__ = ~new_new_n26331__ & ~new_new_n26641__;
  assign new_new_n26645__ = ~new_new_n26643__ & ~new_new_n26644__;
  assign new_new_n26646__ = ys__n602 & ~new_new_n26645__;
  assign ys__n25721 = new_new_n26642__ | new_new_n26646__;
  assign new_new_n26648__ = ~ys__n778 & ys__n25657;
  assign new_new_n26649__ = ys__n778 & ys__n25657;
  assign new_new_n26650__ = ~new_new_n26331__ & new_new_n26649__;
  assign new_new_n26651__ = ~new_new_n26648__ & ~new_new_n26650__;
  assign new_new_n26652__ = ~ys__n602 & ~new_new_n26651__;
  assign new_new_n26653__ = ys__n25470 & new_new_n26331__;
  assign new_new_n26654__ = ~new_new_n26331__ & ~new_new_n26651__;
  assign new_new_n26655__ = ~new_new_n26653__ & ~new_new_n26654__;
  assign new_new_n26656__ = ys__n602 & ~new_new_n26655__;
  assign ys__n25723 = new_new_n26652__ | new_new_n26656__;
  assign new_new_n26658__ = ys__n25292 & new_new_n26274__;
  assign new_new_n26659__ = new_new_n15900__ & new_new_n15911__;
  assign new_new_n26660__ = new_new_n26658__ & new_new_n26659__;
  assign new_new_n26661__ = new_new_n26301__ & new_new_n26660__;
  assign new_new_n26662__ = ~ys__n336 & new_new_n12320__;
  assign new_new_n26663__ = new_new_n26329__ & new_new_n26662__;
  assign new_new_n26664__ = ys__n336 & new_new_n16713__;
  assign new_new_n26665__ = ys__n336 & new_new_n16711__;
  assign new_new_n26666__ = ~new_new_n26664__ & ~new_new_n26665__;
  assign new_new_n26667__ = ~new_new_n26663__ & new_new_n26666__;
  assign new_new_n26668__ = new_new_n12313__ & new_new_n26329__;
  assign new_new_n26669__ = ~ys__n336 & new_new_n26668__;
  assign new_new_n26670__ = ~new_new_n26331__ & ~new_new_n26669__;
  assign new_new_n26671__ = ys__n336 & new_new_n16721__;
  assign new_new_n26672__ = ys__n336 & new_new_n16726__;
  assign new_new_n26673__ = ~new_new_n26671__ & ~new_new_n26672__;
  assign new_new_n26674__ = new_new_n26670__ & new_new_n26673__;
  assign new_new_n26675__ = new_new_n26667__ & new_new_n26674__;
  assign new_new_n26676__ = new_new_n12329__ & new_new_n26675__;
  assign new_new_n26677__ = ~ys__n336 & new_new_n12322__;
  assign new_new_n26678__ = new_new_n26329__ & new_new_n26677__;
  assign new_new_n26679__ = ~new_new_n16727__ & ~new_new_n26678__;
  assign new_new_n26680__ = ys__n25980 & ~new_new_n26679__;
  assign new_new_n26681__ = ys__n26425 & ~new_new_n16715__;
  assign new_new_n26682__ = ys__n26359 & new_new_n16722__;
  assign new_new_n26683__ = ~new_new_n26681__ & ~new_new_n26682__;
  assign new_new_n26684__ = ~new_new_n26680__ & new_new_n26683__;
  assign new_new_n26685__ = new_new_n16715__ & ~new_new_n16722__;
  assign new_new_n26686__ = new_new_n26679__ & new_new_n26685__;
  assign new_new_n26687__ = ~new_new_n26684__ & ~new_new_n26686__;
  assign new_new_n26688__ = new_new_n26676__ & new_new_n26687__;
  assign new_new_n26689__ = ys__n25564 & new_new_n26331__;
  assign new_new_n26690__ = ys__n46955 & ~new_new_n12329__;
  assign new_new_n26691__ = ~new_new_n26689__ & ~new_new_n26690__;
  assign new_new_n26692__ = ~new_new_n26676__ & ~new_new_n26691__;
  assign new_new_n26693__ = ~new_new_n26688__ & ~new_new_n26692__;
  assign new_new_n26694__ = ys__n602 & ~new_new_n26693__;
  assign ys__n25725 = new_new_n26661__ | new_new_n26694__;
  assign new_new_n26696__ = ~ys__n25727 & ~ys__n44988;
  assign new_new_n26697__ = ys__n18317 & new_new_n12242__;
  assign new_new_n26698__ = new_new_n14017__ & new_new_n26697__;
  assign new_new_n26699__ = new_new_n14016__ & new_new_n26698__;
  assign new_new_n26700__ = new_new_n14014__ & new_new_n26699__;
  assign new_new_n26701__ = new_new_n12285__ & new_new_n26700__;
  assign new_new_n26702__ = ~new_new_n26696__ & ~new_new_n26701__;
  assign new_new_n26703__ = ~ys__n18208 & ys__n18210;
  assign new_new_n26704__ = ~new_new_n26696__ & ~new_new_n26703__;
  assign new_new_n26705__ = ys__n18448 & new_new_n26703__;
  assign new_new_n26706__ = ~new_new_n26704__ & ~new_new_n26705__;
  assign new_new_n26707__ = new_new_n26701__ & ~new_new_n26706__;
  assign ys__n25830 = new_new_n26702__ | new_new_n26707__;
  assign new_new_n26709__ = ~ys__n25730 & ~ys__n44989;
  assign new_new_n26710__ = ~new_new_n26701__ & ~new_new_n26709__;
  assign new_new_n26711__ = ~new_new_n26703__ & ~new_new_n26709__;
  assign new_new_n26712__ = ys__n18451 & new_new_n26703__;
  assign new_new_n26713__ = ~new_new_n26711__ & ~new_new_n26712__;
  assign new_new_n26714__ = new_new_n26701__ & ~new_new_n26713__;
  assign ys__n25833 = new_new_n26710__ | new_new_n26714__;
  assign new_new_n26716__ = ~ys__n25733 & ~ys__n44990;
  assign new_new_n26717__ = ~new_new_n26701__ & ~new_new_n26716__;
  assign new_new_n26718__ = ~new_new_n26703__ & ~new_new_n26716__;
  assign new_new_n26719__ = ys__n18454 & new_new_n26703__;
  assign new_new_n26720__ = ~new_new_n26718__ & ~new_new_n26719__;
  assign new_new_n26721__ = new_new_n26701__ & ~new_new_n26720__;
  assign ys__n25836 = new_new_n26717__ | new_new_n26721__;
  assign new_new_n26723__ = ~ys__n25736 & ~ys__n44991;
  assign new_new_n26724__ = ~new_new_n26701__ & ~new_new_n26723__;
  assign new_new_n26725__ = ~new_new_n26703__ & ~new_new_n26723__;
  assign new_new_n26726__ = ys__n18457 & new_new_n26703__;
  assign new_new_n26727__ = ~new_new_n26725__ & ~new_new_n26726__;
  assign new_new_n26728__ = new_new_n26701__ & ~new_new_n26727__;
  assign ys__n25839 = new_new_n26724__ | new_new_n26728__;
  assign ys__n25842 = new_new_n13876__ & ~new_new_n13883__;
  assign ys__n25844 = new_new_n13566__ & ~new_new_n13883__;
  assign ys__n25846 = new_new_n13255__ & ~new_new_n13883__;
  assign ys__n25852 = new_new_n12945__ & ~new_new_n13883__;
  assign new_new_n26734__ = ~ys__n25853 & ~ys__n45707;
  assign new_new_n26735__ = ys__n18317 & new_new_n12250__;
  assign new_new_n26736__ = new_new_n14017__ & new_new_n26735__;
  assign new_new_n26737__ = new_new_n14016__ & new_new_n26736__;
  assign new_new_n26738__ = new_new_n14014__ & new_new_n26737__;
  assign new_new_n26739__ = new_new_n12285__ & new_new_n26738__;
  assign new_new_n26740__ = ~new_new_n26734__ & ~new_new_n26739__;
  assign new_new_n26741__ = ~new_new_n26703__ & ~new_new_n26734__;
  assign new_new_n26742__ = ~new_new_n26705__ & ~new_new_n26741__;
  assign new_new_n26743__ = new_new_n26739__ & ~new_new_n26742__;
  assign ys__n25957 = new_new_n26740__ | new_new_n26743__;
  assign new_new_n26745__ = ~ys__n25856 & ~ys__n45708;
  assign new_new_n26746__ = ~new_new_n26739__ & ~new_new_n26745__;
  assign new_new_n26747__ = ~new_new_n26703__ & ~new_new_n26745__;
  assign new_new_n26748__ = ~new_new_n26712__ & ~new_new_n26747__;
  assign new_new_n26749__ = new_new_n26739__ & ~new_new_n26748__;
  assign ys__n25960 = new_new_n26746__ | new_new_n26749__;
  assign new_new_n26751__ = ~ys__n25859 & ~ys__n45709;
  assign new_new_n26752__ = ~new_new_n26739__ & ~new_new_n26751__;
  assign new_new_n26753__ = ~new_new_n26703__ & ~new_new_n26751__;
  assign new_new_n26754__ = ~new_new_n26719__ & ~new_new_n26753__;
  assign new_new_n26755__ = new_new_n26739__ & ~new_new_n26754__;
  assign ys__n25963 = new_new_n26752__ | new_new_n26755__;
  assign new_new_n26757__ = ~ys__n25862 & ~ys__n45710;
  assign new_new_n26758__ = ~new_new_n26739__ & ~new_new_n26757__;
  assign new_new_n26759__ = ~new_new_n26703__ & ~new_new_n26757__;
  assign new_new_n26760__ = ~new_new_n26726__ & ~new_new_n26759__;
  assign new_new_n26761__ = new_new_n26739__ & ~new_new_n26760__;
  assign ys__n25966 = new_new_n26758__ | new_new_n26761__;
  assign new_new_n26763__ = ys__n18317 & new_new_n12240__;
  assign new_new_n26764__ = new_new_n14017__ & new_new_n26763__;
  assign new_new_n26765__ = new_new_n14016__ & new_new_n26764__;
  assign new_new_n26766__ = new_new_n14014__ & new_new_n26765__;
  assign new_new_n26767__ = new_new_n12285__ & new_new_n26766__;
  assign new_new_n26768__ = ~new_new_n12365__ & ~new_new_n26767__;
  assign new_new_n26769__ = ys__n26002 & new_new_n26768__;
  assign new_new_n26770__ = ys__n18041 & new_new_n12356__;
  assign new_new_n26771__ = ys__n18047 & new_new_n12248__;
  assign new_new_n26772__ = ~new_new_n26770__ & ~new_new_n26771__;
  assign new_new_n26773__ = ys__n18053 & new_new_n12245__;
  assign new_new_n26774__ = ys__n18061 & new_new_n12246__;
  assign new_new_n26775__ = ~new_new_n26773__ & ~new_new_n26774__;
  assign new_new_n26776__ = new_new_n26772__ & new_new_n26775__;
  assign new_new_n26777__ = ~new_new_n12248__ & ~new_new_n12356__;
  assign new_new_n26778__ = new_new_n12247__ & new_new_n26777__;
  assign new_new_n26779__ = new_new_n12240__ & ~new_new_n26778__;
  assign new_new_n26780__ = ~new_new_n26776__ & new_new_n26779__;
  assign new_new_n26781__ = ys__n46266 & new_new_n12356__;
  assign new_new_n26782__ = ys__n46442 & new_new_n12248__;
  assign new_new_n26783__ = ~new_new_n26781__ & ~new_new_n26782__;
  assign new_new_n26784__ = ys__n46618 & new_new_n12245__;
  assign new_new_n26785__ = ys__n46794 & new_new_n12246__;
  assign new_new_n26786__ = ~new_new_n26784__ & ~new_new_n26785__;
  assign new_new_n26787__ = new_new_n26783__ & new_new_n26786__;
  assign new_new_n26788__ = new_new_n12242__ & ~new_new_n26778__;
  assign new_new_n26789__ = ~new_new_n26787__ & new_new_n26788__;
  assign new_new_n26790__ = ~new_new_n26780__ & ~new_new_n26789__;
  assign new_new_n26791__ = ys__n46322 & new_new_n12356__;
  assign new_new_n26792__ = ys__n46498 & new_new_n12248__;
  assign new_new_n26793__ = ~new_new_n26791__ & ~new_new_n26792__;
  assign new_new_n26794__ = ys__n46674 & new_new_n12245__;
  assign new_new_n26795__ = ys__n46850 & new_new_n12246__;
  assign new_new_n26796__ = ~new_new_n26794__ & ~new_new_n26795__;
  assign new_new_n26797__ = new_new_n26793__ & new_new_n26796__;
  assign new_new_n26798__ = new_new_n12250__ & ~new_new_n26778__;
  assign new_new_n26799__ = ~new_new_n26797__ & new_new_n26798__;
  assign new_new_n26800__ = ys__n46399 & new_new_n12356__;
  assign new_new_n26801__ = ys__n46575 & new_new_n12248__;
  assign new_new_n26802__ = ~new_new_n26800__ & ~new_new_n26801__;
  assign new_new_n26803__ = ys__n46751 & new_new_n12245__;
  assign new_new_n26804__ = ys__n46927 & new_new_n12246__;
  assign new_new_n26805__ = ~new_new_n26803__ & ~new_new_n26804__;
  assign new_new_n26806__ = new_new_n26802__ & new_new_n26805__;
  assign new_new_n26807__ = new_new_n12241__ & ~new_new_n26778__;
  assign new_new_n26808__ = ~new_new_n26806__ & new_new_n26807__;
  assign new_new_n26809__ = ~new_new_n26799__ & ~new_new_n26808__;
  assign new_new_n26810__ = new_new_n26790__ & new_new_n26809__;
  assign new_new_n26811__ = ~new_new_n12240__ & ~new_new_n12242__;
  assign new_new_n26812__ = new_new_n12354__ & new_new_n26811__;
  assign new_new_n26813__ = new_new_n12246__ & new_new_n12259__;
  assign new_new_n26814__ = ~new_new_n12260__ & ~new_new_n26813__;
  assign new_new_n26815__ = ~new_new_n26813__ & ~new_new_n26814__;
  assign new_new_n26816__ = ~new_new_n26812__ & new_new_n26815__;
  assign new_new_n26817__ = new_new_n12365__ & new_new_n26816__;
  assign new_new_n26818__ = ~new_new_n26768__ & new_new_n26817__;
  assign new_new_n26819__ = ~new_new_n26810__ & new_new_n26818__;
  assign new_new_n26820__ = ~new_new_n26769__ & ~new_new_n26819__;
  assign new_new_n26821__ = ~new_new_n12286__ & ~new_new_n26701__;
  assign new_new_n26822__ = ~new_new_n26820__ & new_new_n26821__;
  assign new_new_n26823__ = ys__n45648 & new_new_n12356__;
  assign new_new_n26824__ = ys__n45484 & new_new_n12248__;
  assign new_new_n26825__ = ~new_new_n26823__ & ~new_new_n26824__;
  assign new_new_n26826__ = ys__n45320 & new_new_n12245__;
  assign new_new_n26827__ = ys__n45134 & new_new_n12246__;
  assign new_new_n26828__ = ~new_new_n26826__ & ~new_new_n26827__;
  assign new_new_n26829__ = new_new_n26825__ & new_new_n26828__;
  assign new_new_n26830__ = new_new_n26779__ & ~new_new_n26829__;
  assign new_new_n26831__ = ys__n45609 & new_new_n12356__;
  assign new_new_n26832__ = ys__n45445 & new_new_n12248__;
  assign new_new_n26833__ = ~new_new_n26831__ & ~new_new_n26832__;
  assign new_new_n26834__ = ys__n45281 & new_new_n12245__;
  assign new_new_n26835__ = ys__n45087 & new_new_n12246__;
  assign new_new_n26836__ = ~new_new_n26834__ & ~new_new_n26835__;
  assign new_new_n26837__ = new_new_n26833__ & new_new_n26836__;
  assign new_new_n26838__ = new_new_n26788__ & ~new_new_n26837__;
  assign new_new_n26839__ = ~new_new_n26830__ & ~new_new_n26838__;
  assign new_new_n26840__ = ys__n45701 & new_new_n12356__;
  assign new_new_n26841__ = ys__n45537 & new_new_n12248__;
  assign new_new_n26842__ = ~new_new_n26840__ & ~new_new_n26841__;
  assign new_new_n26843__ = ys__n45373 & new_new_n12245__;
  assign new_new_n26844__ = ys__n45211 & new_new_n12246__;
  assign new_new_n26845__ = ~new_new_n26843__ & ~new_new_n26844__;
  assign new_new_n26846__ = new_new_n26842__ & new_new_n26845__;
  assign new_new_n26847__ = new_new_n26798__ & ~new_new_n26846__;
  assign new_new_n26848__ = ys__n45554 & new_new_n12356__;
  assign new_new_n26849__ = ys__n45390 & new_new_n12248__;
  assign new_new_n26850__ = ~new_new_n26848__ & ~new_new_n26849__;
  assign new_new_n26851__ = ys__n45226 & new_new_n12245__;
  assign new_new_n26852__ = ys__n45008 & new_new_n12246__;
  assign new_new_n26853__ = ~new_new_n26851__ & ~new_new_n26852__;
  assign new_new_n26854__ = new_new_n26850__ & new_new_n26853__;
  assign new_new_n26855__ = new_new_n26807__ & ~new_new_n26854__;
  assign new_new_n26856__ = ~new_new_n26847__ & ~new_new_n26855__;
  assign new_new_n26857__ = new_new_n26839__ & new_new_n26856__;
  assign new_new_n26858__ = new_new_n12286__ & new_new_n26816__;
  assign new_new_n26859__ = ~new_new_n26821__ & new_new_n26858__;
  assign new_new_n26860__ = ~new_new_n26857__ & new_new_n26859__;
  assign new_new_n26861__ = ~new_new_n26822__ & ~new_new_n26860__;
  assign new_new_n26862__ = ~new_new_n12395__ & ~new_new_n26739__;
  assign new_new_n26863__ = ~new_new_n26861__ & new_new_n26862__;
  assign new_new_n26864__ = ys__n46102 & new_new_n12356__;
  assign new_new_n26865__ = ys__n46004 & new_new_n12248__;
  assign new_new_n26866__ = ~new_new_n26864__ & ~new_new_n26865__;
  assign new_new_n26867__ = ys__n45906 & new_new_n12245__;
  assign new_new_n26868__ = ys__n45810 & new_new_n12246__;
  assign new_new_n26869__ = ~new_new_n26867__ & ~new_new_n26868__;
  assign new_new_n26870__ = new_new_n26866__ & new_new_n26869__;
  assign new_new_n26871__ = new_new_n26788__ & ~new_new_n26870__;
  assign new_new_n26872__ = ys__n46046 & new_new_n12356__;
  assign new_new_n26873__ = ys__n45948 & new_new_n12248__;
  assign new_new_n26874__ = ~new_new_n26872__ & ~new_new_n26873__;
  assign new_new_n26875__ = ys__n45850 & new_new_n12245__;
  assign new_new_n26876__ = ys__n45730 & new_new_n12246__;
  assign new_new_n26877__ = ~new_new_n26875__ & ~new_new_n26876__;
  assign new_new_n26878__ = new_new_n26874__ & new_new_n26877__;
  assign new_new_n26879__ = new_new_n26807__ & ~new_new_n26878__;
  assign new_new_n26880__ = ~new_new_n26871__ & ~new_new_n26879__;
  assign new_new_n26881__ = ~new_new_n12243__ & new_new_n26815__;
  assign new_new_n26882__ = new_new_n12395__ & new_new_n26881__;
  assign new_new_n26883__ = ~new_new_n26880__ & new_new_n26882__;
  assign new_new_n26884__ = ~new_new_n26862__ & new_new_n26883__;
  assign ys__n26118 = new_new_n26863__ | new_new_n26884__;
  assign new_new_n26886__ = ys__n26005 & new_new_n26768__;
  assign new_new_n26887__ = ys__n47110 & new_new_n12356__;
  assign new_new_n26888__ = ys__n47113 & new_new_n12248__;
  assign new_new_n26889__ = ~new_new_n26887__ & ~new_new_n26888__;
  assign new_new_n26890__ = ys__n47116 & new_new_n12245__;
  assign new_new_n26891__ = ys__n47119 & new_new_n12246__;
  assign new_new_n26892__ = ~new_new_n26890__ & ~new_new_n26891__;
  assign new_new_n26893__ = new_new_n26889__ & new_new_n26892__;
  assign new_new_n26894__ = new_new_n26779__ & ~new_new_n26893__;
  assign new_new_n26895__ = ys__n46268 & new_new_n12356__;
  assign new_new_n26896__ = ys__n46444 & new_new_n12248__;
  assign new_new_n26897__ = ~new_new_n26895__ & ~new_new_n26896__;
  assign new_new_n26898__ = ys__n46620 & new_new_n12245__;
  assign new_new_n26899__ = ys__n46796 & new_new_n12246__;
  assign new_new_n26900__ = ~new_new_n26898__ & ~new_new_n26899__;
  assign new_new_n26901__ = new_new_n26897__ & new_new_n26900__;
  assign new_new_n26902__ = new_new_n26788__ & ~new_new_n26901__;
  assign new_new_n26903__ = ~new_new_n26894__ & ~new_new_n26902__;
  assign new_new_n26904__ = ys__n46323 & new_new_n12356__;
  assign new_new_n26905__ = ys__n46499 & new_new_n12248__;
  assign new_new_n26906__ = ~new_new_n26904__ & ~new_new_n26905__;
  assign new_new_n26907__ = ys__n46675 & new_new_n12245__;
  assign new_new_n26908__ = ys__n46851 & new_new_n12246__;
  assign new_new_n26909__ = ~new_new_n26907__ & ~new_new_n26908__;
  assign new_new_n26910__ = new_new_n26906__ & new_new_n26909__;
  assign new_new_n26911__ = new_new_n26798__ & ~new_new_n26910__;
  assign new_new_n26912__ = ys__n46400 & new_new_n12356__;
  assign new_new_n26913__ = ys__n46576 & new_new_n12248__;
  assign new_new_n26914__ = ~new_new_n26912__ & ~new_new_n26913__;
  assign new_new_n26915__ = ys__n46752 & new_new_n12245__;
  assign new_new_n26916__ = ys__n46928 & new_new_n12246__;
  assign new_new_n26917__ = ~new_new_n26915__ & ~new_new_n26916__;
  assign new_new_n26918__ = new_new_n26914__ & new_new_n26917__;
  assign new_new_n26919__ = new_new_n26807__ & ~new_new_n26918__;
  assign new_new_n26920__ = ~new_new_n26911__ & ~new_new_n26919__;
  assign new_new_n26921__ = new_new_n26903__ & new_new_n26920__;
  assign new_new_n26922__ = new_new_n26818__ & ~new_new_n26921__;
  assign new_new_n26923__ = ~new_new_n26886__ & ~new_new_n26922__;
  assign new_new_n26924__ = new_new_n26821__ & ~new_new_n26923__;
  assign new_new_n26925__ = ys__n45556 & new_new_n12356__;
  assign new_new_n26926__ = ys__n45392 & new_new_n12248__;
  assign new_new_n26927__ = ~new_new_n26925__ & ~new_new_n26926__;
  assign new_new_n26928__ = ys__n45228 & new_new_n12245__;
  assign new_new_n26929__ = ys__n45011 & new_new_n12246__;
  assign new_new_n26930__ = ~new_new_n26928__ & ~new_new_n26929__;
  assign new_new_n26931__ = new_new_n26927__ & new_new_n26930__;
  assign new_new_n26932__ = new_new_n26807__ & ~new_new_n26931__;
  assign new_new_n26933__ = ys__n45650 & new_new_n12356__;
  assign new_new_n26934__ = ys__n45486 & new_new_n12248__;
  assign new_new_n26935__ = ~new_new_n26933__ & ~new_new_n26934__;
  assign new_new_n26936__ = ys__n45322 & new_new_n12245__;
  assign new_new_n26937__ = ys__n45137 & new_new_n12246__;
  assign new_new_n26938__ = ~new_new_n26936__ & ~new_new_n26937__;
  assign new_new_n26939__ = new_new_n26935__ & new_new_n26938__;
  assign new_new_n26940__ = new_new_n26779__ & ~new_new_n26939__;
  assign new_new_n26941__ = ys__n45610 & new_new_n12356__;
  assign new_new_n26942__ = ys__n45446 & new_new_n12248__;
  assign new_new_n26943__ = ~new_new_n26941__ & ~new_new_n26942__;
  assign new_new_n26944__ = ys__n45282 & new_new_n12245__;
  assign new_new_n26945__ = ys__n45088 & new_new_n12246__;
  assign new_new_n26946__ = ~new_new_n26944__ & ~new_new_n26945__;
  assign new_new_n26947__ = new_new_n26943__ & new_new_n26946__;
  assign new_new_n26948__ = new_new_n26788__ & ~new_new_n26947__;
  assign new_new_n26949__ = ~new_new_n26940__ & ~new_new_n26948__;
  assign new_new_n26950__ = ~new_new_n26932__ & new_new_n26949__;
  assign new_new_n26951__ = new_new_n26859__ & ~new_new_n26950__;
  assign new_new_n26952__ = ~new_new_n26924__ & ~new_new_n26951__;
  assign new_new_n26953__ = new_new_n26862__ & ~new_new_n26952__;
  assign new_new_n26954__ = ys__n46103 & new_new_n12356__;
  assign new_new_n26955__ = ys__n46005 & new_new_n12248__;
  assign new_new_n26956__ = ~new_new_n26954__ & ~new_new_n26955__;
  assign new_new_n26957__ = ys__n45907 & new_new_n12245__;
  assign new_new_n26958__ = ys__n45811 & new_new_n12246__;
  assign new_new_n26959__ = ~new_new_n26957__ & ~new_new_n26958__;
  assign new_new_n26960__ = new_new_n26956__ & new_new_n26959__;
  assign new_new_n26961__ = new_new_n26788__ & ~new_new_n26960__;
  assign new_new_n26962__ = ys__n46048 & new_new_n12356__;
  assign new_new_n26963__ = ys__n45950 & new_new_n12248__;
  assign new_new_n26964__ = ~new_new_n26962__ & ~new_new_n26963__;
  assign new_new_n26965__ = ys__n45852 & new_new_n12245__;
  assign new_new_n26966__ = ys__n45733 & new_new_n12246__;
  assign new_new_n26967__ = ~new_new_n26965__ & ~new_new_n26966__;
  assign new_new_n26968__ = new_new_n26964__ & new_new_n26967__;
  assign new_new_n26969__ = new_new_n26807__ & ~new_new_n26968__;
  assign new_new_n26970__ = ~new_new_n26961__ & ~new_new_n26969__;
  assign new_new_n26971__ = new_new_n26882__ & ~new_new_n26970__;
  assign new_new_n26972__ = ~new_new_n26862__ & new_new_n26971__;
  assign ys__n26119 = new_new_n26953__ | new_new_n26972__;
  assign new_new_n26974__ = ys__n26008 & new_new_n26768__;
  assign new_new_n26975__ = ys__n46348 & new_new_n12356__;
  assign new_new_n26976__ = ys__n46524 & new_new_n12248__;
  assign new_new_n26977__ = ~new_new_n26975__ & ~new_new_n26976__;
  assign new_new_n26978__ = ys__n46700 & new_new_n12245__;
  assign new_new_n26979__ = ys__n46876 & new_new_n12246__;
  assign new_new_n26980__ = ~new_new_n26978__ & ~new_new_n26979__;
  assign new_new_n26981__ = new_new_n26977__ & new_new_n26980__;
  assign new_new_n26982__ = new_new_n26779__ & ~new_new_n26981__;
  assign new_new_n26983__ = ys__n46270 & new_new_n12356__;
  assign new_new_n26984__ = ys__n46446 & new_new_n12248__;
  assign new_new_n26985__ = ~new_new_n26983__ & ~new_new_n26984__;
  assign new_new_n26986__ = ys__n46622 & new_new_n12245__;
  assign new_new_n26987__ = ys__n46798 & new_new_n12246__;
  assign new_new_n26988__ = ~new_new_n26986__ & ~new_new_n26987__;
  assign new_new_n26989__ = new_new_n26985__ & new_new_n26988__;
  assign new_new_n26990__ = new_new_n26788__ & ~new_new_n26989__;
  assign new_new_n26991__ = ~new_new_n26982__ & ~new_new_n26990__;
  assign new_new_n26992__ = ys__n46324 & new_new_n12356__;
  assign new_new_n26993__ = ys__n46500 & new_new_n12248__;
  assign new_new_n26994__ = ~new_new_n26992__ & ~new_new_n26993__;
  assign new_new_n26995__ = ys__n46676 & new_new_n12245__;
  assign new_new_n26996__ = ys__n46852 & new_new_n12246__;
  assign new_new_n26997__ = ~new_new_n26995__ & ~new_new_n26996__;
  assign new_new_n26998__ = new_new_n26994__ & new_new_n26997__;
  assign new_new_n26999__ = new_new_n26798__ & ~new_new_n26998__;
  assign new_new_n27000__ = ys__n46401 & new_new_n12356__;
  assign new_new_n27001__ = ys__n46577 & new_new_n12248__;
  assign new_new_n27002__ = ~new_new_n27000__ & ~new_new_n27001__;
  assign new_new_n27003__ = ys__n46753 & new_new_n12245__;
  assign new_new_n27004__ = ys__n46929 & new_new_n12246__;
  assign new_new_n27005__ = ~new_new_n27003__ & ~new_new_n27004__;
  assign new_new_n27006__ = new_new_n27002__ & new_new_n27005__;
  assign new_new_n27007__ = new_new_n26807__ & ~new_new_n27006__;
  assign new_new_n27008__ = ~new_new_n26999__ & ~new_new_n27007__;
  assign new_new_n27009__ = new_new_n26991__ & new_new_n27008__;
  assign new_new_n27010__ = new_new_n26818__ & ~new_new_n27009__;
  assign new_new_n27011__ = ~new_new_n26974__ & ~new_new_n27010__;
  assign new_new_n27012__ = new_new_n26821__ & ~new_new_n27011__;
  assign new_new_n27013__ = ys__n45558 & new_new_n12356__;
  assign new_new_n27014__ = ys__n45394 & new_new_n12248__;
  assign new_new_n27015__ = ~new_new_n27013__ & ~new_new_n27014__;
  assign new_new_n27016__ = ys__n45230 & new_new_n12245__;
  assign new_new_n27017__ = ys__n45014 & new_new_n12246__;
  assign new_new_n27018__ = ~new_new_n27016__ & ~new_new_n27017__;
  assign new_new_n27019__ = new_new_n27015__ & new_new_n27018__;
  assign new_new_n27020__ = new_new_n26807__ & ~new_new_n27019__;
  assign new_new_n27021__ = ys__n45652 & new_new_n12356__;
  assign new_new_n27022__ = ys__n45488 & new_new_n12248__;
  assign new_new_n27023__ = ~new_new_n27021__ & ~new_new_n27022__;
  assign new_new_n27024__ = ys__n45324 & new_new_n12245__;
  assign new_new_n27025__ = ys__n45140 & new_new_n12246__;
  assign new_new_n27026__ = ~new_new_n27024__ & ~new_new_n27025__;
  assign new_new_n27027__ = new_new_n27023__ & new_new_n27026__;
  assign new_new_n27028__ = new_new_n26779__ & ~new_new_n27027__;
  assign new_new_n27029__ = ys__n45611 & new_new_n12356__;
  assign new_new_n27030__ = ys__n45447 & new_new_n12248__;
  assign new_new_n27031__ = ~new_new_n27029__ & ~new_new_n27030__;
  assign new_new_n27032__ = ys__n45283 & new_new_n12245__;
  assign new_new_n27033__ = ys__n45089 & new_new_n12246__;
  assign new_new_n27034__ = ~new_new_n27032__ & ~new_new_n27033__;
  assign new_new_n27035__ = new_new_n27031__ & new_new_n27034__;
  assign new_new_n27036__ = new_new_n26788__ & ~new_new_n27035__;
  assign new_new_n27037__ = ~new_new_n27028__ & ~new_new_n27036__;
  assign new_new_n27038__ = ~new_new_n27020__ & new_new_n27037__;
  assign new_new_n27039__ = new_new_n26859__ & ~new_new_n27038__;
  assign new_new_n27040__ = ~new_new_n27012__ & ~new_new_n27039__;
  assign new_new_n27041__ = new_new_n26862__ & ~new_new_n27040__;
  assign new_new_n27042__ = ys__n46104 & new_new_n12356__;
  assign new_new_n27043__ = ys__n46006 & new_new_n12248__;
  assign new_new_n27044__ = ~new_new_n27042__ & ~new_new_n27043__;
  assign new_new_n27045__ = ys__n45908 & new_new_n12245__;
  assign new_new_n27046__ = ys__n45812 & new_new_n12246__;
  assign new_new_n27047__ = ~new_new_n27045__ & ~new_new_n27046__;
  assign new_new_n27048__ = new_new_n27044__ & new_new_n27047__;
  assign new_new_n27049__ = new_new_n26788__ & ~new_new_n27048__;
  assign new_new_n27050__ = ys__n46050 & new_new_n12356__;
  assign new_new_n27051__ = ys__n45952 & new_new_n12248__;
  assign new_new_n27052__ = ~new_new_n27050__ & ~new_new_n27051__;
  assign new_new_n27053__ = ys__n45854 & new_new_n12245__;
  assign new_new_n27054__ = ys__n45736 & new_new_n12246__;
  assign new_new_n27055__ = ~new_new_n27053__ & ~new_new_n27054__;
  assign new_new_n27056__ = new_new_n27052__ & new_new_n27055__;
  assign new_new_n27057__ = new_new_n26807__ & ~new_new_n27056__;
  assign new_new_n27058__ = ~new_new_n27049__ & ~new_new_n27057__;
  assign new_new_n27059__ = new_new_n26882__ & ~new_new_n27058__;
  assign new_new_n27060__ = ~new_new_n26862__ & new_new_n27059__;
  assign ys__n26120 = new_new_n27041__ | new_new_n27060__;
  assign new_new_n27062__ = ys__n26011 & new_new_n26768__;
  assign new_new_n27063__ = ys__n46350 & new_new_n12356__;
  assign new_new_n27064__ = ys__n46526 & new_new_n12248__;
  assign new_new_n27065__ = ~new_new_n27063__ & ~new_new_n27064__;
  assign new_new_n27066__ = ys__n46702 & new_new_n12245__;
  assign new_new_n27067__ = ys__n46878 & new_new_n12246__;
  assign new_new_n27068__ = ~new_new_n27066__ & ~new_new_n27067__;
  assign new_new_n27069__ = new_new_n27065__ & new_new_n27068__;
  assign new_new_n27070__ = new_new_n26779__ & ~new_new_n27069__;
  assign new_new_n27071__ = ys__n46272 & new_new_n12356__;
  assign new_new_n27072__ = ys__n46448 & new_new_n12248__;
  assign new_new_n27073__ = ~new_new_n27071__ & ~new_new_n27072__;
  assign new_new_n27074__ = ys__n46624 & new_new_n12245__;
  assign new_new_n27075__ = ys__n46800 & new_new_n12246__;
  assign new_new_n27076__ = ~new_new_n27074__ & ~new_new_n27075__;
  assign new_new_n27077__ = new_new_n27073__ & new_new_n27076__;
  assign new_new_n27078__ = new_new_n26788__ & ~new_new_n27077__;
  assign new_new_n27079__ = ~new_new_n27070__ & ~new_new_n27078__;
  assign new_new_n27080__ = ys__n46325 & new_new_n12356__;
  assign new_new_n27081__ = ys__n46501 & new_new_n12248__;
  assign new_new_n27082__ = ~new_new_n27080__ & ~new_new_n27081__;
  assign new_new_n27083__ = ys__n46677 & new_new_n12245__;
  assign new_new_n27084__ = ys__n46853 & new_new_n12246__;
  assign new_new_n27085__ = ~new_new_n27083__ & ~new_new_n27084__;
  assign new_new_n27086__ = new_new_n27082__ & new_new_n27085__;
  assign new_new_n27087__ = new_new_n26798__ & ~new_new_n27086__;
  assign new_new_n27088__ = ys__n46402 & new_new_n12356__;
  assign new_new_n27089__ = ys__n46578 & new_new_n12248__;
  assign new_new_n27090__ = ~new_new_n27088__ & ~new_new_n27089__;
  assign new_new_n27091__ = ys__n46754 & new_new_n12245__;
  assign new_new_n27092__ = ys__n46930 & new_new_n12246__;
  assign new_new_n27093__ = ~new_new_n27091__ & ~new_new_n27092__;
  assign new_new_n27094__ = new_new_n27090__ & new_new_n27093__;
  assign new_new_n27095__ = new_new_n26807__ & ~new_new_n27094__;
  assign new_new_n27096__ = ~new_new_n27087__ & ~new_new_n27095__;
  assign new_new_n27097__ = new_new_n27079__ & new_new_n27096__;
  assign new_new_n27098__ = new_new_n26818__ & ~new_new_n27097__;
  assign new_new_n27099__ = ~new_new_n27062__ & ~new_new_n27098__;
  assign new_new_n27100__ = new_new_n26821__ & ~new_new_n27099__;
  assign new_new_n27101__ = ys__n45560 & new_new_n12356__;
  assign new_new_n27102__ = ys__n45396 & new_new_n12248__;
  assign new_new_n27103__ = ~new_new_n27101__ & ~new_new_n27102__;
  assign new_new_n27104__ = ys__n45232 & new_new_n12245__;
  assign new_new_n27105__ = ys__n45017 & new_new_n12246__;
  assign new_new_n27106__ = ~new_new_n27104__ & ~new_new_n27105__;
  assign new_new_n27107__ = new_new_n27103__ & new_new_n27106__;
  assign new_new_n27108__ = new_new_n26807__ & ~new_new_n27107__;
  assign new_new_n27109__ = ys__n45654 & new_new_n12356__;
  assign new_new_n27110__ = ys__n45490 & new_new_n12248__;
  assign new_new_n27111__ = ~new_new_n27109__ & ~new_new_n27110__;
  assign new_new_n27112__ = ys__n45326 & new_new_n12245__;
  assign new_new_n27113__ = ys__n45143 & new_new_n12246__;
  assign new_new_n27114__ = ~new_new_n27112__ & ~new_new_n27113__;
  assign new_new_n27115__ = new_new_n27111__ & new_new_n27114__;
  assign new_new_n27116__ = new_new_n26779__ & ~new_new_n27115__;
  assign new_new_n27117__ = ys__n45612 & new_new_n12356__;
  assign new_new_n27118__ = ys__n45448 & new_new_n12248__;
  assign new_new_n27119__ = ~new_new_n27117__ & ~new_new_n27118__;
  assign new_new_n27120__ = ys__n45284 & new_new_n12245__;
  assign new_new_n27121__ = ys__n45090 & new_new_n12246__;
  assign new_new_n27122__ = ~new_new_n27120__ & ~new_new_n27121__;
  assign new_new_n27123__ = new_new_n27119__ & new_new_n27122__;
  assign new_new_n27124__ = new_new_n26788__ & ~new_new_n27123__;
  assign new_new_n27125__ = ~new_new_n27116__ & ~new_new_n27124__;
  assign new_new_n27126__ = ~new_new_n27108__ & new_new_n27125__;
  assign new_new_n27127__ = new_new_n26859__ & ~new_new_n27126__;
  assign new_new_n27128__ = ~new_new_n27100__ & ~new_new_n27127__;
  assign new_new_n27129__ = new_new_n26862__ & ~new_new_n27128__;
  assign new_new_n27130__ = ys__n46105 & new_new_n12356__;
  assign new_new_n27131__ = ys__n46007 & new_new_n12248__;
  assign new_new_n27132__ = ~new_new_n27130__ & ~new_new_n27131__;
  assign new_new_n27133__ = ys__n45909 & new_new_n12245__;
  assign new_new_n27134__ = ys__n45813 & new_new_n12246__;
  assign new_new_n27135__ = ~new_new_n27133__ & ~new_new_n27134__;
  assign new_new_n27136__ = new_new_n27132__ & new_new_n27135__;
  assign new_new_n27137__ = new_new_n26788__ & ~new_new_n27136__;
  assign new_new_n27138__ = ys__n46052 & new_new_n12356__;
  assign new_new_n27139__ = ys__n45954 & new_new_n12248__;
  assign new_new_n27140__ = ~new_new_n27138__ & ~new_new_n27139__;
  assign new_new_n27141__ = ys__n45856 & new_new_n12245__;
  assign new_new_n27142__ = ys__n45739 & new_new_n12246__;
  assign new_new_n27143__ = ~new_new_n27141__ & ~new_new_n27142__;
  assign new_new_n27144__ = new_new_n27140__ & new_new_n27143__;
  assign new_new_n27145__ = new_new_n26807__ & ~new_new_n27144__;
  assign new_new_n27146__ = ~new_new_n27137__ & ~new_new_n27145__;
  assign new_new_n27147__ = new_new_n26882__ & ~new_new_n27146__;
  assign new_new_n27148__ = ~new_new_n26862__ & new_new_n27147__;
  assign ys__n26121 = new_new_n27129__ | new_new_n27148__;
  assign new_new_n27150__ = ys__n26014 & new_new_n26768__;
  assign new_new_n27151__ = ys__n46352 & new_new_n12356__;
  assign new_new_n27152__ = ys__n46528 & new_new_n12248__;
  assign new_new_n27153__ = ~new_new_n27151__ & ~new_new_n27152__;
  assign new_new_n27154__ = ys__n46704 & new_new_n12245__;
  assign new_new_n27155__ = ys__n46880 & new_new_n12246__;
  assign new_new_n27156__ = ~new_new_n27154__ & ~new_new_n27155__;
  assign new_new_n27157__ = new_new_n27153__ & new_new_n27156__;
  assign new_new_n27158__ = new_new_n26779__ & ~new_new_n27157__;
  assign new_new_n27159__ = ys__n46274 & new_new_n12356__;
  assign new_new_n27160__ = ys__n46450 & new_new_n12248__;
  assign new_new_n27161__ = ~new_new_n27159__ & ~new_new_n27160__;
  assign new_new_n27162__ = ys__n46626 & new_new_n12245__;
  assign new_new_n27163__ = ys__n46802 & new_new_n12246__;
  assign new_new_n27164__ = ~new_new_n27162__ & ~new_new_n27163__;
  assign new_new_n27165__ = new_new_n27161__ & new_new_n27164__;
  assign new_new_n27166__ = new_new_n26788__ & ~new_new_n27165__;
  assign new_new_n27167__ = ~new_new_n27158__ & ~new_new_n27166__;
  assign new_new_n27168__ = ys__n46326 & new_new_n12356__;
  assign new_new_n27169__ = ys__n46502 & new_new_n12248__;
  assign new_new_n27170__ = ~new_new_n27168__ & ~new_new_n27169__;
  assign new_new_n27171__ = ys__n46678 & new_new_n12245__;
  assign new_new_n27172__ = ys__n46854 & new_new_n12246__;
  assign new_new_n27173__ = ~new_new_n27171__ & ~new_new_n27172__;
  assign new_new_n27174__ = new_new_n27170__ & new_new_n27173__;
  assign new_new_n27175__ = new_new_n26798__ & ~new_new_n27174__;
  assign new_new_n27176__ = ys__n46403 & new_new_n12356__;
  assign new_new_n27177__ = ys__n46579 & new_new_n12248__;
  assign new_new_n27178__ = ~new_new_n27176__ & ~new_new_n27177__;
  assign new_new_n27179__ = ys__n46755 & new_new_n12245__;
  assign new_new_n27180__ = ys__n46931 & new_new_n12246__;
  assign new_new_n27181__ = ~new_new_n27179__ & ~new_new_n27180__;
  assign new_new_n27182__ = new_new_n27178__ & new_new_n27181__;
  assign new_new_n27183__ = new_new_n26807__ & ~new_new_n27182__;
  assign new_new_n27184__ = ~new_new_n27175__ & ~new_new_n27183__;
  assign new_new_n27185__ = new_new_n27167__ & new_new_n27184__;
  assign new_new_n27186__ = new_new_n26818__ & ~new_new_n27185__;
  assign new_new_n27187__ = ~new_new_n27150__ & ~new_new_n27186__;
  assign new_new_n27188__ = new_new_n26821__ & ~new_new_n27187__;
  assign new_new_n27189__ = ys__n45562 & new_new_n12356__;
  assign new_new_n27190__ = ys__n45398 & new_new_n12248__;
  assign new_new_n27191__ = ~new_new_n27189__ & ~new_new_n27190__;
  assign new_new_n27192__ = ys__n45234 & new_new_n12245__;
  assign new_new_n27193__ = ys__n45020 & new_new_n12246__;
  assign new_new_n27194__ = ~new_new_n27192__ & ~new_new_n27193__;
  assign new_new_n27195__ = new_new_n27191__ & new_new_n27194__;
  assign new_new_n27196__ = new_new_n26807__ & ~new_new_n27195__;
  assign new_new_n27197__ = ys__n45656 & new_new_n12356__;
  assign new_new_n27198__ = ys__n45492 & new_new_n12248__;
  assign new_new_n27199__ = ~new_new_n27197__ & ~new_new_n27198__;
  assign new_new_n27200__ = ys__n45328 & new_new_n12245__;
  assign new_new_n27201__ = ys__n45146 & new_new_n12246__;
  assign new_new_n27202__ = ~new_new_n27200__ & ~new_new_n27201__;
  assign new_new_n27203__ = new_new_n27199__ & new_new_n27202__;
  assign new_new_n27204__ = new_new_n26779__ & ~new_new_n27203__;
  assign new_new_n27205__ = ys__n45613 & new_new_n12356__;
  assign new_new_n27206__ = ys__n45449 & new_new_n12248__;
  assign new_new_n27207__ = ~new_new_n27205__ & ~new_new_n27206__;
  assign new_new_n27208__ = ys__n45285 & new_new_n12245__;
  assign new_new_n27209__ = ys__n45091 & new_new_n12246__;
  assign new_new_n27210__ = ~new_new_n27208__ & ~new_new_n27209__;
  assign new_new_n27211__ = new_new_n27207__ & new_new_n27210__;
  assign new_new_n27212__ = new_new_n26788__ & ~new_new_n27211__;
  assign new_new_n27213__ = ~new_new_n27204__ & ~new_new_n27212__;
  assign new_new_n27214__ = ~new_new_n27196__ & new_new_n27213__;
  assign new_new_n27215__ = new_new_n26859__ & ~new_new_n27214__;
  assign new_new_n27216__ = ~new_new_n27188__ & ~new_new_n27215__;
  assign new_new_n27217__ = new_new_n26862__ & ~new_new_n27216__;
  assign new_new_n27218__ = ys__n46106 & new_new_n12356__;
  assign new_new_n27219__ = ys__n46008 & new_new_n12248__;
  assign new_new_n27220__ = ~new_new_n27218__ & ~new_new_n27219__;
  assign new_new_n27221__ = ys__n45910 & new_new_n12245__;
  assign new_new_n27222__ = ys__n45814 & new_new_n12246__;
  assign new_new_n27223__ = ~new_new_n27221__ & ~new_new_n27222__;
  assign new_new_n27224__ = new_new_n27220__ & new_new_n27223__;
  assign new_new_n27225__ = new_new_n26788__ & ~new_new_n27224__;
  assign new_new_n27226__ = ys__n46054 & new_new_n12356__;
  assign new_new_n27227__ = ys__n45956 & new_new_n12248__;
  assign new_new_n27228__ = ~new_new_n27226__ & ~new_new_n27227__;
  assign new_new_n27229__ = ys__n45858 & new_new_n12245__;
  assign new_new_n27230__ = ys__n45742 & new_new_n12246__;
  assign new_new_n27231__ = ~new_new_n27229__ & ~new_new_n27230__;
  assign new_new_n27232__ = new_new_n27228__ & new_new_n27231__;
  assign new_new_n27233__ = new_new_n26807__ & ~new_new_n27232__;
  assign new_new_n27234__ = ~new_new_n27225__ & ~new_new_n27233__;
  assign new_new_n27235__ = new_new_n26882__ & ~new_new_n27234__;
  assign new_new_n27236__ = ~new_new_n26862__ & new_new_n27235__;
  assign ys__n26122 = new_new_n27217__ | new_new_n27236__;
  assign new_new_n27238__ = ys__n26017 & new_new_n26768__;
  assign new_new_n27239__ = ys__n46354 & new_new_n12356__;
  assign new_new_n27240__ = ys__n46530 & new_new_n12248__;
  assign new_new_n27241__ = ~new_new_n27239__ & ~new_new_n27240__;
  assign new_new_n27242__ = ys__n46706 & new_new_n12245__;
  assign new_new_n27243__ = ys__n46882 & new_new_n12246__;
  assign new_new_n27244__ = ~new_new_n27242__ & ~new_new_n27243__;
  assign new_new_n27245__ = new_new_n27241__ & new_new_n27244__;
  assign new_new_n27246__ = new_new_n26779__ & ~new_new_n27245__;
  assign new_new_n27247__ = ys__n46276 & new_new_n12356__;
  assign new_new_n27248__ = ys__n46452 & new_new_n12248__;
  assign new_new_n27249__ = ~new_new_n27247__ & ~new_new_n27248__;
  assign new_new_n27250__ = ys__n46628 & new_new_n12245__;
  assign new_new_n27251__ = ys__n46804 & new_new_n12246__;
  assign new_new_n27252__ = ~new_new_n27250__ & ~new_new_n27251__;
  assign new_new_n27253__ = new_new_n27249__ & new_new_n27252__;
  assign new_new_n27254__ = new_new_n26788__ & ~new_new_n27253__;
  assign new_new_n27255__ = ~new_new_n27246__ & ~new_new_n27254__;
  assign new_new_n27256__ = ys__n46327 & new_new_n12356__;
  assign new_new_n27257__ = ys__n46503 & new_new_n12248__;
  assign new_new_n27258__ = ~new_new_n27256__ & ~new_new_n27257__;
  assign new_new_n27259__ = ys__n46679 & new_new_n12245__;
  assign new_new_n27260__ = ys__n46855 & new_new_n12246__;
  assign new_new_n27261__ = ~new_new_n27259__ & ~new_new_n27260__;
  assign new_new_n27262__ = new_new_n27258__ & new_new_n27261__;
  assign new_new_n27263__ = new_new_n26798__ & ~new_new_n27262__;
  assign new_new_n27264__ = ys__n46404 & new_new_n12356__;
  assign new_new_n27265__ = ys__n46580 & new_new_n12248__;
  assign new_new_n27266__ = ~new_new_n27264__ & ~new_new_n27265__;
  assign new_new_n27267__ = ys__n46756 & new_new_n12245__;
  assign new_new_n27268__ = ys__n46932 & new_new_n12246__;
  assign new_new_n27269__ = ~new_new_n27267__ & ~new_new_n27268__;
  assign new_new_n27270__ = new_new_n27266__ & new_new_n27269__;
  assign new_new_n27271__ = new_new_n26807__ & ~new_new_n27270__;
  assign new_new_n27272__ = ~new_new_n27263__ & ~new_new_n27271__;
  assign new_new_n27273__ = new_new_n27255__ & new_new_n27272__;
  assign new_new_n27274__ = new_new_n26818__ & ~new_new_n27273__;
  assign new_new_n27275__ = ~new_new_n27238__ & ~new_new_n27274__;
  assign new_new_n27276__ = new_new_n26821__ & ~new_new_n27275__;
  assign new_new_n27277__ = ys__n45564 & new_new_n12356__;
  assign new_new_n27278__ = ys__n45400 & new_new_n12248__;
  assign new_new_n27279__ = ~new_new_n27277__ & ~new_new_n27278__;
  assign new_new_n27280__ = ys__n45236 & new_new_n12245__;
  assign new_new_n27281__ = ys__n45023 & new_new_n12246__;
  assign new_new_n27282__ = ~new_new_n27280__ & ~new_new_n27281__;
  assign new_new_n27283__ = new_new_n27279__ & new_new_n27282__;
  assign new_new_n27284__ = new_new_n26807__ & ~new_new_n27283__;
  assign new_new_n27285__ = ys__n45658 & new_new_n12356__;
  assign new_new_n27286__ = ys__n45494 & new_new_n12248__;
  assign new_new_n27287__ = ~new_new_n27285__ & ~new_new_n27286__;
  assign new_new_n27288__ = ys__n45330 & new_new_n12245__;
  assign new_new_n27289__ = ys__n45149 & new_new_n12246__;
  assign new_new_n27290__ = ~new_new_n27288__ & ~new_new_n27289__;
  assign new_new_n27291__ = new_new_n27287__ & new_new_n27290__;
  assign new_new_n27292__ = new_new_n26779__ & ~new_new_n27291__;
  assign new_new_n27293__ = ys__n45614 & new_new_n12356__;
  assign new_new_n27294__ = ys__n45450 & new_new_n12248__;
  assign new_new_n27295__ = ~new_new_n27293__ & ~new_new_n27294__;
  assign new_new_n27296__ = ys__n45286 & new_new_n12245__;
  assign new_new_n27297__ = ys__n45092 & new_new_n12246__;
  assign new_new_n27298__ = ~new_new_n27296__ & ~new_new_n27297__;
  assign new_new_n27299__ = new_new_n27295__ & new_new_n27298__;
  assign new_new_n27300__ = new_new_n26788__ & ~new_new_n27299__;
  assign new_new_n27301__ = ~new_new_n27292__ & ~new_new_n27300__;
  assign new_new_n27302__ = ~new_new_n27284__ & new_new_n27301__;
  assign new_new_n27303__ = new_new_n26859__ & ~new_new_n27302__;
  assign new_new_n27304__ = ~new_new_n27276__ & ~new_new_n27303__;
  assign new_new_n27305__ = new_new_n26862__ & ~new_new_n27304__;
  assign new_new_n27306__ = ys__n46107 & new_new_n12356__;
  assign new_new_n27307__ = ys__n46009 & new_new_n12248__;
  assign new_new_n27308__ = ~new_new_n27306__ & ~new_new_n27307__;
  assign new_new_n27309__ = ys__n45911 & new_new_n12245__;
  assign new_new_n27310__ = ys__n45815 & new_new_n12246__;
  assign new_new_n27311__ = ~new_new_n27309__ & ~new_new_n27310__;
  assign new_new_n27312__ = new_new_n27308__ & new_new_n27311__;
  assign new_new_n27313__ = new_new_n26788__ & ~new_new_n27312__;
  assign new_new_n27314__ = ys__n46056 & new_new_n12356__;
  assign new_new_n27315__ = ys__n45958 & new_new_n12248__;
  assign new_new_n27316__ = ~new_new_n27314__ & ~new_new_n27315__;
  assign new_new_n27317__ = ys__n45860 & new_new_n12245__;
  assign new_new_n27318__ = ys__n45745 & new_new_n12246__;
  assign new_new_n27319__ = ~new_new_n27317__ & ~new_new_n27318__;
  assign new_new_n27320__ = new_new_n27316__ & new_new_n27319__;
  assign new_new_n27321__ = new_new_n26807__ & ~new_new_n27320__;
  assign new_new_n27322__ = ~new_new_n27313__ & ~new_new_n27321__;
  assign new_new_n27323__ = new_new_n26882__ & ~new_new_n27322__;
  assign new_new_n27324__ = ~new_new_n26862__ & new_new_n27323__;
  assign ys__n26123 = new_new_n27305__ | new_new_n27324__;
  assign new_new_n27326__ = ys__n26020 & new_new_n26768__;
  assign new_new_n27327__ = ys__n46356 & new_new_n12356__;
  assign new_new_n27328__ = ys__n46532 & new_new_n12248__;
  assign new_new_n27329__ = ~new_new_n27327__ & ~new_new_n27328__;
  assign new_new_n27330__ = ys__n46708 & new_new_n12245__;
  assign new_new_n27331__ = ys__n46884 & new_new_n12246__;
  assign new_new_n27332__ = ~new_new_n27330__ & ~new_new_n27331__;
  assign new_new_n27333__ = new_new_n27329__ & new_new_n27332__;
  assign new_new_n27334__ = new_new_n26779__ & ~new_new_n27333__;
  assign new_new_n27335__ = ys__n46278 & new_new_n12356__;
  assign new_new_n27336__ = ys__n46454 & new_new_n12248__;
  assign new_new_n27337__ = ~new_new_n27335__ & ~new_new_n27336__;
  assign new_new_n27338__ = ys__n46630 & new_new_n12245__;
  assign new_new_n27339__ = ys__n46806 & new_new_n12246__;
  assign new_new_n27340__ = ~new_new_n27338__ & ~new_new_n27339__;
  assign new_new_n27341__ = new_new_n27337__ & new_new_n27340__;
  assign new_new_n27342__ = new_new_n26788__ & ~new_new_n27341__;
  assign new_new_n27343__ = ~new_new_n27334__ & ~new_new_n27342__;
  assign new_new_n27344__ = ys__n46328 & new_new_n12356__;
  assign new_new_n27345__ = ys__n46504 & new_new_n12248__;
  assign new_new_n27346__ = ~new_new_n27344__ & ~new_new_n27345__;
  assign new_new_n27347__ = ys__n46680 & new_new_n12245__;
  assign new_new_n27348__ = ys__n46856 & new_new_n12246__;
  assign new_new_n27349__ = ~new_new_n27347__ & ~new_new_n27348__;
  assign new_new_n27350__ = new_new_n27346__ & new_new_n27349__;
  assign new_new_n27351__ = new_new_n26798__ & ~new_new_n27350__;
  assign new_new_n27352__ = ys__n46405 & new_new_n12356__;
  assign new_new_n27353__ = ys__n46581 & new_new_n12248__;
  assign new_new_n27354__ = ~new_new_n27352__ & ~new_new_n27353__;
  assign new_new_n27355__ = ys__n46757 & new_new_n12245__;
  assign new_new_n27356__ = ys__n46933 & new_new_n12246__;
  assign new_new_n27357__ = ~new_new_n27355__ & ~new_new_n27356__;
  assign new_new_n27358__ = new_new_n27354__ & new_new_n27357__;
  assign new_new_n27359__ = new_new_n26807__ & ~new_new_n27358__;
  assign new_new_n27360__ = ~new_new_n27351__ & ~new_new_n27359__;
  assign new_new_n27361__ = new_new_n27343__ & new_new_n27360__;
  assign new_new_n27362__ = new_new_n26818__ & ~new_new_n27361__;
  assign new_new_n27363__ = ~new_new_n27326__ & ~new_new_n27362__;
  assign new_new_n27364__ = new_new_n26821__ & ~new_new_n27363__;
  assign new_new_n27365__ = ys__n45566 & new_new_n12356__;
  assign new_new_n27366__ = ys__n45402 & new_new_n12248__;
  assign new_new_n27367__ = ~new_new_n27365__ & ~new_new_n27366__;
  assign new_new_n27368__ = ys__n45238 & new_new_n12245__;
  assign new_new_n27369__ = ys__n45026 & new_new_n12246__;
  assign new_new_n27370__ = ~new_new_n27368__ & ~new_new_n27369__;
  assign new_new_n27371__ = new_new_n27367__ & new_new_n27370__;
  assign new_new_n27372__ = new_new_n26807__ & ~new_new_n27371__;
  assign new_new_n27373__ = ys__n45660 & new_new_n12356__;
  assign new_new_n27374__ = ys__n45496 & new_new_n12248__;
  assign new_new_n27375__ = ~new_new_n27373__ & ~new_new_n27374__;
  assign new_new_n27376__ = ys__n45332 & new_new_n12245__;
  assign new_new_n27377__ = ys__n45152 & new_new_n12246__;
  assign new_new_n27378__ = ~new_new_n27376__ & ~new_new_n27377__;
  assign new_new_n27379__ = new_new_n27375__ & new_new_n27378__;
  assign new_new_n27380__ = new_new_n26779__ & ~new_new_n27379__;
  assign new_new_n27381__ = ys__n45615 & new_new_n12356__;
  assign new_new_n27382__ = ys__n45451 & new_new_n12248__;
  assign new_new_n27383__ = ~new_new_n27381__ & ~new_new_n27382__;
  assign new_new_n27384__ = ys__n45287 & new_new_n12245__;
  assign new_new_n27385__ = ys__n45093 & new_new_n12246__;
  assign new_new_n27386__ = ~new_new_n27384__ & ~new_new_n27385__;
  assign new_new_n27387__ = new_new_n27383__ & new_new_n27386__;
  assign new_new_n27388__ = new_new_n26788__ & ~new_new_n27387__;
  assign new_new_n27389__ = ~new_new_n27380__ & ~new_new_n27388__;
  assign new_new_n27390__ = ~new_new_n27372__ & new_new_n27389__;
  assign new_new_n27391__ = new_new_n26859__ & ~new_new_n27390__;
  assign new_new_n27392__ = ~new_new_n27364__ & ~new_new_n27391__;
  assign new_new_n27393__ = new_new_n26862__ & ~new_new_n27392__;
  assign new_new_n27394__ = ys__n46108 & new_new_n12356__;
  assign new_new_n27395__ = ys__n46010 & new_new_n12248__;
  assign new_new_n27396__ = ~new_new_n27394__ & ~new_new_n27395__;
  assign new_new_n27397__ = ys__n45912 & new_new_n12245__;
  assign new_new_n27398__ = ys__n45816 & new_new_n12246__;
  assign new_new_n27399__ = ~new_new_n27397__ & ~new_new_n27398__;
  assign new_new_n27400__ = new_new_n27396__ & new_new_n27399__;
  assign new_new_n27401__ = new_new_n26788__ & ~new_new_n27400__;
  assign new_new_n27402__ = ys__n46058 & new_new_n12356__;
  assign new_new_n27403__ = ys__n45960 & new_new_n12248__;
  assign new_new_n27404__ = ~new_new_n27402__ & ~new_new_n27403__;
  assign new_new_n27405__ = ys__n45862 & new_new_n12245__;
  assign new_new_n27406__ = ys__n45748 & new_new_n12246__;
  assign new_new_n27407__ = ~new_new_n27405__ & ~new_new_n27406__;
  assign new_new_n27408__ = new_new_n27404__ & new_new_n27407__;
  assign new_new_n27409__ = new_new_n26807__ & ~new_new_n27408__;
  assign new_new_n27410__ = ~new_new_n27401__ & ~new_new_n27409__;
  assign new_new_n27411__ = new_new_n26882__ & ~new_new_n27410__;
  assign new_new_n27412__ = ~new_new_n26862__ & new_new_n27411__;
  assign ys__n26124 = new_new_n27393__ | new_new_n27412__;
  assign new_new_n27414__ = ys__n26023 & new_new_n26768__;
  assign new_new_n27415__ = ys__n46358 & new_new_n12356__;
  assign new_new_n27416__ = ys__n46534 & new_new_n12248__;
  assign new_new_n27417__ = ~new_new_n27415__ & ~new_new_n27416__;
  assign new_new_n27418__ = ys__n46710 & new_new_n12245__;
  assign new_new_n27419__ = ys__n46886 & new_new_n12246__;
  assign new_new_n27420__ = ~new_new_n27418__ & ~new_new_n27419__;
  assign new_new_n27421__ = new_new_n27417__ & new_new_n27420__;
  assign new_new_n27422__ = new_new_n26779__ & ~new_new_n27421__;
  assign new_new_n27423__ = ys__n46280 & new_new_n12356__;
  assign new_new_n27424__ = ys__n46456 & new_new_n12248__;
  assign new_new_n27425__ = ~new_new_n27423__ & ~new_new_n27424__;
  assign new_new_n27426__ = ys__n46632 & new_new_n12245__;
  assign new_new_n27427__ = ys__n46808 & new_new_n12246__;
  assign new_new_n27428__ = ~new_new_n27426__ & ~new_new_n27427__;
  assign new_new_n27429__ = new_new_n27425__ & new_new_n27428__;
  assign new_new_n27430__ = new_new_n26788__ & ~new_new_n27429__;
  assign new_new_n27431__ = ~new_new_n27422__ & ~new_new_n27430__;
  assign new_new_n27432__ = ys__n46329 & new_new_n12356__;
  assign new_new_n27433__ = ys__n46505 & new_new_n12248__;
  assign new_new_n27434__ = ~new_new_n27432__ & ~new_new_n27433__;
  assign new_new_n27435__ = ys__n46681 & new_new_n12245__;
  assign new_new_n27436__ = ys__n46857 & new_new_n12246__;
  assign new_new_n27437__ = ~new_new_n27435__ & ~new_new_n27436__;
  assign new_new_n27438__ = new_new_n27434__ & new_new_n27437__;
  assign new_new_n27439__ = new_new_n26798__ & ~new_new_n27438__;
  assign new_new_n27440__ = ys__n46406 & new_new_n12356__;
  assign new_new_n27441__ = ys__n46582 & new_new_n12248__;
  assign new_new_n27442__ = ~new_new_n27440__ & ~new_new_n27441__;
  assign new_new_n27443__ = ys__n46758 & new_new_n12245__;
  assign new_new_n27444__ = ys__n46934 & new_new_n12246__;
  assign new_new_n27445__ = ~new_new_n27443__ & ~new_new_n27444__;
  assign new_new_n27446__ = new_new_n27442__ & new_new_n27445__;
  assign new_new_n27447__ = new_new_n26807__ & ~new_new_n27446__;
  assign new_new_n27448__ = ~new_new_n27439__ & ~new_new_n27447__;
  assign new_new_n27449__ = new_new_n27431__ & new_new_n27448__;
  assign new_new_n27450__ = new_new_n26818__ & ~new_new_n27449__;
  assign new_new_n27451__ = ~new_new_n27414__ & ~new_new_n27450__;
  assign new_new_n27452__ = new_new_n26821__ & ~new_new_n27451__;
  assign new_new_n27453__ = ys__n45568 & new_new_n12356__;
  assign new_new_n27454__ = ys__n45404 & new_new_n12248__;
  assign new_new_n27455__ = ~new_new_n27453__ & ~new_new_n27454__;
  assign new_new_n27456__ = ys__n45240 & new_new_n12245__;
  assign new_new_n27457__ = ys__n45029 & new_new_n12246__;
  assign new_new_n27458__ = ~new_new_n27456__ & ~new_new_n27457__;
  assign new_new_n27459__ = new_new_n27455__ & new_new_n27458__;
  assign new_new_n27460__ = new_new_n26807__ & ~new_new_n27459__;
  assign new_new_n27461__ = ys__n45662 & new_new_n12356__;
  assign new_new_n27462__ = ys__n45498 & new_new_n12248__;
  assign new_new_n27463__ = ~new_new_n27461__ & ~new_new_n27462__;
  assign new_new_n27464__ = ys__n45334 & new_new_n12245__;
  assign new_new_n27465__ = ys__n45155 & new_new_n12246__;
  assign new_new_n27466__ = ~new_new_n27464__ & ~new_new_n27465__;
  assign new_new_n27467__ = new_new_n27463__ & new_new_n27466__;
  assign new_new_n27468__ = new_new_n26779__ & ~new_new_n27467__;
  assign new_new_n27469__ = ys__n45616 & new_new_n12356__;
  assign new_new_n27470__ = ys__n45452 & new_new_n12248__;
  assign new_new_n27471__ = ~new_new_n27469__ & ~new_new_n27470__;
  assign new_new_n27472__ = ys__n45288 & new_new_n12245__;
  assign new_new_n27473__ = ys__n45094 & new_new_n12246__;
  assign new_new_n27474__ = ~new_new_n27472__ & ~new_new_n27473__;
  assign new_new_n27475__ = new_new_n27471__ & new_new_n27474__;
  assign new_new_n27476__ = new_new_n26788__ & ~new_new_n27475__;
  assign new_new_n27477__ = ~new_new_n27468__ & ~new_new_n27476__;
  assign new_new_n27478__ = ~new_new_n27460__ & new_new_n27477__;
  assign new_new_n27479__ = new_new_n26859__ & ~new_new_n27478__;
  assign new_new_n27480__ = ~new_new_n27452__ & ~new_new_n27479__;
  assign new_new_n27481__ = new_new_n26862__ & ~new_new_n27480__;
  assign new_new_n27482__ = ys__n46109 & new_new_n12356__;
  assign new_new_n27483__ = ys__n46011 & new_new_n12248__;
  assign new_new_n27484__ = ~new_new_n27482__ & ~new_new_n27483__;
  assign new_new_n27485__ = ys__n45913 & new_new_n12245__;
  assign new_new_n27486__ = ys__n45817 & new_new_n12246__;
  assign new_new_n27487__ = ~new_new_n27485__ & ~new_new_n27486__;
  assign new_new_n27488__ = new_new_n27484__ & new_new_n27487__;
  assign new_new_n27489__ = new_new_n26788__ & ~new_new_n27488__;
  assign new_new_n27490__ = ys__n46060 & new_new_n12356__;
  assign new_new_n27491__ = ys__n45962 & new_new_n12248__;
  assign new_new_n27492__ = ~new_new_n27490__ & ~new_new_n27491__;
  assign new_new_n27493__ = ys__n45864 & new_new_n12245__;
  assign new_new_n27494__ = ys__n45751 & new_new_n12246__;
  assign new_new_n27495__ = ~new_new_n27493__ & ~new_new_n27494__;
  assign new_new_n27496__ = new_new_n27492__ & new_new_n27495__;
  assign new_new_n27497__ = new_new_n26807__ & ~new_new_n27496__;
  assign new_new_n27498__ = ~new_new_n27489__ & ~new_new_n27497__;
  assign new_new_n27499__ = new_new_n26882__ & ~new_new_n27498__;
  assign new_new_n27500__ = ~new_new_n26862__ & new_new_n27499__;
  assign ys__n26125 = new_new_n27481__ | new_new_n27500__;
  assign new_new_n27502__ = ys__n26026 & new_new_n26768__;
  assign new_new_n27503__ = ys__n46360 & new_new_n12356__;
  assign new_new_n27504__ = ys__n46536 & new_new_n12248__;
  assign new_new_n27505__ = ~new_new_n27503__ & ~new_new_n27504__;
  assign new_new_n27506__ = ys__n46712 & new_new_n12245__;
  assign new_new_n27507__ = ys__n46888 & new_new_n12246__;
  assign new_new_n27508__ = ~new_new_n27506__ & ~new_new_n27507__;
  assign new_new_n27509__ = new_new_n27505__ & new_new_n27508__;
  assign new_new_n27510__ = new_new_n26779__ & ~new_new_n27509__;
  assign new_new_n27511__ = ys__n46282 & new_new_n12356__;
  assign new_new_n27512__ = ys__n46458 & new_new_n12248__;
  assign new_new_n27513__ = ~new_new_n27511__ & ~new_new_n27512__;
  assign new_new_n27514__ = ys__n46634 & new_new_n12245__;
  assign new_new_n27515__ = ys__n46810 & new_new_n12246__;
  assign new_new_n27516__ = ~new_new_n27514__ & ~new_new_n27515__;
  assign new_new_n27517__ = new_new_n27513__ & new_new_n27516__;
  assign new_new_n27518__ = new_new_n26788__ & ~new_new_n27517__;
  assign new_new_n27519__ = ~new_new_n27510__ & ~new_new_n27518__;
  assign new_new_n27520__ = ys__n46330 & new_new_n12356__;
  assign new_new_n27521__ = ys__n46506 & new_new_n12248__;
  assign new_new_n27522__ = ~new_new_n27520__ & ~new_new_n27521__;
  assign new_new_n27523__ = ys__n46682 & new_new_n12245__;
  assign new_new_n27524__ = ys__n46858 & new_new_n12246__;
  assign new_new_n27525__ = ~new_new_n27523__ & ~new_new_n27524__;
  assign new_new_n27526__ = new_new_n27522__ & new_new_n27525__;
  assign new_new_n27527__ = new_new_n26798__ & ~new_new_n27526__;
  assign new_new_n27528__ = ys__n46407 & new_new_n12356__;
  assign new_new_n27529__ = ys__n46583 & new_new_n12248__;
  assign new_new_n27530__ = ~new_new_n27528__ & ~new_new_n27529__;
  assign new_new_n27531__ = ys__n46759 & new_new_n12245__;
  assign new_new_n27532__ = ys__n46935 & new_new_n12246__;
  assign new_new_n27533__ = ~new_new_n27531__ & ~new_new_n27532__;
  assign new_new_n27534__ = new_new_n27530__ & new_new_n27533__;
  assign new_new_n27535__ = new_new_n26807__ & ~new_new_n27534__;
  assign new_new_n27536__ = ~new_new_n27527__ & ~new_new_n27535__;
  assign new_new_n27537__ = new_new_n27519__ & new_new_n27536__;
  assign new_new_n27538__ = new_new_n26818__ & ~new_new_n27537__;
  assign new_new_n27539__ = ~new_new_n27502__ & ~new_new_n27538__;
  assign new_new_n27540__ = new_new_n26821__ & ~new_new_n27539__;
  assign new_new_n27541__ = ys__n45570 & new_new_n12356__;
  assign new_new_n27542__ = ys__n45406 & new_new_n12248__;
  assign new_new_n27543__ = ~new_new_n27541__ & ~new_new_n27542__;
  assign new_new_n27544__ = ys__n45242 & new_new_n12245__;
  assign new_new_n27545__ = ys__n45032 & new_new_n12246__;
  assign new_new_n27546__ = ~new_new_n27544__ & ~new_new_n27545__;
  assign new_new_n27547__ = new_new_n27543__ & new_new_n27546__;
  assign new_new_n27548__ = new_new_n26807__ & ~new_new_n27547__;
  assign new_new_n27549__ = ys__n45664 & new_new_n12356__;
  assign new_new_n27550__ = ys__n45500 & new_new_n12248__;
  assign new_new_n27551__ = ~new_new_n27549__ & ~new_new_n27550__;
  assign new_new_n27552__ = ys__n45336 & new_new_n12245__;
  assign new_new_n27553__ = ys__n45158 & new_new_n12246__;
  assign new_new_n27554__ = ~new_new_n27552__ & ~new_new_n27553__;
  assign new_new_n27555__ = new_new_n27551__ & new_new_n27554__;
  assign new_new_n27556__ = new_new_n26779__ & ~new_new_n27555__;
  assign new_new_n27557__ = ys__n45617 & new_new_n12356__;
  assign new_new_n27558__ = ys__n45453 & new_new_n12248__;
  assign new_new_n27559__ = ~new_new_n27557__ & ~new_new_n27558__;
  assign new_new_n27560__ = ys__n45289 & new_new_n12245__;
  assign new_new_n27561__ = ys__n45095 & new_new_n12246__;
  assign new_new_n27562__ = ~new_new_n27560__ & ~new_new_n27561__;
  assign new_new_n27563__ = new_new_n27559__ & new_new_n27562__;
  assign new_new_n27564__ = new_new_n26788__ & ~new_new_n27563__;
  assign new_new_n27565__ = ~new_new_n27556__ & ~new_new_n27564__;
  assign new_new_n27566__ = ~new_new_n27548__ & new_new_n27565__;
  assign new_new_n27567__ = new_new_n26859__ & ~new_new_n27566__;
  assign new_new_n27568__ = ~new_new_n27540__ & ~new_new_n27567__;
  assign new_new_n27569__ = new_new_n26862__ & ~new_new_n27568__;
  assign new_new_n27570__ = ys__n46110 & new_new_n12356__;
  assign new_new_n27571__ = ys__n46012 & new_new_n12248__;
  assign new_new_n27572__ = ~new_new_n27570__ & ~new_new_n27571__;
  assign new_new_n27573__ = ys__n45914 & new_new_n12245__;
  assign new_new_n27574__ = ys__n45818 & new_new_n12246__;
  assign new_new_n27575__ = ~new_new_n27573__ & ~new_new_n27574__;
  assign new_new_n27576__ = new_new_n27572__ & new_new_n27575__;
  assign new_new_n27577__ = new_new_n26788__ & ~new_new_n27576__;
  assign new_new_n27578__ = ys__n46062 & new_new_n12356__;
  assign new_new_n27579__ = ys__n45964 & new_new_n12248__;
  assign new_new_n27580__ = ~new_new_n27578__ & ~new_new_n27579__;
  assign new_new_n27581__ = ys__n45866 & new_new_n12245__;
  assign new_new_n27582__ = ys__n45754 & new_new_n12246__;
  assign new_new_n27583__ = ~new_new_n27581__ & ~new_new_n27582__;
  assign new_new_n27584__ = new_new_n27580__ & new_new_n27583__;
  assign new_new_n27585__ = new_new_n26807__ & ~new_new_n27584__;
  assign new_new_n27586__ = ~new_new_n27577__ & ~new_new_n27585__;
  assign new_new_n27587__ = new_new_n26882__ & ~new_new_n27586__;
  assign new_new_n27588__ = ~new_new_n26862__ & new_new_n27587__;
  assign ys__n26126 = new_new_n27569__ | new_new_n27588__;
  assign new_new_n27590__ = ys__n26029 & new_new_n26768__;
  assign new_new_n27591__ = ys__n46362 & new_new_n12356__;
  assign new_new_n27592__ = ys__n46538 & new_new_n12248__;
  assign new_new_n27593__ = ~new_new_n27591__ & ~new_new_n27592__;
  assign new_new_n27594__ = ys__n46714 & new_new_n12245__;
  assign new_new_n27595__ = ys__n46890 & new_new_n12246__;
  assign new_new_n27596__ = ~new_new_n27594__ & ~new_new_n27595__;
  assign new_new_n27597__ = new_new_n27593__ & new_new_n27596__;
  assign new_new_n27598__ = new_new_n26779__ & ~new_new_n27597__;
  assign new_new_n27599__ = ys__n46284 & new_new_n12356__;
  assign new_new_n27600__ = ys__n46460 & new_new_n12248__;
  assign new_new_n27601__ = ~new_new_n27599__ & ~new_new_n27600__;
  assign new_new_n27602__ = ys__n46636 & new_new_n12245__;
  assign new_new_n27603__ = ys__n46812 & new_new_n12246__;
  assign new_new_n27604__ = ~new_new_n27602__ & ~new_new_n27603__;
  assign new_new_n27605__ = new_new_n27601__ & new_new_n27604__;
  assign new_new_n27606__ = new_new_n26788__ & ~new_new_n27605__;
  assign new_new_n27607__ = ~new_new_n27598__ & ~new_new_n27606__;
  assign new_new_n27608__ = ys__n46331 & new_new_n12356__;
  assign new_new_n27609__ = ys__n46507 & new_new_n12248__;
  assign new_new_n27610__ = ~new_new_n27608__ & ~new_new_n27609__;
  assign new_new_n27611__ = ys__n46683 & new_new_n12245__;
  assign new_new_n27612__ = ys__n46859 & new_new_n12246__;
  assign new_new_n27613__ = ~new_new_n27611__ & ~new_new_n27612__;
  assign new_new_n27614__ = new_new_n27610__ & new_new_n27613__;
  assign new_new_n27615__ = new_new_n26798__ & ~new_new_n27614__;
  assign new_new_n27616__ = ys__n46408 & new_new_n12356__;
  assign new_new_n27617__ = ys__n46584 & new_new_n12248__;
  assign new_new_n27618__ = ~new_new_n27616__ & ~new_new_n27617__;
  assign new_new_n27619__ = ys__n46760 & new_new_n12245__;
  assign new_new_n27620__ = ys__n46936 & new_new_n12246__;
  assign new_new_n27621__ = ~new_new_n27619__ & ~new_new_n27620__;
  assign new_new_n27622__ = new_new_n27618__ & new_new_n27621__;
  assign new_new_n27623__ = new_new_n26807__ & ~new_new_n27622__;
  assign new_new_n27624__ = ~new_new_n27615__ & ~new_new_n27623__;
  assign new_new_n27625__ = new_new_n27607__ & new_new_n27624__;
  assign new_new_n27626__ = new_new_n26818__ & ~new_new_n27625__;
  assign new_new_n27627__ = ~new_new_n27590__ & ~new_new_n27626__;
  assign new_new_n27628__ = new_new_n26821__ & ~new_new_n27627__;
  assign new_new_n27629__ = ys__n45572 & new_new_n12356__;
  assign new_new_n27630__ = ys__n45408 & new_new_n12248__;
  assign new_new_n27631__ = ~new_new_n27629__ & ~new_new_n27630__;
  assign new_new_n27632__ = ys__n45244 & new_new_n12245__;
  assign new_new_n27633__ = ys__n45035 & new_new_n12246__;
  assign new_new_n27634__ = ~new_new_n27632__ & ~new_new_n27633__;
  assign new_new_n27635__ = new_new_n27631__ & new_new_n27634__;
  assign new_new_n27636__ = new_new_n26807__ & ~new_new_n27635__;
  assign new_new_n27637__ = ys__n45666 & new_new_n12356__;
  assign new_new_n27638__ = ys__n45502 & new_new_n12248__;
  assign new_new_n27639__ = ~new_new_n27637__ & ~new_new_n27638__;
  assign new_new_n27640__ = ys__n45338 & new_new_n12245__;
  assign new_new_n27641__ = ys__n45161 & new_new_n12246__;
  assign new_new_n27642__ = ~new_new_n27640__ & ~new_new_n27641__;
  assign new_new_n27643__ = new_new_n27639__ & new_new_n27642__;
  assign new_new_n27644__ = new_new_n26779__ & ~new_new_n27643__;
  assign new_new_n27645__ = ys__n45618 & new_new_n12356__;
  assign new_new_n27646__ = ys__n45454 & new_new_n12248__;
  assign new_new_n27647__ = ~new_new_n27645__ & ~new_new_n27646__;
  assign new_new_n27648__ = ys__n45290 & new_new_n12245__;
  assign new_new_n27649__ = ys__n45096 & new_new_n12246__;
  assign new_new_n27650__ = ~new_new_n27648__ & ~new_new_n27649__;
  assign new_new_n27651__ = new_new_n27647__ & new_new_n27650__;
  assign new_new_n27652__ = new_new_n26788__ & ~new_new_n27651__;
  assign new_new_n27653__ = ~new_new_n27644__ & ~new_new_n27652__;
  assign new_new_n27654__ = ~new_new_n27636__ & new_new_n27653__;
  assign new_new_n27655__ = new_new_n26859__ & ~new_new_n27654__;
  assign new_new_n27656__ = ~new_new_n27628__ & ~new_new_n27655__;
  assign new_new_n27657__ = new_new_n26862__ & ~new_new_n27656__;
  assign new_new_n27658__ = ys__n46111 & new_new_n12356__;
  assign new_new_n27659__ = ys__n46013 & new_new_n12248__;
  assign new_new_n27660__ = ~new_new_n27658__ & ~new_new_n27659__;
  assign new_new_n27661__ = ys__n45915 & new_new_n12245__;
  assign new_new_n27662__ = ys__n45819 & new_new_n12246__;
  assign new_new_n27663__ = ~new_new_n27661__ & ~new_new_n27662__;
  assign new_new_n27664__ = new_new_n27660__ & new_new_n27663__;
  assign new_new_n27665__ = new_new_n26788__ & ~new_new_n27664__;
  assign new_new_n27666__ = ys__n46064 & new_new_n12356__;
  assign new_new_n27667__ = ys__n45966 & new_new_n12248__;
  assign new_new_n27668__ = ~new_new_n27666__ & ~new_new_n27667__;
  assign new_new_n27669__ = ys__n45868 & new_new_n12245__;
  assign new_new_n27670__ = ys__n45757 & new_new_n12246__;
  assign new_new_n27671__ = ~new_new_n27669__ & ~new_new_n27670__;
  assign new_new_n27672__ = new_new_n27668__ & new_new_n27671__;
  assign new_new_n27673__ = new_new_n26807__ & ~new_new_n27672__;
  assign new_new_n27674__ = ~new_new_n27665__ & ~new_new_n27673__;
  assign new_new_n27675__ = new_new_n26882__ & ~new_new_n27674__;
  assign new_new_n27676__ = ~new_new_n26862__ & new_new_n27675__;
  assign ys__n26127 = new_new_n27657__ | new_new_n27676__;
  assign new_new_n27678__ = ys__n26032 & new_new_n26768__;
  assign new_new_n27679__ = ys__n46364 & new_new_n12356__;
  assign new_new_n27680__ = ys__n46540 & new_new_n12248__;
  assign new_new_n27681__ = ~new_new_n27679__ & ~new_new_n27680__;
  assign new_new_n27682__ = ys__n46716 & new_new_n12245__;
  assign new_new_n27683__ = ys__n46892 & new_new_n12246__;
  assign new_new_n27684__ = ~new_new_n27682__ & ~new_new_n27683__;
  assign new_new_n27685__ = new_new_n27681__ & new_new_n27684__;
  assign new_new_n27686__ = new_new_n26779__ & ~new_new_n27685__;
  assign new_new_n27687__ = ys__n46286 & new_new_n12356__;
  assign new_new_n27688__ = ys__n46462 & new_new_n12248__;
  assign new_new_n27689__ = ~new_new_n27687__ & ~new_new_n27688__;
  assign new_new_n27690__ = ys__n46638 & new_new_n12245__;
  assign new_new_n27691__ = ys__n46814 & new_new_n12246__;
  assign new_new_n27692__ = ~new_new_n27690__ & ~new_new_n27691__;
  assign new_new_n27693__ = new_new_n27689__ & new_new_n27692__;
  assign new_new_n27694__ = new_new_n26788__ & ~new_new_n27693__;
  assign new_new_n27695__ = ~new_new_n27686__ & ~new_new_n27694__;
  assign new_new_n27696__ = ys__n46332 & new_new_n12356__;
  assign new_new_n27697__ = ys__n46508 & new_new_n12248__;
  assign new_new_n27698__ = ~new_new_n27696__ & ~new_new_n27697__;
  assign new_new_n27699__ = ys__n46684 & new_new_n12245__;
  assign new_new_n27700__ = ys__n46860 & new_new_n12246__;
  assign new_new_n27701__ = ~new_new_n27699__ & ~new_new_n27700__;
  assign new_new_n27702__ = new_new_n27698__ & new_new_n27701__;
  assign new_new_n27703__ = new_new_n26798__ & ~new_new_n27702__;
  assign new_new_n27704__ = ys__n46409 & new_new_n12356__;
  assign new_new_n27705__ = ys__n46585 & new_new_n12248__;
  assign new_new_n27706__ = ~new_new_n27704__ & ~new_new_n27705__;
  assign new_new_n27707__ = ys__n46761 & new_new_n12245__;
  assign new_new_n27708__ = ys__n46937 & new_new_n12246__;
  assign new_new_n27709__ = ~new_new_n27707__ & ~new_new_n27708__;
  assign new_new_n27710__ = new_new_n27706__ & new_new_n27709__;
  assign new_new_n27711__ = new_new_n26807__ & ~new_new_n27710__;
  assign new_new_n27712__ = ~new_new_n27703__ & ~new_new_n27711__;
  assign new_new_n27713__ = new_new_n27695__ & new_new_n27712__;
  assign new_new_n27714__ = new_new_n26818__ & ~new_new_n27713__;
  assign new_new_n27715__ = ~new_new_n27678__ & ~new_new_n27714__;
  assign new_new_n27716__ = new_new_n26821__ & ~new_new_n27715__;
  assign new_new_n27717__ = ys__n45574 & new_new_n12356__;
  assign new_new_n27718__ = ys__n45410 & new_new_n12248__;
  assign new_new_n27719__ = ~new_new_n27717__ & ~new_new_n27718__;
  assign new_new_n27720__ = ys__n45246 & new_new_n12245__;
  assign new_new_n27721__ = ys__n45038 & new_new_n12246__;
  assign new_new_n27722__ = ~new_new_n27720__ & ~new_new_n27721__;
  assign new_new_n27723__ = new_new_n27719__ & new_new_n27722__;
  assign new_new_n27724__ = new_new_n26807__ & ~new_new_n27723__;
  assign new_new_n27725__ = ys__n45668 & new_new_n12356__;
  assign new_new_n27726__ = ys__n45504 & new_new_n12248__;
  assign new_new_n27727__ = ~new_new_n27725__ & ~new_new_n27726__;
  assign new_new_n27728__ = ys__n45340 & new_new_n12245__;
  assign new_new_n27729__ = ys__n45164 & new_new_n12246__;
  assign new_new_n27730__ = ~new_new_n27728__ & ~new_new_n27729__;
  assign new_new_n27731__ = new_new_n27727__ & new_new_n27730__;
  assign new_new_n27732__ = new_new_n26779__ & ~new_new_n27731__;
  assign new_new_n27733__ = ys__n45619 & new_new_n12356__;
  assign new_new_n27734__ = ys__n45455 & new_new_n12248__;
  assign new_new_n27735__ = ~new_new_n27733__ & ~new_new_n27734__;
  assign new_new_n27736__ = ys__n45291 & new_new_n12245__;
  assign new_new_n27737__ = ys__n45097 & new_new_n12246__;
  assign new_new_n27738__ = ~new_new_n27736__ & ~new_new_n27737__;
  assign new_new_n27739__ = new_new_n27735__ & new_new_n27738__;
  assign new_new_n27740__ = new_new_n26788__ & ~new_new_n27739__;
  assign new_new_n27741__ = ~new_new_n27732__ & ~new_new_n27740__;
  assign new_new_n27742__ = ~new_new_n27724__ & new_new_n27741__;
  assign new_new_n27743__ = new_new_n26859__ & ~new_new_n27742__;
  assign new_new_n27744__ = ~new_new_n27716__ & ~new_new_n27743__;
  assign new_new_n27745__ = new_new_n26862__ & ~new_new_n27744__;
  assign new_new_n27746__ = ys__n46112 & new_new_n12356__;
  assign new_new_n27747__ = ys__n46014 & new_new_n12248__;
  assign new_new_n27748__ = ~new_new_n27746__ & ~new_new_n27747__;
  assign new_new_n27749__ = ys__n45916 & new_new_n12245__;
  assign new_new_n27750__ = ys__n45820 & new_new_n12246__;
  assign new_new_n27751__ = ~new_new_n27749__ & ~new_new_n27750__;
  assign new_new_n27752__ = new_new_n27748__ & new_new_n27751__;
  assign new_new_n27753__ = new_new_n26788__ & ~new_new_n27752__;
  assign new_new_n27754__ = ys__n46066 & new_new_n12356__;
  assign new_new_n27755__ = ys__n45968 & new_new_n12248__;
  assign new_new_n27756__ = ~new_new_n27754__ & ~new_new_n27755__;
  assign new_new_n27757__ = ys__n45870 & new_new_n12245__;
  assign new_new_n27758__ = ys__n45760 & new_new_n12246__;
  assign new_new_n27759__ = ~new_new_n27757__ & ~new_new_n27758__;
  assign new_new_n27760__ = new_new_n27756__ & new_new_n27759__;
  assign new_new_n27761__ = new_new_n26807__ & ~new_new_n27760__;
  assign new_new_n27762__ = ~new_new_n27753__ & ~new_new_n27761__;
  assign new_new_n27763__ = new_new_n26882__ & ~new_new_n27762__;
  assign new_new_n27764__ = ~new_new_n26862__ & new_new_n27763__;
  assign ys__n26128 = new_new_n27745__ | new_new_n27764__;
  assign new_new_n27766__ = ys__n26035 & new_new_n26768__;
  assign new_new_n27767__ = ys__n46366 & new_new_n12356__;
  assign new_new_n27768__ = ys__n46542 & new_new_n12248__;
  assign new_new_n27769__ = ~new_new_n27767__ & ~new_new_n27768__;
  assign new_new_n27770__ = ys__n46718 & new_new_n12245__;
  assign new_new_n27771__ = ys__n46894 & new_new_n12246__;
  assign new_new_n27772__ = ~new_new_n27770__ & ~new_new_n27771__;
  assign new_new_n27773__ = new_new_n27769__ & new_new_n27772__;
  assign new_new_n27774__ = new_new_n26779__ & ~new_new_n27773__;
  assign new_new_n27775__ = ys__n46288 & new_new_n12356__;
  assign new_new_n27776__ = ys__n46464 & new_new_n12248__;
  assign new_new_n27777__ = ~new_new_n27775__ & ~new_new_n27776__;
  assign new_new_n27778__ = ys__n46640 & new_new_n12245__;
  assign new_new_n27779__ = ys__n46816 & new_new_n12246__;
  assign new_new_n27780__ = ~new_new_n27778__ & ~new_new_n27779__;
  assign new_new_n27781__ = new_new_n27777__ & new_new_n27780__;
  assign new_new_n27782__ = new_new_n26788__ & ~new_new_n27781__;
  assign new_new_n27783__ = ~new_new_n27774__ & ~new_new_n27782__;
  assign new_new_n27784__ = ys__n46333 & new_new_n12356__;
  assign new_new_n27785__ = ys__n46509 & new_new_n12248__;
  assign new_new_n27786__ = ~new_new_n27784__ & ~new_new_n27785__;
  assign new_new_n27787__ = ys__n46685 & new_new_n12245__;
  assign new_new_n27788__ = ys__n46861 & new_new_n12246__;
  assign new_new_n27789__ = ~new_new_n27787__ & ~new_new_n27788__;
  assign new_new_n27790__ = new_new_n27786__ & new_new_n27789__;
  assign new_new_n27791__ = new_new_n26798__ & ~new_new_n27790__;
  assign new_new_n27792__ = ys__n46410 & new_new_n12356__;
  assign new_new_n27793__ = ys__n46586 & new_new_n12248__;
  assign new_new_n27794__ = ~new_new_n27792__ & ~new_new_n27793__;
  assign new_new_n27795__ = ys__n46762 & new_new_n12245__;
  assign new_new_n27796__ = ys__n46938 & new_new_n12246__;
  assign new_new_n27797__ = ~new_new_n27795__ & ~new_new_n27796__;
  assign new_new_n27798__ = new_new_n27794__ & new_new_n27797__;
  assign new_new_n27799__ = new_new_n26807__ & ~new_new_n27798__;
  assign new_new_n27800__ = ~new_new_n27791__ & ~new_new_n27799__;
  assign new_new_n27801__ = new_new_n27783__ & new_new_n27800__;
  assign new_new_n27802__ = new_new_n26818__ & ~new_new_n27801__;
  assign new_new_n27803__ = ~new_new_n27766__ & ~new_new_n27802__;
  assign new_new_n27804__ = new_new_n26821__ & ~new_new_n27803__;
  assign new_new_n27805__ = ys__n45576 & new_new_n12356__;
  assign new_new_n27806__ = ys__n45412 & new_new_n12248__;
  assign new_new_n27807__ = ~new_new_n27805__ & ~new_new_n27806__;
  assign new_new_n27808__ = ys__n45248 & new_new_n12245__;
  assign new_new_n27809__ = ys__n45041 & new_new_n12246__;
  assign new_new_n27810__ = ~new_new_n27808__ & ~new_new_n27809__;
  assign new_new_n27811__ = new_new_n27807__ & new_new_n27810__;
  assign new_new_n27812__ = new_new_n26807__ & ~new_new_n27811__;
  assign new_new_n27813__ = ys__n45670 & new_new_n12356__;
  assign new_new_n27814__ = ys__n45506 & new_new_n12248__;
  assign new_new_n27815__ = ~new_new_n27813__ & ~new_new_n27814__;
  assign new_new_n27816__ = ys__n45342 & new_new_n12245__;
  assign new_new_n27817__ = ys__n45167 & new_new_n12246__;
  assign new_new_n27818__ = ~new_new_n27816__ & ~new_new_n27817__;
  assign new_new_n27819__ = new_new_n27815__ & new_new_n27818__;
  assign new_new_n27820__ = new_new_n26779__ & ~new_new_n27819__;
  assign new_new_n27821__ = ys__n45620 & new_new_n12356__;
  assign new_new_n27822__ = ys__n45456 & new_new_n12248__;
  assign new_new_n27823__ = ~new_new_n27821__ & ~new_new_n27822__;
  assign new_new_n27824__ = ys__n45292 & new_new_n12245__;
  assign new_new_n27825__ = ys__n45098 & new_new_n12246__;
  assign new_new_n27826__ = ~new_new_n27824__ & ~new_new_n27825__;
  assign new_new_n27827__ = new_new_n27823__ & new_new_n27826__;
  assign new_new_n27828__ = new_new_n26788__ & ~new_new_n27827__;
  assign new_new_n27829__ = ~new_new_n27820__ & ~new_new_n27828__;
  assign new_new_n27830__ = ~new_new_n27812__ & new_new_n27829__;
  assign new_new_n27831__ = new_new_n26859__ & ~new_new_n27830__;
  assign new_new_n27832__ = ~new_new_n27804__ & ~new_new_n27831__;
  assign new_new_n27833__ = new_new_n26862__ & ~new_new_n27832__;
  assign new_new_n27834__ = ys__n46113 & new_new_n12356__;
  assign new_new_n27835__ = ys__n46015 & new_new_n12248__;
  assign new_new_n27836__ = ~new_new_n27834__ & ~new_new_n27835__;
  assign new_new_n27837__ = ys__n45917 & new_new_n12245__;
  assign new_new_n27838__ = ys__n45821 & new_new_n12246__;
  assign new_new_n27839__ = ~new_new_n27837__ & ~new_new_n27838__;
  assign new_new_n27840__ = new_new_n27836__ & new_new_n27839__;
  assign new_new_n27841__ = new_new_n26788__ & ~new_new_n27840__;
  assign new_new_n27842__ = ys__n46068 & new_new_n12356__;
  assign new_new_n27843__ = ys__n45970 & new_new_n12248__;
  assign new_new_n27844__ = ~new_new_n27842__ & ~new_new_n27843__;
  assign new_new_n27845__ = ys__n45872 & new_new_n12245__;
  assign new_new_n27846__ = ys__n45763 & new_new_n12246__;
  assign new_new_n27847__ = ~new_new_n27845__ & ~new_new_n27846__;
  assign new_new_n27848__ = new_new_n27844__ & new_new_n27847__;
  assign new_new_n27849__ = new_new_n26807__ & ~new_new_n27848__;
  assign new_new_n27850__ = ~new_new_n27841__ & ~new_new_n27849__;
  assign new_new_n27851__ = new_new_n26882__ & ~new_new_n27850__;
  assign new_new_n27852__ = ~new_new_n26862__ & new_new_n27851__;
  assign ys__n26129 = new_new_n27833__ | new_new_n27852__;
  assign new_new_n27854__ = ys__n26038 & new_new_n26768__;
  assign new_new_n27855__ = ys__n46368 & new_new_n12356__;
  assign new_new_n27856__ = ys__n46544 & new_new_n12248__;
  assign new_new_n27857__ = ~new_new_n27855__ & ~new_new_n27856__;
  assign new_new_n27858__ = ys__n46720 & new_new_n12245__;
  assign new_new_n27859__ = ys__n46896 & new_new_n12246__;
  assign new_new_n27860__ = ~new_new_n27858__ & ~new_new_n27859__;
  assign new_new_n27861__ = new_new_n27857__ & new_new_n27860__;
  assign new_new_n27862__ = new_new_n26779__ & ~new_new_n27861__;
  assign new_new_n27863__ = ys__n46290 & new_new_n12356__;
  assign new_new_n27864__ = ys__n46466 & new_new_n12248__;
  assign new_new_n27865__ = ~new_new_n27863__ & ~new_new_n27864__;
  assign new_new_n27866__ = ys__n46642 & new_new_n12245__;
  assign new_new_n27867__ = ys__n46818 & new_new_n12246__;
  assign new_new_n27868__ = ~new_new_n27866__ & ~new_new_n27867__;
  assign new_new_n27869__ = new_new_n27865__ & new_new_n27868__;
  assign new_new_n27870__ = new_new_n26788__ & ~new_new_n27869__;
  assign new_new_n27871__ = ~new_new_n27862__ & ~new_new_n27870__;
  assign new_new_n27872__ = ys__n46334 & new_new_n12356__;
  assign new_new_n27873__ = ys__n46510 & new_new_n12248__;
  assign new_new_n27874__ = ~new_new_n27872__ & ~new_new_n27873__;
  assign new_new_n27875__ = ys__n46686 & new_new_n12245__;
  assign new_new_n27876__ = ys__n46862 & new_new_n12246__;
  assign new_new_n27877__ = ~new_new_n27875__ & ~new_new_n27876__;
  assign new_new_n27878__ = new_new_n27874__ & new_new_n27877__;
  assign new_new_n27879__ = new_new_n26798__ & ~new_new_n27878__;
  assign new_new_n27880__ = ys__n46411 & new_new_n12356__;
  assign new_new_n27881__ = ys__n46587 & new_new_n12248__;
  assign new_new_n27882__ = ~new_new_n27880__ & ~new_new_n27881__;
  assign new_new_n27883__ = ys__n46763 & new_new_n12245__;
  assign new_new_n27884__ = ys__n46939 & new_new_n12246__;
  assign new_new_n27885__ = ~new_new_n27883__ & ~new_new_n27884__;
  assign new_new_n27886__ = new_new_n27882__ & new_new_n27885__;
  assign new_new_n27887__ = new_new_n26807__ & ~new_new_n27886__;
  assign new_new_n27888__ = ~new_new_n27879__ & ~new_new_n27887__;
  assign new_new_n27889__ = new_new_n27871__ & new_new_n27888__;
  assign new_new_n27890__ = new_new_n26818__ & ~new_new_n27889__;
  assign new_new_n27891__ = ~new_new_n27854__ & ~new_new_n27890__;
  assign new_new_n27892__ = new_new_n26821__ & ~new_new_n27891__;
  assign new_new_n27893__ = ys__n45578 & new_new_n12356__;
  assign new_new_n27894__ = ys__n45414 & new_new_n12248__;
  assign new_new_n27895__ = ~new_new_n27893__ & ~new_new_n27894__;
  assign new_new_n27896__ = ys__n45250 & new_new_n12245__;
  assign new_new_n27897__ = ys__n45044 & new_new_n12246__;
  assign new_new_n27898__ = ~new_new_n27896__ & ~new_new_n27897__;
  assign new_new_n27899__ = new_new_n27895__ & new_new_n27898__;
  assign new_new_n27900__ = new_new_n26807__ & ~new_new_n27899__;
  assign new_new_n27901__ = ys__n45672 & new_new_n12356__;
  assign new_new_n27902__ = ys__n45508 & new_new_n12248__;
  assign new_new_n27903__ = ~new_new_n27901__ & ~new_new_n27902__;
  assign new_new_n27904__ = ys__n45344 & new_new_n12245__;
  assign new_new_n27905__ = ys__n45170 & new_new_n12246__;
  assign new_new_n27906__ = ~new_new_n27904__ & ~new_new_n27905__;
  assign new_new_n27907__ = new_new_n27903__ & new_new_n27906__;
  assign new_new_n27908__ = new_new_n26779__ & ~new_new_n27907__;
  assign new_new_n27909__ = ys__n45621 & new_new_n12356__;
  assign new_new_n27910__ = ys__n45457 & new_new_n12248__;
  assign new_new_n27911__ = ~new_new_n27909__ & ~new_new_n27910__;
  assign new_new_n27912__ = ys__n45293 & new_new_n12245__;
  assign new_new_n27913__ = ys__n45099 & new_new_n12246__;
  assign new_new_n27914__ = ~new_new_n27912__ & ~new_new_n27913__;
  assign new_new_n27915__ = new_new_n27911__ & new_new_n27914__;
  assign new_new_n27916__ = new_new_n26788__ & ~new_new_n27915__;
  assign new_new_n27917__ = ~new_new_n27908__ & ~new_new_n27916__;
  assign new_new_n27918__ = ~new_new_n27900__ & new_new_n27917__;
  assign new_new_n27919__ = new_new_n26859__ & ~new_new_n27918__;
  assign new_new_n27920__ = ~new_new_n27892__ & ~new_new_n27919__;
  assign new_new_n27921__ = new_new_n26862__ & ~new_new_n27920__;
  assign new_new_n27922__ = ys__n46114 & new_new_n12356__;
  assign new_new_n27923__ = ys__n46016 & new_new_n12248__;
  assign new_new_n27924__ = ~new_new_n27922__ & ~new_new_n27923__;
  assign new_new_n27925__ = ys__n45918 & new_new_n12245__;
  assign new_new_n27926__ = ys__n45822 & new_new_n12246__;
  assign new_new_n27927__ = ~new_new_n27925__ & ~new_new_n27926__;
  assign new_new_n27928__ = new_new_n27924__ & new_new_n27927__;
  assign new_new_n27929__ = new_new_n26788__ & ~new_new_n27928__;
  assign new_new_n27930__ = ys__n46070 & new_new_n12356__;
  assign new_new_n27931__ = ys__n45972 & new_new_n12248__;
  assign new_new_n27932__ = ~new_new_n27930__ & ~new_new_n27931__;
  assign new_new_n27933__ = ys__n45874 & new_new_n12245__;
  assign new_new_n27934__ = ys__n45766 & new_new_n12246__;
  assign new_new_n27935__ = ~new_new_n27933__ & ~new_new_n27934__;
  assign new_new_n27936__ = new_new_n27932__ & new_new_n27935__;
  assign new_new_n27937__ = new_new_n26807__ & ~new_new_n27936__;
  assign new_new_n27938__ = ~new_new_n27929__ & ~new_new_n27937__;
  assign new_new_n27939__ = new_new_n26882__ & ~new_new_n27938__;
  assign new_new_n27940__ = ~new_new_n26862__ & new_new_n27939__;
  assign ys__n26130 = new_new_n27921__ | new_new_n27940__;
  assign new_new_n27942__ = ys__n26041 & new_new_n26768__;
  assign new_new_n27943__ = ys__n46370 & new_new_n12356__;
  assign new_new_n27944__ = ys__n46546 & new_new_n12248__;
  assign new_new_n27945__ = ~new_new_n27943__ & ~new_new_n27944__;
  assign new_new_n27946__ = ys__n46722 & new_new_n12245__;
  assign new_new_n27947__ = ys__n46898 & new_new_n12246__;
  assign new_new_n27948__ = ~new_new_n27946__ & ~new_new_n27947__;
  assign new_new_n27949__ = new_new_n27945__ & new_new_n27948__;
  assign new_new_n27950__ = new_new_n26779__ & ~new_new_n27949__;
  assign new_new_n27951__ = ys__n46292 & new_new_n12356__;
  assign new_new_n27952__ = ys__n46468 & new_new_n12248__;
  assign new_new_n27953__ = ~new_new_n27951__ & ~new_new_n27952__;
  assign new_new_n27954__ = ys__n46644 & new_new_n12245__;
  assign new_new_n27955__ = ys__n46820 & new_new_n12246__;
  assign new_new_n27956__ = ~new_new_n27954__ & ~new_new_n27955__;
  assign new_new_n27957__ = new_new_n27953__ & new_new_n27956__;
  assign new_new_n27958__ = new_new_n26788__ & ~new_new_n27957__;
  assign new_new_n27959__ = ~new_new_n27950__ & ~new_new_n27958__;
  assign new_new_n27960__ = ys__n46335 & new_new_n12356__;
  assign new_new_n27961__ = ys__n46511 & new_new_n12248__;
  assign new_new_n27962__ = ~new_new_n27960__ & ~new_new_n27961__;
  assign new_new_n27963__ = ys__n46687 & new_new_n12245__;
  assign new_new_n27964__ = ys__n46863 & new_new_n12246__;
  assign new_new_n27965__ = ~new_new_n27963__ & ~new_new_n27964__;
  assign new_new_n27966__ = new_new_n27962__ & new_new_n27965__;
  assign new_new_n27967__ = new_new_n26798__ & ~new_new_n27966__;
  assign new_new_n27968__ = ys__n46412 & new_new_n12356__;
  assign new_new_n27969__ = ys__n46588 & new_new_n12248__;
  assign new_new_n27970__ = ~new_new_n27968__ & ~new_new_n27969__;
  assign new_new_n27971__ = ys__n46764 & new_new_n12245__;
  assign new_new_n27972__ = ys__n46940 & new_new_n12246__;
  assign new_new_n27973__ = ~new_new_n27971__ & ~new_new_n27972__;
  assign new_new_n27974__ = new_new_n27970__ & new_new_n27973__;
  assign new_new_n27975__ = new_new_n26807__ & ~new_new_n27974__;
  assign new_new_n27976__ = ~new_new_n27967__ & ~new_new_n27975__;
  assign new_new_n27977__ = new_new_n27959__ & new_new_n27976__;
  assign new_new_n27978__ = new_new_n26818__ & ~new_new_n27977__;
  assign new_new_n27979__ = ~new_new_n27942__ & ~new_new_n27978__;
  assign new_new_n27980__ = new_new_n26821__ & ~new_new_n27979__;
  assign new_new_n27981__ = ys__n45580 & new_new_n12356__;
  assign new_new_n27982__ = ys__n45416 & new_new_n12248__;
  assign new_new_n27983__ = ~new_new_n27981__ & ~new_new_n27982__;
  assign new_new_n27984__ = ys__n45252 & new_new_n12245__;
  assign new_new_n27985__ = ys__n45047 & new_new_n12246__;
  assign new_new_n27986__ = ~new_new_n27984__ & ~new_new_n27985__;
  assign new_new_n27987__ = new_new_n27983__ & new_new_n27986__;
  assign new_new_n27988__ = new_new_n26807__ & ~new_new_n27987__;
  assign new_new_n27989__ = ys__n45674 & new_new_n12356__;
  assign new_new_n27990__ = ys__n45510 & new_new_n12248__;
  assign new_new_n27991__ = ~new_new_n27989__ & ~new_new_n27990__;
  assign new_new_n27992__ = ys__n45346 & new_new_n12245__;
  assign new_new_n27993__ = ys__n45173 & new_new_n12246__;
  assign new_new_n27994__ = ~new_new_n27992__ & ~new_new_n27993__;
  assign new_new_n27995__ = new_new_n27991__ & new_new_n27994__;
  assign new_new_n27996__ = new_new_n26779__ & ~new_new_n27995__;
  assign new_new_n27997__ = ys__n45622 & new_new_n12356__;
  assign new_new_n27998__ = ys__n45458 & new_new_n12248__;
  assign new_new_n27999__ = ~new_new_n27997__ & ~new_new_n27998__;
  assign new_new_n28000__ = ys__n45294 & new_new_n12245__;
  assign new_new_n28001__ = ys__n45100 & new_new_n12246__;
  assign new_new_n28002__ = ~new_new_n28000__ & ~new_new_n28001__;
  assign new_new_n28003__ = new_new_n27999__ & new_new_n28002__;
  assign new_new_n28004__ = new_new_n26788__ & ~new_new_n28003__;
  assign new_new_n28005__ = ~new_new_n27996__ & ~new_new_n28004__;
  assign new_new_n28006__ = ~new_new_n27988__ & new_new_n28005__;
  assign new_new_n28007__ = new_new_n26859__ & ~new_new_n28006__;
  assign new_new_n28008__ = ~new_new_n27980__ & ~new_new_n28007__;
  assign new_new_n28009__ = new_new_n26862__ & ~new_new_n28008__;
  assign new_new_n28010__ = ys__n46115 & new_new_n12356__;
  assign new_new_n28011__ = ys__n46017 & new_new_n12248__;
  assign new_new_n28012__ = ~new_new_n28010__ & ~new_new_n28011__;
  assign new_new_n28013__ = ys__n45919 & new_new_n12245__;
  assign new_new_n28014__ = ys__n45823 & new_new_n12246__;
  assign new_new_n28015__ = ~new_new_n28013__ & ~new_new_n28014__;
  assign new_new_n28016__ = new_new_n28012__ & new_new_n28015__;
  assign new_new_n28017__ = new_new_n26788__ & ~new_new_n28016__;
  assign new_new_n28018__ = ys__n46072 & new_new_n12356__;
  assign new_new_n28019__ = ys__n45974 & new_new_n12248__;
  assign new_new_n28020__ = ~new_new_n28018__ & ~new_new_n28019__;
  assign new_new_n28021__ = ys__n45876 & new_new_n12245__;
  assign new_new_n28022__ = ys__n45769 & new_new_n12246__;
  assign new_new_n28023__ = ~new_new_n28021__ & ~new_new_n28022__;
  assign new_new_n28024__ = new_new_n28020__ & new_new_n28023__;
  assign new_new_n28025__ = new_new_n26807__ & ~new_new_n28024__;
  assign new_new_n28026__ = ~new_new_n28017__ & ~new_new_n28025__;
  assign new_new_n28027__ = new_new_n26882__ & ~new_new_n28026__;
  assign new_new_n28028__ = ~new_new_n26862__ & new_new_n28027__;
  assign ys__n26131 = new_new_n28009__ | new_new_n28028__;
  assign new_new_n28030__ = ys__n26044 & new_new_n26768__;
  assign new_new_n28031__ = ys__n46372 & new_new_n12356__;
  assign new_new_n28032__ = ys__n46548 & new_new_n12248__;
  assign new_new_n28033__ = ~new_new_n28031__ & ~new_new_n28032__;
  assign new_new_n28034__ = ys__n46724 & new_new_n12245__;
  assign new_new_n28035__ = ys__n46900 & new_new_n12246__;
  assign new_new_n28036__ = ~new_new_n28034__ & ~new_new_n28035__;
  assign new_new_n28037__ = new_new_n28033__ & new_new_n28036__;
  assign new_new_n28038__ = new_new_n26779__ & ~new_new_n28037__;
  assign new_new_n28039__ = ys__n46294 & new_new_n12356__;
  assign new_new_n28040__ = ys__n46470 & new_new_n12248__;
  assign new_new_n28041__ = ~new_new_n28039__ & ~new_new_n28040__;
  assign new_new_n28042__ = ys__n46646 & new_new_n12245__;
  assign new_new_n28043__ = ys__n46822 & new_new_n12246__;
  assign new_new_n28044__ = ~new_new_n28042__ & ~new_new_n28043__;
  assign new_new_n28045__ = new_new_n28041__ & new_new_n28044__;
  assign new_new_n28046__ = new_new_n26788__ & ~new_new_n28045__;
  assign new_new_n28047__ = ~new_new_n28038__ & ~new_new_n28046__;
  assign new_new_n28048__ = ys__n46336 & new_new_n12356__;
  assign new_new_n28049__ = ys__n46512 & new_new_n12248__;
  assign new_new_n28050__ = ~new_new_n28048__ & ~new_new_n28049__;
  assign new_new_n28051__ = ys__n46688 & new_new_n12245__;
  assign new_new_n28052__ = ys__n46864 & new_new_n12246__;
  assign new_new_n28053__ = ~new_new_n28051__ & ~new_new_n28052__;
  assign new_new_n28054__ = new_new_n28050__ & new_new_n28053__;
  assign new_new_n28055__ = new_new_n26798__ & ~new_new_n28054__;
  assign new_new_n28056__ = ys__n46413 & new_new_n12356__;
  assign new_new_n28057__ = ys__n46589 & new_new_n12248__;
  assign new_new_n28058__ = ~new_new_n28056__ & ~new_new_n28057__;
  assign new_new_n28059__ = ys__n46765 & new_new_n12245__;
  assign new_new_n28060__ = ys__n46941 & new_new_n12246__;
  assign new_new_n28061__ = ~new_new_n28059__ & ~new_new_n28060__;
  assign new_new_n28062__ = new_new_n28058__ & new_new_n28061__;
  assign new_new_n28063__ = new_new_n26807__ & ~new_new_n28062__;
  assign new_new_n28064__ = ~new_new_n28055__ & ~new_new_n28063__;
  assign new_new_n28065__ = new_new_n28047__ & new_new_n28064__;
  assign new_new_n28066__ = new_new_n26818__ & ~new_new_n28065__;
  assign new_new_n28067__ = ~new_new_n28030__ & ~new_new_n28066__;
  assign new_new_n28068__ = new_new_n26821__ & ~new_new_n28067__;
  assign new_new_n28069__ = ys__n45582 & new_new_n12356__;
  assign new_new_n28070__ = ys__n45418 & new_new_n12248__;
  assign new_new_n28071__ = ~new_new_n28069__ & ~new_new_n28070__;
  assign new_new_n28072__ = ys__n45254 & new_new_n12245__;
  assign new_new_n28073__ = ys__n45050 & new_new_n12246__;
  assign new_new_n28074__ = ~new_new_n28072__ & ~new_new_n28073__;
  assign new_new_n28075__ = new_new_n28071__ & new_new_n28074__;
  assign new_new_n28076__ = new_new_n26807__ & ~new_new_n28075__;
  assign new_new_n28077__ = ys__n45676 & new_new_n12356__;
  assign new_new_n28078__ = ys__n45512 & new_new_n12248__;
  assign new_new_n28079__ = ~new_new_n28077__ & ~new_new_n28078__;
  assign new_new_n28080__ = ys__n45348 & new_new_n12245__;
  assign new_new_n28081__ = ys__n45176 & new_new_n12246__;
  assign new_new_n28082__ = ~new_new_n28080__ & ~new_new_n28081__;
  assign new_new_n28083__ = new_new_n28079__ & new_new_n28082__;
  assign new_new_n28084__ = new_new_n26779__ & ~new_new_n28083__;
  assign new_new_n28085__ = ys__n45623 & new_new_n12356__;
  assign new_new_n28086__ = ys__n45459 & new_new_n12248__;
  assign new_new_n28087__ = ~new_new_n28085__ & ~new_new_n28086__;
  assign new_new_n28088__ = ys__n45295 & new_new_n12245__;
  assign new_new_n28089__ = ys__n45101 & new_new_n12246__;
  assign new_new_n28090__ = ~new_new_n28088__ & ~new_new_n28089__;
  assign new_new_n28091__ = new_new_n28087__ & new_new_n28090__;
  assign new_new_n28092__ = new_new_n26788__ & ~new_new_n28091__;
  assign new_new_n28093__ = ~new_new_n28084__ & ~new_new_n28092__;
  assign new_new_n28094__ = ~new_new_n28076__ & new_new_n28093__;
  assign new_new_n28095__ = new_new_n26859__ & ~new_new_n28094__;
  assign new_new_n28096__ = ~new_new_n28068__ & ~new_new_n28095__;
  assign new_new_n28097__ = new_new_n26862__ & ~new_new_n28096__;
  assign new_new_n28098__ = ys__n46116 & new_new_n12356__;
  assign new_new_n28099__ = ys__n46018 & new_new_n12248__;
  assign new_new_n28100__ = ~new_new_n28098__ & ~new_new_n28099__;
  assign new_new_n28101__ = ys__n45920 & new_new_n12245__;
  assign new_new_n28102__ = ys__n45824 & new_new_n12246__;
  assign new_new_n28103__ = ~new_new_n28101__ & ~new_new_n28102__;
  assign new_new_n28104__ = new_new_n28100__ & new_new_n28103__;
  assign new_new_n28105__ = new_new_n26788__ & ~new_new_n28104__;
  assign new_new_n28106__ = ys__n46074 & new_new_n12356__;
  assign new_new_n28107__ = ys__n45976 & new_new_n12248__;
  assign new_new_n28108__ = ~new_new_n28106__ & ~new_new_n28107__;
  assign new_new_n28109__ = ys__n45878 & new_new_n12245__;
  assign new_new_n28110__ = ys__n45772 & new_new_n12246__;
  assign new_new_n28111__ = ~new_new_n28109__ & ~new_new_n28110__;
  assign new_new_n28112__ = new_new_n28108__ & new_new_n28111__;
  assign new_new_n28113__ = new_new_n26807__ & ~new_new_n28112__;
  assign new_new_n28114__ = ~new_new_n28105__ & ~new_new_n28113__;
  assign new_new_n28115__ = new_new_n26882__ & ~new_new_n28114__;
  assign new_new_n28116__ = ~new_new_n26862__ & new_new_n28115__;
  assign ys__n26132 = new_new_n28097__ | new_new_n28116__;
  assign new_new_n28118__ = ys__n26047 & new_new_n26768__;
  assign new_new_n28119__ = ys__n46374 & new_new_n12356__;
  assign new_new_n28120__ = ys__n46550 & new_new_n12248__;
  assign new_new_n28121__ = ~new_new_n28119__ & ~new_new_n28120__;
  assign new_new_n28122__ = ys__n46726 & new_new_n12245__;
  assign new_new_n28123__ = ys__n46902 & new_new_n12246__;
  assign new_new_n28124__ = ~new_new_n28122__ & ~new_new_n28123__;
  assign new_new_n28125__ = new_new_n28121__ & new_new_n28124__;
  assign new_new_n28126__ = new_new_n26779__ & ~new_new_n28125__;
  assign new_new_n28127__ = ys__n46296 & new_new_n12356__;
  assign new_new_n28128__ = ys__n46472 & new_new_n12248__;
  assign new_new_n28129__ = ~new_new_n28127__ & ~new_new_n28128__;
  assign new_new_n28130__ = ys__n46648 & new_new_n12245__;
  assign new_new_n28131__ = ys__n46824 & new_new_n12246__;
  assign new_new_n28132__ = ~new_new_n28130__ & ~new_new_n28131__;
  assign new_new_n28133__ = new_new_n28129__ & new_new_n28132__;
  assign new_new_n28134__ = new_new_n26788__ & ~new_new_n28133__;
  assign new_new_n28135__ = ~new_new_n28126__ & ~new_new_n28134__;
  assign new_new_n28136__ = ys__n46337 & new_new_n12356__;
  assign new_new_n28137__ = ys__n46513 & new_new_n12248__;
  assign new_new_n28138__ = ~new_new_n28136__ & ~new_new_n28137__;
  assign new_new_n28139__ = ys__n46689 & new_new_n12245__;
  assign new_new_n28140__ = ys__n46865 & new_new_n12246__;
  assign new_new_n28141__ = ~new_new_n28139__ & ~new_new_n28140__;
  assign new_new_n28142__ = new_new_n28138__ & new_new_n28141__;
  assign new_new_n28143__ = new_new_n26798__ & ~new_new_n28142__;
  assign new_new_n28144__ = ys__n46414 & new_new_n12356__;
  assign new_new_n28145__ = ys__n46590 & new_new_n12248__;
  assign new_new_n28146__ = ~new_new_n28144__ & ~new_new_n28145__;
  assign new_new_n28147__ = ys__n46766 & new_new_n12245__;
  assign new_new_n28148__ = ys__n46942 & new_new_n12246__;
  assign new_new_n28149__ = ~new_new_n28147__ & ~new_new_n28148__;
  assign new_new_n28150__ = new_new_n28146__ & new_new_n28149__;
  assign new_new_n28151__ = new_new_n26807__ & ~new_new_n28150__;
  assign new_new_n28152__ = ~new_new_n28143__ & ~new_new_n28151__;
  assign new_new_n28153__ = new_new_n28135__ & new_new_n28152__;
  assign new_new_n28154__ = new_new_n26818__ & ~new_new_n28153__;
  assign new_new_n28155__ = ~new_new_n28118__ & ~new_new_n28154__;
  assign new_new_n28156__ = new_new_n26821__ & ~new_new_n28155__;
  assign new_new_n28157__ = ys__n45584 & new_new_n12356__;
  assign new_new_n28158__ = ys__n45420 & new_new_n12248__;
  assign new_new_n28159__ = ~new_new_n28157__ & ~new_new_n28158__;
  assign new_new_n28160__ = ys__n45256 & new_new_n12245__;
  assign new_new_n28161__ = ys__n45053 & new_new_n12246__;
  assign new_new_n28162__ = ~new_new_n28160__ & ~new_new_n28161__;
  assign new_new_n28163__ = new_new_n28159__ & new_new_n28162__;
  assign new_new_n28164__ = new_new_n26807__ & ~new_new_n28163__;
  assign new_new_n28165__ = ys__n45678 & new_new_n12356__;
  assign new_new_n28166__ = ys__n45514 & new_new_n12248__;
  assign new_new_n28167__ = ~new_new_n28165__ & ~new_new_n28166__;
  assign new_new_n28168__ = ys__n45350 & new_new_n12245__;
  assign new_new_n28169__ = ys__n45179 & new_new_n12246__;
  assign new_new_n28170__ = ~new_new_n28168__ & ~new_new_n28169__;
  assign new_new_n28171__ = new_new_n28167__ & new_new_n28170__;
  assign new_new_n28172__ = new_new_n26779__ & ~new_new_n28171__;
  assign new_new_n28173__ = ys__n45624 & new_new_n12356__;
  assign new_new_n28174__ = ys__n45460 & new_new_n12248__;
  assign new_new_n28175__ = ~new_new_n28173__ & ~new_new_n28174__;
  assign new_new_n28176__ = ys__n45296 & new_new_n12245__;
  assign new_new_n28177__ = ys__n45102 & new_new_n12246__;
  assign new_new_n28178__ = ~new_new_n28176__ & ~new_new_n28177__;
  assign new_new_n28179__ = new_new_n28175__ & new_new_n28178__;
  assign new_new_n28180__ = new_new_n26788__ & ~new_new_n28179__;
  assign new_new_n28181__ = ~new_new_n28172__ & ~new_new_n28180__;
  assign new_new_n28182__ = ~new_new_n28164__ & new_new_n28181__;
  assign new_new_n28183__ = new_new_n26859__ & ~new_new_n28182__;
  assign new_new_n28184__ = ~new_new_n28156__ & ~new_new_n28183__;
  assign new_new_n28185__ = new_new_n26862__ & ~new_new_n28184__;
  assign new_new_n28186__ = ys__n46117 & new_new_n12356__;
  assign new_new_n28187__ = ys__n46019 & new_new_n12248__;
  assign new_new_n28188__ = ~new_new_n28186__ & ~new_new_n28187__;
  assign new_new_n28189__ = ys__n45921 & new_new_n12245__;
  assign new_new_n28190__ = ys__n45825 & new_new_n12246__;
  assign new_new_n28191__ = ~new_new_n28189__ & ~new_new_n28190__;
  assign new_new_n28192__ = new_new_n28188__ & new_new_n28191__;
  assign new_new_n28193__ = new_new_n26788__ & ~new_new_n28192__;
  assign new_new_n28194__ = ys__n46076 & new_new_n12356__;
  assign new_new_n28195__ = ys__n45978 & new_new_n12248__;
  assign new_new_n28196__ = ~new_new_n28194__ & ~new_new_n28195__;
  assign new_new_n28197__ = ys__n45880 & new_new_n12245__;
  assign new_new_n28198__ = ys__n45775 & new_new_n12246__;
  assign new_new_n28199__ = ~new_new_n28197__ & ~new_new_n28198__;
  assign new_new_n28200__ = new_new_n28196__ & new_new_n28199__;
  assign new_new_n28201__ = new_new_n26807__ & ~new_new_n28200__;
  assign new_new_n28202__ = ~new_new_n28193__ & ~new_new_n28201__;
  assign new_new_n28203__ = new_new_n26882__ & ~new_new_n28202__;
  assign new_new_n28204__ = ~new_new_n26862__ & new_new_n28203__;
  assign ys__n26133 = new_new_n28185__ | new_new_n28204__;
  assign new_new_n28206__ = ys__n26050 & new_new_n26768__;
  assign new_new_n28207__ = ys__n46376 & new_new_n12356__;
  assign new_new_n28208__ = ys__n46552 & new_new_n12248__;
  assign new_new_n28209__ = ~new_new_n28207__ & ~new_new_n28208__;
  assign new_new_n28210__ = ys__n46728 & new_new_n12245__;
  assign new_new_n28211__ = ys__n46904 & new_new_n12246__;
  assign new_new_n28212__ = ~new_new_n28210__ & ~new_new_n28211__;
  assign new_new_n28213__ = new_new_n28209__ & new_new_n28212__;
  assign new_new_n28214__ = new_new_n26779__ & ~new_new_n28213__;
  assign new_new_n28215__ = ys__n46298 & new_new_n12356__;
  assign new_new_n28216__ = ys__n46474 & new_new_n12248__;
  assign new_new_n28217__ = ~new_new_n28215__ & ~new_new_n28216__;
  assign new_new_n28218__ = ys__n46650 & new_new_n12245__;
  assign new_new_n28219__ = ys__n46826 & new_new_n12246__;
  assign new_new_n28220__ = ~new_new_n28218__ & ~new_new_n28219__;
  assign new_new_n28221__ = new_new_n28217__ & new_new_n28220__;
  assign new_new_n28222__ = new_new_n26788__ & ~new_new_n28221__;
  assign new_new_n28223__ = ~new_new_n28214__ & ~new_new_n28222__;
  assign new_new_n28224__ = ys__n46338 & new_new_n12356__;
  assign new_new_n28225__ = ys__n46514 & new_new_n12248__;
  assign new_new_n28226__ = ~new_new_n28224__ & ~new_new_n28225__;
  assign new_new_n28227__ = ys__n46690 & new_new_n12245__;
  assign new_new_n28228__ = ys__n46866 & new_new_n12246__;
  assign new_new_n28229__ = ~new_new_n28227__ & ~new_new_n28228__;
  assign new_new_n28230__ = new_new_n28226__ & new_new_n28229__;
  assign new_new_n28231__ = new_new_n26798__ & ~new_new_n28230__;
  assign new_new_n28232__ = ys__n46415 & new_new_n12356__;
  assign new_new_n28233__ = ys__n46591 & new_new_n12248__;
  assign new_new_n28234__ = ~new_new_n28232__ & ~new_new_n28233__;
  assign new_new_n28235__ = ys__n46767 & new_new_n12245__;
  assign new_new_n28236__ = ys__n46943 & new_new_n12246__;
  assign new_new_n28237__ = ~new_new_n28235__ & ~new_new_n28236__;
  assign new_new_n28238__ = new_new_n28234__ & new_new_n28237__;
  assign new_new_n28239__ = new_new_n26807__ & ~new_new_n28238__;
  assign new_new_n28240__ = ~new_new_n28231__ & ~new_new_n28239__;
  assign new_new_n28241__ = new_new_n28223__ & new_new_n28240__;
  assign new_new_n28242__ = new_new_n26818__ & ~new_new_n28241__;
  assign new_new_n28243__ = ~new_new_n28206__ & ~new_new_n28242__;
  assign new_new_n28244__ = new_new_n26821__ & ~new_new_n28243__;
  assign new_new_n28245__ = ys__n45586 & new_new_n12356__;
  assign new_new_n28246__ = ys__n45422 & new_new_n12248__;
  assign new_new_n28247__ = ~new_new_n28245__ & ~new_new_n28246__;
  assign new_new_n28248__ = ys__n45258 & new_new_n12245__;
  assign new_new_n28249__ = ys__n45056 & new_new_n12246__;
  assign new_new_n28250__ = ~new_new_n28248__ & ~new_new_n28249__;
  assign new_new_n28251__ = new_new_n28247__ & new_new_n28250__;
  assign new_new_n28252__ = new_new_n26807__ & ~new_new_n28251__;
  assign new_new_n28253__ = ys__n45680 & new_new_n12356__;
  assign new_new_n28254__ = ys__n45516 & new_new_n12248__;
  assign new_new_n28255__ = ~new_new_n28253__ & ~new_new_n28254__;
  assign new_new_n28256__ = ys__n45352 & new_new_n12245__;
  assign new_new_n28257__ = ys__n45182 & new_new_n12246__;
  assign new_new_n28258__ = ~new_new_n28256__ & ~new_new_n28257__;
  assign new_new_n28259__ = new_new_n28255__ & new_new_n28258__;
  assign new_new_n28260__ = new_new_n26779__ & ~new_new_n28259__;
  assign new_new_n28261__ = ys__n45625 & new_new_n12356__;
  assign new_new_n28262__ = ys__n45461 & new_new_n12248__;
  assign new_new_n28263__ = ~new_new_n28261__ & ~new_new_n28262__;
  assign new_new_n28264__ = ys__n45297 & new_new_n12245__;
  assign new_new_n28265__ = ys__n45103 & new_new_n12246__;
  assign new_new_n28266__ = ~new_new_n28264__ & ~new_new_n28265__;
  assign new_new_n28267__ = new_new_n28263__ & new_new_n28266__;
  assign new_new_n28268__ = new_new_n26788__ & ~new_new_n28267__;
  assign new_new_n28269__ = ~new_new_n28260__ & ~new_new_n28268__;
  assign new_new_n28270__ = ~new_new_n28252__ & new_new_n28269__;
  assign new_new_n28271__ = new_new_n26859__ & ~new_new_n28270__;
  assign new_new_n28272__ = ~new_new_n28244__ & ~new_new_n28271__;
  assign new_new_n28273__ = new_new_n26862__ & ~new_new_n28272__;
  assign new_new_n28274__ = ys__n46118 & new_new_n12356__;
  assign new_new_n28275__ = ys__n46020 & new_new_n12248__;
  assign new_new_n28276__ = ~new_new_n28274__ & ~new_new_n28275__;
  assign new_new_n28277__ = ys__n45922 & new_new_n12245__;
  assign new_new_n28278__ = ys__n45826 & new_new_n12246__;
  assign new_new_n28279__ = ~new_new_n28277__ & ~new_new_n28278__;
  assign new_new_n28280__ = new_new_n28276__ & new_new_n28279__;
  assign new_new_n28281__ = new_new_n26788__ & ~new_new_n28280__;
  assign new_new_n28282__ = ys__n46078 & new_new_n12356__;
  assign new_new_n28283__ = ys__n45980 & new_new_n12248__;
  assign new_new_n28284__ = ~new_new_n28282__ & ~new_new_n28283__;
  assign new_new_n28285__ = ys__n45882 & new_new_n12245__;
  assign new_new_n28286__ = ys__n45778 & new_new_n12246__;
  assign new_new_n28287__ = ~new_new_n28285__ & ~new_new_n28286__;
  assign new_new_n28288__ = new_new_n28284__ & new_new_n28287__;
  assign new_new_n28289__ = new_new_n26807__ & ~new_new_n28288__;
  assign new_new_n28290__ = ~new_new_n28281__ & ~new_new_n28289__;
  assign new_new_n28291__ = new_new_n26882__ & ~new_new_n28290__;
  assign new_new_n28292__ = ~new_new_n26862__ & new_new_n28291__;
  assign ys__n26134 = new_new_n28273__ | new_new_n28292__;
  assign new_new_n28294__ = ys__n26053 & new_new_n26768__;
  assign new_new_n28295__ = ys__n46378 & new_new_n12356__;
  assign new_new_n28296__ = ys__n46554 & new_new_n12248__;
  assign new_new_n28297__ = ~new_new_n28295__ & ~new_new_n28296__;
  assign new_new_n28298__ = ys__n46730 & new_new_n12245__;
  assign new_new_n28299__ = ys__n46906 & new_new_n12246__;
  assign new_new_n28300__ = ~new_new_n28298__ & ~new_new_n28299__;
  assign new_new_n28301__ = new_new_n28297__ & new_new_n28300__;
  assign new_new_n28302__ = new_new_n26779__ & ~new_new_n28301__;
  assign new_new_n28303__ = ys__n46300 & new_new_n12356__;
  assign new_new_n28304__ = ys__n46476 & new_new_n12248__;
  assign new_new_n28305__ = ~new_new_n28303__ & ~new_new_n28304__;
  assign new_new_n28306__ = ys__n46652 & new_new_n12245__;
  assign new_new_n28307__ = ys__n46828 & new_new_n12246__;
  assign new_new_n28308__ = ~new_new_n28306__ & ~new_new_n28307__;
  assign new_new_n28309__ = new_new_n28305__ & new_new_n28308__;
  assign new_new_n28310__ = new_new_n26788__ & ~new_new_n28309__;
  assign new_new_n28311__ = ~new_new_n28302__ & ~new_new_n28310__;
  assign new_new_n28312__ = ys__n46339 & new_new_n12356__;
  assign new_new_n28313__ = ys__n46515 & new_new_n12248__;
  assign new_new_n28314__ = ~new_new_n28312__ & ~new_new_n28313__;
  assign new_new_n28315__ = ys__n46691 & new_new_n12245__;
  assign new_new_n28316__ = ys__n46867 & new_new_n12246__;
  assign new_new_n28317__ = ~new_new_n28315__ & ~new_new_n28316__;
  assign new_new_n28318__ = new_new_n28314__ & new_new_n28317__;
  assign new_new_n28319__ = new_new_n26798__ & ~new_new_n28318__;
  assign new_new_n28320__ = ys__n46416 & new_new_n12356__;
  assign new_new_n28321__ = ys__n46592 & new_new_n12248__;
  assign new_new_n28322__ = ~new_new_n28320__ & ~new_new_n28321__;
  assign new_new_n28323__ = ys__n46768 & new_new_n12245__;
  assign new_new_n28324__ = ys__n46944 & new_new_n12246__;
  assign new_new_n28325__ = ~new_new_n28323__ & ~new_new_n28324__;
  assign new_new_n28326__ = new_new_n28322__ & new_new_n28325__;
  assign new_new_n28327__ = new_new_n26807__ & ~new_new_n28326__;
  assign new_new_n28328__ = ~new_new_n28319__ & ~new_new_n28327__;
  assign new_new_n28329__ = new_new_n28311__ & new_new_n28328__;
  assign new_new_n28330__ = new_new_n26818__ & ~new_new_n28329__;
  assign new_new_n28331__ = ~new_new_n28294__ & ~new_new_n28330__;
  assign new_new_n28332__ = new_new_n26821__ & ~new_new_n28331__;
  assign new_new_n28333__ = ys__n45588 & new_new_n12356__;
  assign new_new_n28334__ = ys__n45424 & new_new_n12248__;
  assign new_new_n28335__ = ~new_new_n28333__ & ~new_new_n28334__;
  assign new_new_n28336__ = ys__n45260 & new_new_n12245__;
  assign new_new_n28337__ = ys__n45059 & new_new_n12246__;
  assign new_new_n28338__ = ~new_new_n28336__ & ~new_new_n28337__;
  assign new_new_n28339__ = new_new_n28335__ & new_new_n28338__;
  assign new_new_n28340__ = new_new_n26807__ & ~new_new_n28339__;
  assign new_new_n28341__ = ys__n45682 & new_new_n12356__;
  assign new_new_n28342__ = ys__n45518 & new_new_n12248__;
  assign new_new_n28343__ = ~new_new_n28341__ & ~new_new_n28342__;
  assign new_new_n28344__ = ys__n45354 & new_new_n12245__;
  assign new_new_n28345__ = ys__n45185 & new_new_n12246__;
  assign new_new_n28346__ = ~new_new_n28344__ & ~new_new_n28345__;
  assign new_new_n28347__ = new_new_n28343__ & new_new_n28346__;
  assign new_new_n28348__ = new_new_n26779__ & ~new_new_n28347__;
  assign new_new_n28349__ = ys__n45626 & new_new_n12356__;
  assign new_new_n28350__ = ys__n45462 & new_new_n12248__;
  assign new_new_n28351__ = ~new_new_n28349__ & ~new_new_n28350__;
  assign new_new_n28352__ = ys__n45298 & new_new_n12245__;
  assign new_new_n28353__ = ys__n45104 & new_new_n12246__;
  assign new_new_n28354__ = ~new_new_n28352__ & ~new_new_n28353__;
  assign new_new_n28355__ = new_new_n28351__ & new_new_n28354__;
  assign new_new_n28356__ = new_new_n26788__ & ~new_new_n28355__;
  assign new_new_n28357__ = ~new_new_n28348__ & ~new_new_n28356__;
  assign new_new_n28358__ = ~new_new_n28340__ & new_new_n28357__;
  assign new_new_n28359__ = new_new_n26859__ & ~new_new_n28358__;
  assign new_new_n28360__ = ~new_new_n28332__ & ~new_new_n28359__;
  assign new_new_n28361__ = new_new_n26862__ & ~new_new_n28360__;
  assign new_new_n28362__ = ys__n46119 & new_new_n12356__;
  assign new_new_n28363__ = ys__n46021 & new_new_n12248__;
  assign new_new_n28364__ = ~new_new_n28362__ & ~new_new_n28363__;
  assign new_new_n28365__ = ys__n45923 & new_new_n12245__;
  assign new_new_n28366__ = ys__n45827 & new_new_n12246__;
  assign new_new_n28367__ = ~new_new_n28365__ & ~new_new_n28366__;
  assign new_new_n28368__ = new_new_n28364__ & new_new_n28367__;
  assign new_new_n28369__ = new_new_n26788__ & ~new_new_n28368__;
  assign new_new_n28370__ = ys__n46080 & new_new_n12356__;
  assign new_new_n28371__ = ys__n45982 & new_new_n12248__;
  assign new_new_n28372__ = ~new_new_n28370__ & ~new_new_n28371__;
  assign new_new_n28373__ = ys__n45884 & new_new_n12245__;
  assign new_new_n28374__ = ys__n45781 & new_new_n12246__;
  assign new_new_n28375__ = ~new_new_n28373__ & ~new_new_n28374__;
  assign new_new_n28376__ = new_new_n28372__ & new_new_n28375__;
  assign new_new_n28377__ = new_new_n26807__ & ~new_new_n28376__;
  assign new_new_n28378__ = ~new_new_n28369__ & ~new_new_n28377__;
  assign new_new_n28379__ = new_new_n26882__ & ~new_new_n28378__;
  assign new_new_n28380__ = ~new_new_n26862__ & new_new_n28379__;
  assign ys__n26135 = new_new_n28361__ | new_new_n28380__;
  assign new_new_n28382__ = ys__n26056 & new_new_n26768__;
  assign new_new_n28383__ = ys__n46380 & new_new_n12356__;
  assign new_new_n28384__ = ys__n46556 & new_new_n12248__;
  assign new_new_n28385__ = ~new_new_n28383__ & ~new_new_n28384__;
  assign new_new_n28386__ = ys__n46732 & new_new_n12245__;
  assign new_new_n28387__ = ys__n46908 & new_new_n12246__;
  assign new_new_n28388__ = ~new_new_n28386__ & ~new_new_n28387__;
  assign new_new_n28389__ = new_new_n28385__ & new_new_n28388__;
  assign new_new_n28390__ = new_new_n26779__ & ~new_new_n28389__;
  assign new_new_n28391__ = ys__n46302 & new_new_n12356__;
  assign new_new_n28392__ = ys__n46478 & new_new_n12248__;
  assign new_new_n28393__ = ~new_new_n28391__ & ~new_new_n28392__;
  assign new_new_n28394__ = ys__n46654 & new_new_n12245__;
  assign new_new_n28395__ = ys__n46830 & new_new_n12246__;
  assign new_new_n28396__ = ~new_new_n28394__ & ~new_new_n28395__;
  assign new_new_n28397__ = new_new_n28393__ & new_new_n28396__;
  assign new_new_n28398__ = new_new_n26788__ & ~new_new_n28397__;
  assign new_new_n28399__ = ~new_new_n28390__ & ~new_new_n28398__;
  assign new_new_n28400__ = ys__n46340 & new_new_n12356__;
  assign new_new_n28401__ = ys__n46516 & new_new_n12248__;
  assign new_new_n28402__ = ~new_new_n28400__ & ~new_new_n28401__;
  assign new_new_n28403__ = ys__n46692 & new_new_n12245__;
  assign new_new_n28404__ = ys__n46868 & new_new_n12246__;
  assign new_new_n28405__ = ~new_new_n28403__ & ~new_new_n28404__;
  assign new_new_n28406__ = new_new_n28402__ & new_new_n28405__;
  assign new_new_n28407__ = new_new_n26798__ & ~new_new_n28406__;
  assign new_new_n28408__ = ys__n46417 & new_new_n12356__;
  assign new_new_n28409__ = ys__n46593 & new_new_n12248__;
  assign new_new_n28410__ = ~new_new_n28408__ & ~new_new_n28409__;
  assign new_new_n28411__ = ys__n46769 & new_new_n12245__;
  assign new_new_n28412__ = ys__n46945 & new_new_n12246__;
  assign new_new_n28413__ = ~new_new_n28411__ & ~new_new_n28412__;
  assign new_new_n28414__ = new_new_n28410__ & new_new_n28413__;
  assign new_new_n28415__ = new_new_n26807__ & ~new_new_n28414__;
  assign new_new_n28416__ = ~new_new_n28407__ & ~new_new_n28415__;
  assign new_new_n28417__ = new_new_n28399__ & new_new_n28416__;
  assign new_new_n28418__ = new_new_n26818__ & ~new_new_n28417__;
  assign new_new_n28419__ = ~new_new_n28382__ & ~new_new_n28418__;
  assign new_new_n28420__ = new_new_n26821__ & ~new_new_n28419__;
  assign new_new_n28421__ = ys__n45590 & new_new_n12356__;
  assign new_new_n28422__ = ys__n45426 & new_new_n12248__;
  assign new_new_n28423__ = ~new_new_n28421__ & ~new_new_n28422__;
  assign new_new_n28424__ = ys__n45262 & new_new_n12245__;
  assign new_new_n28425__ = ys__n45062 & new_new_n12246__;
  assign new_new_n28426__ = ~new_new_n28424__ & ~new_new_n28425__;
  assign new_new_n28427__ = new_new_n28423__ & new_new_n28426__;
  assign new_new_n28428__ = new_new_n26807__ & ~new_new_n28427__;
  assign new_new_n28429__ = ys__n45684 & new_new_n12356__;
  assign new_new_n28430__ = ys__n45520 & new_new_n12248__;
  assign new_new_n28431__ = ~new_new_n28429__ & ~new_new_n28430__;
  assign new_new_n28432__ = ys__n45356 & new_new_n12245__;
  assign new_new_n28433__ = ys__n45188 & new_new_n12246__;
  assign new_new_n28434__ = ~new_new_n28432__ & ~new_new_n28433__;
  assign new_new_n28435__ = new_new_n28431__ & new_new_n28434__;
  assign new_new_n28436__ = new_new_n26779__ & ~new_new_n28435__;
  assign new_new_n28437__ = ys__n45627 & new_new_n12356__;
  assign new_new_n28438__ = ys__n45463 & new_new_n12248__;
  assign new_new_n28439__ = ~new_new_n28437__ & ~new_new_n28438__;
  assign new_new_n28440__ = ys__n45299 & new_new_n12245__;
  assign new_new_n28441__ = ys__n45105 & new_new_n12246__;
  assign new_new_n28442__ = ~new_new_n28440__ & ~new_new_n28441__;
  assign new_new_n28443__ = new_new_n28439__ & new_new_n28442__;
  assign new_new_n28444__ = new_new_n26788__ & ~new_new_n28443__;
  assign new_new_n28445__ = ~new_new_n28436__ & ~new_new_n28444__;
  assign new_new_n28446__ = ~new_new_n28428__ & new_new_n28445__;
  assign new_new_n28447__ = new_new_n26859__ & ~new_new_n28446__;
  assign new_new_n28448__ = ~new_new_n28420__ & ~new_new_n28447__;
  assign new_new_n28449__ = new_new_n26862__ & ~new_new_n28448__;
  assign new_new_n28450__ = ys__n46120 & new_new_n12356__;
  assign new_new_n28451__ = ys__n46022 & new_new_n12248__;
  assign new_new_n28452__ = ~new_new_n28450__ & ~new_new_n28451__;
  assign new_new_n28453__ = ys__n45924 & new_new_n12245__;
  assign new_new_n28454__ = ys__n45828 & new_new_n12246__;
  assign new_new_n28455__ = ~new_new_n28453__ & ~new_new_n28454__;
  assign new_new_n28456__ = new_new_n28452__ & new_new_n28455__;
  assign new_new_n28457__ = new_new_n26788__ & ~new_new_n28456__;
  assign new_new_n28458__ = ys__n46082 & new_new_n12356__;
  assign new_new_n28459__ = ys__n45984 & new_new_n12248__;
  assign new_new_n28460__ = ~new_new_n28458__ & ~new_new_n28459__;
  assign new_new_n28461__ = ys__n45886 & new_new_n12245__;
  assign new_new_n28462__ = ys__n45784 & new_new_n12246__;
  assign new_new_n28463__ = ~new_new_n28461__ & ~new_new_n28462__;
  assign new_new_n28464__ = new_new_n28460__ & new_new_n28463__;
  assign new_new_n28465__ = new_new_n26807__ & ~new_new_n28464__;
  assign new_new_n28466__ = ~new_new_n28457__ & ~new_new_n28465__;
  assign new_new_n28467__ = new_new_n26882__ & ~new_new_n28466__;
  assign new_new_n28468__ = ~new_new_n26862__ & new_new_n28467__;
  assign ys__n26136 = new_new_n28449__ | new_new_n28468__;
  assign new_new_n28470__ = ys__n26059 & new_new_n26768__;
  assign new_new_n28471__ = ys__n46382 & new_new_n12356__;
  assign new_new_n28472__ = ys__n46558 & new_new_n12248__;
  assign new_new_n28473__ = ~new_new_n28471__ & ~new_new_n28472__;
  assign new_new_n28474__ = ys__n46734 & new_new_n12245__;
  assign new_new_n28475__ = ys__n46910 & new_new_n12246__;
  assign new_new_n28476__ = ~new_new_n28474__ & ~new_new_n28475__;
  assign new_new_n28477__ = new_new_n28473__ & new_new_n28476__;
  assign new_new_n28478__ = new_new_n26779__ & ~new_new_n28477__;
  assign new_new_n28479__ = ys__n46304 & new_new_n12356__;
  assign new_new_n28480__ = ys__n46480 & new_new_n12248__;
  assign new_new_n28481__ = ~new_new_n28479__ & ~new_new_n28480__;
  assign new_new_n28482__ = ys__n46656 & new_new_n12245__;
  assign new_new_n28483__ = ys__n46832 & new_new_n12246__;
  assign new_new_n28484__ = ~new_new_n28482__ & ~new_new_n28483__;
  assign new_new_n28485__ = new_new_n28481__ & new_new_n28484__;
  assign new_new_n28486__ = new_new_n26788__ & ~new_new_n28485__;
  assign new_new_n28487__ = ~new_new_n28478__ & ~new_new_n28486__;
  assign new_new_n28488__ = ys__n46341 & new_new_n12356__;
  assign new_new_n28489__ = ys__n46517 & new_new_n12248__;
  assign new_new_n28490__ = ~new_new_n28488__ & ~new_new_n28489__;
  assign new_new_n28491__ = ys__n46693 & new_new_n12245__;
  assign new_new_n28492__ = ys__n46869 & new_new_n12246__;
  assign new_new_n28493__ = ~new_new_n28491__ & ~new_new_n28492__;
  assign new_new_n28494__ = new_new_n28490__ & new_new_n28493__;
  assign new_new_n28495__ = new_new_n26798__ & ~new_new_n28494__;
  assign new_new_n28496__ = ys__n46418 & new_new_n12356__;
  assign new_new_n28497__ = ys__n46594 & new_new_n12248__;
  assign new_new_n28498__ = ~new_new_n28496__ & ~new_new_n28497__;
  assign new_new_n28499__ = ys__n46770 & new_new_n12245__;
  assign new_new_n28500__ = ys__n46946 & new_new_n12246__;
  assign new_new_n28501__ = ~new_new_n28499__ & ~new_new_n28500__;
  assign new_new_n28502__ = new_new_n28498__ & new_new_n28501__;
  assign new_new_n28503__ = new_new_n26807__ & ~new_new_n28502__;
  assign new_new_n28504__ = ~new_new_n28495__ & ~new_new_n28503__;
  assign new_new_n28505__ = new_new_n28487__ & new_new_n28504__;
  assign new_new_n28506__ = new_new_n26817__ & ~new_new_n28505__;
  assign new_new_n28507__ = new_new_n12365__ & ~new_new_n28506__;
  assign new_new_n28508__ = ~new_new_n26768__ & ~new_new_n28507__;
  assign new_new_n28509__ = ~new_new_n28470__ & ~new_new_n28508__;
  assign new_new_n28510__ = new_new_n26821__ & ~new_new_n28509__;
  assign new_new_n28511__ = ys__n45592 & new_new_n12356__;
  assign new_new_n28512__ = ys__n45428 & new_new_n12248__;
  assign new_new_n28513__ = ~new_new_n28511__ & ~new_new_n28512__;
  assign new_new_n28514__ = ys__n45264 & new_new_n12245__;
  assign new_new_n28515__ = ys__n45065 & new_new_n12246__;
  assign new_new_n28516__ = ~new_new_n28514__ & ~new_new_n28515__;
  assign new_new_n28517__ = new_new_n28513__ & new_new_n28516__;
  assign new_new_n28518__ = new_new_n26807__ & ~new_new_n28517__;
  assign new_new_n28519__ = ys__n45686 & new_new_n12356__;
  assign new_new_n28520__ = ys__n45522 & new_new_n12248__;
  assign new_new_n28521__ = ~new_new_n28519__ & ~new_new_n28520__;
  assign new_new_n28522__ = ys__n45358 & new_new_n12245__;
  assign new_new_n28523__ = ys__n45191 & new_new_n12246__;
  assign new_new_n28524__ = ~new_new_n28522__ & ~new_new_n28523__;
  assign new_new_n28525__ = new_new_n28521__ & new_new_n28524__;
  assign new_new_n28526__ = new_new_n26779__ & ~new_new_n28525__;
  assign new_new_n28527__ = ys__n45628 & new_new_n12356__;
  assign new_new_n28528__ = ys__n45464 & new_new_n12248__;
  assign new_new_n28529__ = ~new_new_n28527__ & ~new_new_n28528__;
  assign new_new_n28530__ = ys__n45300 & new_new_n12245__;
  assign new_new_n28531__ = ys__n45106 & new_new_n12246__;
  assign new_new_n28532__ = ~new_new_n28530__ & ~new_new_n28531__;
  assign new_new_n28533__ = new_new_n28529__ & new_new_n28532__;
  assign new_new_n28534__ = new_new_n26788__ & ~new_new_n28533__;
  assign new_new_n28535__ = ~new_new_n28526__ & ~new_new_n28534__;
  assign new_new_n28536__ = ~new_new_n28518__ & new_new_n28535__;
  assign new_new_n28537__ = new_new_n26858__ & ~new_new_n28536__;
  assign new_new_n28538__ = new_new_n12286__ & ~new_new_n28537__;
  assign new_new_n28539__ = ~new_new_n26821__ & ~new_new_n28538__;
  assign new_new_n28540__ = ~new_new_n28510__ & ~new_new_n28539__;
  assign new_new_n28541__ = new_new_n26862__ & ~new_new_n28540__;
  assign new_new_n28542__ = ys__n46121 & new_new_n12356__;
  assign new_new_n28543__ = ys__n46023 & new_new_n12248__;
  assign new_new_n28544__ = ~new_new_n28542__ & ~new_new_n28543__;
  assign new_new_n28545__ = ys__n45925 & new_new_n12245__;
  assign new_new_n28546__ = ys__n45829 & new_new_n12246__;
  assign new_new_n28547__ = ~new_new_n28545__ & ~new_new_n28546__;
  assign new_new_n28548__ = new_new_n28544__ & new_new_n28547__;
  assign new_new_n28549__ = new_new_n26788__ & ~new_new_n28548__;
  assign new_new_n28550__ = ys__n46084 & new_new_n12356__;
  assign new_new_n28551__ = ys__n45986 & new_new_n12248__;
  assign new_new_n28552__ = ~new_new_n28550__ & ~new_new_n28551__;
  assign new_new_n28553__ = ys__n45888 & new_new_n12245__;
  assign new_new_n28554__ = ys__n45787 & new_new_n12246__;
  assign new_new_n28555__ = ~new_new_n28553__ & ~new_new_n28554__;
  assign new_new_n28556__ = new_new_n28552__ & new_new_n28555__;
  assign new_new_n28557__ = new_new_n26807__ & ~new_new_n28556__;
  assign new_new_n28558__ = ~new_new_n28549__ & ~new_new_n28557__;
  assign new_new_n28559__ = new_new_n26882__ & ~new_new_n28558__;
  assign new_new_n28560__ = new_new_n12395__ & ~new_new_n28559__;
  assign new_new_n28561__ = ~new_new_n26862__ & ~new_new_n28560__;
  assign ys__n26137 = new_new_n28541__ | new_new_n28561__;
  assign new_new_n28563__ = ys__n26062 & new_new_n26768__;
  assign new_new_n28564__ = ys__n46384 & new_new_n12356__;
  assign new_new_n28565__ = ys__n46560 & new_new_n12248__;
  assign new_new_n28566__ = ~new_new_n28564__ & ~new_new_n28565__;
  assign new_new_n28567__ = ys__n46736 & new_new_n12245__;
  assign new_new_n28568__ = ys__n46912 & new_new_n12246__;
  assign new_new_n28569__ = ~new_new_n28567__ & ~new_new_n28568__;
  assign new_new_n28570__ = new_new_n28566__ & new_new_n28569__;
  assign new_new_n28571__ = new_new_n26779__ & ~new_new_n28570__;
  assign new_new_n28572__ = ys__n46306 & new_new_n12356__;
  assign new_new_n28573__ = ys__n46482 & new_new_n12248__;
  assign new_new_n28574__ = ~new_new_n28572__ & ~new_new_n28573__;
  assign new_new_n28575__ = ys__n46658 & new_new_n12245__;
  assign new_new_n28576__ = ys__n46834 & new_new_n12246__;
  assign new_new_n28577__ = ~new_new_n28575__ & ~new_new_n28576__;
  assign new_new_n28578__ = new_new_n28574__ & new_new_n28577__;
  assign new_new_n28579__ = new_new_n26788__ & ~new_new_n28578__;
  assign new_new_n28580__ = ~new_new_n28571__ & ~new_new_n28579__;
  assign new_new_n28581__ = ys__n46342 & new_new_n12356__;
  assign new_new_n28582__ = ys__n46518 & new_new_n12248__;
  assign new_new_n28583__ = ~new_new_n28581__ & ~new_new_n28582__;
  assign new_new_n28584__ = ys__n46694 & new_new_n12245__;
  assign new_new_n28585__ = ys__n46870 & new_new_n12246__;
  assign new_new_n28586__ = ~new_new_n28584__ & ~new_new_n28585__;
  assign new_new_n28587__ = new_new_n28583__ & new_new_n28586__;
  assign new_new_n28588__ = new_new_n26798__ & ~new_new_n28587__;
  assign new_new_n28589__ = ys__n46419 & new_new_n12356__;
  assign new_new_n28590__ = ys__n46595 & new_new_n12248__;
  assign new_new_n28591__ = ~new_new_n28589__ & ~new_new_n28590__;
  assign new_new_n28592__ = ys__n46771 & new_new_n12245__;
  assign new_new_n28593__ = ys__n46947 & new_new_n12246__;
  assign new_new_n28594__ = ~new_new_n28592__ & ~new_new_n28593__;
  assign new_new_n28595__ = new_new_n28591__ & new_new_n28594__;
  assign new_new_n28596__ = new_new_n26807__ & ~new_new_n28595__;
  assign new_new_n28597__ = ~new_new_n28588__ & ~new_new_n28596__;
  assign new_new_n28598__ = new_new_n28580__ & new_new_n28597__;
  assign new_new_n28599__ = new_new_n26818__ & ~new_new_n28598__;
  assign new_new_n28600__ = ~new_new_n28563__ & ~new_new_n28599__;
  assign new_new_n28601__ = new_new_n26821__ & ~new_new_n28600__;
  assign new_new_n28602__ = ys__n45594 & new_new_n12356__;
  assign new_new_n28603__ = ys__n45430 & new_new_n12248__;
  assign new_new_n28604__ = ~new_new_n28602__ & ~new_new_n28603__;
  assign new_new_n28605__ = ys__n45266 & new_new_n12245__;
  assign new_new_n28606__ = ys__n45068 & new_new_n12246__;
  assign new_new_n28607__ = ~new_new_n28605__ & ~new_new_n28606__;
  assign new_new_n28608__ = new_new_n28604__ & new_new_n28607__;
  assign new_new_n28609__ = new_new_n26807__ & ~new_new_n28608__;
  assign new_new_n28610__ = ys__n45688 & new_new_n12356__;
  assign new_new_n28611__ = ys__n45524 & new_new_n12248__;
  assign new_new_n28612__ = ~new_new_n28610__ & ~new_new_n28611__;
  assign new_new_n28613__ = ys__n45360 & new_new_n12245__;
  assign new_new_n28614__ = ys__n45194 & new_new_n12246__;
  assign new_new_n28615__ = ~new_new_n28613__ & ~new_new_n28614__;
  assign new_new_n28616__ = new_new_n28612__ & new_new_n28615__;
  assign new_new_n28617__ = new_new_n26779__ & ~new_new_n28616__;
  assign new_new_n28618__ = ys__n45629 & new_new_n12356__;
  assign new_new_n28619__ = ys__n45465 & new_new_n12248__;
  assign new_new_n28620__ = ~new_new_n28618__ & ~new_new_n28619__;
  assign new_new_n28621__ = ys__n45301 & new_new_n12245__;
  assign new_new_n28622__ = ys__n45107 & new_new_n12246__;
  assign new_new_n28623__ = ~new_new_n28621__ & ~new_new_n28622__;
  assign new_new_n28624__ = new_new_n28620__ & new_new_n28623__;
  assign new_new_n28625__ = new_new_n26788__ & ~new_new_n28624__;
  assign new_new_n28626__ = ~new_new_n28617__ & ~new_new_n28625__;
  assign new_new_n28627__ = ~new_new_n28609__ & new_new_n28626__;
  assign new_new_n28628__ = new_new_n26859__ & ~new_new_n28627__;
  assign new_new_n28629__ = ~new_new_n28601__ & ~new_new_n28628__;
  assign new_new_n28630__ = new_new_n26862__ & ~new_new_n28629__;
  assign new_new_n28631__ = ys__n46122 & new_new_n12356__;
  assign new_new_n28632__ = ys__n46024 & new_new_n12248__;
  assign new_new_n28633__ = ~new_new_n28631__ & ~new_new_n28632__;
  assign new_new_n28634__ = ys__n45926 & new_new_n12245__;
  assign new_new_n28635__ = ys__n45830 & new_new_n12246__;
  assign new_new_n28636__ = ~new_new_n28634__ & ~new_new_n28635__;
  assign new_new_n28637__ = new_new_n28633__ & new_new_n28636__;
  assign new_new_n28638__ = new_new_n26788__ & ~new_new_n28637__;
  assign new_new_n28639__ = ys__n46086 & new_new_n12356__;
  assign new_new_n28640__ = ys__n45988 & new_new_n12248__;
  assign new_new_n28641__ = ~new_new_n28639__ & ~new_new_n28640__;
  assign new_new_n28642__ = ys__n45890 & new_new_n12245__;
  assign new_new_n28643__ = ys__n45790 & new_new_n12246__;
  assign new_new_n28644__ = ~new_new_n28642__ & ~new_new_n28643__;
  assign new_new_n28645__ = new_new_n28641__ & new_new_n28644__;
  assign new_new_n28646__ = new_new_n26807__ & ~new_new_n28645__;
  assign new_new_n28647__ = ~new_new_n28638__ & ~new_new_n28646__;
  assign new_new_n28648__ = new_new_n26882__ & ~new_new_n28647__;
  assign new_new_n28649__ = ~new_new_n26862__ & new_new_n28648__;
  assign ys__n26138 = new_new_n28630__ | new_new_n28649__;
  assign new_new_n28651__ = ys__n26065 & new_new_n26768__;
  assign new_new_n28652__ = ys__n46386 & new_new_n12356__;
  assign new_new_n28653__ = ys__n46562 & new_new_n12248__;
  assign new_new_n28654__ = ~new_new_n28652__ & ~new_new_n28653__;
  assign new_new_n28655__ = ys__n46738 & new_new_n12245__;
  assign new_new_n28656__ = ys__n46914 & new_new_n12246__;
  assign new_new_n28657__ = ~new_new_n28655__ & ~new_new_n28656__;
  assign new_new_n28658__ = new_new_n28654__ & new_new_n28657__;
  assign new_new_n28659__ = new_new_n26779__ & ~new_new_n28658__;
  assign new_new_n28660__ = ys__n46308 & new_new_n12356__;
  assign new_new_n28661__ = ys__n46484 & new_new_n12248__;
  assign new_new_n28662__ = ~new_new_n28660__ & ~new_new_n28661__;
  assign new_new_n28663__ = ys__n46660 & new_new_n12245__;
  assign new_new_n28664__ = ys__n46836 & new_new_n12246__;
  assign new_new_n28665__ = ~new_new_n28663__ & ~new_new_n28664__;
  assign new_new_n28666__ = new_new_n28662__ & new_new_n28665__;
  assign new_new_n28667__ = new_new_n26788__ & ~new_new_n28666__;
  assign new_new_n28668__ = ~new_new_n28659__ & ~new_new_n28667__;
  assign new_new_n28669__ = ys__n46343 & new_new_n12356__;
  assign new_new_n28670__ = ys__n46519 & new_new_n12248__;
  assign new_new_n28671__ = ~new_new_n28669__ & ~new_new_n28670__;
  assign new_new_n28672__ = ys__n46695 & new_new_n12245__;
  assign new_new_n28673__ = ys__n46871 & new_new_n12246__;
  assign new_new_n28674__ = ~new_new_n28672__ & ~new_new_n28673__;
  assign new_new_n28675__ = new_new_n28671__ & new_new_n28674__;
  assign new_new_n28676__ = new_new_n26798__ & ~new_new_n28675__;
  assign new_new_n28677__ = ys__n46420 & new_new_n12356__;
  assign new_new_n28678__ = ys__n46596 & new_new_n12248__;
  assign new_new_n28679__ = ~new_new_n28677__ & ~new_new_n28678__;
  assign new_new_n28680__ = ys__n46772 & new_new_n12245__;
  assign new_new_n28681__ = ys__n46948 & new_new_n12246__;
  assign new_new_n28682__ = ~new_new_n28680__ & ~new_new_n28681__;
  assign new_new_n28683__ = new_new_n28679__ & new_new_n28682__;
  assign new_new_n28684__ = new_new_n26807__ & ~new_new_n28683__;
  assign new_new_n28685__ = ~new_new_n28676__ & ~new_new_n28684__;
  assign new_new_n28686__ = new_new_n28668__ & new_new_n28685__;
  assign new_new_n28687__ = new_new_n26818__ & ~new_new_n28686__;
  assign new_new_n28688__ = ~new_new_n28651__ & ~new_new_n28687__;
  assign new_new_n28689__ = new_new_n26821__ & ~new_new_n28688__;
  assign new_new_n28690__ = ys__n45596 & new_new_n12356__;
  assign new_new_n28691__ = ys__n45432 & new_new_n12248__;
  assign new_new_n28692__ = ~new_new_n28690__ & ~new_new_n28691__;
  assign new_new_n28693__ = ys__n45268 & new_new_n12245__;
  assign new_new_n28694__ = ys__n45071 & new_new_n12246__;
  assign new_new_n28695__ = ~new_new_n28693__ & ~new_new_n28694__;
  assign new_new_n28696__ = new_new_n28692__ & new_new_n28695__;
  assign new_new_n28697__ = new_new_n26807__ & ~new_new_n28696__;
  assign new_new_n28698__ = ys__n45690 & new_new_n12356__;
  assign new_new_n28699__ = ys__n45526 & new_new_n12248__;
  assign new_new_n28700__ = ~new_new_n28698__ & ~new_new_n28699__;
  assign new_new_n28701__ = ys__n45362 & new_new_n12245__;
  assign new_new_n28702__ = ys__n45197 & new_new_n12246__;
  assign new_new_n28703__ = ~new_new_n28701__ & ~new_new_n28702__;
  assign new_new_n28704__ = new_new_n28700__ & new_new_n28703__;
  assign new_new_n28705__ = new_new_n26779__ & ~new_new_n28704__;
  assign new_new_n28706__ = ys__n45630 & new_new_n12356__;
  assign new_new_n28707__ = ys__n45466 & new_new_n12248__;
  assign new_new_n28708__ = ~new_new_n28706__ & ~new_new_n28707__;
  assign new_new_n28709__ = ys__n45302 & new_new_n12245__;
  assign new_new_n28710__ = ys__n45108 & new_new_n12246__;
  assign new_new_n28711__ = ~new_new_n28709__ & ~new_new_n28710__;
  assign new_new_n28712__ = new_new_n28708__ & new_new_n28711__;
  assign new_new_n28713__ = new_new_n26788__ & ~new_new_n28712__;
  assign new_new_n28714__ = ~new_new_n28705__ & ~new_new_n28713__;
  assign new_new_n28715__ = ~new_new_n28697__ & new_new_n28714__;
  assign new_new_n28716__ = new_new_n26859__ & ~new_new_n28715__;
  assign new_new_n28717__ = ~new_new_n28689__ & ~new_new_n28716__;
  assign new_new_n28718__ = new_new_n26862__ & ~new_new_n28717__;
  assign new_new_n28719__ = ys__n46123 & new_new_n12356__;
  assign new_new_n28720__ = ys__n46025 & new_new_n12248__;
  assign new_new_n28721__ = ~new_new_n28719__ & ~new_new_n28720__;
  assign new_new_n28722__ = ys__n45927 & new_new_n12245__;
  assign new_new_n28723__ = ys__n45831 & new_new_n12246__;
  assign new_new_n28724__ = ~new_new_n28722__ & ~new_new_n28723__;
  assign new_new_n28725__ = new_new_n28721__ & new_new_n28724__;
  assign new_new_n28726__ = new_new_n26788__ & ~new_new_n28725__;
  assign new_new_n28727__ = ys__n46088 & new_new_n12356__;
  assign new_new_n28728__ = ys__n45990 & new_new_n12248__;
  assign new_new_n28729__ = ~new_new_n28727__ & ~new_new_n28728__;
  assign new_new_n28730__ = ys__n45892 & new_new_n12245__;
  assign new_new_n28731__ = ys__n45793 & new_new_n12246__;
  assign new_new_n28732__ = ~new_new_n28730__ & ~new_new_n28731__;
  assign new_new_n28733__ = new_new_n28729__ & new_new_n28732__;
  assign new_new_n28734__ = new_new_n26807__ & ~new_new_n28733__;
  assign new_new_n28735__ = ~new_new_n28726__ & ~new_new_n28734__;
  assign new_new_n28736__ = new_new_n26882__ & ~new_new_n28735__;
  assign new_new_n28737__ = ~new_new_n26862__ & new_new_n28736__;
  assign ys__n26139 = new_new_n28718__ | new_new_n28737__;
  assign new_new_n28739__ = ys__n26071 & new_new_n26768__;
  assign new_new_n28740__ = ys__n46390 & new_new_n12356__;
  assign new_new_n28741__ = ys__n46566 & new_new_n12248__;
  assign new_new_n28742__ = ~new_new_n28740__ & ~new_new_n28741__;
  assign new_new_n28743__ = ys__n46742 & new_new_n12245__;
  assign new_new_n28744__ = ys__n46918 & new_new_n12246__;
  assign new_new_n28745__ = ~new_new_n28743__ & ~new_new_n28744__;
  assign new_new_n28746__ = new_new_n28742__ & new_new_n28745__;
  assign new_new_n28747__ = new_new_n26779__ & ~new_new_n28746__;
  assign new_new_n28748__ = ys__n46312 & new_new_n12356__;
  assign new_new_n28749__ = ys__n46488 & new_new_n12248__;
  assign new_new_n28750__ = ~new_new_n28748__ & ~new_new_n28749__;
  assign new_new_n28751__ = ys__n46664 & new_new_n12245__;
  assign new_new_n28752__ = ys__n46840 & new_new_n12246__;
  assign new_new_n28753__ = ~new_new_n28751__ & ~new_new_n28752__;
  assign new_new_n28754__ = new_new_n28750__ & new_new_n28753__;
  assign new_new_n28755__ = new_new_n26788__ & ~new_new_n28754__;
  assign new_new_n28756__ = ~new_new_n28747__ & ~new_new_n28755__;
  assign new_new_n28757__ = ys__n46345 & new_new_n12356__;
  assign new_new_n28758__ = ys__n46521 & new_new_n12248__;
  assign new_new_n28759__ = ~new_new_n28757__ & ~new_new_n28758__;
  assign new_new_n28760__ = ys__n46697 & new_new_n12245__;
  assign new_new_n28761__ = ys__n46873 & new_new_n12246__;
  assign new_new_n28762__ = ~new_new_n28760__ & ~new_new_n28761__;
  assign new_new_n28763__ = new_new_n28759__ & new_new_n28762__;
  assign new_new_n28764__ = new_new_n26798__ & ~new_new_n28763__;
  assign new_new_n28765__ = ys__n46422 & new_new_n12356__;
  assign new_new_n28766__ = ys__n46598 & new_new_n12248__;
  assign new_new_n28767__ = ~new_new_n28765__ & ~new_new_n28766__;
  assign new_new_n28768__ = ys__n46774 & new_new_n12245__;
  assign new_new_n28769__ = ys__n46950 & new_new_n12246__;
  assign new_new_n28770__ = ~new_new_n28768__ & ~new_new_n28769__;
  assign new_new_n28771__ = new_new_n28767__ & new_new_n28770__;
  assign new_new_n28772__ = new_new_n26807__ & ~new_new_n28771__;
  assign new_new_n28773__ = ~new_new_n28764__ & ~new_new_n28772__;
  assign new_new_n28774__ = new_new_n28756__ & new_new_n28773__;
  assign new_new_n28775__ = new_new_n26818__ & ~new_new_n28774__;
  assign new_new_n28776__ = ~new_new_n28739__ & ~new_new_n28775__;
  assign new_new_n28777__ = new_new_n26821__ & ~new_new_n28776__;
  assign new_new_n28778__ = ys__n45600 & new_new_n12356__;
  assign new_new_n28779__ = ys__n45436 & new_new_n12248__;
  assign new_new_n28780__ = ~new_new_n28778__ & ~new_new_n28779__;
  assign new_new_n28781__ = ys__n45272 & new_new_n12245__;
  assign new_new_n28782__ = ys__n45077 & new_new_n12246__;
  assign new_new_n28783__ = ~new_new_n28781__ & ~new_new_n28782__;
  assign new_new_n28784__ = new_new_n28780__ & new_new_n28783__;
  assign new_new_n28785__ = new_new_n26807__ & ~new_new_n28784__;
  assign new_new_n28786__ = ys__n45694 & new_new_n12356__;
  assign new_new_n28787__ = ys__n45530 & new_new_n12248__;
  assign new_new_n28788__ = ~new_new_n28786__ & ~new_new_n28787__;
  assign new_new_n28789__ = ys__n45366 & new_new_n12245__;
  assign new_new_n28790__ = ys__n45203 & new_new_n12246__;
  assign new_new_n28791__ = ~new_new_n28789__ & ~new_new_n28790__;
  assign new_new_n28792__ = new_new_n28788__ & new_new_n28791__;
  assign new_new_n28793__ = new_new_n26779__ & ~new_new_n28792__;
  assign new_new_n28794__ = ys__n45632 & new_new_n12356__;
  assign new_new_n28795__ = ys__n45468 & new_new_n12248__;
  assign new_new_n28796__ = ~new_new_n28794__ & ~new_new_n28795__;
  assign new_new_n28797__ = ys__n45304 & new_new_n12245__;
  assign new_new_n28798__ = ys__n45110 & new_new_n12246__;
  assign new_new_n28799__ = ~new_new_n28797__ & ~new_new_n28798__;
  assign new_new_n28800__ = new_new_n28796__ & new_new_n28799__;
  assign new_new_n28801__ = new_new_n26788__ & ~new_new_n28800__;
  assign new_new_n28802__ = ~new_new_n28793__ & ~new_new_n28801__;
  assign new_new_n28803__ = ~new_new_n28785__ & new_new_n28802__;
  assign new_new_n28804__ = new_new_n26859__ & ~new_new_n28803__;
  assign new_new_n28805__ = ~new_new_n28777__ & ~new_new_n28804__;
  assign new_new_n28806__ = new_new_n26862__ & ~new_new_n28805__;
  assign new_new_n28807__ = ys__n46125 & new_new_n12356__;
  assign new_new_n28808__ = ys__n46027 & new_new_n12248__;
  assign new_new_n28809__ = ~new_new_n28807__ & ~new_new_n28808__;
  assign new_new_n28810__ = ys__n45929 & new_new_n12245__;
  assign new_new_n28811__ = ys__n45833 & new_new_n12246__;
  assign new_new_n28812__ = ~new_new_n28810__ & ~new_new_n28811__;
  assign new_new_n28813__ = new_new_n28809__ & new_new_n28812__;
  assign new_new_n28814__ = new_new_n26788__ & ~new_new_n28813__;
  assign new_new_n28815__ = ys__n46092 & new_new_n12356__;
  assign new_new_n28816__ = ys__n45994 & new_new_n12248__;
  assign new_new_n28817__ = ~new_new_n28815__ & ~new_new_n28816__;
  assign new_new_n28818__ = ys__n45896 & new_new_n12245__;
  assign new_new_n28819__ = ys__n45799 & new_new_n12246__;
  assign new_new_n28820__ = ~new_new_n28818__ & ~new_new_n28819__;
  assign new_new_n28821__ = new_new_n28817__ & new_new_n28820__;
  assign new_new_n28822__ = new_new_n26807__ & ~new_new_n28821__;
  assign new_new_n28823__ = ~new_new_n28814__ & ~new_new_n28822__;
  assign new_new_n28824__ = new_new_n26882__ & ~new_new_n28823__;
  assign new_new_n28825__ = ~new_new_n26862__ & new_new_n28824__;
  assign ys__n26141 = new_new_n28806__ | new_new_n28825__;
  assign new_new_n28827__ = ys__n25980 & new_new_n26768__;
  assign new_new_n28828__ = ys__n26766 & ~new_new_n12365__;
  assign new_new_n28829__ = ys__n46315 & new_new_n12356__;
  assign new_new_n28830__ = ys__n46491 & new_new_n12248__;
  assign new_new_n28831__ = ~new_new_n28829__ & ~new_new_n28830__;
  assign new_new_n28832__ = ys__n46667 & new_new_n12245__;
  assign new_new_n28833__ = ys__n46843 & new_new_n12246__;
  assign new_new_n28834__ = ~new_new_n28832__ & ~new_new_n28833__;
  assign new_new_n28835__ = new_new_n28831__ & new_new_n28834__;
  assign new_new_n28836__ = new_new_n26798__ & ~new_new_n28835__;
  assign new_new_n28837__ = ys__n27518 & new_new_n12356__;
  assign new_new_n28838__ = ys__n27507 & new_new_n12248__;
  assign new_new_n28839__ = ~new_new_n28837__ & ~new_new_n28838__;
  assign new_new_n28840__ = ys__n27496 & new_new_n12245__;
  assign new_new_n28841__ = ys__n27481 & new_new_n12246__;
  assign new_new_n28842__ = ~new_new_n28840__ & ~new_new_n28841__;
  assign new_new_n28843__ = new_new_n28839__ & new_new_n28842__;
  assign new_new_n28844__ = new_new_n26779__ & ~new_new_n28843__;
  assign new_new_n28845__ = ys__n46252 & new_new_n12356__;
  assign new_new_n28846__ = ys__n46428 & new_new_n12248__;
  assign new_new_n28847__ = ~new_new_n28845__ & ~new_new_n28846__;
  assign new_new_n28848__ = ys__n46604 & new_new_n12245__;
  assign new_new_n28849__ = ys__n46780 & new_new_n12246__;
  assign new_new_n28850__ = ~new_new_n28848__ & ~new_new_n28849__;
  assign new_new_n28851__ = new_new_n28847__ & new_new_n28850__;
  assign new_new_n28852__ = new_new_n26788__ & ~new_new_n28851__;
  assign new_new_n28853__ = ~new_new_n28844__ & ~new_new_n28852__;
  assign new_new_n28854__ = ~new_new_n28836__ & new_new_n28853__;
  assign new_new_n28855__ = new_new_n26817__ & ~new_new_n28854__;
  assign new_new_n28856__ = ~new_new_n28828__ & ~new_new_n28855__;
  assign new_new_n28857__ = ~new_new_n26768__ & ~new_new_n28856__;
  assign new_new_n28858__ = ~new_new_n28827__ & ~new_new_n28857__;
  assign new_new_n28859__ = new_new_n26821__ & ~new_new_n28858__;
  assign new_new_n28860__ = ys__n25727 & ~new_new_n12286__;
  assign new_new_n28861__ = ys__n45634 & new_new_n12356__;
  assign new_new_n28862__ = ys__n45470 & new_new_n12248__;
  assign new_new_n28863__ = ~new_new_n28861__ & ~new_new_n28862__;
  assign new_new_n28864__ = ys__n45306 & new_new_n12245__;
  assign new_new_n28865__ = ys__n45113 & new_new_n12246__;
  assign new_new_n28866__ = ~new_new_n28864__ & ~new_new_n28865__;
  assign new_new_n28867__ = new_new_n28863__ & new_new_n28866__;
  assign new_new_n28868__ = new_new_n26779__ & ~new_new_n28867__;
  assign new_new_n28869__ = ys__n45702 & new_new_n12356__;
  assign new_new_n28870__ = ys__n45538 & new_new_n12248__;
  assign new_new_n28871__ = ~new_new_n28869__ & ~new_new_n28870__;
  assign new_new_n28872__ = ys__n45374 & new_new_n12245__;
  assign new_new_n28873__ = ys__n45212 & new_new_n12246__;
  assign new_new_n28874__ = ~new_new_n28872__ & ~new_new_n28873__;
  assign new_new_n28875__ = new_new_n28871__ & new_new_n28874__;
  assign new_new_n28876__ = new_new_n26798__ & ~new_new_n28875__;
  assign new_new_n28877__ = ~new_new_n28868__ & ~new_new_n28876__;
  assign new_new_n28878__ = new_new_n12244__ & ~new_new_n12250__;
  assign new_new_n28879__ = new_new_n26815__ & ~new_new_n28878__;
  assign new_new_n28880__ = new_new_n12286__ & new_new_n28879__;
  assign new_new_n28881__ = ~new_new_n28877__ & new_new_n28880__;
  assign new_new_n28882__ = ~new_new_n28860__ & ~new_new_n28881__;
  assign new_new_n28883__ = ~new_new_n26821__ & ~new_new_n28882__;
  assign new_new_n28884__ = ~new_new_n28859__ & ~new_new_n28883__;
  assign new_new_n28885__ = new_new_n26862__ & ~new_new_n28884__;
  assign new_new_n28886__ = ys__n25853 & ~new_new_n12395__;
  assign new_new_n28887__ = ys__n46127 & new_new_n12356__;
  assign new_new_n28888__ = ys__n46029 & new_new_n12248__;
  assign new_new_n28889__ = ~new_new_n28887__ & ~new_new_n28888__;
  assign new_new_n28890__ = ys__n45931 & new_new_n12245__;
  assign new_new_n28891__ = ys__n45835 & new_new_n12246__;
  assign new_new_n28892__ = ~new_new_n28890__ & ~new_new_n28891__;
  assign new_new_n28893__ = new_new_n28889__ & new_new_n28892__;
  assign new_new_n28894__ = new_new_n26798__ & new_new_n26815__;
  assign new_new_n28895__ = ~new_new_n28893__ & new_new_n28894__;
  assign new_new_n28896__ = new_new_n12395__ & new_new_n28895__;
  assign new_new_n28897__ = ~new_new_n28886__ & ~new_new_n28896__;
  assign new_new_n28898__ = ~new_new_n26862__ & ~new_new_n28897__;
  assign new_new_n28899__ = ~new_new_n28885__ & ~new_new_n28898__;
  assign new_new_n28900__ = ~new_new_n14022__ & ~new_new_n28899__;
  assign new_new_n28901__ = ys__n26143 & new_new_n14022__;
  assign ys__n26144 = new_new_n28900__ | new_new_n28901__;
  assign new_new_n28903__ = ys__n25984 & new_new_n26768__;
  assign new_new_n28904__ = ys__n26768 & ~new_new_n12365__;
  assign new_new_n28905__ = ys__n47108 & new_new_n12356__;
  assign new_new_n28906__ = ys__n47111 & new_new_n12248__;
  assign new_new_n28907__ = ~new_new_n28905__ & ~new_new_n28906__;
  assign new_new_n28908__ = ys__n47114 & new_new_n12245__;
  assign new_new_n28909__ = ys__n47117 & new_new_n12246__;
  assign new_new_n28910__ = ~new_new_n28908__ & ~new_new_n28909__;
  assign new_new_n28911__ = new_new_n28907__ & new_new_n28910__;
  assign new_new_n28912__ = new_new_n26779__ & ~new_new_n28911__;
  assign new_new_n28913__ = ys__n46254 & new_new_n12356__;
  assign new_new_n28914__ = ys__n46430 & new_new_n12248__;
  assign new_new_n28915__ = ~new_new_n28913__ & ~new_new_n28914__;
  assign new_new_n28916__ = ys__n46606 & new_new_n12245__;
  assign new_new_n28917__ = ys__n46782 & new_new_n12246__;
  assign new_new_n28918__ = ~new_new_n28916__ & ~new_new_n28917__;
  assign new_new_n28919__ = new_new_n28915__ & new_new_n28918__;
  assign new_new_n28920__ = new_new_n26788__ & ~new_new_n28919__;
  assign new_new_n28921__ = ~new_new_n28912__ & ~new_new_n28920__;
  assign new_new_n28922__ = ys__n46316 & new_new_n12356__;
  assign new_new_n28923__ = ys__n46492 & new_new_n12248__;
  assign new_new_n28924__ = ~new_new_n28922__ & ~new_new_n28923__;
  assign new_new_n28925__ = ys__n46668 & new_new_n12245__;
  assign new_new_n28926__ = ys__n46844 & new_new_n12246__;
  assign new_new_n28927__ = ~new_new_n28925__ & ~new_new_n28926__;
  assign new_new_n28928__ = new_new_n28924__ & new_new_n28927__;
  assign new_new_n28929__ = new_new_n26798__ & ~new_new_n28928__;
  assign new_new_n28930__ = ys__n46393 & new_new_n12356__;
  assign new_new_n28931__ = ys__n46569 & new_new_n12248__;
  assign new_new_n28932__ = ~new_new_n28930__ & ~new_new_n28931__;
  assign new_new_n28933__ = ys__n46745 & new_new_n12245__;
  assign new_new_n28934__ = ys__n46921 & new_new_n12246__;
  assign new_new_n28935__ = ~new_new_n28933__ & ~new_new_n28934__;
  assign new_new_n28936__ = new_new_n28932__ & new_new_n28935__;
  assign new_new_n28937__ = new_new_n26807__ & ~new_new_n28936__;
  assign new_new_n28938__ = ~new_new_n28929__ & ~new_new_n28937__;
  assign new_new_n28939__ = new_new_n28921__ & new_new_n28938__;
  assign new_new_n28940__ = new_new_n26817__ & ~new_new_n28939__;
  assign new_new_n28941__ = ~new_new_n28904__ & ~new_new_n28940__;
  assign new_new_n28942__ = ~new_new_n26768__ & ~new_new_n28941__;
  assign new_new_n28943__ = ~new_new_n28903__ & ~new_new_n28942__;
  assign new_new_n28944__ = new_new_n26821__ & ~new_new_n28943__;
  assign new_new_n28945__ = ys__n25730 & ~new_new_n12286__;
  assign new_new_n28946__ = new_new_n26779__ & new_new_n26815__;
  assign new_new_n28947__ = ys__n45636 & new_new_n12356__;
  assign new_new_n28948__ = ys__n45472 & new_new_n12248__;
  assign new_new_n28949__ = ~new_new_n28947__ & ~new_new_n28948__;
  assign new_new_n28950__ = ys__n45308 & new_new_n12245__;
  assign new_new_n28951__ = ys__n45116 & new_new_n12246__;
  assign new_new_n28952__ = ~new_new_n28950__ & ~new_new_n28951__;
  assign new_new_n28953__ = new_new_n28949__ & new_new_n28952__;
  assign new_new_n28954__ = ~new_new_n12240__ & new_new_n12355__;
  assign new_new_n28955__ = ~new_new_n28953__ & ~new_new_n28954__;
  assign new_new_n28956__ = new_new_n28946__ & new_new_n28955__;
  assign new_new_n28957__ = new_new_n12286__ & new_new_n28956__;
  assign new_new_n28958__ = ~new_new_n28945__ & ~new_new_n28957__;
  assign new_new_n28959__ = ~new_new_n26821__ & ~new_new_n28958__;
  assign new_new_n28960__ = ~new_new_n28944__ & ~new_new_n28959__;
  assign new_new_n28961__ = new_new_n26862__ & ~new_new_n28960__;
  assign new_new_n28962__ = ys__n25856 & ~new_new_n12395__;
  assign new_new_n28963__ = ys__n46096 & new_new_n12356__;
  assign new_new_n28964__ = ys__n45998 & new_new_n12248__;
  assign new_new_n28965__ = ~new_new_n28963__ & ~new_new_n28964__;
  assign new_new_n28966__ = ys__n45900 & new_new_n12245__;
  assign new_new_n28967__ = ys__n45804 & new_new_n12246__;
  assign new_new_n28968__ = ~new_new_n28966__ & ~new_new_n28967__;
  assign new_new_n28969__ = new_new_n28965__ & new_new_n28968__;
  assign new_new_n28970__ = new_new_n26788__ & ~new_new_n28969__;
  assign new_new_n28971__ = ys__n46034 & new_new_n12356__;
  assign new_new_n28972__ = ys__n45936 & new_new_n12248__;
  assign new_new_n28973__ = ~new_new_n28971__ & ~new_new_n28972__;
  assign new_new_n28974__ = ys__n45838 & new_new_n12245__;
  assign new_new_n28975__ = ys__n45712 & new_new_n12246__;
  assign new_new_n28976__ = ~new_new_n28974__ & ~new_new_n28975__;
  assign new_new_n28977__ = new_new_n28973__ & new_new_n28976__;
  assign new_new_n28978__ = new_new_n26807__ & ~new_new_n28977__;
  assign new_new_n28979__ = ~new_new_n28970__ & ~new_new_n28978__;
  assign new_new_n28980__ = new_new_n26882__ & ~new_new_n28979__;
  assign new_new_n28981__ = ~new_new_n28962__ & ~new_new_n28980__;
  assign new_new_n28982__ = ~new_new_n26862__ & ~new_new_n28981__;
  assign new_new_n28983__ = ~new_new_n28961__ & ~new_new_n28982__;
  assign new_new_n28984__ = ~new_new_n14022__ & ~new_new_n28983__;
  assign new_new_n28985__ = ys__n26145 & new_new_n14022__;
  assign ys__n26146 = new_new_n28984__ | new_new_n28985__;
  assign new_new_n28987__ = ys__n25987 & new_new_n26768__;
  assign new_new_n28988__ = ys__n26770 & ~new_new_n12365__;
  assign new_new_n28989__ = ys__n27520 & new_new_n12356__;
  assign new_new_n28990__ = ys__n27509 & new_new_n12248__;
  assign new_new_n28991__ = ~new_new_n28989__ & ~new_new_n28990__;
  assign new_new_n28992__ = ys__n27498 & new_new_n12245__;
  assign new_new_n28993__ = ys__n27485 & new_new_n12246__;
  assign new_new_n28994__ = ~new_new_n28992__ & ~new_new_n28993__;
  assign new_new_n28995__ = new_new_n28991__ & new_new_n28994__;
  assign new_new_n28996__ = new_new_n26779__ & ~new_new_n28995__;
  assign new_new_n28997__ = ys__n46256 & new_new_n12356__;
  assign new_new_n28998__ = ys__n46432 & new_new_n12248__;
  assign new_new_n28999__ = ~new_new_n28997__ & ~new_new_n28998__;
  assign new_new_n29000__ = ys__n46608 & new_new_n12245__;
  assign new_new_n29001__ = ys__n46784 & new_new_n12246__;
  assign new_new_n29002__ = ~new_new_n29000__ & ~new_new_n29001__;
  assign new_new_n29003__ = new_new_n28999__ & new_new_n29002__;
  assign new_new_n29004__ = new_new_n26788__ & ~new_new_n29003__;
  assign new_new_n29005__ = ~new_new_n28996__ & ~new_new_n29004__;
  assign new_new_n29006__ = ys__n46317 & new_new_n12356__;
  assign new_new_n29007__ = ys__n46493 & new_new_n12248__;
  assign new_new_n29008__ = ~new_new_n29006__ & ~new_new_n29007__;
  assign new_new_n29009__ = ys__n46669 & new_new_n12245__;
  assign new_new_n29010__ = ys__n46845 & new_new_n12246__;
  assign new_new_n29011__ = ~new_new_n29009__ & ~new_new_n29010__;
  assign new_new_n29012__ = new_new_n29008__ & new_new_n29011__;
  assign new_new_n29013__ = new_new_n26798__ & ~new_new_n29012__;
  assign new_new_n29014__ = ys__n46394 & new_new_n12356__;
  assign new_new_n29015__ = ys__n46570 & new_new_n12248__;
  assign new_new_n29016__ = ~new_new_n29014__ & ~new_new_n29015__;
  assign new_new_n29017__ = ys__n46746 & new_new_n12245__;
  assign new_new_n29018__ = ys__n46922 & new_new_n12246__;
  assign new_new_n29019__ = ~new_new_n29017__ & ~new_new_n29018__;
  assign new_new_n29020__ = new_new_n29016__ & new_new_n29019__;
  assign new_new_n29021__ = new_new_n26807__ & ~new_new_n29020__;
  assign new_new_n29022__ = ~new_new_n29013__ & ~new_new_n29021__;
  assign new_new_n29023__ = new_new_n29005__ & new_new_n29022__;
  assign new_new_n29024__ = new_new_n26817__ & ~new_new_n29023__;
  assign new_new_n29025__ = ~new_new_n28988__ & ~new_new_n29024__;
  assign new_new_n29026__ = ~new_new_n26768__ & ~new_new_n29025__;
  assign new_new_n29027__ = ~new_new_n28987__ & ~new_new_n29026__;
  assign new_new_n29028__ = new_new_n26821__ & ~new_new_n29027__;
  assign new_new_n29029__ = ys__n25733 & ~new_new_n12286__;
  assign new_new_n29030__ = ys__n45638 & new_new_n12356__;
  assign new_new_n29031__ = ys__n45474 & new_new_n12248__;
  assign new_new_n29032__ = ~new_new_n29030__ & ~new_new_n29031__;
  assign new_new_n29033__ = ys__n45310 & new_new_n12245__;
  assign new_new_n29034__ = ys__n45119 & new_new_n12246__;
  assign new_new_n29035__ = ~new_new_n29033__ & ~new_new_n29034__;
  assign new_new_n29036__ = new_new_n29032__ & new_new_n29035__;
  assign new_new_n29037__ = new_new_n26779__ & ~new_new_n29036__;
  assign new_new_n29038__ = ys__n45604 & new_new_n12356__;
  assign new_new_n29039__ = ys__n45440 & new_new_n12248__;
  assign new_new_n29040__ = ~new_new_n29038__ & ~new_new_n29039__;
  assign new_new_n29041__ = ys__n45276 & new_new_n12245__;
  assign new_new_n29042__ = ys__n45082 & new_new_n12246__;
  assign new_new_n29043__ = ~new_new_n29041__ & ~new_new_n29042__;
  assign new_new_n29044__ = new_new_n29040__ & new_new_n29043__;
  assign new_new_n29045__ = new_new_n26788__ & ~new_new_n29044__;
  assign new_new_n29046__ = ~new_new_n29037__ & ~new_new_n29045__;
  assign new_new_n29047__ = ys__n45704 & new_new_n12356__;
  assign new_new_n29048__ = ys__n45541 & new_new_n12248__;
  assign new_new_n29049__ = ~new_new_n29047__ & ~new_new_n29048__;
  assign new_new_n29050__ = ys__n45377 & new_new_n12245__;
  assign new_new_n29051__ = ys__n45214 & new_new_n12246__;
  assign new_new_n29052__ = ~new_new_n29050__ & ~new_new_n29051__;
  assign new_new_n29053__ = new_new_n29049__ & new_new_n29052__;
  assign new_new_n29054__ = new_new_n26798__ & ~new_new_n29053__;
  assign new_new_n29055__ = ys__n45544 & new_new_n12356__;
  assign new_new_n29056__ = ys__n45380 & new_new_n12248__;
  assign new_new_n29057__ = ~new_new_n29055__ & ~new_new_n29056__;
  assign new_new_n29058__ = ys__n45216 & new_new_n12245__;
  assign new_new_n29059__ = ys__n44993 & new_new_n12246__;
  assign new_new_n29060__ = ~new_new_n29058__ & ~new_new_n29059__;
  assign new_new_n29061__ = new_new_n29057__ & new_new_n29060__;
  assign new_new_n29062__ = new_new_n26807__ & ~new_new_n29061__;
  assign new_new_n29063__ = ~new_new_n29054__ & ~new_new_n29062__;
  assign new_new_n29064__ = new_new_n29046__ & new_new_n29063__;
  assign new_new_n29065__ = new_new_n26858__ & ~new_new_n29064__;
  assign new_new_n29066__ = ~new_new_n29029__ & ~new_new_n29065__;
  assign new_new_n29067__ = ~new_new_n26821__ & ~new_new_n29066__;
  assign new_new_n29068__ = ~new_new_n29028__ & ~new_new_n29067__;
  assign new_new_n29069__ = new_new_n26862__ & ~new_new_n29068__;
  assign new_new_n29070__ = ys__n25859 & ~new_new_n12395__;
  assign new_new_n29071__ = ys__n46036 & new_new_n12356__;
  assign new_new_n29072__ = ys__n45938 & new_new_n12248__;
  assign new_new_n29073__ = ~new_new_n29071__ & ~new_new_n29072__;
  assign new_new_n29074__ = ys__n45840 & new_new_n12245__;
  assign new_new_n29075__ = ys__n45715 & new_new_n12246__;
  assign new_new_n29076__ = ~new_new_n29074__ & ~new_new_n29075__;
  assign new_new_n29077__ = new_new_n29073__ & new_new_n29076__;
  assign new_new_n29078__ = new_new_n26807__ & ~new_new_n29077__;
  assign new_new_n29079__ = ys__n46097 & new_new_n12356__;
  assign new_new_n29080__ = ys__n45999 & new_new_n12248__;
  assign new_new_n29081__ = ~new_new_n29079__ & ~new_new_n29080__;
  assign new_new_n29082__ = ys__n45901 & new_new_n12245__;
  assign new_new_n29083__ = ys__n45805 & new_new_n12246__;
  assign new_new_n29084__ = ~new_new_n29082__ & ~new_new_n29083__;
  assign new_new_n29085__ = new_new_n29081__ & new_new_n29084__;
  assign new_new_n29086__ = new_new_n26788__ & ~new_new_n29085__;
  assign new_new_n29087__ = ys__n46128 & new_new_n12356__;
  assign new_new_n29088__ = ys__n46031 & new_new_n12248__;
  assign new_new_n29089__ = ~new_new_n29087__ & ~new_new_n29088__;
  assign new_new_n29090__ = ys__n45933 & new_new_n12245__;
  assign new_new_n29091__ = ys__n45836 & new_new_n12246__;
  assign new_new_n29092__ = ~new_new_n29090__ & ~new_new_n29091__;
  assign new_new_n29093__ = new_new_n29089__ & new_new_n29092__;
  assign new_new_n29094__ = new_new_n26798__ & ~new_new_n29093__;
  assign new_new_n29095__ = ~new_new_n29086__ & ~new_new_n29094__;
  assign new_new_n29096__ = ~new_new_n29078__ & new_new_n29095__;
  assign new_new_n29097__ = ~new_new_n12241__ & new_new_n12377__;
  assign new_new_n29098__ = new_new_n26815__ & ~new_new_n29097__;
  assign new_new_n29099__ = new_new_n12395__ & new_new_n29098__;
  assign new_new_n29100__ = ~new_new_n29096__ & new_new_n29099__;
  assign new_new_n29101__ = ~new_new_n29070__ & ~new_new_n29100__;
  assign new_new_n29102__ = ~new_new_n26862__ & ~new_new_n29101__;
  assign new_new_n29103__ = ~new_new_n29069__ & ~new_new_n29102__;
  assign new_new_n29104__ = ~new_new_n14022__ & ~new_new_n29103__;
  assign new_new_n29105__ = ys__n26147 & new_new_n14022__;
  assign ys__n26148 = new_new_n29104__ | new_new_n29105__;
  assign new_new_n29107__ = ys__n25990 & new_new_n26768__;
  assign new_new_n29108__ = ys__n26772 & ~new_new_n12365__;
  assign new_new_n29109__ = ys__n47109 & new_new_n12356__;
  assign new_new_n29110__ = ys__n47112 & new_new_n12248__;
  assign new_new_n29111__ = ~new_new_n29109__ & ~new_new_n29110__;
  assign new_new_n29112__ = ys__n47115 & new_new_n12245__;
  assign new_new_n29113__ = ys__n47118 & new_new_n12246__;
  assign new_new_n29114__ = ~new_new_n29112__ & ~new_new_n29113__;
  assign new_new_n29115__ = new_new_n29111__ & new_new_n29114__;
  assign new_new_n29116__ = new_new_n26779__ & ~new_new_n29115__;
  assign new_new_n29117__ = ys__n46258 & new_new_n12356__;
  assign new_new_n29118__ = ys__n46434 & new_new_n12248__;
  assign new_new_n29119__ = ~new_new_n29117__ & ~new_new_n29118__;
  assign new_new_n29120__ = ys__n46610 & new_new_n12245__;
  assign new_new_n29121__ = ys__n46786 & new_new_n12246__;
  assign new_new_n29122__ = ~new_new_n29120__ & ~new_new_n29121__;
  assign new_new_n29123__ = new_new_n29119__ & new_new_n29122__;
  assign new_new_n29124__ = new_new_n26788__ & ~new_new_n29123__;
  assign new_new_n29125__ = ~new_new_n29116__ & ~new_new_n29124__;
  assign new_new_n29126__ = ys__n46318 & new_new_n12356__;
  assign new_new_n29127__ = ys__n46494 & new_new_n12248__;
  assign new_new_n29128__ = ~new_new_n29126__ & ~new_new_n29127__;
  assign new_new_n29129__ = ys__n46670 & new_new_n12245__;
  assign new_new_n29130__ = ys__n46846 & new_new_n12246__;
  assign new_new_n29131__ = ~new_new_n29129__ & ~new_new_n29130__;
  assign new_new_n29132__ = new_new_n29128__ & new_new_n29131__;
  assign new_new_n29133__ = new_new_n26798__ & ~new_new_n29132__;
  assign new_new_n29134__ = ys__n46395 & new_new_n12356__;
  assign new_new_n29135__ = ys__n46571 & new_new_n12248__;
  assign new_new_n29136__ = ~new_new_n29134__ & ~new_new_n29135__;
  assign new_new_n29137__ = ys__n46747 & new_new_n12245__;
  assign new_new_n29138__ = ys__n46923 & new_new_n12246__;
  assign new_new_n29139__ = ~new_new_n29137__ & ~new_new_n29138__;
  assign new_new_n29140__ = new_new_n29136__ & new_new_n29139__;
  assign new_new_n29141__ = new_new_n26807__ & ~new_new_n29140__;
  assign new_new_n29142__ = ~new_new_n29133__ & ~new_new_n29141__;
  assign new_new_n29143__ = new_new_n29125__ & new_new_n29142__;
  assign new_new_n29144__ = new_new_n26817__ & ~new_new_n29143__;
  assign new_new_n29145__ = ~new_new_n29108__ & ~new_new_n29144__;
  assign new_new_n29146__ = ~new_new_n26768__ & ~new_new_n29145__;
  assign new_new_n29147__ = ~new_new_n29107__ & ~new_new_n29146__;
  assign new_new_n29148__ = new_new_n26821__ & ~new_new_n29147__;
  assign new_new_n29149__ = ys__n25736 & ~new_new_n12286__;
  assign new_new_n29150__ = ys__n45546 & new_new_n12356__;
  assign new_new_n29151__ = ys__n45382 & new_new_n12248__;
  assign new_new_n29152__ = ~new_new_n29150__ & ~new_new_n29151__;
  assign new_new_n29153__ = ys__n45218 & new_new_n12245__;
  assign new_new_n29154__ = ys__n44996 & new_new_n12246__;
  assign new_new_n29155__ = ~new_new_n29153__ & ~new_new_n29154__;
  assign new_new_n29156__ = new_new_n29152__ & new_new_n29155__;
  assign new_new_n29157__ = new_new_n26807__ & ~new_new_n29156__;
  assign new_new_n29158__ = ys__n45640 & new_new_n12356__;
  assign new_new_n29159__ = ys__n45476 & new_new_n12248__;
  assign new_new_n29160__ = ~new_new_n29158__ & ~new_new_n29159__;
  assign new_new_n29161__ = ys__n45312 & new_new_n12245__;
  assign new_new_n29162__ = ys__n45122 & new_new_n12246__;
  assign new_new_n29163__ = ~new_new_n29161__ & ~new_new_n29162__;
  assign new_new_n29164__ = new_new_n29160__ & new_new_n29163__;
  assign new_new_n29165__ = new_new_n26779__ & ~new_new_n29164__;
  assign new_new_n29166__ = ys__n45605 & new_new_n12356__;
  assign new_new_n29167__ = ys__n45441 & new_new_n12248__;
  assign new_new_n29168__ = ~new_new_n29166__ & ~new_new_n29167__;
  assign new_new_n29169__ = ys__n45277 & new_new_n12245__;
  assign new_new_n29170__ = ys__n45083 & new_new_n12246__;
  assign new_new_n29171__ = ~new_new_n29169__ & ~new_new_n29170__;
  assign new_new_n29172__ = new_new_n29168__ & new_new_n29171__;
  assign new_new_n29173__ = new_new_n26788__ & ~new_new_n29172__;
  assign new_new_n29174__ = ~new_new_n29165__ & ~new_new_n29173__;
  assign new_new_n29175__ = ~new_new_n29157__ & new_new_n29174__;
  assign new_new_n29176__ = new_new_n26858__ & ~new_new_n29175__;
  assign new_new_n29177__ = ~new_new_n29149__ & ~new_new_n29176__;
  assign new_new_n29178__ = ~new_new_n26821__ & ~new_new_n29177__;
  assign new_new_n29179__ = ~new_new_n29148__ & ~new_new_n29178__;
  assign new_new_n29180__ = new_new_n26862__ & ~new_new_n29179__;
  assign new_new_n29181__ = ys__n25862 & ~new_new_n12395__;
  assign new_new_n29182__ = ys__n46098 & new_new_n12356__;
  assign new_new_n29183__ = ys__n46000 & new_new_n12248__;
  assign new_new_n29184__ = ~new_new_n29182__ & ~new_new_n29183__;
  assign new_new_n29185__ = ys__n45902 & new_new_n12245__;
  assign new_new_n29186__ = ys__n45806 & new_new_n12246__;
  assign new_new_n29187__ = ~new_new_n29185__ & ~new_new_n29186__;
  assign new_new_n29188__ = new_new_n29184__ & new_new_n29187__;
  assign new_new_n29189__ = new_new_n26788__ & ~new_new_n29188__;
  assign new_new_n29190__ = ys__n46038 & new_new_n12356__;
  assign new_new_n29191__ = ys__n45940 & new_new_n12248__;
  assign new_new_n29192__ = ~new_new_n29190__ & ~new_new_n29191__;
  assign new_new_n29193__ = ys__n45842 & new_new_n12245__;
  assign new_new_n29194__ = ys__n45718 & new_new_n12246__;
  assign new_new_n29195__ = ~new_new_n29193__ & ~new_new_n29194__;
  assign new_new_n29196__ = new_new_n29192__ & new_new_n29195__;
  assign new_new_n29197__ = new_new_n26807__ & ~new_new_n29196__;
  assign new_new_n29198__ = ~new_new_n29189__ & ~new_new_n29197__;
  assign new_new_n29199__ = new_new_n26882__ & ~new_new_n29198__;
  assign new_new_n29200__ = ~new_new_n29181__ & ~new_new_n29199__;
  assign new_new_n29201__ = ~new_new_n26862__ & ~new_new_n29200__;
  assign new_new_n29202__ = ~new_new_n29180__ & ~new_new_n29201__;
  assign new_new_n29203__ = ~new_new_n14022__ & ~new_new_n29202__;
  assign new_new_n29204__ = ys__n26149 & new_new_n14022__;
  assign ys__n26150 = new_new_n29203__ | new_new_n29204__;
  assign new_new_n29206__ = ys__n25993 & new_new_n26768__;
  assign new_new_n29207__ = ys__n27510 & new_new_n12356__;
  assign new_new_n29208__ = ys__n27499 & new_new_n12248__;
  assign new_new_n29209__ = ~new_new_n29207__ & ~new_new_n29208__;
  assign new_new_n29210__ = ys__n27488 & new_new_n12245__;
  assign new_new_n29211__ = ys__n27479 & new_new_n12246__;
  assign new_new_n29212__ = ~new_new_n29210__ & ~new_new_n29211__;
  assign new_new_n29213__ = new_new_n29209__ & new_new_n29212__;
  assign new_new_n29214__ = new_new_n26779__ & ~new_new_n29213__;
  assign new_new_n29215__ = ys__n46260 & new_new_n12356__;
  assign new_new_n29216__ = ys__n46436 & new_new_n12248__;
  assign new_new_n29217__ = ~new_new_n29215__ & ~new_new_n29216__;
  assign new_new_n29218__ = ys__n46612 & new_new_n12245__;
  assign new_new_n29219__ = ys__n46788 & new_new_n12246__;
  assign new_new_n29220__ = ~new_new_n29218__ & ~new_new_n29219__;
  assign new_new_n29221__ = new_new_n29217__ & new_new_n29220__;
  assign new_new_n29222__ = new_new_n26788__ & ~new_new_n29221__;
  assign new_new_n29223__ = ~new_new_n29214__ & ~new_new_n29222__;
  assign new_new_n29224__ = ys__n46319 & new_new_n12356__;
  assign new_new_n29225__ = ys__n46495 & new_new_n12248__;
  assign new_new_n29226__ = ~new_new_n29224__ & ~new_new_n29225__;
  assign new_new_n29227__ = ys__n46671 & new_new_n12245__;
  assign new_new_n29228__ = ys__n46847 & new_new_n12246__;
  assign new_new_n29229__ = ~new_new_n29227__ & ~new_new_n29228__;
  assign new_new_n29230__ = new_new_n29226__ & new_new_n29229__;
  assign new_new_n29231__ = new_new_n26798__ & ~new_new_n29230__;
  assign new_new_n29232__ = ys__n46396 & new_new_n12356__;
  assign new_new_n29233__ = ys__n46572 & new_new_n12248__;
  assign new_new_n29234__ = ~new_new_n29232__ & ~new_new_n29233__;
  assign new_new_n29235__ = ys__n46748 & new_new_n12245__;
  assign new_new_n29236__ = ys__n46924 & new_new_n12246__;
  assign new_new_n29237__ = ~new_new_n29235__ & ~new_new_n29236__;
  assign new_new_n29238__ = new_new_n29234__ & new_new_n29237__;
  assign new_new_n29239__ = new_new_n26807__ & ~new_new_n29238__;
  assign new_new_n29240__ = ~new_new_n29231__ & ~new_new_n29239__;
  assign new_new_n29241__ = new_new_n29223__ & new_new_n29240__;
  assign new_new_n29242__ = new_new_n26818__ & ~new_new_n29241__;
  assign new_new_n29243__ = ~new_new_n29206__ & ~new_new_n29242__;
  assign new_new_n29244__ = new_new_n26821__ & ~new_new_n29243__;
  assign new_new_n29245__ = ys__n45642 & new_new_n12356__;
  assign new_new_n29246__ = ys__n45478 & new_new_n12248__;
  assign new_new_n29247__ = ~new_new_n29245__ & ~new_new_n29246__;
  assign new_new_n29248__ = ys__n45314 & new_new_n12245__;
  assign new_new_n29249__ = ys__n45125 & new_new_n12246__;
  assign new_new_n29250__ = ~new_new_n29248__ & ~new_new_n29249__;
  assign new_new_n29251__ = new_new_n29247__ & new_new_n29250__;
  assign new_new_n29252__ = new_new_n26779__ & ~new_new_n29251__;
  assign new_new_n29253__ = ys__n45606 & new_new_n12356__;
  assign new_new_n29254__ = ys__n45442 & new_new_n12248__;
  assign new_new_n29255__ = ~new_new_n29253__ & ~new_new_n29254__;
  assign new_new_n29256__ = ys__n45278 & new_new_n12245__;
  assign new_new_n29257__ = ys__n45084 & new_new_n12246__;
  assign new_new_n29258__ = ~new_new_n29256__ & ~new_new_n29257__;
  assign new_new_n29259__ = new_new_n29255__ & new_new_n29258__;
  assign new_new_n29260__ = new_new_n26788__ & ~new_new_n29259__;
  assign new_new_n29261__ = ~new_new_n29252__ & ~new_new_n29260__;
  assign new_new_n29262__ = ys__n45698 & new_new_n12356__;
  assign new_new_n29263__ = ys__n45534 & new_new_n12248__;
  assign new_new_n29264__ = ~new_new_n29262__ & ~new_new_n29263__;
  assign new_new_n29265__ = ys__n45370 & new_new_n12245__;
  assign new_new_n29266__ = ys__n45208 & new_new_n12246__;
  assign new_new_n29267__ = ~new_new_n29265__ & ~new_new_n29266__;
  assign new_new_n29268__ = new_new_n29264__ & new_new_n29267__;
  assign new_new_n29269__ = new_new_n26798__ & ~new_new_n29268__;
  assign new_new_n29270__ = ys__n45548 & new_new_n12356__;
  assign new_new_n29271__ = ys__n45384 & new_new_n12248__;
  assign new_new_n29272__ = ~new_new_n29270__ & ~new_new_n29271__;
  assign new_new_n29273__ = ys__n45220 & new_new_n12245__;
  assign new_new_n29274__ = ys__n44999 & new_new_n12246__;
  assign new_new_n29275__ = ~new_new_n29273__ & ~new_new_n29274__;
  assign new_new_n29276__ = new_new_n29272__ & new_new_n29275__;
  assign new_new_n29277__ = new_new_n26807__ & ~new_new_n29276__;
  assign new_new_n29278__ = ~new_new_n29269__ & ~new_new_n29277__;
  assign new_new_n29279__ = new_new_n29261__ & new_new_n29278__;
  assign new_new_n29280__ = new_new_n26859__ & ~new_new_n29279__;
  assign new_new_n29281__ = ~new_new_n29244__ & ~new_new_n29280__;
  assign new_new_n29282__ = new_new_n26862__ & ~new_new_n29281__;
  assign new_new_n29283__ = ys__n46099 & new_new_n12356__;
  assign new_new_n29284__ = ys__n46001 & new_new_n12248__;
  assign new_new_n29285__ = ~new_new_n29283__ & ~new_new_n29284__;
  assign new_new_n29286__ = ys__n45903 & new_new_n12245__;
  assign new_new_n29287__ = ys__n45807 & new_new_n12246__;
  assign new_new_n29288__ = ~new_new_n29286__ & ~new_new_n29287__;
  assign new_new_n29289__ = new_new_n29285__ & new_new_n29288__;
  assign new_new_n29290__ = new_new_n26788__ & ~new_new_n29289__;
  assign new_new_n29291__ = ys__n46040 & new_new_n12356__;
  assign new_new_n29292__ = ys__n45942 & new_new_n12248__;
  assign new_new_n29293__ = ~new_new_n29291__ & ~new_new_n29292__;
  assign new_new_n29294__ = ys__n45844 & new_new_n12245__;
  assign new_new_n29295__ = ys__n45721 & new_new_n12246__;
  assign new_new_n29296__ = ~new_new_n29294__ & ~new_new_n29295__;
  assign new_new_n29297__ = new_new_n29293__ & new_new_n29296__;
  assign new_new_n29298__ = new_new_n26807__ & ~new_new_n29297__;
  assign new_new_n29299__ = ~new_new_n29290__ & ~new_new_n29298__;
  assign new_new_n29300__ = new_new_n26882__ & ~new_new_n29299__;
  assign new_new_n29301__ = ~new_new_n26862__ & new_new_n29300__;
  assign new_new_n29302__ = ~new_new_n29282__ & ~new_new_n29301__;
  assign new_new_n29303__ = ~new_new_n14022__ & ~new_new_n29302__;
  assign new_new_n29304__ = ys__n26151 & new_new_n14022__;
  assign ys__n26152 = new_new_n29303__ | new_new_n29304__;
  assign new_new_n29306__ = ys__n25996 & new_new_n26768__;
  assign new_new_n29307__ = ys__n18045 & new_new_n12356__;
  assign new_new_n29308__ = ys__n18051 & new_new_n12248__;
  assign new_new_n29309__ = ~new_new_n29307__ & ~new_new_n29308__;
  assign new_new_n29310__ = ys__n18057 & new_new_n12245__;
  assign new_new_n29311__ = ys__n18067 & new_new_n12246__;
  assign new_new_n29312__ = ~new_new_n29310__ & ~new_new_n29311__;
  assign new_new_n29313__ = new_new_n29309__ & new_new_n29312__;
  assign new_new_n29314__ = new_new_n26779__ & ~new_new_n29313__;
  assign new_new_n29315__ = ys__n46262 & new_new_n12356__;
  assign new_new_n29316__ = ys__n46438 & new_new_n12248__;
  assign new_new_n29317__ = ~new_new_n29315__ & ~new_new_n29316__;
  assign new_new_n29318__ = ys__n46614 & new_new_n12245__;
  assign new_new_n29319__ = ys__n46790 & new_new_n12246__;
  assign new_new_n29320__ = ~new_new_n29318__ & ~new_new_n29319__;
  assign new_new_n29321__ = new_new_n29317__ & new_new_n29320__;
  assign new_new_n29322__ = new_new_n26788__ & ~new_new_n29321__;
  assign new_new_n29323__ = ~new_new_n29314__ & ~new_new_n29322__;
  assign new_new_n29324__ = ys__n46320 & new_new_n12356__;
  assign new_new_n29325__ = ys__n46496 & new_new_n12248__;
  assign new_new_n29326__ = ~new_new_n29324__ & ~new_new_n29325__;
  assign new_new_n29327__ = ys__n46672 & new_new_n12245__;
  assign new_new_n29328__ = ys__n46848 & new_new_n12246__;
  assign new_new_n29329__ = ~new_new_n29327__ & ~new_new_n29328__;
  assign new_new_n29330__ = new_new_n29326__ & new_new_n29329__;
  assign new_new_n29331__ = new_new_n26798__ & ~new_new_n29330__;
  assign new_new_n29332__ = ys__n46397 & new_new_n12356__;
  assign new_new_n29333__ = ys__n46573 & new_new_n12248__;
  assign new_new_n29334__ = ~new_new_n29332__ & ~new_new_n29333__;
  assign new_new_n29335__ = ys__n46749 & new_new_n12245__;
  assign new_new_n29336__ = ys__n46925 & new_new_n12246__;
  assign new_new_n29337__ = ~new_new_n29335__ & ~new_new_n29336__;
  assign new_new_n29338__ = new_new_n29334__ & new_new_n29337__;
  assign new_new_n29339__ = new_new_n26807__ & ~new_new_n29338__;
  assign new_new_n29340__ = ~new_new_n29331__ & ~new_new_n29339__;
  assign new_new_n29341__ = new_new_n29323__ & new_new_n29340__;
  assign new_new_n29342__ = new_new_n26818__ & ~new_new_n29341__;
  assign new_new_n29343__ = ~new_new_n29306__ & ~new_new_n29342__;
  assign new_new_n29344__ = new_new_n26821__ & ~new_new_n29343__;
  assign new_new_n29345__ = ys__n45644 & new_new_n12356__;
  assign new_new_n29346__ = ys__n45480 & new_new_n12248__;
  assign new_new_n29347__ = ~new_new_n29345__ & ~new_new_n29346__;
  assign new_new_n29348__ = ys__n45316 & new_new_n12245__;
  assign new_new_n29349__ = ys__n45128 & new_new_n12246__;
  assign new_new_n29350__ = ~new_new_n29348__ & ~new_new_n29349__;
  assign new_new_n29351__ = new_new_n29347__ & new_new_n29350__;
  assign new_new_n29352__ = new_new_n26779__ & ~new_new_n29351__;
  assign new_new_n29353__ = ys__n45607 & new_new_n12356__;
  assign new_new_n29354__ = ys__n45443 & new_new_n12248__;
  assign new_new_n29355__ = ~new_new_n29353__ & ~new_new_n29354__;
  assign new_new_n29356__ = ys__n45279 & new_new_n12245__;
  assign new_new_n29357__ = ys__n45085 & new_new_n12246__;
  assign new_new_n29358__ = ~new_new_n29356__ & ~new_new_n29357__;
  assign new_new_n29359__ = new_new_n29355__ & new_new_n29358__;
  assign new_new_n29360__ = new_new_n26788__ & ~new_new_n29359__;
  assign new_new_n29361__ = ~new_new_n29352__ & ~new_new_n29360__;
  assign new_new_n29362__ = ys__n45699 & new_new_n12356__;
  assign new_new_n29363__ = ys__n45535 & new_new_n12248__;
  assign new_new_n29364__ = ~new_new_n29362__ & ~new_new_n29363__;
  assign new_new_n29365__ = ys__n45371 & new_new_n12245__;
  assign new_new_n29366__ = ys__n45209 & new_new_n12246__;
  assign new_new_n29367__ = ~new_new_n29365__ & ~new_new_n29366__;
  assign new_new_n29368__ = new_new_n29364__ & new_new_n29367__;
  assign new_new_n29369__ = new_new_n26798__ & ~new_new_n29368__;
  assign new_new_n29370__ = ys__n45550 & new_new_n12356__;
  assign new_new_n29371__ = ys__n45386 & new_new_n12248__;
  assign new_new_n29372__ = ~new_new_n29370__ & ~new_new_n29371__;
  assign new_new_n29373__ = ys__n45222 & new_new_n12245__;
  assign new_new_n29374__ = ys__n45002 & new_new_n12246__;
  assign new_new_n29375__ = ~new_new_n29373__ & ~new_new_n29374__;
  assign new_new_n29376__ = new_new_n29372__ & new_new_n29375__;
  assign new_new_n29377__ = new_new_n26807__ & ~new_new_n29376__;
  assign new_new_n29378__ = ~new_new_n29369__ & ~new_new_n29377__;
  assign new_new_n29379__ = new_new_n29361__ & new_new_n29378__;
  assign new_new_n29380__ = new_new_n26859__ & ~new_new_n29379__;
  assign new_new_n29381__ = ~new_new_n29344__ & ~new_new_n29380__;
  assign new_new_n29382__ = new_new_n26862__ & ~new_new_n29381__;
  assign new_new_n29383__ = ys__n46100 & new_new_n12356__;
  assign new_new_n29384__ = ys__n46002 & new_new_n12248__;
  assign new_new_n29385__ = ~new_new_n29383__ & ~new_new_n29384__;
  assign new_new_n29386__ = ys__n45904 & new_new_n12245__;
  assign new_new_n29387__ = ys__n45808 & new_new_n12246__;
  assign new_new_n29388__ = ~new_new_n29386__ & ~new_new_n29387__;
  assign new_new_n29389__ = new_new_n29385__ & new_new_n29388__;
  assign new_new_n29390__ = new_new_n26788__ & ~new_new_n29389__;
  assign new_new_n29391__ = ys__n46042 & new_new_n12356__;
  assign new_new_n29392__ = ys__n45944 & new_new_n12248__;
  assign new_new_n29393__ = ~new_new_n29391__ & ~new_new_n29392__;
  assign new_new_n29394__ = ys__n45846 & new_new_n12245__;
  assign new_new_n29395__ = ys__n45724 & new_new_n12246__;
  assign new_new_n29396__ = ~new_new_n29394__ & ~new_new_n29395__;
  assign new_new_n29397__ = new_new_n29393__ & new_new_n29396__;
  assign new_new_n29398__ = new_new_n26807__ & ~new_new_n29397__;
  assign new_new_n29399__ = ~new_new_n29390__ & ~new_new_n29398__;
  assign new_new_n29400__ = new_new_n26882__ & ~new_new_n29399__;
  assign new_new_n29401__ = ~new_new_n26862__ & new_new_n29400__;
  assign new_new_n29402__ = ~new_new_n29382__ & ~new_new_n29401__;
  assign new_new_n29403__ = ~new_new_n14022__ & ~new_new_n29402__;
  assign new_new_n29404__ = ys__n26153 & new_new_n14022__;
  assign ys__n26154 = new_new_n29403__ | new_new_n29404__;
  assign new_new_n29406__ = ys__n25999 & new_new_n26768__;
  assign new_new_n29407__ = ys__n18043 & new_new_n12356__;
  assign new_new_n29408__ = ys__n18049 & new_new_n12248__;
  assign new_new_n29409__ = ~new_new_n29407__ & ~new_new_n29408__;
  assign new_new_n29410__ = ys__n18055 & new_new_n12245__;
  assign new_new_n29411__ = ys__n18063 & new_new_n12246__;
  assign new_new_n29412__ = ~new_new_n29410__ & ~new_new_n29411__;
  assign new_new_n29413__ = new_new_n29409__ & new_new_n29412__;
  assign new_new_n29414__ = new_new_n26779__ & ~new_new_n29413__;
  assign new_new_n29415__ = ys__n46264 & new_new_n12356__;
  assign new_new_n29416__ = ys__n46440 & new_new_n12248__;
  assign new_new_n29417__ = ~new_new_n29415__ & ~new_new_n29416__;
  assign new_new_n29418__ = ys__n46616 & new_new_n12245__;
  assign new_new_n29419__ = ys__n46792 & new_new_n12246__;
  assign new_new_n29420__ = ~new_new_n29418__ & ~new_new_n29419__;
  assign new_new_n29421__ = new_new_n29417__ & new_new_n29420__;
  assign new_new_n29422__ = new_new_n26788__ & ~new_new_n29421__;
  assign new_new_n29423__ = ~new_new_n29414__ & ~new_new_n29422__;
  assign new_new_n29424__ = ys__n46321 & new_new_n12356__;
  assign new_new_n29425__ = ys__n46497 & new_new_n12248__;
  assign new_new_n29426__ = ~new_new_n29424__ & ~new_new_n29425__;
  assign new_new_n29427__ = ys__n46673 & new_new_n12245__;
  assign new_new_n29428__ = ys__n46849 & new_new_n12246__;
  assign new_new_n29429__ = ~new_new_n29427__ & ~new_new_n29428__;
  assign new_new_n29430__ = new_new_n29426__ & new_new_n29429__;
  assign new_new_n29431__ = new_new_n26798__ & ~new_new_n29430__;
  assign new_new_n29432__ = ys__n46398 & new_new_n12356__;
  assign new_new_n29433__ = ys__n46574 & new_new_n12248__;
  assign new_new_n29434__ = ~new_new_n29432__ & ~new_new_n29433__;
  assign new_new_n29435__ = ys__n46750 & new_new_n12245__;
  assign new_new_n29436__ = ys__n46926 & new_new_n12246__;
  assign new_new_n29437__ = ~new_new_n29435__ & ~new_new_n29436__;
  assign new_new_n29438__ = new_new_n29434__ & new_new_n29437__;
  assign new_new_n29439__ = new_new_n26807__ & ~new_new_n29438__;
  assign new_new_n29440__ = ~new_new_n29431__ & ~new_new_n29439__;
  assign new_new_n29441__ = new_new_n29423__ & new_new_n29440__;
  assign new_new_n29442__ = new_new_n26818__ & ~new_new_n29441__;
  assign new_new_n29443__ = ~new_new_n29406__ & ~new_new_n29442__;
  assign new_new_n29444__ = new_new_n26821__ & ~new_new_n29443__;
  assign new_new_n29445__ = ys__n45646 & new_new_n12356__;
  assign new_new_n29446__ = ys__n45482 & new_new_n12248__;
  assign new_new_n29447__ = ~new_new_n29445__ & ~new_new_n29446__;
  assign new_new_n29448__ = ys__n45318 & new_new_n12245__;
  assign new_new_n29449__ = ys__n45131 & new_new_n12246__;
  assign new_new_n29450__ = ~new_new_n29448__ & ~new_new_n29449__;
  assign new_new_n29451__ = new_new_n29447__ & new_new_n29450__;
  assign new_new_n29452__ = new_new_n26779__ & ~new_new_n29451__;
  assign new_new_n29453__ = ys__n45608 & new_new_n12356__;
  assign new_new_n29454__ = ys__n45444 & new_new_n12248__;
  assign new_new_n29455__ = ~new_new_n29453__ & ~new_new_n29454__;
  assign new_new_n29456__ = ys__n45280 & new_new_n12245__;
  assign new_new_n29457__ = ys__n45086 & new_new_n12246__;
  assign new_new_n29458__ = ~new_new_n29456__ & ~new_new_n29457__;
  assign new_new_n29459__ = new_new_n29455__ & new_new_n29458__;
  assign new_new_n29460__ = new_new_n26788__ & ~new_new_n29459__;
  assign new_new_n29461__ = ~new_new_n29452__ & ~new_new_n29460__;
  assign new_new_n29462__ = ys__n45700 & new_new_n12356__;
  assign new_new_n29463__ = ys__n45536 & new_new_n12248__;
  assign new_new_n29464__ = ~new_new_n29462__ & ~new_new_n29463__;
  assign new_new_n29465__ = ys__n45372 & new_new_n12245__;
  assign new_new_n29466__ = ys__n45210 & new_new_n12246__;
  assign new_new_n29467__ = ~new_new_n29465__ & ~new_new_n29466__;
  assign new_new_n29468__ = new_new_n29464__ & new_new_n29467__;
  assign new_new_n29469__ = new_new_n26798__ & ~new_new_n29468__;
  assign new_new_n29470__ = ys__n45552 & new_new_n12356__;
  assign new_new_n29471__ = ys__n45388 & new_new_n12248__;
  assign new_new_n29472__ = ~new_new_n29470__ & ~new_new_n29471__;
  assign new_new_n29473__ = ys__n45224 & new_new_n12245__;
  assign new_new_n29474__ = ys__n45005 & new_new_n12246__;
  assign new_new_n29475__ = ~new_new_n29473__ & ~new_new_n29474__;
  assign new_new_n29476__ = new_new_n29472__ & new_new_n29475__;
  assign new_new_n29477__ = new_new_n26807__ & ~new_new_n29476__;
  assign new_new_n29478__ = ~new_new_n29469__ & ~new_new_n29477__;
  assign new_new_n29479__ = new_new_n29461__ & new_new_n29478__;
  assign new_new_n29480__ = new_new_n26859__ & ~new_new_n29479__;
  assign new_new_n29481__ = ~new_new_n29444__ & ~new_new_n29480__;
  assign new_new_n29482__ = new_new_n26862__ & ~new_new_n29481__;
  assign new_new_n29483__ = ys__n46101 & new_new_n12356__;
  assign new_new_n29484__ = ys__n46003 & new_new_n12248__;
  assign new_new_n29485__ = ~new_new_n29483__ & ~new_new_n29484__;
  assign new_new_n29486__ = ys__n45905 & new_new_n12245__;
  assign new_new_n29487__ = ys__n45809 & new_new_n12246__;
  assign new_new_n29488__ = ~new_new_n29486__ & ~new_new_n29487__;
  assign new_new_n29489__ = new_new_n29485__ & new_new_n29488__;
  assign new_new_n29490__ = new_new_n26788__ & ~new_new_n29489__;
  assign new_new_n29491__ = ys__n46044 & new_new_n12356__;
  assign new_new_n29492__ = ys__n45946 & new_new_n12248__;
  assign new_new_n29493__ = ~new_new_n29491__ & ~new_new_n29492__;
  assign new_new_n29494__ = ys__n45848 & new_new_n12245__;
  assign new_new_n29495__ = ys__n45727 & new_new_n12246__;
  assign new_new_n29496__ = ~new_new_n29494__ & ~new_new_n29495__;
  assign new_new_n29497__ = new_new_n29493__ & new_new_n29496__;
  assign new_new_n29498__ = new_new_n26807__ & ~new_new_n29497__;
  assign new_new_n29499__ = ~new_new_n29490__ & ~new_new_n29498__;
  assign new_new_n29500__ = new_new_n26882__ & ~new_new_n29499__;
  assign new_new_n29501__ = ~new_new_n26862__ & new_new_n29500__;
  assign new_new_n29502__ = ~new_new_n29482__ & ~new_new_n29501__;
  assign new_new_n29503__ = ~new_new_n14022__ & ~new_new_n29502__;
  assign new_new_n29504__ = ys__n26155 & new_new_n14022__;
  assign ys__n26156 = new_new_n29503__ | new_new_n29504__;
  assign new_new_n29506__ = ys__n26068 & new_new_n26768__;
  assign new_new_n29507__ = ys__n46388 & new_new_n12356__;
  assign new_new_n29508__ = ys__n46564 & new_new_n12248__;
  assign new_new_n29509__ = ~new_new_n29507__ & ~new_new_n29508__;
  assign new_new_n29510__ = ys__n46740 & new_new_n12245__;
  assign new_new_n29511__ = ys__n46916 & new_new_n12246__;
  assign new_new_n29512__ = ~new_new_n29510__ & ~new_new_n29511__;
  assign new_new_n29513__ = new_new_n29509__ & new_new_n29512__;
  assign new_new_n29514__ = new_new_n26779__ & ~new_new_n29513__;
  assign new_new_n29515__ = ys__n46310 & new_new_n12356__;
  assign new_new_n29516__ = ys__n46486 & new_new_n12248__;
  assign new_new_n29517__ = ~new_new_n29515__ & ~new_new_n29516__;
  assign new_new_n29518__ = ys__n46662 & new_new_n12245__;
  assign new_new_n29519__ = ys__n46838 & new_new_n12246__;
  assign new_new_n29520__ = ~new_new_n29518__ & ~new_new_n29519__;
  assign new_new_n29521__ = new_new_n29517__ & new_new_n29520__;
  assign new_new_n29522__ = new_new_n26788__ & ~new_new_n29521__;
  assign new_new_n29523__ = ~new_new_n29514__ & ~new_new_n29522__;
  assign new_new_n29524__ = ys__n46344 & new_new_n12356__;
  assign new_new_n29525__ = ys__n46520 & new_new_n12248__;
  assign new_new_n29526__ = ~new_new_n29524__ & ~new_new_n29525__;
  assign new_new_n29527__ = ys__n46696 & new_new_n12245__;
  assign new_new_n29528__ = ys__n46872 & new_new_n12246__;
  assign new_new_n29529__ = ~new_new_n29527__ & ~new_new_n29528__;
  assign new_new_n29530__ = new_new_n29526__ & new_new_n29529__;
  assign new_new_n29531__ = new_new_n26798__ & ~new_new_n29530__;
  assign new_new_n29532__ = ys__n46421 & new_new_n12356__;
  assign new_new_n29533__ = ys__n46597 & new_new_n12248__;
  assign new_new_n29534__ = ~new_new_n29532__ & ~new_new_n29533__;
  assign new_new_n29535__ = ys__n46773 & new_new_n12245__;
  assign new_new_n29536__ = ys__n46949 & new_new_n12246__;
  assign new_new_n29537__ = ~new_new_n29535__ & ~new_new_n29536__;
  assign new_new_n29538__ = new_new_n29534__ & new_new_n29537__;
  assign new_new_n29539__ = new_new_n26807__ & ~new_new_n29538__;
  assign new_new_n29540__ = ~new_new_n29531__ & ~new_new_n29539__;
  assign new_new_n29541__ = new_new_n29523__ & new_new_n29540__;
  assign new_new_n29542__ = new_new_n26818__ & ~new_new_n29541__;
  assign new_new_n29543__ = ~new_new_n29506__ & ~new_new_n29542__;
  assign new_new_n29544__ = new_new_n26821__ & ~new_new_n29543__;
  assign new_new_n29545__ = ys__n45598 & new_new_n12356__;
  assign new_new_n29546__ = ys__n45434 & new_new_n12248__;
  assign new_new_n29547__ = ~new_new_n29545__ & ~new_new_n29546__;
  assign new_new_n29548__ = ys__n45270 & new_new_n12245__;
  assign new_new_n29549__ = ys__n45074 & new_new_n12246__;
  assign new_new_n29550__ = ~new_new_n29548__ & ~new_new_n29549__;
  assign new_new_n29551__ = new_new_n29547__ & new_new_n29550__;
  assign new_new_n29552__ = new_new_n26807__ & ~new_new_n29551__;
  assign new_new_n29553__ = ys__n45692 & new_new_n12356__;
  assign new_new_n29554__ = ys__n45528 & new_new_n12248__;
  assign new_new_n29555__ = ~new_new_n29553__ & ~new_new_n29554__;
  assign new_new_n29556__ = ys__n45364 & new_new_n12245__;
  assign new_new_n29557__ = ys__n45200 & new_new_n12246__;
  assign new_new_n29558__ = ~new_new_n29556__ & ~new_new_n29557__;
  assign new_new_n29559__ = new_new_n29555__ & new_new_n29558__;
  assign new_new_n29560__ = new_new_n26779__ & ~new_new_n29559__;
  assign new_new_n29561__ = ys__n45631 & new_new_n12356__;
  assign new_new_n29562__ = ys__n45467 & new_new_n12248__;
  assign new_new_n29563__ = ~new_new_n29561__ & ~new_new_n29562__;
  assign new_new_n29564__ = ys__n45303 & new_new_n12245__;
  assign new_new_n29565__ = ys__n45109 & new_new_n12246__;
  assign new_new_n29566__ = ~new_new_n29564__ & ~new_new_n29565__;
  assign new_new_n29567__ = new_new_n29563__ & new_new_n29566__;
  assign new_new_n29568__ = new_new_n26788__ & ~new_new_n29567__;
  assign new_new_n29569__ = ~new_new_n29560__ & ~new_new_n29568__;
  assign new_new_n29570__ = ~new_new_n29552__ & new_new_n29569__;
  assign new_new_n29571__ = new_new_n26859__ & ~new_new_n29570__;
  assign new_new_n29572__ = ~new_new_n29544__ & ~new_new_n29571__;
  assign new_new_n29573__ = new_new_n26862__ & ~new_new_n29572__;
  assign new_new_n29574__ = ys__n46124 & new_new_n12356__;
  assign new_new_n29575__ = ys__n46026 & new_new_n12248__;
  assign new_new_n29576__ = ~new_new_n29574__ & ~new_new_n29575__;
  assign new_new_n29577__ = ys__n45928 & new_new_n12245__;
  assign new_new_n29578__ = ys__n45832 & new_new_n12246__;
  assign new_new_n29579__ = ~new_new_n29577__ & ~new_new_n29578__;
  assign new_new_n29580__ = new_new_n29576__ & new_new_n29579__;
  assign new_new_n29581__ = new_new_n26788__ & ~new_new_n29580__;
  assign new_new_n29582__ = ys__n46090 & new_new_n12356__;
  assign new_new_n29583__ = ys__n45992 & new_new_n12248__;
  assign new_new_n29584__ = ~new_new_n29582__ & ~new_new_n29583__;
  assign new_new_n29585__ = ys__n45894 & new_new_n12245__;
  assign new_new_n29586__ = ys__n45796 & new_new_n12246__;
  assign new_new_n29587__ = ~new_new_n29585__ & ~new_new_n29586__;
  assign new_new_n29588__ = new_new_n29584__ & new_new_n29587__;
  assign new_new_n29589__ = new_new_n26807__ & ~new_new_n29588__;
  assign new_new_n29590__ = ~new_new_n29581__ & ~new_new_n29589__;
  assign new_new_n29591__ = new_new_n26882__ & ~new_new_n29590__;
  assign new_new_n29592__ = ~new_new_n26862__ & new_new_n29591__;
  assign new_new_n29593__ = ~new_new_n29573__ & ~new_new_n29592__;
  assign new_new_n29594__ = ~new_new_n14022__ & ~new_new_n29593__;
  assign new_new_n29595__ = ys__n26157 & new_new_n14022__;
  assign ys__n26158 = new_new_n29594__ | new_new_n29595__;
  assign new_new_n29597__ = ys__n26074 & new_new_n26768__;
  assign new_new_n29598__ = ys__n46392 & new_new_n12356__;
  assign new_new_n29599__ = ys__n46568 & new_new_n12248__;
  assign new_new_n29600__ = ~new_new_n29598__ & ~new_new_n29599__;
  assign new_new_n29601__ = ys__n46744 & new_new_n12245__;
  assign new_new_n29602__ = ys__n46920 & new_new_n12246__;
  assign new_new_n29603__ = ~new_new_n29601__ & ~new_new_n29602__;
  assign new_new_n29604__ = new_new_n29600__ & new_new_n29603__;
  assign new_new_n29605__ = new_new_n26779__ & ~new_new_n29604__;
  assign new_new_n29606__ = ys__n46314 & new_new_n12356__;
  assign new_new_n29607__ = ys__n46490 & new_new_n12248__;
  assign new_new_n29608__ = ~new_new_n29606__ & ~new_new_n29607__;
  assign new_new_n29609__ = ys__n46666 & new_new_n12245__;
  assign new_new_n29610__ = ys__n46842 & new_new_n12246__;
  assign new_new_n29611__ = ~new_new_n29609__ & ~new_new_n29610__;
  assign new_new_n29612__ = new_new_n29608__ & new_new_n29611__;
  assign new_new_n29613__ = new_new_n26788__ & ~new_new_n29612__;
  assign new_new_n29614__ = ~new_new_n29605__ & ~new_new_n29613__;
  assign new_new_n29615__ = ys__n46346 & new_new_n12356__;
  assign new_new_n29616__ = ys__n46522 & new_new_n12248__;
  assign new_new_n29617__ = ~new_new_n29615__ & ~new_new_n29616__;
  assign new_new_n29618__ = ys__n46698 & new_new_n12245__;
  assign new_new_n29619__ = ys__n46874 & new_new_n12246__;
  assign new_new_n29620__ = ~new_new_n29618__ & ~new_new_n29619__;
  assign new_new_n29621__ = new_new_n29617__ & new_new_n29620__;
  assign new_new_n29622__ = new_new_n26798__ & ~new_new_n29621__;
  assign new_new_n29623__ = ys__n46423 & new_new_n12356__;
  assign new_new_n29624__ = ys__n46599 & new_new_n12248__;
  assign new_new_n29625__ = ~new_new_n29623__ & ~new_new_n29624__;
  assign new_new_n29626__ = ys__n46775 & new_new_n12245__;
  assign new_new_n29627__ = ys__n46951 & new_new_n12246__;
  assign new_new_n29628__ = ~new_new_n29626__ & ~new_new_n29627__;
  assign new_new_n29629__ = new_new_n29625__ & new_new_n29628__;
  assign new_new_n29630__ = new_new_n26807__ & ~new_new_n29629__;
  assign new_new_n29631__ = ~new_new_n29622__ & ~new_new_n29630__;
  assign new_new_n29632__ = new_new_n29614__ & new_new_n29631__;
  assign new_new_n29633__ = new_new_n26818__ & ~new_new_n29632__;
  assign new_new_n29634__ = ~new_new_n29597__ & ~new_new_n29633__;
  assign new_new_n29635__ = new_new_n26821__ & ~new_new_n29634__;
  assign new_new_n29636__ = ys__n45602 & new_new_n12356__;
  assign new_new_n29637__ = ys__n45438 & new_new_n12248__;
  assign new_new_n29638__ = ~new_new_n29636__ & ~new_new_n29637__;
  assign new_new_n29639__ = ys__n45274 & new_new_n12245__;
  assign new_new_n29640__ = ys__n45080 & new_new_n12246__;
  assign new_new_n29641__ = ~new_new_n29639__ & ~new_new_n29640__;
  assign new_new_n29642__ = new_new_n29638__ & new_new_n29641__;
  assign new_new_n29643__ = new_new_n26807__ & ~new_new_n29642__;
  assign new_new_n29644__ = ys__n45696 & new_new_n12356__;
  assign new_new_n29645__ = ys__n45532 & new_new_n12248__;
  assign new_new_n29646__ = ~new_new_n29644__ & ~new_new_n29645__;
  assign new_new_n29647__ = ys__n45368 & new_new_n12245__;
  assign new_new_n29648__ = ys__n45206 & new_new_n12246__;
  assign new_new_n29649__ = ~new_new_n29647__ & ~new_new_n29648__;
  assign new_new_n29650__ = new_new_n29646__ & new_new_n29649__;
  assign new_new_n29651__ = new_new_n26779__ & ~new_new_n29650__;
  assign new_new_n29652__ = ys__n45633 & new_new_n12356__;
  assign new_new_n29653__ = ys__n45469 & new_new_n12248__;
  assign new_new_n29654__ = ~new_new_n29652__ & ~new_new_n29653__;
  assign new_new_n29655__ = ys__n45305 & new_new_n12245__;
  assign new_new_n29656__ = ys__n45111 & new_new_n12246__;
  assign new_new_n29657__ = ~new_new_n29655__ & ~new_new_n29656__;
  assign new_new_n29658__ = new_new_n29654__ & new_new_n29657__;
  assign new_new_n29659__ = new_new_n26788__ & ~new_new_n29658__;
  assign new_new_n29660__ = ~new_new_n29651__ & ~new_new_n29659__;
  assign new_new_n29661__ = ~new_new_n29643__ & new_new_n29660__;
  assign new_new_n29662__ = new_new_n26859__ & ~new_new_n29661__;
  assign new_new_n29663__ = ~new_new_n29635__ & ~new_new_n29662__;
  assign new_new_n29664__ = new_new_n26862__ & ~new_new_n29663__;
  assign new_new_n29665__ = ys__n46126 & new_new_n12356__;
  assign new_new_n29666__ = ys__n46028 & new_new_n12248__;
  assign new_new_n29667__ = ~new_new_n29665__ & ~new_new_n29666__;
  assign new_new_n29668__ = ys__n45930 & new_new_n12245__;
  assign new_new_n29669__ = ys__n45834 & new_new_n12246__;
  assign new_new_n29670__ = ~new_new_n29668__ & ~new_new_n29669__;
  assign new_new_n29671__ = new_new_n29667__ & new_new_n29670__;
  assign new_new_n29672__ = new_new_n26788__ & ~new_new_n29671__;
  assign new_new_n29673__ = ys__n46094 & new_new_n12356__;
  assign new_new_n29674__ = ys__n45996 & new_new_n12248__;
  assign new_new_n29675__ = ~new_new_n29673__ & ~new_new_n29674__;
  assign new_new_n29676__ = ys__n45898 & new_new_n12245__;
  assign new_new_n29677__ = ys__n45802 & new_new_n12246__;
  assign new_new_n29678__ = ~new_new_n29676__ & ~new_new_n29677__;
  assign new_new_n29679__ = new_new_n29675__ & new_new_n29678__;
  assign new_new_n29680__ = new_new_n26807__ & ~new_new_n29679__;
  assign new_new_n29681__ = ~new_new_n29672__ & ~new_new_n29680__;
  assign new_new_n29682__ = new_new_n26882__ & ~new_new_n29681__;
  assign new_new_n29683__ = ~new_new_n26862__ & new_new_n29682__;
  assign new_new_n29684__ = ~new_new_n29664__ & ~new_new_n29683__;
  assign new_new_n29685__ = ~new_new_n14022__ & ~new_new_n29684__;
  assign new_new_n29686__ = ys__n26159 & new_new_n14022__;
  assign ys__n26160 = new_new_n29685__ | new_new_n29686__;
  assign new_new_n29688__ = ys__n18833 & ~ys__n18174;
  assign new_new_n29689__ = ys__n26161 & ys__n18174;
  assign new_new_n29690__ = ~new_new_n29688__ & ~new_new_n29689__;
  assign new_new_n29691__ = ys__n18169 & ys__n18170;
  assign new_new_n29692__ = ~new_new_n29690__ & ~new_new_n29691__;
  assign new_new_n29693__ = new_new_n29690__ & new_new_n29691__;
  assign ys__n26220 = new_new_n29692__ | new_new_n29693__;
  assign new_new_n29695__ = ys__n18835 & ~ys__n18174;
  assign new_new_n29696__ = ys__n26162 & ys__n18174;
  assign new_new_n29697__ = ~new_new_n29695__ & ~new_new_n29696__;
  assign new_new_n29698__ = ~new_new_n29691__ & ~new_new_n29697__;
  assign new_new_n29699__ = ~new_new_n29690__ & new_new_n29697__;
  assign new_new_n29700__ = new_new_n29690__ & ~new_new_n29697__;
  assign new_new_n29701__ = ~new_new_n29699__ & ~new_new_n29700__;
  assign new_new_n29702__ = new_new_n29691__ & ~new_new_n29701__;
  assign ys__n26222 = new_new_n29698__ | new_new_n29702__;
  assign new_new_n29704__ = ys__n18837 & ~ys__n18174;
  assign new_new_n29705__ = ys__n26164 & ys__n18174;
  assign new_new_n29706__ = ~new_new_n29704__ & ~new_new_n29705__;
  assign new_new_n29707__ = ~new_new_n29691__ & ~new_new_n29706__;
  assign new_new_n29708__ = ~new_new_n29690__ & ~new_new_n29697__;
  assign new_new_n29709__ = new_new_n29706__ & new_new_n29708__;
  assign new_new_n29710__ = ~new_new_n29706__ & ~new_new_n29708__;
  assign new_new_n29711__ = ~new_new_n29709__ & ~new_new_n29710__;
  assign new_new_n29712__ = new_new_n29691__ & ~new_new_n29711__;
  assign ys__n26224 = new_new_n29707__ | new_new_n29712__;
  assign new_new_n29714__ = ys__n18839 & ~ys__n18174;
  assign new_new_n29715__ = ys__n26166 & ys__n18174;
  assign new_new_n29716__ = ~new_new_n29714__ & ~new_new_n29715__;
  assign new_new_n29717__ = ~new_new_n29691__ & ~new_new_n29716__;
  assign new_new_n29718__ = ~new_new_n29706__ & new_new_n29708__;
  assign new_new_n29719__ = new_new_n29716__ & new_new_n29718__;
  assign new_new_n29720__ = ~new_new_n29716__ & ~new_new_n29718__;
  assign new_new_n29721__ = ~new_new_n29719__ & ~new_new_n29720__;
  assign new_new_n29722__ = new_new_n29691__ & ~new_new_n29721__;
  assign ys__n26226 = new_new_n29717__ | new_new_n29722__;
  assign new_new_n29724__ = ys__n18841 & ~ys__n18174;
  assign new_new_n29725__ = ys__n26168 & ys__n18174;
  assign new_new_n29726__ = ~new_new_n29724__ & ~new_new_n29725__;
  assign new_new_n29727__ = ~new_new_n29691__ & ~new_new_n29726__;
  assign new_new_n29728__ = ~new_new_n29706__ & ~new_new_n29716__;
  assign new_new_n29729__ = new_new_n29708__ & new_new_n29728__;
  assign new_new_n29730__ = new_new_n29726__ & new_new_n29729__;
  assign new_new_n29731__ = ~new_new_n29726__ & ~new_new_n29729__;
  assign new_new_n29732__ = ~new_new_n29730__ & ~new_new_n29731__;
  assign new_new_n29733__ = new_new_n29691__ & ~new_new_n29732__;
  assign ys__n26228 = new_new_n29727__ | new_new_n29733__;
  assign new_new_n29735__ = ys__n18843 & ~ys__n18174;
  assign new_new_n29736__ = ys__n26170 & ys__n18174;
  assign new_new_n29737__ = ~new_new_n29735__ & ~new_new_n29736__;
  assign new_new_n29738__ = ~new_new_n29691__ & ~new_new_n29737__;
  assign new_new_n29739__ = ~new_new_n29726__ & new_new_n29729__;
  assign new_new_n29740__ = new_new_n29737__ & new_new_n29739__;
  assign new_new_n29741__ = ~new_new_n29737__ & ~new_new_n29739__;
  assign new_new_n29742__ = ~new_new_n29740__ & ~new_new_n29741__;
  assign new_new_n29743__ = new_new_n29691__ & ~new_new_n29742__;
  assign ys__n26230 = new_new_n29738__ | new_new_n29743__;
  assign new_new_n29745__ = ys__n18845 & ~ys__n18174;
  assign new_new_n29746__ = ys__n26172 & ys__n18174;
  assign new_new_n29747__ = ~new_new_n29745__ & ~new_new_n29746__;
  assign new_new_n29748__ = ~new_new_n29691__ & ~new_new_n29747__;
  assign new_new_n29749__ = ~new_new_n29726__ & ~new_new_n29737__;
  assign new_new_n29750__ = new_new_n29708__ & new_new_n29749__;
  assign new_new_n29751__ = new_new_n29728__ & new_new_n29750__;
  assign new_new_n29752__ = new_new_n29747__ & new_new_n29751__;
  assign new_new_n29753__ = ~new_new_n29747__ & ~new_new_n29751__;
  assign new_new_n29754__ = ~new_new_n29752__ & ~new_new_n29753__;
  assign new_new_n29755__ = new_new_n29691__ & ~new_new_n29754__;
  assign ys__n26232 = new_new_n29748__ | new_new_n29755__;
  assign new_new_n29757__ = ys__n18847 & ~ys__n18174;
  assign new_new_n29758__ = ys__n26174 & ys__n18174;
  assign new_new_n29759__ = ~new_new_n29757__ & ~new_new_n29758__;
  assign new_new_n29760__ = ~new_new_n29691__ & ~new_new_n29759__;
  assign new_new_n29761__ = ~new_new_n29747__ & new_new_n29751__;
  assign new_new_n29762__ = new_new_n29759__ & new_new_n29761__;
  assign new_new_n29763__ = ~new_new_n29759__ & ~new_new_n29761__;
  assign new_new_n29764__ = ~new_new_n29762__ & ~new_new_n29763__;
  assign new_new_n29765__ = new_new_n29691__ & ~new_new_n29764__;
  assign ys__n26234 = new_new_n29760__ | new_new_n29765__;
  assign new_new_n29767__ = ys__n18849 & ~ys__n18174;
  assign new_new_n29768__ = ys__n26176 & ys__n18174;
  assign new_new_n29769__ = ~new_new_n29767__ & ~new_new_n29768__;
  assign new_new_n29770__ = ~new_new_n29691__ & ~new_new_n29769__;
  assign new_new_n29771__ = ~new_new_n29747__ & ~new_new_n29759__;
  assign new_new_n29772__ = new_new_n29751__ & new_new_n29771__;
  assign new_new_n29773__ = new_new_n29769__ & new_new_n29772__;
  assign new_new_n29774__ = ~new_new_n29769__ & ~new_new_n29772__;
  assign new_new_n29775__ = ~new_new_n29773__ & ~new_new_n29774__;
  assign new_new_n29776__ = new_new_n29691__ & ~new_new_n29775__;
  assign ys__n26236 = new_new_n29770__ | new_new_n29776__;
  assign new_new_n29778__ = ys__n18851 & ~ys__n18174;
  assign new_new_n29779__ = ys__n26178 & ys__n18174;
  assign new_new_n29780__ = ~new_new_n29778__ & ~new_new_n29779__;
  assign new_new_n29781__ = ~new_new_n29691__ & ~new_new_n29780__;
  assign new_new_n29782__ = ~new_new_n29769__ & new_new_n29772__;
  assign new_new_n29783__ = new_new_n29780__ & new_new_n29782__;
  assign new_new_n29784__ = ~new_new_n29780__ & ~new_new_n29782__;
  assign new_new_n29785__ = ~new_new_n29783__ & ~new_new_n29784__;
  assign new_new_n29786__ = new_new_n29691__ & ~new_new_n29785__;
  assign ys__n26238 = new_new_n29781__ | new_new_n29786__;
  assign new_new_n29788__ = ys__n18853 & ~ys__n18174;
  assign new_new_n29789__ = ys__n26180 & ys__n18174;
  assign new_new_n29790__ = ~new_new_n29788__ & ~new_new_n29789__;
  assign new_new_n29791__ = ~new_new_n29691__ & ~new_new_n29790__;
  assign new_new_n29792__ = ~new_new_n29769__ & ~new_new_n29780__;
  assign new_new_n29793__ = new_new_n29771__ & new_new_n29792__;
  assign new_new_n29794__ = new_new_n29751__ & new_new_n29793__;
  assign new_new_n29795__ = new_new_n29790__ & new_new_n29794__;
  assign new_new_n29796__ = ~new_new_n29790__ & ~new_new_n29794__;
  assign new_new_n29797__ = ~new_new_n29795__ & ~new_new_n29796__;
  assign new_new_n29798__ = new_new_n29691__ & ~new_new_n29797__;
  assign ys__n26240 = new_new_n29791__ | new_new_n29798__;
  assign new_new_n29800__ = ys__n18855 & ~ys__n18174;
  assign new_new_n29801__ = ys__n26182 & ys__n18174;
  assign new_new_n29802__ = ~new_new_n29800__ & ~new_new_n29801__;
  assign new_new_n29803__ = ~new_new_n29691__ & ~new_new_n29802__;
  assign new_new_n29804__ = ~new_new_n29790__ & new_new_n29794__;
  assign new_new_n29805__ = new_new_n29802__ & new_new_n29804__;
  assign new_new_n29806__ = ~new_new_n29802__ & ~new_new_n29804__;
  assign new_new_n29807__ = ~new_new_n29805__ & ~new_new_n29806__;
  assign new_new_n29808__ = new_new_n29691__ & ~new_new_n29807__;
  assign ys__n26242 = new_new_n29803__ | new_new_n29808__;
  assign new_new_n29810__ = ys__n18857 & ~ys__n18174;
  assign new_new_n29811__ = ys__n26184 & ys__n18174;
  assign new_new_n29812__ = ~new_new_n29810__ & ~new_new_n29811__;
  assign new_new_n29813__ = ~new_new_n29691__ & ~new_new_n29812__;
  assign new_new_n29814__ = ~new_new_n29790__ & ~new_new_n29802__;
  assign new_new_n29815__ = new_new_n29794__ & new_new_n29814__;
  assign new_new_n29816__ = new_new_n29812__ & new_new_n29815__;
  assign new_new_n29817__ = ~new_new_n29812__ & ~new_new_n29815__;
  assign new_new_n29818__ = ~new_new_n29816__ & ~new_new_n29817__;
  assign new_new_n29819__ = new_new_n29691__ & ~new_new_n29818__;
  assign ys__n26244 = new_new_n29813__ | new_new_n29819__;
  assign new_new_n29821__ = ys__n18859 & ~ys__n18174;
  assign new_new_n29822__ = ys__n26186 & ys__n18174;
  assign new_new_n29823__ = ~new_new_n29821__ & ~new_new_n29822__;
  assign new_new_n29824__ = ~new_new_n29691__ & ~new_new_n29823__;
  assign new_new_n29825__ = ~new_new_n29812__ & new_new_n29815__;
  assign new_new_n29826__ = new_new_n29823__ & new_new_n29825__;
  assign new_new_n29827__ = ~new_new_n29823__ & ~new_new_n29825__;
  assign new_new_n29828__ = ~new_new_n29826__ & ~new_new_n29827__;
  assign new_new_n29829__ = new_new_n29691__ & ~new_new_n29828__;
  assign ys__n26246 = new_new_n29824__ | new_new_n29829__;
  assign new_new_n29831__ = ys__n18861 & ~ys__n18174;
  assign new_new_n29832__ = ys__n26188 & ys__n18174;
  assign new_new_n29833__ = ~new_new_n29831__ & ~new_new_n29832__;
  assign new_new_n29834__ = ~new_new_n29691__ & ~new_new_n29833__;
  assign new_new_n29835__ = ~new_new_n29812__ & ~new_new_n29823__;
  assign new_new_n29836__ = new_new_n29814__ & new_new_n29835__;
  assign new_new_n29837__ = new_new_n29793__ & new_new_n29836__;
  assign new_new_n29838__ = new_new_n29751__ & new_new_n29837__;
  assign new_new_n29839__ = new_new_n29833__ & new_new_n29838__;
  assign new_new_n29840__ = ~new_new_n29833__ & ~new_new_n29838__;
  assign new_new_n29841__ = ~new_new_n29839__ & ~new_new_n29840__;
  assign new_new_n29842__ = new_new_n29691__ & ~new_new_n29841__;
  assign ys__n26248 = new_new_n29834__ | new_new_n29842__;
  assign new_new_n29844__ = ys__n18863 & ~ys__n18174;
  assign new_new_n29845__ = ys__n26190 & ys__n18174;
  assign new_new_n29846__ = ~new_new_n29844__ & ~new_new_n29845__;
  assign new_new_n29847__ = ~new_new_n29691__ & ~new_new_n29846__;
  assign new_new_n29848__ = ~new_new_n29833__ & new_new_n29838__;
  assign new_new_n29849__ = new_new_n29846__ & new_new_n29848__;
  assign new_new_n29850__ = ~new_new_n29846__ & ~new_new_n29848__;
  assign new_new_n29851__ = ~new_new_n29849__ & ~new_new_n29850__;
  assign new_new_n29852__ = new_new_n29691__ & ~new_new_n29851__;
  assign ys__n26250 = new_new_n29847__ | new_new_n29852__;
  assign new_new_n29854__ = ys__n18865 & ~ys__n18174;
  assign new_new_n29855__ = ys__n26192 & ys__n18174;
  assign new_new_n29856__ = ~new_new_n29854__ & ~new_new_n29855__;
  assign new_new_n29857__ = ~new_new_n29691__ & ~new_new_n29856__;
  assign new_new_n29858__ = ~new_new_n29833__ & ~new_new_n29846__;
  assign new_new_n29859__ = new_new_n29838__ & new_new_n29858__;
  assign new_new_n29860__ = new_new_n29856__ & new_new_n29859__;
  assign new_new_n29861__ = ~new_new_n29856__ & ~new_new_n29859__;
  assign new_new_n29862__ = ~new_new_n29860__ & ~new_new_n29861__;
  assign new_new_n29863__ = new_new_n29691__ & ~new_new_n29862__;
  assign ys__n26252 = new_new_n29857__ | new_new_n29863__;
  assign new_new_n29865__ = ys__n18867 & ~ys__n18174;
  assign new_new_n29866__ = ys__n26194 & ys__n18174;
  assign new_new_n29867__ = ~new_new_n29865__ & ~new_new_n29866__;
  assign new_new_n29868__ = ~new_new_n29691__ & ~new_new_n29867__;
  assign new_new_n29869__ = ~new_new_n29856__ & new_new_n29859__;
  assign new_new_n29870__ = new_new_n29867__ & new_new_n29869__;
  assign new_new_n29871__ = ~new_new_n29867__ & ~new_new_n29869__;
  assign new_new_n29872__ = ~new_new_n29870__ & ~new_new_n29871__;
  assign new_new_n29873__ = new_new_n29691__ & ~new_new_n29872__;
  assign ys__n26254 = new_new_n29868__ | new_new_n29873__;
  assign new_new_n29875__ = ys__n18869 & ~ys__n18174;
  assign new_new_n29876__ = ys__n26196 & ys__n18174;
  assign new_new_n29877__ = ~new_new_n29875__ & ~new_new_n29876__;
  assign new_new_n29878__ = ~new_new_n29691__ & ~new_new_n29877__;
  assign new_new_n29879__ = ~new_new_n29856__ & ~new_new_n29867__;
  assign new_new_n29880__ = new_new_n29858__ & new_new_n29879__;
  assign new_new_n29881__ = new_new_n29838__ & new_new_n29880__;
  assign new_new_n29882__ = new_new_n29877__ & new_new_n29881__;
  assign new_new_n29883__ = ~new_new_n29877__ & ~new_new_n29881__;
  assign new_new_n29884__ = ~new_new_n29882__ & ~new_new_n29883__;
  assign new_new_n29885__ = new_new_n29691__ & ~new_new_n29884__;
  assign ys__n26256 = new_new_n29878__ | new_new_n29885__;
  assign new_new_n29887__ = ys__n18871 & ~ys__n18174;
  assign new_new_n29888__ = ys__n26198 & ys__n18174;
  assign new_new_n29889__ = ~new_new_n29887__ & ~new_new_n29888__;
  assign new_new_n29890__ = ~new_new_n29691__ & ~new_new_n29889__;
  assign new_new_n29891__ = ~new_new_n29877__ & new_new_n29881__;
  assign new_new_n29892__ = new_new_n29889__ & new_new_n29891__;
  assign new_new_n29893__ = ~new_new_n29889__ & ~new_new_n29891__;
  assign new_new_n29894__ = ~new_new_n29892__ & ~new_new_n29893__;
  assign new_new_n29895__ = new_new_n29691__ & ~new_new_n29894__;
  assign ys__n26258 = new_new_n29890__ | new_new_n29895__;
  assign new_new_n29897__ = ys__n18873 & ~ys__n18174;
  assign new_new_n29898__ = ys__n26200 & ys__n18174;
  assign new_new_n29899__ = ~new_new_n29897__ & ~new_new_n29898__;
  assign new_new_n29900__ = ~new_new_n29691__ & ~new_new_n29899__;
  assign new_new_n29901__ = ~new_new_n29877__ & ~new_new_n29889__;
  assign new_new_n29902__ = new_new_n29881__ & new_new_n29901__;
  assign new_new_n29903__ = new_new_n29899__ & new_new_n29902__;
  assign new_new_n29904__ = ~new_new_n29899__ & ~new_new_n29902__;
  assign new_new_n29905__ = ~new_new_n29903__ & ~new_new_n29904__;
  assign new_new_n29906__ = new_new_n29691__ & ~new_new_n29905__;
  assign ys__n26260 = new_new_n29900__ | new_new_n29906__;
  assign new_new_n29908__ = ys__n18875 & ~ys__n18174;
  assign new_new_n29909__ = ys__n26202 & ys__n18174;
  assign new_new_n29910__ = ~new_new_n29908__ & ~new_new_n29909__;
  assign new_new_n29911__ = ~new_new_n29691__ & ~new_new_n29910__;
  assign new_new_n29912__ = ~new_new_n29899__ & new_new_n29902__;
  assign new_new_n29913__ = new_new_n29910__ & new_new_n29912__;
  assign new_new_n29914__ = ~new_new_n29910__ & ~new_new_n29912__;
  assign new_new_n29915__ = ~new_new_n29913__ & ~new_new_n29914__;
  assign new_new_n29916__ = new_new_n29691__ & ~new_new_n29915__;
  assign ys__n26262 = new_new_n29911__ | new_new_n29916__;
  assign new_new_n29918__ = ys__n18877 & ~ys__n18174;
  assign new_new_n29919__ = ys__n26204 & ys__n18174;
  assign new_new_n29920__ = ~new_new_n29918__ & ~new_new_n29919__;
  assign new_new_n29921__ = ~new_new_n29691__ & ~new_new_n29920__;
  assign new_new_n29922__ = ~new_new_n29899__ & ~new_new_n29910__;
  assign new_new_n29923__ = new_new_n29901__ & new_new_n29922__;
  assign new_new_n29924__ = new_new_n29880__ & new_new_n29923__;
  assign new_new_n29925__ = new_new_n29838__ & new_new_n29924__;
  assign new_new_n29926__ = new_new_n29920__ & new_new_n29925__;
  assign new_new_n29927__ = ~new_new_n29920__ & ~new_new_n29925__;
  assign new_new_n29928__ = ~new_new_n29926__ & ~new_new_n29927__;
  assign new_new_n29929__ = new_new_n29691__ & ~new_new_n29928__;
  assign ys__n26264 = new_new_n29921__ | new_new_n29929__;
  assign new_new_n29931__ = ys__n18879 & ~ys__n18174;
  assign new_new_n29932__ = ys__n26206 & ys__n18174;
  assign new_new_n29933__ = ~new_new_n29931__ & ~new_new_n29932__;
  assign new_new_n29934__ = ~new_new_n29691__ & ~new_new_n29933__;
  assign new_new_n29935__ = ~new_new_n29920__ & new_new_n29925__;
  assign new_new_n29936__ = new_new_n29933__ & new_new_n29935__;
  assign new_new_n29937__ = ~new_new_n29933__ & ~new_new_n29935__;
  assign new_new_n29938__ = ~new_new_n29936__ & ~new_new_n29937__;
  assign new_new_n29939__ = new_new_n29691__ & ~new_new_n29938__;
  assign ys__n26266 = new_new_n29934__ | new_new_n29939__;
  assign new_new_n29941__ = ys__n18881 & ~ys__n18174;
  assign new_new_n29942__ = ys__n26208 & ys__n18174;
  assign new_new_n29943__ = ~new_new_n29941__ & ~new_new_n29942__;
  assign new_new_n29944__ = ~new_new_n29691__ & ~new_new_n29943__;
  assign new_new_n29945__ = ~new_new_n29920__ & ~new_new_n29933__;
  assign new_new_n29946__ = new_new_n29925__ & new_new_n29945__;
  assign new_new_n29947__ = new_new_n29943__ & new_new_n29946__;
  assign new_new_n29948__ = ~new_new_n29943__ & ~new_new_n29946__;
  assign new_new_n29949__ = ~new_new_n29947__ & ~new_new_n29948__;
  assign new_new_n29950__ = new_new_n29691__ & ~new_new_n29949__;
  assign ys__n26268 = new_new_n29944__ | new_new_n29950__;
  assign new_new_n29952__ = ys__n18883 & ~ys__n18174;
  assign new_new_n29953__ = ys__n26210 & ys__n18174;
  assign new_new_n29954__ = ~new_new_n29952__ & ~new_new_n29953__;
  assign new_new_n29955__ = ~new_new_n29691__ & ~new_new_n29954__;
  assign new_new_n29956__ = ~new_new_n29943__ & new_new_n29946__;
  assign new_new_n29957__ = new_new_n29954__ & new_new_n29956__;
  assign new_new_n29958__ = ~new_new_n29954__ & ~new_new_n29956__;
  assign new_new_n29959__ = ~new_new_n29957__ & ~new_new_n29958__;
  assign new_new_n29960__ = new_new_n29691__ & ~new_new_n29959__;
  assign ys__n26270 = new_new_n29955__ | new_new_n29960__;
  assign new_new_n29962__ = ys__n18885 & ~ys__n18174;
  assign new_new_n29963__ = ys__n26212 & ys__n18174;
  assign new_new_n29964__ = ~new_new_n29962__ & ~new_new_n29963__;
  assign new_new_n29965__ = ~new_new_n29691__ & ~new_new_n29964__;
  assign new_new_n29966__ = ~new_new_n29943__ & ~new_new_n29954__;
  assign new_new_n29967__ = new_new_n29945__ & new_new_n29966__;
  assign new_new_n29968__ = new_new_n29925__ & new_new_n29967__;
  assign new_new_n29969__ = new_new_n29964__ & new_new_n29968__;
  assign new_new_n29970__ = ~new_new_n29964__ & ~new_new_n29968__;
  assign new_new_n29971__ = ~new_new_n29969__ & ~new_new_n29970__;
  assign new_new_n29972__ = new_new_n29691__ & ~new_new_n29971__;
  assign ys__n26272 = new_new_n29965__ | new_new_n29972__;
  assign new_new_n29974__ = ys__n18887 & ~ys__n18174;
  assign new_new_n29975__ = ys__n26214 & ys__n18174;
  assign new_new_n29976__ = ~new_new_n29974__ & ~new_new_n29975__;
  assign new_new_n29977__ = ~new_new_n29691__ & ~new_new_n29976__;
  assign new_new_n29978__ = ~new_new_n29964__ & new_new_n29968__;
  assign new_new_n29979__ = new_new_n29976__ & new_new_n29978__;
  assign new_new_n29980__ = ~new_new_n29976__ & ~new_new_n29978__;
  assign new_new_n29981__ = ~new_new_n29979__ & ~new_new_n29980__;
  assign new_new_n29982__ = new_new_n29691__ & ~new_new_n29981__;
  assign ys__n26274 = new_new_n29977__ | new_new_n29982__;
  assign new_new_n29984__ = ys__n18889 & ~ys__n18174;
  assign new_new_n29985__ = ys__n26216 & ys__n18174;
  assign new_new_n29986__ = ~new_new_n29984__ & ~new_new_n29985__;
  assign new_new_n29987__ = ~new_new_n29691__ & ~new_new_n29986__;
  assign new_new_n29988__ = ~new_new_n29964__ & ~new_new_n29976__;
  assign new_new_n29989__ = new_new_n29968__ & new_new_n29988__;
  assign new_new_n29990__ = new_new_n29986__ & new_new_n29989__;
  assign new_new_n29991__ = ~new_new_n29986__ & ~new_new_n29989__;
  assign new_new_n29992__ = ~new_new_n29990__ & ~new_new_n29991__;
  assign new_new_n29993__ = new_new_n29691__ & ~new_new_n29992__;
  assign ys__n26276 = new_new_n29987__ | new_new_n29993__;
  assign new_new_n29995__ = ys__n18891 & ~ys__n18174;
  assign new_new_n29996__ = ys__n26218 & ys__n18174;
  assign new_new_n29997__ = ~new_new_n29995__ & ~new_new_n29996__;
  assign new_new_n29998__ = ~new_new_n29691__ & ~new_new_n29997__;
  assign new_new_n29999__ = ~new_new_n29986__ & new_new_n29989__;
  assign new_new_n30000__ = new_new_n29997__ & new_new_n29999__;
  assign new_new_n30001__ = ~new_new_n29997__ & ~new_new_n29999__;
  assign new_new_n30002__ = ~new_new_n30000__ & ~new_new_n30001__;
  assign new_new_n30003__ = new_new_n29691__ & ~new_new_n30002__;
  assign ys__n26278 = new_new_n29998__ | new_new_n30003__;
  assign new_new_n30005__ = ~ys__n26428 & ~ys__n30941;
  assign ys__n26282 = ys__n18169 & new_new_n30005__;
  assign new_new_n30007__ = ys__n26431 & ~ys__n30941;
  assign ys__n26284 = ys__n18169 & new_new_n30007__;
  assign ys__n26286 = ys__n26285 & ys__n18169;
  assign new_new_n30010__ = ys__n26460 & ~ys__n30941;
  assign ys__n26288 = ys__n18169 & new_new_n30010__;
  assign new_new_n30012__ = ys__n336 & ys__n776;
  assign ys__n26573 = new_new_n26668__ & new_new_n30012__;
  assign new_new_n30014__ = ys__n26569 & ~ys__n26573;
  assign new_new_n30015__ = ~ys__n18169 & new_new_n30014__;
  assign new_new_n30016__ = ~ys__n26478 & ys__n26493;
  assign new_new_n30017__ = ys__n35031 & new_new_n30016__;
  assign new_new_n30018__ = ys__n18169 & new_new_n30017__;
  assign ys__n26291 = new_new_n30015__ | new_new_n30018__;
  assign ys__n26293 = ~ys__n18466 & ys__n18178;
  assign ys__n26294 = ys__n18463 & ys__n18178;
  assign new_new_n30022__ = ~ys__n18208 & ~ys__n26565;
  assign new_new_n30023__ = ys__n26565 & ys__n30962;
  assign ys__n26566 = new_new_n30022__ | new_new_n30023__;
  assign new_new_n30025__ = ~ys__n778 & ys__n25980;
  assign new_new_n30026__ = new_new_n16728__ & ~new_new_n26678__;
  assign new_new_n30027__ = ys__n25980 & new_new_n30026__;
  assign new_new_n30028__ = ~ys__n18173 & ys__n18448;
  assign new_new_n30029__ = ys__n18173 & ys__n30877;
  assign new_new_n30030__ = ~new_new_n30028__ & ~new_new_n30029__;
  assign new_new_n30031__ = ~new_new_n16728__ & ~new_new_n30030__;
  assign new_new_n30032__ = ~new_new_n30026__ & new_new_n30031__;
  assign new_new_n30033__ = ~new_new_n30027__ & ~new_new_n30032__;
  assign new_new_n30034__ = ys__n778 & ~new_new_n30033__;
  assign new_new_n30035__ = ~new_new_n30025__ & ~new_new_n30034__;
  assign new_new_n30036__ = ~ys__n602 & ~new_new_n30035__;
  assign new_new_n30037__ = ~new_new_n16712__ & new_new_n26679__;
  assign new_new_n30038__ = ~new_new_n30035__ & new_new_n30037__;
  assign new_new_n30039__ = ys__n25984 & new_new_n16712__;
  assign new_new_n30040__ = ys__n25984 & ~new_new_n26679__;
  assign new_new_n30041__ = ~new_new_n30039__ & ~new_new_n30040__;
  assign new_new_n30042__ = ~new_new_n30037__ & ~new_new_n30041__;
  assign new_new_n30043__ = ~new_new_n30038__ & ~new_new_n30042__;
  assign new_new_n30044__ = ys__n602 & ~new_new_n30043__;
  assign ys__n26607 = new_new_n30036__ | new_new_n30044__;
  assign new_new_n30046__ = ~ys__n778 & ys__n25984;
  assign new_new_n30047__ = ys__n25984 & new_new_n30026__;
  assign new_new_n30048__ = ~ys__n18173 & ys__n18451;
  assign new_new_n30049__ = ys__n18173 & ys__n30879;
  assign new_new_n30050__ = ~new_new_n30048__ & ~new_new_n30049__;
  assign new_new_n30051__ = ~new_new_n16728__ & ~new_new_n30050__;
  assign new_new_n30052__ = ~new_new_n30026__ & new_new_n30051__;
  assign new_new_n30053__ = ~new_new_n30047__ & ~new_new_n30052__;
  assign new_new_n30054__ = ys__n778 & ~new_new_n30053__;
  assign new_new_n30055__ = ~new_new_n30046__ & ~new_new_n30054__;
  assign new_new_n30056__ = ~ys__n602 & ~new_new_n30055__;
  assign new_new_n30057__ = new_new_n30037__ & ~new_new_n30055__;
  assign new_new_n30058__ = ys__n25987 & new_new_n16712__;
  assign new_new_n30059__ = ys__n25987 & ~new_new_n26679__;
  assign new_new_n30060__ = ~new_new_n30058__ & ~new_new_n30059__;
  assign new_new_n30061__ = ~new_new_n30037__ & ~new_new_n30060__;
  assign new_new_n30062__ = ~new_new_n30057__ & ~new_new_n30061__;
  assign new_new_n30063__ = ys__n602 & ~new_new_n30062__;
  assign ys__n26609 = new_new_n30056__ | new_new_n30063__;
  assign new_new_n30065__ = ~ys__n778 & ys__n25987;
  assign new_new_n30066__ = ys__n25987 & new_new_n30026__;
  assign new_new_n30067__ = ~ys__n18173 & ys__n18454;
  assign new_new_n30068__ = ys__n18173 & ys__n30881;
  assign new_new_n30069__ = ~new_new_n30067__ & ~new_new_n30068__;
  assign new_new_n30070__ = ~new_new_n16728__ & ~new_new_n30069__;
  assign new_new_n30071__ = ~new_new_n30026__ & new_new_n30070__;
  assign new_new_n30072__ = ~new_new_n30066__ & ~new_new_n30071__;
  assign new_new_n30073__ = ys__n778 & ~new_new_n30072__;
  assign new_new_n30074__ = ~new_new_n30065__ & ~new_new_n30073__;
  assign new_new_n30075__ = ~ys__n602 & ~new_new_n30074__;
  assign new_new_n30076__ = new_new_n30037__ & ~new_new_n30074__;
  assign new_new_n30077__ = ys__n25990 & new_new_n16712__;
  assign new_new_n30078__ = ys__n25990 & ~new_new_n26679__;
  assign new_new_n30079__ = ~new_new_n30077__ & ~new_new_n30078__;
  assign new_new_n30080__ = ~new_new_n30037__ & ~new_new_n30079__;
  assign new_new_n30081__ = ~new_new_n30076__ & ~new_new_n30080__;
  assign new_new_n30082__ = ys__n602 & ~new_new_n30081__;
  assign ys__n26611 = new_new_n30075__ | new_new_n30082__;
  assign new_new_n30084__ = ~ys__n778 & ys__n25990;
  assign new_new_n30085__ = ys__n25990 & new_new_n30026__;
  assign new_new_n30086__ = ~ys__n18173 & ys__n18457;
  assign new_new_n30087__ = ys__n18173 & ys__n30883;
  assign new_new_n30088__ = ~new_new_n30086__ & ~new_new_n30087__;
  assign new_new_n30089__ = ~new_new_n16728__ & ~new_new_n30088__;
  assign new_new_n30090__ = ~new_new_n30026__ & new_new_n30089__;
  assign new_new_n30091__ = ~new_new_n30085__ & ~new_new_n30090__;
  assign new_new_n30092__ = ys__n778 & ~new_new_n30091__;
  assign new_new_n30093__ = ~new_new_n30084__ & ~new_new_n30092__;
  assign new_new_n30094__ = ~ys__n602 & ~new_new_n30093__;
  assign new_new_n30095__ = new_new_n30037__ & ~new_new_n30093__;
  assign new_new_n30096__ = ys__n25993 & new_new_n16712__;
  assign new_new_n30097__ = ys__n25993 & ~new_new_n26679__;
  assign new_new_n30098__ = ~new_new_n30096__ & ~new_new_n30097__;
  assign new_new_n30099__ = ~new_new_n30037__ & ~new_new_n30098__;
  assign new_new_n30100__ = ~new_new_n30095__ & ~new_new_n30099__;
  assign new_new_n30101__ = ys__n602 & ~new_new_n30100__;
  assign ys__n26613 = new_new_n30094__ | new_new_n30101__;
  assign new_new_n30103__ = ~ys__n778 & ys__n25993;
  assign new_new_n30104__ = ys__n25993 & new_new_n30026__;
  assign new_new_n30105__ = ~ys__n18173 & ys__n18460;
  assign new_new_n30106__ = ys__n18173 & ys__n30885;
  assign new_new_n30107__ = ~new_new_n30105__ & ~new_new_n30106__;
  assign new_new_n30108__ = ~new_new_n16728__ & ~new_new_n30107__;
  assign new_new_n30109__ = ~new_new_n30026__ & new_new_n30108__;
  assign new_new_n30110__ = ~new_new_n30104__ & ~new_new_n30109__;
  assign new_new_n30111__ = ys__n778 & ~new_new_n30110__;
  assign new_new_n30112__ = ~new_new_n30103__ & ~new_new_n30111__;
  assign new_new_n30113__ = ~ys__n602 & ~new_new_n30112__;
  assign new_new_n30114__ = new_new_n30037__ & ~new_new_n30112__;
  assign new_new_n30115__ = ys__n25996 & new_new_n16712__;
  assign new_new_n30116__ = ys__n25996 & ~new_new_n26679__;
  assign new_new_n30117__ = ~new_new_n30115__ & ~new_new_n30116__;
  assign new_new_n30118__ = ~new_new_n30037__ & ~new_new_n30117__;
  assign new_new_n30119__ = ~new_new_n30114__ & ~new_new_n30118__;
  assign new_new_n30120__ = ys__n602 & ~new_new_n30119__;
  assign ys__n26615 = new_new_n30113__ | new_new_n30120__;
  assign new_new_n30122__ = ~ys__n778 & ys__n25996;
  assign new_new_n30123__ = ys__n25996 & new_new_n30026__;
  assign new_new_n30124__ = ~ys__n18173 & ys__n18463;
  assign new_new_n30125__ = ys__n18173 & ys__n30887;
  assign new_new_n30126__ = ~new_new_n30124__ & ~new_new_n30125__;
  assign new_new_n30127__ = ~new_new_n16728__ & ~new_new_n30126__;
  assign new_new_n30128__ = ~new_new_n30026__ & new_new_n30127__;
  assign new_new_n30129__ = ~new_new_n30123__ & ~new_new_n30128__;
  assign new_new_n30130__ = ys__n778 & ~new_new_n30129__;
  assign new_new_n30131__ = ~new_new_n30122__ & ~new_new_n30130__;
  assign new_new_n30132__ = ~ys__n602 & ~new_new_n30131__;
  assign new_new_n30133__ = new_new_n30037__ & ~new_new_n30131__;
  assign new_new_n30134__ = ys__n25999 & new_new_n16712__;
  assign new_new_n30135__ = ys__n25999 & ~new_new_n26679__;
  assign new_new_n30136__ = ~new_new_n30134__ & ~new_new_n30135__;
  assign new_new_n30137__ = ~new_new_n30037__ & ~new_new_n30136__;
  assign new_new_n30138__ = ~new_new_n30133__ & ~new_new_n30137__;
  assign new_new_n30139__ = ys__n602 & ~new_new_n30138__;
  assign ys__n26617 = new_new_n30132__ | new_new_n30139__;
  assign new_new_n30141__ = ~ys__n778 & ys__n25999;
  assign new_new_n30142__ = ys__n25999 & new_new_n30026__;
  assign new_new_n30143__ = ~ys__n18173 & ys__n18466;
  assign new_new_n30144__ = ys__n18173 & ys__n30889;
  assign new_new_n30145__ = ~new_new_n30143__ & ~new_new_n30144__;
  assign new_new_n30146__ = ~new_new_n16728__ & ~new_new_n30145__;
  assign new_new_n30147__ = ~new_new_n30026__ & new_new_n30146__;
  assign new_new_n30148__ = ~new_new_n30142__ & ~new_new_n30147__;
  assign new_new_n30149__ = ys__n778 & ~new_new_n30148__;
  assign new_new_n30150__ = ~new_new_n30141__ & ~new_new_n30149__;
  assign new_new_n30151__ = ~ys__n602 & ~new_new_n30150__;
  assign new_new_n30152__ = new_new_n30037__ & ~new_new_n30150__;
  assign new_new_n30153__ = ys__n26002 & new_new_n16712__;
  assign new_new_n30154__ = ys__n26002 & ~new_new_n26679__;
  assign new_new_n30155__ = ~new_new_n30153__ & ~new_new_n30154__;
  assign new_new_n30156__ = ~new_new_n30037__ & ~new_new_n30155__;
  assign new_new_n30157__ = ~new_new_n30152__ & ~new_new_n30156__;
  assign new_new_n30158__ = ys__n602 & ~new_new_n30157__;
  assign ys__n26619 = new_new_n30151__ | new_new_n30158__;
  assign new_new_n30160__ = ~ys__n778 & ys__n26002;
  assign new_new_n30161__ = ys__n26002 & new_new_n30026__;
  assign new_new_n30162__ = ~ys__n18173 & ys__n18469;
  assign new_new_n30163__ = ys__n18173 & ys__n30891;
  assign new_new_n30164__ = ~new_new_n30162__ & ~new_new_n30163__;
  assign new_new_n30165__ = ~new_new_n16728__ & ~new_new_n30164__;
  assign new_new_n30166__ = ~new_new_n30026__ & new_new_n30165__;
  assign new_new_n30167__ = ~new_new_n30161__ & ~new_new_n30166__;
  assign new_new_n30168__ = ys__n778 & ~new_new_n30167__;
  assign new_new_n30169__ = ~new_new_n30160__ & ~new_new_n30168__;
  assign new_new_n30170__ = ~ys__n602 & ~new_new_n30169__;
  assign new_new_n30171__ = new_new_n30037__ & ~new_new_n30169__;
  assign new_new_n30172__ = ys__n26005 & new_new_n16712__;
  assign new_new_n30173__ = ys__n26005 & ~new_new_n26679__;
  assign new_new_n30174__ = ~new_new_n30172__ & ~new_new_n30173__;
  assign new_new_n30175__ = ~new_new_n30037__ & ~new_new_n30174__;
  assign new_new_n30176__ = ~new_new_n30171__ & ~new_new_n30175__;
  assign new_new_n30177__ = ys__n602 & ~new_new_n30176__;
  assign ys__n26621 = new_new_n30170__ | new_new_n30177__;
  assign new_new_n30179__ = ~ys__n778 & ys__n26005;
  assign new_new_n30180__ = ys__n26005 & new_new_n30026__;
  assign new_new_n30181__ = ys__n35059 & new_new_n26678__;
  assign new_new_n30182__ = ~ys__n18173 & ys__n18472;
  assign new_new_n30183__ = ys__n18173 & ys__n30893;
  assign new_new_n30184__ = ~new_new_n30182__ & ~new_new_n30183__;
  assign new_new_n30185__ = ~new_new_n16728__ & ~new_new_n30184__;
  assign new_new_n30186__ = ~new_new_n30181__ & ~new_new_n30185__;
  assign new_new_n30187__ = ~new_new_n30026__ & ~new_new_n30186__;
  assign new_new_n30188__ = ~new_new_n30180__ & ~new_new_n30187__;
  assign new_new_n30189__ = ys__n778 & ~new_new_n30188__;
  assign new_new_n30190__ = ~new_new_n30179__ & ~new_new_n30189__;
  assign new_new_n30191__ = ~ys__n602 & ~new_new_n30190__;
  assign new_new_n30192__ = new_new_n30037__ & ~new_new_n30190__;
  assign new_new_n30193__ = ys__n26008 & new_new_n16712__;
  assign new_new_n30194__ = ys__n26008 & ~new_new_n26679__;
  assign new_new_n30195__ = ~new_new_n30193__ & ~new_new_n30194__;
  assign new_new_n30196__ = ~new_new_n30037__ & ~new_new_n30195__;
  assign new_new_n30197__ = ~new_new_n30192__ & ~new_new_n30196__;
  assign new_new_n30198__ = ys__n602 & ~new_new_n30197__;
  assign ys__n26623 = new_new_n30191__ | new_new_n30198__;
  assign new_new_n30200__ = ~ys__n778 & ys__n26008;
  assign new_new_n30201__ = ys__n26008 & new_new_n30026__;
  assign new_new_n30202__ = ys__n35057 & new_new_n26678__;
  assign new_new_n30203__ = ~ys__n18173 & ys__n18475;
  assign new_new_n30204__ = ys__n18173 & ys__n30895;
  assign new_new_n30205__ = ~new_new_n30203__ & ~new_new_n30204__;
  assign new_new_n30206__ = ~new_new_n16728__ & ~new_new_n30205__;
  assign new_new_n30207__ = ~new_new_n30202__ & ~new_new_n30206__;
  assign new_new_n30208__ = ~new_new_n30026__ & ~new_new_n30207__;
  assign new_new_n30209__ = ~new_new_n30201__ & ~new_new_n30208__;
  assign new_new_n30210__ = ys__n778 & ~new_new_n30209__;
  assign new_new_n30211__ = ~new_new_n30200__ & ~new_new_n30210__;
  assign new_new_n30212__ = ~ys__n602 & ~new_new_n30211__;
  assign new_new_n30213__ = new_new_n30037__ & ~new_new_n30211__;
  assign new_new_n30214__ = ys__n26011 & new_new_n16712__;
  assign new_new_n30215__ = ys__n26011 & ~new_new_n26679__;
  assign new_new_n30216__ = ~new_new_n30214__ & ~new_new_n30215__;
  assign new_new_n30217__ = ~new_new_n30037__ & ~new_new_n30216__;
  assign new_new_n30218__ = ~new_new_n30213__ & ~new_new_n30217__;
  assign new_new_n30219__ = ys__n602 & ~new_new_n30218__;
  assign ys__n26625 = new_new_n30212__ | new_new_n30219__;
  assign new_new_n30221__ = ~ys__n778 & ys__n26011;
  assign new_new_n30222__ = ys__n26011 & new_new_n30026__;
  assign new_new_n30223__ = ~ys__n18173 & ys__n18478;
  assign new_new_n30224__ = ys__n18173 & ys__n30897;
  assign new_new_n30225__ = ~new_new_n30223__ & ~new_new_n30224__;
  assign new_new_n30226__ = ~new_new_n16728__ & ~new_new_n30225__;
  assign new_new_n30227__ = ~new_new_n30026__ & new_new_n30226__;
  assign new_new_n30228__ = ~new_new_n30222__ & ~new_new_n30227__;
  assign new_new_n30229__ = ys__n778 & ~new_new_n30228__;
  assign new_new_n30230__ = ~new_new_n30221__ & ~new_new_n30229__;
  assign new_new_n30231__ = ~ys__n602 & ~new_new_n30230__;
  assign new_new_n30232__ = new_new_n30037__ & ~new_new_n30230__;
  assign new_new_n30233__ = ys__n26014 & new_new_n16712__;
  assign new_new_n30234__ = ys__n26014 & ~new_new_n26679__;
  assign new_new_n30235__ = ~new_new_n30233__ & ~new_new_n30234__;
  assign new_new_n30236__ = ~new_new_n30037__ & ~new_new_n30235__;
  assign new_new_n30237__ = ~new_new_n30232__ & ~new_new_n30236__;
  assign new_new_n30238__ = ys__n602 & ~new_new_n30237__;
  assign ys__n26627 = new_new_n30231__ | new_new_n30238__;
  assign new_new_n30240__ = ~ys__n778 & ys__n26014;
  assign new_new_n30241__ = ys__n26014 & new_new_n30026__;
  assign new_new_n30242__ = ys__n184 & new_new_n26678__;
  assign new_new_n30243__ = ~ys__n18173 & ys__n18481;
  assign new_new_n30244__ = ys__n18173 & ys__n30899;
  assign new_new_n30245__ = ~new_new_n30243__ & ~new_new_n30244__;
  assign new_new_n30246__ = ~new_new_n16728__ & ~new_new_n30245__;
  assign new_new_n30247__ = ~new_new_n30242__ & ~new_new_n30246__;
  assign new_new_n30248__ = ~new_new_n30026__ & ~new_new_n30247__;
  assign new_new_n30249__ = ~new_new_n30241__ & ~new_new_n30248__;
  assign new_new_n30250__ = ys__n778 & ~new_new_n30249__;
  assign new_new_n30251__ = ~new_new_n30240__ & ~new_new_n30250__;
  assign new_new_n30252__ = ~ys__n602 & ~new_new_n30251__;
  assign new_new_n30253__ = new_new_n30037__ & ~new_new_n30251__;
  assign new_new_n30254__ = ys__n26017 & new_new_n16712__;
  assign new_new_n30255__ = ys__n26017 & ~new_new_n26679__;
  assign new_new_n30256__ = ~new_new_n30254__ & ~new_new_n30255__;
  assign new_new_n30257__ = ~new_new_n30037__ & ~new_new_n30256__;
  assign new_new_n30258__ = ~new_new_n30253__ & ~new_new_n30257__;
  assign new_new_n30259__ = ys__n602 & ~new_new_n30258__;
  assign ys__n26629 = new_new_n30252__ | new_new_n30259__;
  assign new_new_n30261__ = ~ys__n778 & ys__n26017;
  assign new_new_n30262__ = ys__n26017 & new_new_n30026__;
  assign new_new_n30263__ = ys__n182 & new_new_n26678__;
  assign new_new_n30264__ = ~ys__n18173 & ys__n18484;
  assign new_new_n30265__ = ys__n18173 & ys__n30901;
  assign new_new_n30266__ = ~new_new_n30264__ & ~new_new_n30265__;
  assign new_new_n30267__ = ~new_new_n16728__ & ~new_new_n30266__;
  assign new_new_n30268__ = ~new_new_n30263__ & ~new_new_n30267__;
  assign new_new_n30269__ = ~new_new_n30026__ & ~new_new_n30268__;
  assign new_new_n30270__ = ~new_new_n30262__ & ~new_new_n30269__;
  assign new_new_n30271__ = ys__n778 & ~new_new_n30270__;
  assign new_new_n30272__ = ~new_new_n30261__ & ~new_new_n30271__;
  assign new_new_n30273__ = ~ys__n602 & ~new_new_n30272__;
  assign new_new_n30274__ = new_new_n30037__ & ~new_new_n30272__;
  assign new_new_n30275__ = ys__n26020 & new_new_n16712__;
  assign new_new_n30276__ = ys__n26020 & ~new_new_n26679__;
  assign new_new_n30277__ = ~new_new_n30275__ & ~new_new_n30276__;
  assign new_new_n30278__ = ~new_new_n30037__ & ~new_new_n30277__;
  assign new_new_n30279__ = ~new_new_n30274__ & ~new_new_n30278__;
  assign new_new_n30280__ = ys__n602 & ~new_new_n30279__;
  assign ys__n26631 = new_new_n30273__ | new_new_n30280__;
  assign new_new_n30282__ = ~ys__n778 & ys__n26020;
  assign new_new_n30283__ = ys__n26020 & new_new_n30026__;
  assign new_new_n30284__ = ~ys__n18173 & ys__n18487;
  assign new_new_n30285__ = ys__n18173 & ys__n30903;
  assign new_new_n30286__ = ~new_new_n30284__ & ~new_new_n30285__;
  assign new_new_n30287__ = ~new_new_n16728__ & ~new_new_n30286__;
  assign new_new_n30288__ = ~new_new_n30026__ & new_new_n30287__;
  assign new_new_n30289__ = ~new_new_n30283__ & ~new_new_n30288__;
  assign new_new_n30290__ = ys__n778 & ~new_new_n30289__;
  assign new_new_n30291__ = ~new_new_n30282__ & ~new_new_n30290__;
  assign new_new_n30292__ = ~ys__n602 & ~new_new_n30291__;
  assign new_new_n30293__ = new_new_n30037__ & ~new_new_n30291__;
  assign new_new_n30294__ = ys__n26023 & new_new_n16712__;
  assign new_new_n30295__ = ys__n26023 & ~new_new_n26679__;
  assign new_new_n30296__ = ~new_new_n30294__ & ~new_new_n30295__;
  assign new_new_n30297__ = ~new_new_n30037__ & ~new_new_n30296__;
  assign new_new_n30298__ = ~new_new_n30293__ & ~new_new_n30297__;
  assign new_new_n30299__ = ys__n602 & ~new_new_n30298__;
  assign ys__n26633 = new_new_n30292__ | new_new_n30299__;
  assign new_new_n30301__ = ~ys__n778 & ys__n26023;
  assign new_new_n30302__ = ys__n26023 & new_new_n30026__;
  assign new_new_n30303__ = ~ys__n18173 & ys__n18490;
  assign new_new_n30304__ = ys__n18173 & ys__n30905;
  assign new_new_n30305__ = ~new_new_n30303__ & ~new_new_n30304__;
  assign new_new_n30306__ = ~new_new_n16728__ & ~new_new_n30305__;
  assign new_new_n30307__ = ~new_new_n30026__ & new_new_n30306__;
  assign new_new_n30308__ = ~new_new_n30302__ & ~new_new_n30307__;
  assign new_new_n30309__ = ys__n778 & ~new_new_n30308__;
  assign new_new_n30310__ = ~new_new_n30301__ & ~new_new_n30309__;
  assign new_new_n30311__ = ~ys__n602 & ~new_new_n30310__;
  assign new_new_n30312__ = new_new_n30037__ & ~new_new_n30310__;
  assign new_new_n30313__ = ys__n26026 & new_new_n16712__;
  assign new_new_n30314__ = ys__n26026 & ~new_new_n26679__;
  assign new_new_n30315__ = ~new_new_n30313__ & ~new_new_n30314__;
  assign new_new_n30316__ = ~new_new_n30037__ & ~new_new_n30315__;
  assign new_new_n30317__ = ~new_new_n30312__ & ~new_new_n30316__;
  assign new_new_n30318__ = ys__n602 & ~new_new_n30317__;
  assign ys__n26635 = new_new_n30311__ | new_new_n30318__;
  assign new_new_n30320__ = ~ys__n778 & ys__n26026;
  assign new_new_n30321__ = ys__n26026 & new_new_n30026__;
  assign new_new_n30322__ = ~ys__n18173 & ys__n18493;
  assign new_new_n30323__ = ys__n18173 & ys__n30907;
  assign new_new_n30324__ = ~new_new_n30322__ & ~new_new_n30323__;
  assign new_new_n30325__ = ~new_new_n16728__ & ~new_new_n30324__;
  assign new_new_n30326__ = ~new_new_n30026__ & new_new_n30325__;
  assign new_new_n30327__ = ~new_new_n30321__ & ~new_new_n30326__;
  assign new_new_n30328__ = ys__n778 & ~new_new_n30327__;
  assign new_new_n30329__ = ~new_new_n30320__ & ~new_new_n30328__;
  assign new_new_n30330__ = ~ys__n602 & ~new_new_n30329__;
  assign new_new_n30331__ = new_new_n30037__ & ~new_new_n30329__;
  assign new_new_n30332__ = ys__n26029 & new_new_n16712__;
  assign new_new_n30333__ = ys__n26029 & ~new_new_n26679__;
  assign new_new_n30334__ = ~new_new_n30332__ & ~new_new_n30333__;
  assign new_new_n30335__ = ~new_new_n30037__ & ~new_new_n30334__;
  assign new_new_n30336__ = ~new_new_n30331__ & ~new_new_n30335__;
  assign new_new_n30337__ = ys__n602 & ~new_new_n30336__;
  assign ys__n26637 = new_new_n30330__ | new_new_n30337__;
  assign new_new_n30339__ = ~ys__n778 & ys__n26029;
  assign new_new_n30340__ = ys__n26029 & new_new_n30026__;
  assign new_new_n30341__ = ~ys__n18173 & ys__n18496;
  assign new_new_n30342__ = ys__n18173 & ys__n30909;
  assign new_new_n30343__ = ~new_new_n30341__ & ~new_new_n30342__;
  assign new_new_n30344__ = ~new_new_n16728__ & ~new_new_n30343__;
  assign new_new_n30345__ = ~new_new_n26678__ & ~new_new_n30344__;
  assign new_new_n30346__ = ~new_new_n30026__ & ~new_new_n30345__;
  assign new_new_n30347__ = ~new_new_n30340__ & ~new_new_n30346__;
  assign new_new_n30348__ = ys__n778 & ~new_new_n30347__;
  assign new_new_n30349__ = ~new_new_n30339__ & ~new_new_n30348__;
  assign new_new_n30350__ = ~ys__n602 & ~new_new_n30349__;
  assign new_new_n30351__ = new_new_n30037__ & ~new_new_n30349__;
  assign new_new_n30352__ = ys__n26032 & new_new_n16712__;
  assign new_new_n30353__ = ys__n26032 & ~new_new_n26679__;
  assign new_new_n30354__ = ~new_new_n30352__ & ~new_new_n30353__;
  assign new_new_n30355__ = ~new_new_n30037__ & ~new_new_n30354__;
  assign new_new_n30356__ = ~new_new_n30351__ & ~new_new_n30355__;
  assign new_new_n30357__ = ys__n602 & ~new_new_n30356__;
  assign ys__n26639 = new_new_n30350__ | new_new_n30357__;
  assign new_new_n30359__ = ~ys__n778 & ys__n26032;
  assign new_new_n30360__ = ys__n26032 & new_new_n30026__;
  assign new_new_n30361__ = ~ys__n18173 & ys__n18499;
  assign new_new_n30362__ = ys__n18173 & ys__n30911;
  assign new_new_n30363__ = ~new_new_n30361__ & ~new_new_n30362__;
  assign new_new_n30364__ = ~new_new_n16728__ & ~new_new_n30363__;
  assign new_new_n30365__ = ~new_new_n30026__ & new_new_n30364__;
  assign new_new_n30366__ = ~new_new_n30360__ & ~new_new_n30365__;
  assign new_new_n30367__ = ys__n778 & ~new_new_n30366__;
  assign new_new_n30368__ = ~new_new_n30359__ & ~new_new_n30367__;
  assign new_new_n30369__ = ~ys__n602 & ~new_new_n30368__;
  assign new_new_n30370__ = new_new_n30037__ & ~new_new_n30368__;
  assign new_new_n30371__ = ys__n26035 & new_new_n16712__;
  assign new_new_n30372__ = ys__n26035 & ~new_new_n26679__;
  assign new_new_n30373__ = ~new_new_n30371__ & ~new_new_n30372__;
  assign new_new_n30374__ = ~new_new_n30037__ & ~new_new_n30373__;
  assign new_new_n30375__ = ~new_new_n30370__ & ~new_new_n30374__;
  assign new_new_n30376__ = ys__n602 & ~new_new_n30375__;
  assign ys__n26641 = new_new_n30369__ | new_new_n30376__;
  assign new_new_n30378__ = ~ys__n778 & ys__n26035;
  assign new_new_n30379__ = ys__n26035 & new_new_n30026__;
  assign new_new_n30380__ = ~ys__n18173 & ys__n18502;
  assign new_new_n30381__ = ys__n18173 & ys__n30913;
  assign new_new_n30382__ = ~new_new_n30380__ & ~new_new_n30381__;
  assign new_new_n30383__ = ~new_new_n16728__ & ~new_new_n30382__;
  assign new_new_n30384__ = ~new_new_n30026__ & new_new_n30383__;
  assign new_new_n30385__ = ~new_new_n30379__ & ~new_new_n30384__;
  assign new_new_n30386__ = ys__n778 & ~new_new_n30385__;
  assign new_new_n30387__ = ~new_new_n30378__ & ~new_new_n30386__;
  assign new_new_n30388__ = ~ys__n602 & ~new_new_n30387__;
  assign new_new_n30389__ = new_new_n30037__ & ~new_new_n30387__;
  assign new_new_n30390__ = ys__n26038 & new_new_n16712__;
  assign new_new_n30391__ = ys__n26038 & ~new_new_n26679__;
  assign new_new_n30392__ = ~new_new_n30390__ & ~new_new_n30391__;
  assign new_new_n30393__ = ~new_new_n30037__ & ~new_new_n30392__;
  assign new_new_n30394__ = ~new_new_n30389__ & ~new_new_n30393__;
  assign new_new_n30395__ = ys__n602 & ~new_new_n30394__;
  assign ys__n26643 = new_new_n30388__ | new_new_n30395__;
  assign new_new_n30397__ = ~ys__n778 & ys__n26038;
  assign new_new_n30398__ = ys__n26038 & new_new_n30026__;
  assign new_new_n30399__ = ~ys__n18173 & ys__n18505;
  assign new_new_n30400__ = ys__n18173 & ys__n30915;
  assign new_new_n30401__ = ~new_new_n30399__ & ~new_new_n30400__;
  assign new_new_n30402__ = ~new_new_n16728__ & ~new_new_n30401__;
  assign new_new_n30403__ = ~new_new_n30026__ & new_new_n30402__;
  assign new_new_n30404__ = ~new_new_n30398__ & ~new_new_n30403__;
  assign new_new_n30405__ = ys__n778 & ~new_new_n30404__;
  assign new_new_n30406__ = ~new_new_n30397__ & ~new_new_n30405__;
  assign new_new_n30407__ = ~ys__n602 & ~new_new_n30406__;
  assign new_new_n30408__ = new_new_n30037__ & ~new_new_n30406__;
  assign new_new_n30409__ = ys__n26041 & new_new_n16712__;
  assign new_new_n30410__ = ys__n26041 & ~new_new_n26679__;
  assign new_new_n30411__ = ~new_new_n30409__ & ~new_new_n30410__;
  assign new_new_n30412__ = ~new_new_n30037__ & ~new_new_n30411__;
  assign new_new_n30413__ = ~new_new_n30408__ & ~new_new_n30412__;
  assign new_new_n30414__ = ys__n602 & ~new_new_n30413__;
  assign ys__n26645 = new_new_n30407__ | new_new_n30414__;
  assign new_new_n30416__ = ~ys__n778 & ys__n26041;
  assign new_new_n30417__ = ys__n26041 & new_new_n30026__;
  assign new_new_n30418__ = ~ys__n18173 & ys__n18508;
  assign new_new_n30419__ = ys__n18173 & ys__n30917;
  assign new_new_n30420__ = ~new_new_n30418__ & ~new_new_n30419__;
  assign new_new_n30421__ = ~new_new_n16728__ & ~new_new_n30420__;
  assign new_new_n30422__ = ~new_new_n30026__ & new_new_n30421__;
  assign new_new_n30423__ = ~new_new_n30417__ & ~new_new_n30422__;
  assign new_new_n30424__ = ys__n778 & ~new_new_n30423__;
  assign new_new_n30425__ = ~new_new_n30416__ & ~new_new_n30424__;
  assign new_new_n30426__ = ~ys__n602 & ~new_new_n30425__;
  assign new_new_n30427__ = new_new_n30037__ & ~new_new_n30425__;
  assign new_new_n30428__ = ys__n26044 & new_new_n16712__;
  assign new_new_n30429__ = ys__n26044 & ~new_new_n26679__;
  assign new_new_n30430__ = ~new_new_n30428__ & ~new_new_n30429__;
  assign new_new_n30431__ = ~new_new_n30037__ & ~new_new_n30430__;
  assign new_new_n30432__ = ~new_new_n30427__ & ~new_new_n30431__;
  assign new_new_n30433__ = ys__n602 & ~new_new_n30432__;
  assign ys__n26647 = new_new_n30426__ | new_new_n30433__;
  assign new_new_n30435__ = ~ys__n778 & ys__n26044;
  assign new_new_n30436__ = ys__n26044 & new_new_n30026__;
  assign new_new_n30437__ = ~ys__n18173 & ys__n18511;
  assign new_new_n30438__ = ys__n18173 & ys__n30919;
  assign new_new_n30439__ = ~new_new_n30437__ & ~new_new_n30438__;
  assign new_new_n30440__ = ~new_new_n16728__ & ~new_new_n30439__;
  assign new_new_n30441__ = ~new_new_n30026__ & new_new_n30440__;
  assign new_new_n30442__ = ~new_new_n30436__ & ~new_new_n30441__;
  assign new_new_n30443__ = ys__n778 & ~new_new_n30442__;
  assign new_new_n30444__ = ~new_new_n30435__ & ~new_new_n30443__;
  assign new_new_n30445__ = ~ys__n602 & ~new_new_n30444__;
  assign new_new_n30446__ = new_new_n30037__ & ~new_new_n30444__;
  assign new_new_n30447__ = ys__n26047 & new_new_n16712__;
  assign new_new_n30448__ = ys__n26047 & ~new_new_n26679__;
  assign new_new_n30449__ = ~new_new_n30447__ & ~new_new_n30448__;
  assign new_new_n30450__ = ~new_new_n30037__ & ~new_new_n30449__;
  assign new_new_n30451__ = ~new_new_n30446__ & ~new_new_n30450__;
  assign new_new_n30452__ = ys__n602 & ~new_new_n30451__;
  assign ys__n26649 = new_new_n30445__ | new_new_n30452__;
  assign new_new_n30454__ = ~ys__n778 & ys__n26047;
  assign new_new_n30455__ = ys__n26047 & new_new_n30026__;
  assign new_new_n30456__ = ~ys__n18173 & ys__n18514;
  assign new_new_n30457__ = ys__n18173 & ys__n30921;
  assign new_new_n30458__ = ~new_new_n30456__ & ~new_new_n30457__;
  assign new_new_n30459__ = ~new_new_n16728__ & ~new_new_n30458__;
  assign new_new_n30460__ = ~new_new_n30026__ & new_new_n30459__;
  assign new_new_n30461__ = ~new_new_n30455__ & ~new_new_n30460__;
  assign new_new_n30462__ = ys__n778 & ~new_new_n30461__;
  assign new_new_n30463__ = ~new_new_n30454__ & ~new_new_n30462__;
  assign new_new_n30464__ = ~ys__n602 & ~new_new_n30463__;
  assign new_new_n30465__ = new_new_n30037__ & ~new_new_n30463__;
  assign new_new_n30466__ = ys__n26050 & new_new_n16712__;
  assign new_new_n30467__ = ys__n26050 & ~new_new_n26679__;
  assign new_new_n30468__ = ~new_new_n30466__ & ~new_new_n30467__;
  assign new_new_n30469__ = ~new_new_n30037__ & ~new_new_n30468__;
  assign new_new_n30470__ = ~new_new_n30465__ & ~new_new_n30469__;
  assign new_new_n30471__ = ys__n602 & ~new_new_n30470__;
  assign ys__n26651 = new_new_n30464__ | new_new_n30471__;
  assign new_new_n30473__ = ~ys__n778 & ys__n26050;
  assign new_new_n30474__ = ys__n26050 & new_new_n30026__;
  assign new_new_n30475__ = ~ys__n18173 & ys__n18517;
  assign new_new_n30476__ = ys__n18173 & ys__n30923;
  assign new_new_n30477__ = ~new_new_n30475__ & ~new_new_n30476__;
  assign new_new_n30478__ = ~new_new_n16728__ & ~new_new_n30477__;
  assign new_new_n30479__ = ~new_new_n26678__ & ~new_new_n30478__;
  assign new_new_n30480__ = ~new_new_n30026__ & ~new_new_n30479__;
  assign new_new_n30481__ = ~new_new_n30474__ & ~new_new_n30480__;
  assign new_new_n30482__ = ys__n778 & ~new_new_n30481__;
  assign new_new_n30483__ = ~new_new_n30473__ & ~new_new_n30482__;
  assign new_new_n30484__ = ~ys__n602 & ~new_new_n30483__;
  assign new_new_n30485__ = new_new_n30037__ & ~new_new_n30483__;
  assign new_new_n30486__ = ys__n26053 & new_new_n16712__;
  assign new_new_n30487__ = ys__n26053 & ~new_new_n26679__;
  assign new_new_n30488__ = ~new_new_n30486__ & ~new_new_n30487__;
  assign new_new_n30489__ = ~new_new_n30037__ & ~new_new_n30488__;
  assign new_new_n30490__ = ~new_new_n30485__ & ~new_new_n30489__;
  assign new_new_n30491__ = ys__n602 & ~new_new_n30490__;
  assign ys__n26653 = new_new_n30484__ | new_new_n30491__;
  assign new_new_n30493__ = ~ys__n778 & ys__n26053;
  assign new_new_n30494__ = ys__n26053 & new_new_n30026__;
  assign new_new_n30495__ = ~ys__n18173 & ys__n18520;
  assign new_new_n30496__ = ys__n18173 & ys__n30925;
  assign new_new_n30497__ = ~new_new_n30495__ & ~new_new_n30496__;
  assign new_new_n30498__ = ~new_new_n16728__ & ~new_new_n30497__;
  assign new_new_n30499__ = ~new_new_n30026__ & new_new_n30498__;
  assign new_new_n30500__ = ~new_new_n30494__ & ~new_new_n30499__;
  assign new_new_n30501__ = ys__n778 & ~new_new_n30500__;
  assign new_new_n30502__ = ~new_new_n30493__ & ~new_new_n30501__;
  assign new_new_n30503__ = ~ys__n602 & ~new_new_n30502__;
  assign new_new_n30504__ = new_new_n30037__ & ~new_new_n30502__;
  assign new_new_n30505__ = ys__n26056 & new_new_n16712__;
  assign new_new_n30506__ = ys__n26056 & ~new_new_n26679__;
  assign new_new_n30507__ = ~new_new_n30505__ & ~new_new_n30506__;
  assign new_new_n30508__ = ~new_new_n30037__ & ~new_new_n30507__;
  assign new_new_n30509__ = ~new_new_n30504__ & ~new_new_n30508__;
  assign new_new_n30510__ = ys__n602 & ~new_new_n30509__;
  assign ys__n26655 = new_new_n30503__ | new_new_n30510__;
  assign new_new_n30512__ = ~ys__n778 & ys__n26056;
  assign new_new_n30513__ = ys__n26056 & new_new_n30026__;
  assign new_new_n30514__ = ~ys__n18173 & ys__n18523;
  assign new_new_n30515__ = ys__n18173 & ys__n30927;
  assign new_new_n30516__ = ~new_new_n30514__ & ~new_new_n30515__;
  assign new_new_n30517__ = ~new_new_n16728__ & ~new_new_n30516__;
  assign new_new_n30518__ = ~new_new_n30026__ & new_new_n30517__;
  assign new_new_n30519__ = ~new_new_n30513__ & ~new_new_n30518__;
  assign new_new_n30520__ = ys__n778 & ~new_new_n30519__;
  assign new_new_n30521__ = ~new_new_n30512__ & ~new_new_n30520__;
  assign new_new_n30522__ = ~ys__n602 & ~new_new_n30521__;
  assign new_new_n30523__ = new_new_n30037__ & ~new_new_n30521__;
  assign new_new_n30524__ = ys__n26059 & new_new_n16712__;
  assign new_new_n30525__ = ys__n26059 & ~new_new_n26679__;
  assign new_new_n30526__ = ~new_new_n30524__ & ~new_new_n30525__;
  assign new_new_n30527__ = ~new_new_n30037__ & ~new_new_n30526__;
  assign new_new_n30528__ = ~new_new_n30523__ & ~new_new_n30527__;
  assign new_new_n30529__ = ys__n602 & ~new_new_n30528__;
  assign ys__n26657 = new_new_n30522__ | new_new_n30529__;
  assign new_new_n30531__ = ~ys__n778 & ys__n26059;
  assign new_new_n30532__ = ys__n26059 & new_new_n30026__;
  assign new_new_n30533__ = ys__n30941 & new_new_n26678__;
  assign new_new_n30534__ = ~ys__n18173 & ys__n18526;
  assign new_new_n30535__ = ys__n18173 & ys__n30929;
  assign new_new_n30536__ = ~new_new_n30534__ & ~new_new_n30535__;
  assign new_new_n30537__ = ~new_new_n16728__ & ~new_new_n30536__;
  assign new_new_n30538__ = ~new_new_n30533__ & ~new_new_n30537__;
  assign new_new_n30539__ = ~new_new_n30026__ & ~new_new_n30538__;
  assign new_new_n30540__ = ~new_new_n30532__ & ~new_new_n30539__;
  assign new_new_n30541__ = ys__n778 & ~new_new_n30540__;
  assign new_new_n30542__ = ~new_new_n30531__ & ~new_new_n30541__;
  assign new_new_n30543__ = ~ys__n602 & ~new_new_n30542__;
  assign new_new_n30544__ = new_new_n30037__ & ~new_new_n30542__;
  assign new_new_n30545__ = ys__n26062 & new_new_n16712__;
  assign new_new_n30546__ = ys__n26062 & ~new_new_n26679__;
  assign new_new_n30547__ = ~new_new_n30545__ & ~new_new_n30546__;
  assign new_new_n30548__ = ~new_new_n30037__ & ~new_new_n30547__;
  assign new_new_n30549__ = ~new_new_n30544__ & ~new_new_n30548__;
  assign new_new_n30550__ = ys__n602 & ~new_new_n30549__;
  assign ys__n26659 = new_new_n30543__ | new_new_n30550__;
  assign new_new_n30552__ = ~ys__n778 & ys__n26062;
  assign new_new_n30553__ = ys__n26062 & new_new_n30026__;
  assign new_new_n30554__ = ys__n202 & new_new_n26678__;
  assign new_new_n30555__ = ~ys__n18173 & ys__n18529;
  assign new_new_n30556__ = ys__n18173 & ys__n30931;
  assign new_new_n30557__ = ~new_new_n30555__ & ~new_new_n30556__;
  assign new_new_n30558__ = ~new_new_n16728__ & ~new_new_n30557__;
  assign new_new_n30559__ = ~new_new_n30554__ & ~new_new_n30558__;
  assign new_new_n30560__ = ~new_new_n30026__ & ~new_new_n30559__;
  assign new_new_n30561__ = ~new_new_n30553__ & ~new_new_n30560__;
  assign new_new_n30562__ = ys__n778 & ~new_new_n30561__;
  assign new_new_n30563__ = ~new_new_n30552__ & ~new_new_n30562__;
  assign new_new_n30564__ = ~ys__n602 & ~new_new_n30563__;
  assign new_new_n30565__ = new_new_n30037__ & ~new_new_n30563__;
  assign new_new_n30566__ = ys__n26065 & new_new_n16712__;
  assign new_new_n30567__ = ys__n26065 & ~new_new_n26679__;
  assign new_new_n30568__ = ~new_new_n30566__ & ~new_new_n30567__;
  assign new_new_n30569__ = ~new_new_n30037__ & ~new_new_n30568__;
  assign new_new_n30570__ = ~new_new_n30565__ & ~new_new_n30569__;
  assign new_new_n30571__ = ys__n602 & ~new_new_n30570__;
  assign ys__n26661 = new_new_n30564__ | new_new_n30571__;
  assign new_new_n30573__ = ~ys__n778 & ys__n26065;
  assign new_new_n30574__ = ys__n26065 & new_new_n30026__;
  assign new_new_n30575__ = ~ys__n18173 & ys__n18532;
  assign new_new_n30576__ = ys__n18173 & ys__n30933;
  assign new_new_n30577__ = ~new_new_n30575__ & ~new_new_n30576__;
  assign new_new_n30578__ = ~new_new_n16728__ & ~new_new_n30577__;
  assign new_new_n30579__ = ~new_new_n30026__ & new_new_n30578__;
  assign new_new_n30580__ = ~new_new_n30574__ & ~new_new_n30579__;
  assign new_new_n30581__ = ys__n778 & ~new_new_n30580__;
  assign new_new_n30582__ = ~new_new_n30573__ & ~new_new_n30581__;
  assign new_new_n30583__ = ~ys__n602 & ~new_new_n30582__;
  assign new_new_n30584__ = new_new_n30037__ & ~new_new_n30582__;
  assign new_new_n30585__ = ys__n26068 & new_new_n16712__;
  assign new_new_n30586__ = ys__n26068 & ~new_new_n26679__;
  assign new_new_n30587__ = ~new_new_n30585__ & ~new_new_n30586__;
  assign new_new_n30588__ = ~new_new_n30037__ & ~new_new_n30587__;
  assign new_new_n30589__ = ~new_new_n30584__ & ~new_new_n30588__;
  assign new_new_n30590__ = ys__n602 & ~new_new_n30589__;
  assign ys__n26663 = new_new_n30583__ | new_new_n30590__;
  assign new_new_n30592__ = ~ys__n778 & ys__n26068;
  assign new_new_n30593__ = ys__n26068 & new_new_n30026__;
  assign new_new_n30594__ = ~ys__n18173 & ys__n18535;
  assign new_new_n30595__ = ys__n18173 & ys__n30935;
  assign new_new_n30596__ = ~new_new_n30594__ & ~new_new_n30595__;
  assign new_new_n30597__ = ~new_new_n16728__ & ~new_new_n30596__;
  assign new_new_n30598__ = ~new_new_n30026__ & new_new_n30597__;
  assign new_new_n30599__ = ~new_new_n30593__ & ~new_new_n30598__;
  assign new_new_n30600__ = ys__n778 & ~new_new_n30599__;
  assign new_new_n30601__ = ~new_new_n30592__ & ~new_new_n30600__;
  assign new_new_n30602__ = ~ys__n602 & ~new_new_n30601__;
  assign new_new_n30603__ = new_new_n30037__ & ~new_new_n30601__;
  assign new_new_n30604__ = ys__n26071 & new_new_n16712__;
  assign new_new_n30605__ = ys__n26071 & ~new_new_n26679__;
  assign new_new_n30606__ = ~new_new_n30604__ & ~new_new_n30605__;
  assign new_new_n30607__ = ~new_new_n30037__ & ~new_new_n30606__;
  assign new_new_n30608__ = ~new_new_n30603__ & ~new_new_n30607__;
  assign new_new_n30609__ = ys__n602 & ~new_new_n30608__;
  assign ys__n26665 = new_new_n30602__ | new_new_n30609__;
  assign new_new_n30611__ = ~ys__n778 & ys__n26071;
  assign new_new_n30612__ = ys__n26071 & new_new_n30026__;
  assign new_new_n30613__ = ~ys__n18173 & ys__n18538;
  assign new_new_n30614__ = ys__n18173 & ys__n30937;
  assign new_new_n30615__ = ~new_new_n30613__ & ~new_new_n30614__;
  assign new_new_n30616__ = ~new_new_n16728__ & ~new_new_n30615__;
  assign new_new_n30617__ = ~new_new_n30026__ & new_new_n30616__;
  assign new_new_n30618__ = ~new_new_n30612__ & ~new_new_n30617__;
  assign new_new_n30619__ = ys__n778 & ~new_new_n30618__;
  assign new_new_n30620__ = ~new_new_n30611__ & ~new_new_n30619__;
  assign new_new_n30621__ = ~ys__n602 & ~new_new_n30620__;
  assign new_new_n30622__ = new_new_n30037__ & ~new_new_n30620__;
  assign new_new_n30623__ = ys__n26074 & new_new_n16712__;
  assign new_new_n30624__ = ys__n26074 & ~new_new_n26679__;
  assign new_new_n30625__ = ~new_new_n30623__ & ~new_new_n30624__;
  assign new_new_n30626__ = ~new_new_n30037__ & ~new_new_n30625__;
  assign new_new_n30627__ = ~new_new_n30622__ & ~new_new_n30626__;
  assign new_new_n30628__ = ys__n602 & ~new_new_n30627__;
  assign ys__n26667 = new_new_n30621__ | new_new_n30628__;
  assign new_new_n30630__ = ~ys__n778 & ys__n26074;
  assign new_new_n30631__ = ys__n26074 & new_new_n30026__;
  assign new_new_n30632__ = ~ys__n18173 & ys__n18541;
  assign new_new_n30633__ = ys__n18173 & ys__n30939;
  assign new_new_n30634__ = ~new_new_n30632__ & ~new_new_n30633__;
  assign new_new_n30635__ = ~new_new_n16728__ & ~new_new_n30634__;
  assign new_new_n30636__ = ~new_new_n30026__ & new_new_n30635__;
  assign new_new_n30637__ = ~new_new_n30631__ & ~new_new_n30636__;
  assign new_new_n30638__ = ys__n778 & ~new_new_n30637__;
  assign new_new_n30639__ = ~new_new_n30630__ & ~new_new_n30638__;
  assign new_new_n30640__ = ~ys__n602 & ~new_new_n30639__;
  assign new_new_n30641__ = new_new_n30037__ & ~new_new_n30639__;
  assign new_new_n30642__ = ys__n26359 & new_new_n16712__;
  assign new_new_n30643__ = ys__n25470 & ~new_new_n12328__;
  assign new_new_n30644__ = new_new_n26674__ & new_new_n30643__;
  assign new_new_n30645__ = new_new_n12325__ & new_new_n26667__;
  assign new_new_n30646__ = new_new_n30644__ & new_new_n30645__;
  assign new_new_n30647__ = ~new_new_n26679__ & new_new_n30646__;
  assign new_new_n30648__ = ~new_new_n30642__ & ~new_new_n30647__;
  assign new_new_n30649__ = ~new_new_n30037__ & ~new_new_n30648__;
  assign new_new_n30650__ = ~new_new_n30641__ & ~new_new_n30649__;
  assign new_new_n30651__ = ys__n602 & ~new_new_n30650__;
  assign ys__n26669 = new_new_n30640__ | new_new_n30651__;
  assign new_new_n30653__ = ~ys__n778 & ys__n26425;
  assign new_new_n30654__ = ys__n26425 & new_new_n16715__;
  assign new_new_n30655__ = ys__n26552 & ~new_new_n16715__;
  assign new_new_n30656__ = ~new_new_n30654__ & ~new_new_n30655__;
  assign new_new_n30657__ = ys__n778 & ~new_new_n30656__;
  assign new_new_n30658__ = ~new_new_n30653__ & ~new_new_n30657__;
  assign new_new_n30659__ = ~ys__n602 & ~new_new_n30658__;
  assign new_new_n30660__ = new_new_n16715__ & ~new_new_n30658__;
  assign new_new_n30661__ = ys__n26428 & new_new_n16712__;
  assign new_new_n30662__ = ys__n26428 & new_new_n16714__;
  assign new_new_n30663__ = ~new_new_n30661__ & ~new_new_n30662__;
  assign new_new_n30664__ = ~new_new_n16715__ & ~new_new_n30663__;
  assign new_new_n30665__ = ~new_new_n30660__ & ~new_new_n30664__;
  assign new_new_n30666__ = ys__n602 & ~new_new_n30665__;
  assign ys__n26671 = new_new_n30659__ | new_new_n30666__;
  assign new_new_n30668__ = ~ys__n778 & ys__n26428;
  assign new_new_n30669__ = ys__n26428 & new_new_n16715__;
  assign new_new_n30670__ = ys__n26553 & ~new_new_n16715__;
  assign new_new_n30671__ = ~new_new_n30669__ & ~new_new_n30670__;
  assign new_new_n30672__ = ys__n778 & ~new_new_n30671__;
  assign new_new_n30673__ = ~new_new_n30668__ & ~new_new_n30672__;
  assign new_new_n30674__ = ~ys__n602 & ~new_new_n30673__;
  assign new_new_n30675__ = new_new_n16715__ & ~new_new_n30673__;
  assign new_new_n30676__ = ys__n26431 & new_new_n16712__;
  assign new_new_n30677__ = ys__n26431 & new_new_n16714__;
  assign new_new_n30678__ = ~new_new_n30676__ & ~new_new_n30677__;
  assign new_new_n30679__ = ~new_new_n16715__ & ~new_new_n30678__;
  assign new_new_n30680__ = ~new_new_n30675__ & ~new_new_n30679__;
  assign new_new_n30681__ = ys__n602 & ~new_new_n30680__;
  assign ys__n26673 = new_new_n30674__ | new_new_n30681__;
  assign new_new_n30683__ = ~ys__n778 & ys__n26431;
  assign new_new_n30684__ = ys__n26431 & new_new_n16715__;
  assign new_new_n30685__ = ys__n26554 & ~new_new_n16715__;
  assign new_new_n30686__ = ~new_new_n30684__ & ~new_new_n30685__;
  assign new_new_n30687__ = ys__n778 & ~new_new_n30686__;
  assign new_new_n30688__ = ~new_new_n30683__ & ~new_new_n30687__;
  assign new_new_n30689__ = ~ys__n602 & ~new_new_n30688__;
  assign new_new_n30690__ = new_new_n16715__ & ~new_new_n30688__;
  assign new_new_n30691__ = ys__n26434 & new_new_n16712__;
  assign new_new_n30692__ = ys__n26434 & new_new_n16714__;
  assign new_new_n30693__ = ~new_new_n30691__ & ~new_new_n30692__;
  assign new_new_n30694__ = ~new_new_n16715__ & ~new_new_n30693__;
  assign new_new_n30695__ = ~new_new_n30690__ & ~new_new_n30694__;
  assign new_new_n30696__ = ys__n602 & ~new_new_n30695__;
  assign ys__n26675 = new_new_n30689__ | new_new_n30696__;
  assign new_new_n30698__ = ~ys__n778 & ys__n26434;
  assign new_new_n30699__ = ys__n26434 & new_new_n16715__;
  assign new_new_n30700__ = ys__n26555 & ~new_new_n16715__;
  assign new_new_n30701__ = ~new_new_n30699__ & ~new_new_n30700__;
  assign new_new_n30702__ = ys__n778 & ~new_new_n30701__;
  assign new_new_n30703__ = ~new_new_n30698__ & ~new_new_n30702__;
  assign new_new_n30704__ = ~ys__n602 & ~new_new_n30703__;
  assign new_new_n30705__ = new_new_n16715__ & ~new_new_n30703__;
  assign new_new_n30706__ = ys__n26437 & new_new_n16712__;
  assign new_new_n30707__ = ys__n26437 & new_new_n16714__;
  assign new_new_n30708__ = ~new_new_n30706__ & ~new_new_n30707__;
  assign new_new_n30709__ = ~new_new_n16715__ & ~new_new_n30708__;
  assign new_new_n30710__ = ~new_new_n30705__ & ~new_new_n30709__;
  assign new_new_n30711__ = ys__n602 & ~new_new_n30710__;
  assign ys__n26677 = new_new_n30704__ | new_new_n30711__;
  assign new_new_n30713__ = ~ys__n778 & ys__n26437;
  assign new_new_n30714__ = ys__n26437 & new_new_n16715__;
  assign new_new_n30715__ = ys__n26279 & ~new_new_n16715__;
  assign new_new_n30716__ = ~new_new_n30714__ & ~new_new_n30715__;
  assign new_new_n30717__ = ys__n778 & ~new_new_n30716__;
  assign new_new_n30718__ = ~new_new_n30713__ & ~new_new_n30717__;
  assign new_new_n30719__ = ~ys__n602 & ~new_new_n30718__;
  assign new_new_n30720__ = new_new_n16715__ & ~new_new_n30718__;
  assign new_new_n30721__ = ys__n26440 & new_new_n16712__;
  assign new_new_n30722__ = ys__n26440 & new_new_n16714__;
  assign new_new_n30723__ = ~new_new_n30721__ & ~new_new_n30722__;
  assign new_new_n30724__ = ~new_new_n16715__ & ~new_new_n30723__;
  assign new_new_n30725__ = ~new_new_n30720__ & ~new_new_n30724__;
  assign new_new_n30726__ = ys__n602 & ~new_new_n30725__;
  assign ys__n26679 = new_new_n30719__ | new_new_n30726__;
  assign new_new_n30728__ = ~ys__n778 & ys__n26440;
  assign new_new_n30729__ = ys__n26440 & new_new_n16715__;
  assign new_new_n30730__ = ys__n26556 & ~new_new_n16715__;
  assign new_new_n30731__ = ~new_new_n30729__ & ~new_new_n30730__;
  assign new_new_n30732__ = ys__n778 & ~new_new_n30731__;
  assign new_new_n30733__ = ~new_new_n30728__ & ~new_new_n30732__;
  assign new_new_n30734__ = ~ys__n602 & ~new_new_n30733__;
  assign new_new_n30735__ = new_new_n16715__ & ~new_new_n30733__;
  assign new_new_n30736__ = ys__n26443 & new_new_n16712__;
  assign new_new_n30737__ = ys__n26443 & new_new_n16714__;
  assign new_new_n30738__ = ~new_new_n30736__ & ~new_new_n30737__;
  assign new_new_n30739__ = ~new_new_n16715__ & ~new_new_n30738__;
  assign new_new_n30740__ = ~new_new_n30735__ & ~new_new_n30739__;
  assign new_new_n30741__ = ys__n602 & ~new_new_n30740__;
  assign ys__n26681 = new_new_n30734__ | new_new_n30741__;
  assign new_new_n30743__ = ~ys__n778 & ys__n26443;
  assign new_new_n30744__ = ys__n778 & ys__n26443;
  assign new_new_n30745__ = new_new_n16715__ & new_new_n30744__;
  assign new_new_n30746__ = ~new_new_n30743__ & ~new_new_n30745__;
  assign new_new_n30747__ = ~ys__n602 & ~new_new_n30746__;
  assign new_new_n30748__ = new_new_n16715__ & ~new_new_n30746__;
  assign new_new_n30749__ = ys__n26446 & new_new_n16712__;
  assign new_new_n30750__ = ys__n26446 & new_new_n16714__;
  assign new_new_n30751__ = ~new_new_n30749__ & ~new_new_n30750__;
  assign new_new_n30752__ = ~new_new_n16715__ & ~new_new_n30751__;
  assign new_new_n30753__ = ~new_new_n30748__ & ~new_new_n30752__;
  assign new_new_n30754__ = ys__n602 & ~new_new_n30753__;
  assign ys__n26683 = new_new_n30747__ | new_new_n30754__;
  assign new_new_n30756__ = ~ys__n778 & ys__n26446;
  assign new_new_n30757__ = ys__n26446 & new_new_n16715__;
  assign new_new_n30758__ = ys__n26557 & ~new_new_n16715__;
  assign new_new_n30759__ = ~new_new_n30757__ & ~new_new_n30758__;
  assign new_new_n30760__ = ys__n778 & ~new_new_n30759__;
  assign new_new_n30761__ = ~new_new_n30756__ & ~new_new_n30760__;
  assign new_new_n30762__ = ~ys__n602 & ~new_new_n30761__;
  assign new_new_n30763__ = new_new_n16715__ & ~new_new_n30761__;
  assign new_new_n30764__ = ys__n26449 & new_new_n16712__;
  assign new_new_n30765__ = ys__n26449 & new_new_n16714__;
  assign new_new_n30766__ = ~new_new_n30764__ & ~new_new_n30765__;
  assign new_new_n30767__ = ~new_new_n16715__ & ~new_new_n30766__;
  assign new_new_n30768__ = ~new_new_n30763__ & ~new_new_n30767__;
  assign new_new_n30769__ = ys__n602 & ~new_new_n30768__;
  assign ys__n26685 = new_new_n30762__ | new_new_n30769__;
  assign new_new_n30771__ = ~ys__n778 & ys__n26449;
  assign new_new_n30772__ = ys__n26449 & new_new_n16715__;
  assign new_new_n30773__ = ys__n26558 & ~new_new_n16715__;
  assign new_new_n30774__ = ~new_new_n30772__ & ~new_new_n30773__;
  assign new_new_n30775__ = ys__n778 & ~new_new_n30774__;
  assign new_new_n30776__ = ~new_new_n30771__ & ~new_new_n30775__;
  assign new_new_n30777__ = ~ys__n602 & ~new_new_n30776__;
  assign new_new_n30778__ = new_new_n16715__ & ~new_new_n30776__;
  assign new_new_n30779__ = ys__n26452 & new_new_n16712__;
  assign new_new_n30780__ = ys__n26452 & new_new_n16714__;
  assign new_new_n30781__ = ~new_new_n30779__ & ~new_new_n30780__;
  assign new_new_n30782__ = ~new_new_n16715__ & ~new_new_n30781__;
  assign new_new_n30783__ = ~new_new_n30778__ & ~new_new_n30782__;
  assign new_new_n30784__ = ys__n602 & ~new_new_n30783__;
  assign ys__n26687 = new_new_n30777__ | new_new_n30784__;
  assign new_new_n30786__ = ~ys__n778 & ys__n26452;
  assign new_new_n30787__ = ys__n26452 & new_new_n16715__;
  assign new_new_n30788__ = ys__n26559 & ~new_new_n16715__;
  assign new_new_n30789__ = ~new_new_n30787__ & ~new_new_n30788__;
  assign new_new_n30790__ = ys__n778 & ~new_new_n30789__;
  assign new_new_n30791__ = ~new_new_n30786__ & ~new_new_n30790__;
  assign new_new_n30792__ = ~ys__n602 & ~new_new_n30791__;
  assign new_new_n30793__ = new_new_n16715__ & ~new_new_n30791__;
  assign new_new_n30794__ = ys__n26455 & new_new_n16712__;
  assign new_new_n30795__ = ys__n26455 & new_new_n16714__;
  assign new_new_n30796__ = ~new_new_n30794__ & ~new_new_n30795__;
  assign new_new_n30797__ = ~new_new_n16715__ & ~new_new_n30796__;
  assign new_new_n30798__ = ~new_new_n30793__ & ~new_new_n30797__;
  assign new_new_n30799__ = ys__n602 & ~new_new_n30798__;
  assign ys__n26689 = new_new_n30792__ | new_new_n30799__;
  assign new_new_n30801__ = ~ys__n778 & ys__n26455;
  assign new_new_n30802__ = ys__n778 & ys__n26455;
  assign new_new_n30803__ = new_new_n16715__ & new_new_n30802__;
  assign new_new_n30804__ = ~new_new_n30801__ & ~new_new_n30803__;
  assign new_new_n30805__ = ~ys__n602 & ~new_new_n30804__;
  assign new_new_n30806__ = new_new_n16715__ & ~new_new_n30804__;
  assign new_new_n30807__ = ys__n26285 & new_new_n16712__;
  assign new_new_n30808__ = ys__n26285 & new_new_n16714__;
  assign new_new_n30809__ = ~new_new_n30807__ & ~new_new_n30808__;
  assign new_new_n30810__ = ~new_new_n16715__ & ~new_new_n30809__;
  assign new_new_n30811__ = ~new_new_n30806__ & ~new_new_n30810__;
  assign new_new_n30812__ = ys__n602 & ~new_new_n30811__;
  assign ys__n26691 = new_new_n30805__ | new_new_n30812__;
  assign new_new_n30814__ = ~ys__n778 & ys__n26285;
  assign new_new_n30815__ = ys__n26285 & new_new_n16715__;
  assign new_new_n30816__ = ys__n26560 & ~new_new_n16715__;
  assign new_new_n30817__ = ~new_new_n30815__ & ~new_new_n30816__;
  assign new_new_n30818__ = ys__n778 & ~new_new_n30817__;
  assign new_new_n30819__ = ~new_new_n30814__ & ~new_new_n30818__;
  assign new_new_n30820__ = ~ys__n602 & ~new_new_n30819__;
  assign new_new_n30821__ = new_new_n16715__ & ~new_new_n30819__;
  assign new_new_n30822__ = ys__n26460 & new_new_n16712__;
  assign new_new_n30823__ = ys__n26460 & new_new_n16714__;
  assign new_new_n30824__ = ~new_new_n30822__ & ~new_new_n30823__;
  assign new_new_n30825__ = ~new_new_n16715__ & ~new_new_n30824__;
  assign new_new_n30826__ = ~new_new_n30821__ & ~new_new_n30825__;
  assign new_new_n30827__ = ys__n602 & ~new_new_n30826__;
  assign ys__n26693 = new_new_n30820__ | new_new_n30827__;
  assign new_new_n30829__ = ~ys__n778 & ys__n26460;
  assign new_new_n30830__ = ys__n26460 & new_new_n16715__;
  assign new_new_n30831__ = ys__n26561 & ~new_new_n16715__;
  assign new_new_n30832__ = ~new_new_n30830__ & ~new_new_n30831__;
  assign new_new_n30833__ = ys__n778 & ~new_new_n30832__;
  assign new_new_n30834__ = ~new_new_n30829__ & ~new_new_n30833__;
  assign new_new_n30835__ = ~ys__n602 & ~new_new_n30834__;
  assign new_new_n30836__ = new_new_n16715__ & ~new_new_n30834__;
  assign new_new_n30837__ = ys__n26463 & new_new_n16712__;
  assign new_new_n30838__ = ys__n26463 & new_new_n16714__;
  assign new_new_n30839__ = ~new_new_n30837__ & ~new_new_n30838__;
  assign new_new_n30840__ = ~new_new_n16715__ & ~new_new_n30839__;
  assign new_new_n30841__ = ~new_new_n30836__ & ~new_new_n30840__;
  assign new_new_n30842__ = ys__n602 & ~new_new_n30841__;
  assign ys__n26695 = new_new_n30835__ | new_new_n30842__;
  assign new_new_n30844__ = ~ys__n778 & ys__n26463;
  assign new_new_n30845__ = ys__n778 & ys__n26463;
  assign new_new_n30846__ = new_new_n16715__ & new_new_n30845__;
  assign new_new_n30847__ = ~new_new_n30844__ & ~new_new_n30846__;
  assign new_new_n30848__ = ~ys__n602 & ~new_new_n30847__;
  assign new_new_n30849__ = new_new_n16715__ & ~new_new_n30847__;
  assign new_new_n30850__ = ys__n26466 & new_new_n16712__;
  assign new_new_n30851__ = ys__n26466 & new_new_n16714__;
  assign new_new_n30852__ = ~new_new_n30850__ & ~new_new_n30851__;
  assign new_new_n30853__ = ~new_new_n16715__ & ~new_new_n30852__;
  assign new_new_n30854__ = ~new_new_n30849__ & ~new_new_n30853__;
  assign new_new_n30855__ = ys__n602 & ~new_new_n30854__;
  assign ys__n26697 = new_new_n30848__ | new_new_n30855__;
  assign new_new_n30857__ = ~ys__n778 & ys__n26466;
  assign new_new_n30858__ = ys__n26466 & new_new_n16715__;
  assign new_new_n30859__ = ys__n26562 & ~new_new_n16715__;
  assign new_new_n30860__ = ~new_new_n30858__ & ~new_new_n30859__;
  assign new_new_n30861__ = ys__n778 & ~new_new_n30860__;
  assign new_new_n30862__ = ~new_new_n30857__ & ~new_new_n30861__;
  assign new_new_n30863__ = ~ys__n602 & ~new_new_n30862__;
  assign new_new_n30864__ = new_new_n16715__ & ~new_new_n30862__;
  assign new_new_n30865__ = ys__n26469 & new_new_n16712__;
  assign new_new_n30866__ = ys__n26469 & new_new_n16714__;
  assign new_new_n30867__ = ~new_new_n30865__ & ~new_new_n30866__;
  assign new_new_n30868__ = ~new_new_n16715__ & ~new_new_n30867__;
  assign new_new_n30869__ = ~new_new_n30864__ & ~new_new_n30868__;
  assign new_new_n30870__ = ys__n602 & ~new_new_n30869__;
  assign ys__n26699 = new_new_n30863__ | new_new_n30870__;
  assign new_new_n30872__ = ~ys__n778 & ys__n26469;
  assign new_new_n30873__ = ys__n26469 & new_new_n16715__;
  assign new_new_n30874__ = ys__n26563 & ~new_new_n16715__;
  assign new_new_n30875__ = ~new_new_n30873__ & ~new_new_n30874__;
  assign new_new_n30876__ = ys__n778 & ~new_new_n30875__;
  assign new_new_n30877__ = ~new_new_n30872__ & ~new_new_n30876__;
  assign new_new_n30878__ = ~ys__n602 & ~new_new_n30877__;
  assign new_new_n30879__ = new_new_n16715__ & ~new_new_n30877__;
  assign new_new_n30880__ = ys__n26472 & new_new_n16712__;
  assign new_new_n30881__ = ys__n26472 & new_new_n16714__;
  assign new_new_n30882__ = ~new_new_n30880__ & ~new_new_n30881__;
  assign new_new_n30883__ = ~new_new_n16715__ & ~new_new_n30882__;
  assign new_new_n30884__ = ~new_new_n30879__ & ~new_new_n30883__;
  assign new_new_n30885__ = ys__n602 & ~new_new_n30884__;
  assign ys__n26701 = new_new_n30878__ | new_new_n30885__;
  assign new_new_n30887__ = ~ys__n778 & ys__n26472;
  assign new_new_n30888__ = ys__n26472 & new_new_n16715__;
  assign new_new_n30889__ = ys__n26564 & ~new_new_n16715__;
  assign new_new_n30890__ = ~new_new_n30888__ & ~new_new_n30889__;
  assign new_new_n30891__ = ys__n778 & ~new_new_n30890__;
  assign new_new_n30892__ = ~new_new_n30887__ & ~new_new_n30891__;
  assign new_new_n30893__ = ~ys__n602 & ~new_new_n30892__;
  assign new_new_n30894__ = new_new_n16715__ & ~new_new_n30892__;
  assign new_new_n30895__ = ys__n26475 & new_new_n16712__;
  assign new_new_n30896__ = ys__n26475 & new_new_n16714__;
  assign new_new_n30897__ = ~new_new_n30895__ & ~new_new_n30896__;
  assign new_new_n30898__ = ~new_new_n16715__ & ~new_new_n30897__;
  assign new_new_n30899__ = ~new_new_n30894__ & ~new_new_n30898__;
  assign new_new_n30900__ = ys__n602 & ~new_new_n30899__;
  assign ys__n26703 = new_new_n30893__ | new_new_n30900__;
  assign new_new_n30902__ = ~ys__n778 & ys__n26475;
  assign new_new_n30903__ = ys__n26475 & new_new_n16715__;
  assign new_new_n30904__ = ys__n18173 & ~new_new_n16715__;
  assign new_new_n30905__ = ~new_new_n30903__ & ~new_new_n30904__;
  assign new_new_n30906__ = ys__n778 & ~new_new_n30905__;
  assign new_new_n30907__ = ~new_new_n30902__ & ~new_new_n30906__;
  assign new_new_n30908__ = ~ys__n602 & ~new_new_n30907__;
  assign new_new_n30909__ = new_new_n16715__ & ~new_new_n30907__;
  assign new_new_n30910__ = ys__n26478 & new_new_n16712__;
  assign new_new_n30911__ = ys__n26478 & new_new_n16714__;
  assign new_new_n30912__ = ~new_new_n30910__ & ~new_new_n30911__;
  assign new_new_n30913__ = ~new_new_n16715__ & ~new_new_n30912__;
  assign new_new_n30914__ = ~new_new_n30909__ & ~new_new_n30913__;
  assign new_new_n30915__ = ys__n602 & ~new_new_n30914__;
  assign ys__n26705 = new_new_n30908__ | new_new_n30915__;
  assign new_new_n30917__ = ~ys__n778 & ys__n26478;
  assign new_new_n30918__ = ys__n26478 & new_new_n16715__;
  assign new_new_n30919__ = ys__n26565 & ~new_new_n16715__;
  assign new_new_n30920__ = ~new_new_n30918__ & ~new_new_n30919__;
  assign new_new_n30921__ = ys__n778 & ~new_new_n30920__;
  assign new_new_n30922__ = ~new_new_n30917__ & ~new_new_n30921__;
  assign new_new_n30923__ = ~ys__n602 & ~new_new_n30922__;
  assign new_new_n30924__ = new_new_n16715__ & ~new_new_n30922__;
  assign new_new_n30925__ = ys__n26481 & new_new_n16712__;
  assign new_new_n30926__ = ys__n26481 & new_new_n16714__;
  assign new_new_n30927__ = ~new_new_n30925__ & ~new_new_n30926__;
  assign new_new_n30928__ = ~new_new_n16715__ & ~new_new_n30927__;
  assign new_new_n30929__ = ~new_new_n30924__ & ~new_new_n30928__;
  assign new_new_n30930__ = ys__n602 & ~new_new_n30929__;
  assign ys__n26707 = new_new_n30923__ | new_new_n30930__;
  assign new_new_n30932__ = ~ys__n778 & ys__n26481;
  assign new_new_n30933__ = ys__n26481 & new_new_n16715__;
  assign new_new_n30934__ = ~new_new_n16715__ & ys__n26566;
  assign new_new_n30935__ = ~new_new_n30933__ & ~new_new_n30934__;
  assign new_new_n30936__ = ys__n778 & ~new_new_n30935__;
  assign new_new_n30937__ = ~new_new_n30932__ & ~new_new_n30936__;
  assign new_new_n30938__ = ~ys__n602 & ~new_new_n30937__;
  assign new_new_n30939__ = new_new_n16715__ & ~new_new_n30937__;
  assign new_new_n30940__ = ys__n26484 & new_new_n16712__;
  assign new_new_n30941__ = ys__n26484 & new_new_n16714__;
  assign new_new_n30942__ = ~new_new_n30940__ & ~new_new_n30941__;
  assign new_new_n30943__ = ~new_new_n16715__ & ~new_new_n30942__;
  assign new_new_n30944__ = ~new_new_n30939__ & ~new_new_n30943__;
  assign new_new_n30945__ = ys__n602 & ~new_new_n30944__;
  assign ys__n26709 = new_new_n30938__ | new_new_n30945__;
  assign new_new_n30947__ = ~ys__n778 & ys__n26484;
  assign new_new_n30948__ = ys__n26484 & new_new_n16715__;
  assign new_new_n30949__ = ys__n26567 & ~new_new_n16715__;
  assign new_new_n30950__ = ~new_new_n30948__ & ~new_new_n30949__;
  assign new_new_n30951__ = ys__n778 & ~new_new_n30950__;
  assign new_new_n30952__ = ~new_new_n30947__ & ~new_new_n30951__;
  assign new_new_n30953__ = ~ys__n602 & ~new_new_n30952__;
  assign new_new_n30954__ = new_new_n16715__ & ~new_new_n30952__;
  assign new_new_n30955__ = ys__n26487 & new_new_n16712__;
  assign new_new_n30956__ = ys__n26487 & new_new_n16714__;
  assign new_new_n30957__ = ~new_new_n30955__ & ~new_new_n30956__;
  assign new_new_n30958__ = ~new_new_n16715__ & ~new_new_n30957__;
  assign new_new_n30959__ = ~new_new_n30954__ & ~new_new_n30958__;
  assign new_new_n30960__ = ys__n602 & ~new_new_n30959__;
  assign ys__n26711 = new_new_n30953__ | new_new_n30960__;
  assign new_new_n30962__ = ~ys__n778 & ys__n26487;
  assign new_new_n30963__ = ys__n26487 & new_new_n16715__;
  assign new_new_n30964__ = new_new_n16715__ & ~new_new_n30963__;
  assign new_new_n30965__ = ys__n778 & ~new_new_n30964__;
  assign new_new_n30966__ = ~new_new_n30962__ & ~new_new_n30965__;
  assign new_new_n30967__ = ~ys__n602 & ~new_new_n30966__;
  assign new_new_n30968__ = new_new_n16715__ & ~new_new_n30966__;
  assign new_new_n30969__ = ys__n26490 & new_new_n16712__;
  assign new_new_n30970__ = ys__n26490 & new_new_n16714__;
  assign new_new_n30971__ = ~new_new_n30969__ & ~new_new_n30970__;
  assign new_new_n30972__ = ~new_new_n16715__ & ~new_new_n30971__;
  assign new_new_n30973__ = ~new_new_n30968__ & ~new_new_n30972__;
  assign new_new_n30974__ = ys__n602 & ~new_new_n30973__;
  assign ys__n26713 = new_new_n30967__ | new_new_n30974__;
  assign new_new_n30976__ = ~ys__n778 & ys__n26490;
  assign new_new_n30977__ = ys__n26490 & new_new_n16715__;
  assign new_new_n30978__ = ys__n26568 & ~new_new_n16715__;
  assign new_new_n30979__ = ~new_new_n30977__ & ~new_new_n30978__;
  assign new_new_n30980__ = ys__n778 & ~new_new_n30979__;
  assign new_new_n30981__ = ~new_new_n30976__ & ~new_new_n30980__;
  assign new_new_n30982__ = ~ys__n602 & ~new_new_n30981__;
  assign new_new_n30983__ = new_new_n16715__ & ~new_new_n30981__;
  assign new_new_n30984__ = ys__n26493 & new_new_n16712__;
  assign new_new_n30985__ = ys__n26493 & new_new_n16714__;
  assign new_new_n30986__ = ~new_new_n30984__ & ~new_new_n30985__;
  assign new_new_n30987__ = ~new_new_n16715__ & ~new_new_n30986__;
  assign new_new_n30988__ = ~new_new_n30983__ & ~new_new_n30987__;
  assign new_new_n30989__ = ys__n602 & ~new_new_n30988__;
  assign ys__n26715 = new_new_n30982__ | new_new_n30989__;
  assign new_new_n30991__ = ~ys__n778 & ys__n26493;
  assign new_new_n30992__ = ys__n26493 & new_new_n16715__;
  assign new_new_n30993__ = ys__n26569 & ~new_new_n16715__;
  assign new_new_n30994__ = ~new_new_n30992__ & ~new_new_n30993__;
  assign new_new_n30995__ = ys__n778 & ~new_new_n30994__;
  assign new_new_n30996__ = ~new_new_n30991__ & ~new_new_n30995__;
  assign new_new_n30997__ = ~ys__n602 & ~new_new_n30996__;
  assign new_new_n30998__ = new_new_n16715__ & ~new_new_n30996__;
  assign new_new_n30999__ = ys__n26496 & new_new_n16712__;
  assign new_new_n31000__ = ys__n26496 & new_new_n16714__;
  assign new_new_n31001__ = ~new_new_n30999__ & ~new_new_n31000__;
  assign new_new_n31002__ = ~new_new_n16715__ & ~new_new_n31001__;
  assign new_new_n31003__ = ~new_new_n30998__ & ~new_new_n31002__;
  assign new_new_n31004__ = ys__n602 & ~new_new_n31003__;
  assign ys__n26717 = new_new_n30997__ | new_new_n31004__;
  assign new_new_n31006__ = ~ys__n778 & ys__n26496;
  assign new_new_n31007__ = ys__n26496 & new_new_n16715__;
  assign new_new_n31008__ = ys__n26570 & ~new_new_n16715__;
  assign new_new_n31009__ = ~new_new_n31007__ & ~new_new_n31008__;
  assign new_new_n31010__ = ys__n778 & ~new_new_n31009__;
  assign new_new_n31011__ = ~new_new_n31006__ & ~new_new_n31010__;
  assign new_new_n31012__ = ~ys__n602 & ~new_new_n31011__;
  assign new_new_n31013__ = new_new_n16715__ & ~new_new_n31011__;
  assign new_new_n31014__ = ys__n26499 & new_new_n16712__;
  assign new_new_n31015__ = ys__n26499 & new_new_n16714__;
  assign new_new_n31016__ = ~new_new_n31014__ & ~new_new_n31015__;
  assign new_new_n31017__ = ~new_new_n16715__ & ~new_new_n31016__;
  assign new_new_n31018__ = ~new_new_n31013__ & ~new_new_n31017__;
  assign new_new_n31019__ = ys__n602 & ~new_new_n31018__;
  assign ys__n26719 = new_new_n31012__ | new_new_n31019__;
  assign new_new_n31021__ = ~ys__n778 & ys__n26499;
  assign new_new_n31022__ = ys__n26499 & new_new_n16715__;
  assign new_new_n31023__ = ys__n26571 & ~new_new_n16715__;
  assign new_new_n31024__ = ~new_new_n31022__ & ~new_new_n31023__;
  assign new_new_n31025__ = ys__n778 & ~new_new_n31024__;
  assign new_new_n31026__ = ~new_new_n31021__ & ~new_new_n31025__;
  assign new_new_n31027__ = ~ys__n602 & ~new_new_n31026__;
  assign new_new_n31028__ = new_new_n16715__ & ~new_new_n31026__;
  assign new_new_n31029__ = ys__n26502 & new_new_n16712__;
  assign new_new_n31030__ = ys__n26502 & new_new_n16714__;
  assign new_new_n31031__ = ~new_new_n31029__ & ~new_new_n31030__;
  assign new_new_n31032__ = ~new_new_n16715__ & ~new_new_n31031__;
  assign new_new_n31033__ = ~new_new_n31028__ & ~new_new_n31032__;
  assign new_new_n31034__ = ys__n602 & ~new_new_n31033__;
  assign ys__n26721 = new_new_n31027__ | new_new_n31034__;
  assign new_new_n31036__ = ~ys__n778 & ys__n26502;
  assign new_new_n31037__ = ys__n778 & ys__n26502;
  assign new_new_n31038__ = new_new_n16715__ & new_new_n31037__;
  assign new_new_n31039__ = ~new_new_n31036__ & ~new_new_n31038__;
  assign new_new_n31040__ = ~ys__n602 & ~new_new_n31039__;
  assign new_new_n31041__ = new_new_n16715__ & ~new_new_n31039__;
  assign new_new_n31042__ = ys__n26505 & new_new_n16712__;
  assign new_new_n31043__ = ys__n26505 & new_new_n16714__;
  assign new_new_n31044__ = ~new_new_n31042__ & ~new_new_n31043__;
  assign new_new_n31045__ = ~new_new_n16715__ & ~new_new_n31044__;
  assign new_new_n31046__ = ~new_new_n31041__ & ~new_new_n31045__;
  assign new_new_n31047__ = ys__n602 & ~new_new_n31046__;
  assign ys__n26723 = new_new_n31040__ | new_new_n31047__;
  assign new_new_n31049__ = ~ys__n778 & ys__n26505;
  assign new_new_n31050__ = ys__n778 & ys__n26505;
  assign new_new_n31051__ = new_new_n16715__ & new_new_n31050__;
  assign new_new_n31052__ = ~new_new_n31049__ & ~new_new_n31051__;
  assign new_new_n31053__ = ~ys__n602 & ~new_new_n31052__;
  assign new_new_n31054__ = new_new_n16715__ & ~new_new_n31052__;
  assign new_new_n31055__ = ys__n26508 & new_new_n16712__;
  assign new_new_n31056__ = ys__n26508 & new_new_n16714__;
  assign new_new_n31057__ = ~new_new_n31055__ & ~new_new_n31056__;
  assign new_new_n31058__ = ~new_new_n16715__ & ~new_new_n31057__;
  assign new_new_n31059__ = ~new_new_n31054__ & ~new_new_n31058__;
  assign new_new_n31060__ = ys__n602 & ~new_new_n31059__;
  assign ys__n26725 = new_new_n31053__ | new_new_n31060__;
  assign new_new_n31062__ = ~ys__n778 & ys__n26508;
  assign new_new_n31063__ = ys__n778 & ys__n26508;
  assign new_new_n31064__ = new_new_n16715__ & new_new_n31063__;
  assign new_new_n31065__ = ~new_new_n31062__ & ~new_new_n31064__;
  assign new_new_n31066__ = ~ys__n602 & ~new_new_n31065__;
  assign new_new_n31067__ = new_new_n16715__ & ~new_new_n31065__;
  assign new_new_n31068__ = ys__n26511 & new_new_n16712__;
  assign new_new_n31069__ = ys__n26511 & new_new_n16714__;
  assign new_new_n31070__ = ~new_new_n31068__ & ~new_new_n31069__;
  assign new_new_n31071__ = ~new_new_n16715__ & ~new_new_n31070__;
  assign new_new_n31072__ = ~new_new_n31067__ & ~new_new_n31071__;
  assign new_new_n31073__ = ys__n602 & ~new_new_n31072__;
  assign ys__n26727 = new_new_n31066__ | new_new_n31073__;
  assign new_new_n31075__ = ~ys__n778 & ys__n26511;
  assign new_new_n31076__ = ys__n778 & ys__n26511;
  assign new_new_n31077__ = new_new_n16715__ & new_new_n31076__;
  assign new_new_n31078__ = ~new_new_n31075__ & ~new_new_n31077__;
  assign new_new_n31079__ = ~ys__n602 & ~new_new_n31078__;
  assign new_new_n31080__ = new_new_n16715__ & ~new_new_n31078__;
  assign new_new_n31081__ = ys__n26514 & new_new_n16712__;
  assign new_new_n31082__ = ys__n26514 & new_new_n16714__;
  assign new_new_n31083__ = ~new_new_n31081__ & ~new_new_n31082__;
  assign new_new_n31084__ = ~new_new_n16715__ & ~new_new_n31083__;
  assign new_new_n31085__ = ~new_new_n31080__ & ~new_new_n31084__;
  assign new_new_n31086__ = ys__n602 & ~new_new_n31085__;
  assign ys__n26729 = new_new_n31079__ | new_new_n31086__;
  assign new_new_n31088__ = ~ys__n778 & ys__n26514;
  assign new_new_n31089__ = ys__n778 & ys__n26514;
  assign new_new_n31090__ = new_new_n16715__ & new_new_n31089__;
  assign new_new_n31091__ = ~new_new_n31088__ & ~new_new_n31090__;
  assign new_new_n31092__ = ~ys__n602 & ~new_new_n31091__;
  assign new_new_n31093__ = new_new_n16715__ & ~new_new_n31091__;
  assign new_new_n31094__ = ys__n26517 & new_new_n16712__;
  assign new_new_n31095__ = ys__n26517 & new_new_n16714__;
  assign new_new_n31096__ = ~new_new_n31094__ & ~new_new_n31095__;
  assign new_new_n31097__ = ~new_new_n16715__ & ~new_new_n31096__;
  assign new_new_n31098__ = ~new_new_n31093__ & ~new_new_n31097__;
  assign new_new_n31099__ = ys__n602 & ~new_new_n31098__;
  assign ys__n26731 = new_new_n31092__ | new_new_n31099__;
  assign new_new_n31101__ = ~ys__n778 & ys__n26517;
  assign new_new_n31102__ = ys__n26517 & new_new_n16715__;
  assign new_new_n31103__ = ys__n26572 & ~new_new_n16715__;
  assign new_new_n31104__ = ~new_new_n31102__ & ~new_new_n31103__;
  assign new_new_n31105__ = ys__n778 & ~new_new_n31104__;
  assign new_new_n31106__ = ~new_new_n31101__ & ~new_new_n31105__;
  assign new_new_n31107__ = ~ys__n602 & ~new_new_n31106__;
  assign new_new_n31108__ = new_new_n16715__ & ~new_new_n31106__;
  assign new_new_n31109__ = ys__n25980 & new_new_n16712__;
  assign new_new_n31110__ = new_new_n16714__ & new_new_n30646__;
  assign new_new_n31111__ = ~new_new_n31109__ & ~new_new_n31110__;
  assign new_new_n31112__ = ~new_new_n16715__ & ~new_new_n31111__;
  assign new_new_n31113__ = ~new_new_n31108__ & ~new_new_n31112__;
  assign new_new_n31114__ = ys__n602 & ~new_new_n31113__;
  assign ys__n26733 = new_new_n31107__ | new_new_n31114__;
  assign new_new_n31116__ = ~ys__n778 & ys__n26359;
  assign new_new_n31117__ = ys__n26359 & new_new_n16723__;
  assign new_new_n31118__ = ys__n6112 & ~ys__n18173;
  assign new_new_n31119__ = ys__n18173 & ys__n18829;
  assign new_new_n31120__ = ~new_new_n31118__ & ~new_new_n31119__;
  assign new_new_n31121__ = ~new_new_n16723__ & ~new_new_n31120__;
  assign new_new_n31122__ = ~new_new_n31117__ & ~new_new_n31121__;
  assign new_new_n31123__ = ys__n778 & ~new_new_n31122__;
  assign new_new_n31124__ = ~new_new_n31116__ & ~new_new_n31123__;
  assign new_new_n31125__ = ~ys__n602 & ~new_new_n31124__;
  assign new_new_n31126__ = new_new_n16723__ & ~new_new_n31124__;
  assign new_new_n31127__ = ys__n26362 & ~new_new_n16723__;
  assign new_new_n31128__ = ~new_new_n31126__ & ~new_new_n31127__;
  assign new_new_n31129__ = ys__n602 & ~new_new_n31128__;
  assign ys__n26734 = new_new_n31125__ | new_new_n31129__;
  assign new_new_n31131__ = ~ys__n778 & ys__n26362;
  assign new_new_n31132__ = ys__n26362 & new_new_n16723__;
  assign new_new_n31133__ = ys__n6113 & ~ys__n18173;
  assign new_new_n31134__ = ys__n18173 & ys__n18831;
  assign new_new_n31135__ = ~new_new_n31133__ & ~new_new_n31134__;
  assign new_new_n31136__ = ~new_new_n16723__ & ~new_new_n31135__;
  assign new_new_n31137__ = ~new_new_n31132__ & ~new_new_n31136__;
  assign new_new_n31138__ = ys__n778 & ~new_new_n31137__;
  assign new_new_n31139__ = ~new_new_n31131__ & ~new_new_n31138__;
  assign new_new_n31140__ = ~ys__n602 & ~new_new_n31139__;
  assign new_new_n31141__ = new_new_n16723__ & ~new_new_n31139__;
  assign new_new_n31142__ = ys__n26161 & ~new_new_n16723__;
  assign new_new_n31143__ = ~new_new_n31141__ & ~new_new_n31142__;
  assign new_new_n31144__ = ys__n602 & ~new_new_n31143__;
  assign ys__n26735 = new_new_n31140__ | new_new_n31144__;
  assign new_new_n31146__ = ~ys__n778 & ys__n26161;
  assign new_new_n31147__ = ys__n26161 & new_new_n16723__;
  assign new_new_n31148__ = ys__n172 & ~ys__n18173;
  assign new_new_n31149__ = ys__n18173 & ys__n18833;
  assign new_new_n31150__ = ~new_new_n31148__ & ~new_new_n31149__;
  assign new_new_n31151__ = ~new_new_n16723__ & ~new_new_n31150__;
  assign new_new_n31152__ = ~new_new_n31147__ & ~new_new_n31151__;
  assign new_new_n31153__ = ys__n778 & ~new_new_n31152__;
  assign new_new_n31154__ = ~new_new_n31146__ & ~new_new_n31153__;
  assign new_new_n31155__ = ~ys__n602 & ~new_new_n31154__;
  assign new_new_n31156__ = new_new_n16723__ & ~new_new_n31154__;
  assign new_new_n31157__ = ys__n26162 & ~new_new_n16723__;
  assign new_new_n31158__ = ~new_new_n31156__ & ~new_new_n31157__;
  assign new_new_n31159__ = ys__n602 & ~new_new_n31158__;
  assign ys__n26736 = new_new_n31155__ | new_new_n31159__;
  assign new_new_n31161__ = ~ys__n778 & ys__n26162;
  assign new_new_n31162__ = ys__n26162 & new_new_n16723__;
  assign new_new_n31163__ = ys__n338 & ~ys__n18173;
  assign new_new_n31164__ = ys__n18173 & ys__n18835;
  assign new_new_n31165__ = ~new_new_n31163__ & ~new_new_n31164__;
  assign new_new_n31166__ = ~new_new_n16723__ & ~new_new_n31165__;
  assign new_new_n31167__ = ~new_new_n31162__ & ~new_new_n31166__;
  assign new_new_n31168__ = ys__n778 & ~new_new_n31167__;
  assign new_new_n31169__ = ~new_new_n31161__ & ~new_new_n31168__;
  assign new_new_n31170__ = ~ys__n602 & ~new_new_n31169__;
  assign new_new_n31171__ = new_new_n16723__ & ~new_new_n31169__;
  assign new_new_n31172__ = ys__n26164 & ~new_new_n16723__;
  assign new_new_n31173__ = ~new_new_n31171__ & ~new_new_n31172__;
  assign new_new_n31174__ = ys__n602 & ~new_new_n31173__;
  assign ys__n26737 = new_new_n31170__ | new_new_n31174__;
  assign new_new_n31176__ = ~ys__n778 & ys__n26164;
  assign new_new_n31177__ = ys__n26164 & new_new_n16723__;
  assign new_new_n31178__ = ys__n22 & ~ys__n18173;
  assign new_new_n31179__ = ys__n18173 & ys__n18837;
  assign new_new_n31180__ = ~new_new_n31178__ & ~new_new_n31179__;
  assign new_new_n31181__ = ~new_new_n16723__ & ~new_new_n31180__;
  assign new_new_n31182__ = ~new_new_n31177__ & ~new_new_n31181__;
  assign new_new_n31183__ = ys__n778 & ~new_new_n31182__;
  assign new_new_n31184__ = ~new_new_n31176__ & ~new_new_n31183__;
  assign new_new_n31185__ = ~ys__n602 & ~new_new_n31184__;
  assign new_new_n31186__ = new_new_n16723__ & ~new_new_n31184__;
  assign new_new_n31187__ = ys__n26166 & ~new_new_n16723__;
  assign new_new_n31188__ = ~new_new_n31186__ & ~new_new_n31187__;
  assign new_new_n31189__ = ys__n602 & ~new_new_n31188__;
  assign ys__n26738 = new_new_n31185__ | new_new_n31189__;
  assign new_new_n31191__ = ~ys__n778 & ys__n26166;
  assign new_new_n31192__ = ys__n26166 & new_new_n16723__;
  assign new_new_n31193__ = ys__n316 & ~ys__n18173;
  assign new_new_n31194__ = ys__n18173 & ys__n18839;
  assign new_new_n31195__ = ~new_new_n31193__ & ~new_new_n31194__;
  assign new_new_n31196__ = ~new_new_n16723__ & ~new_new_n31195__;
  assign new_new_n31197__ = ~new_new_n31192__ & ~new_new_n31196__;
  assign new_new_n31198__ = ys__n778 & ~new_new_n31197__;
  assign new_new_n31199__ = ~new_new_n31191__ & ~new_new_n31198__;
  assign new_new_n31200__ = ~ys__n602 & ~new_new_n31199__;
  assign new_new_n31201__ = new_new_n16723__ & ~new_new_n31199__;
  assign new_new_n31202__ = ys__n26168 & ~new_new_n16723__;
  assign new_new_n31203__ = ~new_new_n31201__ & ~new_new_n31202__;
  assign new_new_n31204__ = ys__n602 & ~new_new_n31203__;
  assign ys__n26739 = new_new_n31200__ | new_new_n31204__;
  assign new_new_n31206__ = ~ys__n778 & ys__n26168;
  assign new_new_n31207__ = ys__n26168 & new_new_n16723__;
  assign new_new_n31208__ = ys__n6115 & ~ys__n18173;
  assign new_new_n31209__ = ys__n18173 & ys__n18841;
  assign new_new_n31210__ = ~new_new_n31208__ & ~new_new_n31209__;
  assign new_new_n31211__ = ~new_new_n16723__ & ~new_new_n31210__;
  assign new_new_n31212__ = ~new_new_n31207__ & ~new_new_n31211__;
  assign new_new_n31213__ = ys__n778 & ~new_new_n31212__;
  assign new_new_n31214__ = ~new_new_n31206__ & ~new_new_n31213__;
  assign new_new_n31215__ = ~ys__n602 & ~new_new_n31214__;
  assign new_new_n31216__ = new_new_n16723__ & ~new_new_n31214__;
  assign new_new_n31217__ = ys__n26170 & ~new_new_n16723__;
  assign new_new_n31218__ = ~new_new_n31216__ & ~new_new_n31217__;
  assign new_new_n31219__ = ys__n602 & ~new_new_n31218__;
  assign ys__n26740 = new_new_n31215__ | new_new_n31219__;
  assign new_new_n31221__ = ~ys__n778 & ys__n26170;
  assign new_new_n31222__ = ys__n26170 & new_new_n16723__;
  assign new_new_n31223__ = ys__n44 & ~ys__n18173;
  assign new_new_n31224__ = ys__n18173 & ys__n18843;
  assign new_new_n31225__ = ~new_new_n31223__ & ~new_new_n31224__;
  assign new_new_n31226__ = ~new_new_n16723__ & ~new_new_n31225__;
  assign new_new_n31227__ = ~new_new_n31222__ & ~new_new_n31226__;
  assign new_new_n31228__ = ys__n778 & ~new_new_n31227__;
  assign new_new_n31229__ = ~new_new_n31221__ & ~new_new_n31228__;
  assign new_new_n31230__ = ~ys__n602 & ~new_new_n31229__;
  assign new_new_n31231__ = new_new_n16723__ & ~new_new_n31229__;
  assign new_new_n31232__ = ys__n26172 & ~new_new_n16723__;
  assign new_new_n31233__ = ~new_new_n31231__ & ~new_new_n31232__;
  assign new_new_n31234__ = ys__n602 & ~new_new_n31233__;
  assign ys__n26741 = new_new_n31230__ | new_new_n31234__;
  assign new_new_n31236__ = ~ys__n778 & ys__n26172;
  assign new_new_n31237__ = ys__n26172 & new_new_n16723__;
  assign new_new_n31238__ = ys__n340 & ~ys__n18173;
  assign new_new_n31239__ = ys__n18173 & ys__n18845;
  assign new_new_n31240__ = ~new_new_n31238__ & ~new_new_n31239__;
  assign new_new_n31241__ = ~new_new_n16723__ & ~new_new_n31240__;
  assign new_new_n31242__ = ~new_new_n31237__ & ~new_new_n31241__;
  assign new_new_n31243__ = ys__n778 & ~new_new_n31242__;
  assign new_new_n31244__ = ~new_new_n31236__ & ~new_new_n31243__;
  assign new_new_n31245__ = ~ys__n602 & ~new_new_n31244__;
  assign new_new_n31246__ = new_new_n16723__ & ~new_new_n31244__;
  assign new_new_n31247__ = ys__n26174 & ~new_new_n16723__;
  assign new_new_n31248__ = ~new_new_n31246__ & ~new_new_n31247__;
  assign new_new_n31249__ = ys__n602 & ~new_new_n31248__;
  assign ys__n26742 = new_new_n31245__ | new_new_n31249__;
  assign new_new_n31251__ = ~ys__n778 & ys__n26174;
  assign new_new_n31252__ = ys__n26174 & new_new_n16723__;
  assign new_new_n31253__ = ys__n46 & ~ys__n18173;
  assign new_new_n31254__ = ys__n18173 & ys__n18847;
  assign new_new_n31255__ = ~new_new_n31253__ & ~new_new_n31254__;
  assign new_new_n31256__ = ~new_new_n16723__ & ~new_new_n31255__;
  assign new_new_n31257__ = ~new_new_n31252__ & ~new_new_n31256__;
  assign new_new_n31258__ = ys__n778 & ~new_new_n31257__;
  assign new_new_n31259__ = ~new_new_n31251__ & ~new_new_n31258__;
  assign new_new_n31260__ = ~ys__n602 & ~new_new_n31259__;
  assign new_new_n31261__ = new_new_n16723__ & ~new_new_n31259__;
  assign new_new_n31262__ = ys__n26176 & ~new_new_n16723__;
  assign new_new_n31263__ = ~new_new_n31261__ & ~new_new_n31262__;
  assign new_new_n31264__ = ys__n602 & ~new_new_n31263__;
  assign ys__n26743 = new_new_n31260__ | new_new_n31264__;
  assign new_new_n31266__ = ~ys__n778 & ys__n26176;
  assign new_new_n31267__ = ys__n26176 & new_new_n16723__;
  assign new_new_n31268__ = ys__n6118 & ~ys__n18173;
  assign new_new_n31269__ = ys__n18173 & ys__n18849;
  assign new_new_n31270__ = ~new_new_n31268__ & ~new_new_n31269__;
  assign new_new_n31271__ = ~new_new_n16723__ & ~new_new_n31270__;
  assign new_new_n31272__ = ~new_new_n31267__ & ~new_new_n31271__;
  assign new_new_n31273__ = ys__n778 & ~new_new_n31272__;
  assign new_new_n31274__ = ~new_new_n31266__ & ~new_new_n31273__;
  assign new_new_n31275__ = ~ys__n602 & ~new_new_n31274__;
  assign new_new_n31276__ = new_new_n16723__ & ~new_new_n31274__;
  assign new_new_n31277__ = ys__n26178 & ~new_new_n16723__;
  assign new_new_n31278__ = ~new_new_n31276__ & ~new_new_n31277__;
  assign new_new_n31279__ = ys__n602 & ~new_new_n31278__;
  assign ys__n26744 = new_new_n31275__ | new_new_n31279__;
  assign new_new_n31281__ = ~ys__n778 & ys__n26178;
  assign new_new_n31282__ = ys__n26178 & new_new_n16723__;
  assign new_new_n31283__ = ys__n6119 & ~ys__n18173;
  assign new_new_n31284__ = ys__n18173 & ys__n18851;
  assign new_new_n31285__ = ~new_new_n31283__ & ~new_new_n31284__;
  assign new_new_n31286__ = ~new_new_n16723__ & ~new_new_n31285__;
  assign new_new_n31287__ = ~new_new_n31282__ & ~new_new_n31286__;
  assign new_new_n31288__ = ys__n778 & ~new_new_n31287__;
  assign new_new_n31289__ = ~new_new_n31281__ & ~new_new_n31288__;
  assign new_new_n31290__ = ~ys__n602 & ~new_new_n31289__;
  assign new_new_n31291__ = new_new_n16723__ & ~new_new_n31289__;
  assign new_new_n31292__ = ys__n26180 & ~new_new_n16723__;
  assign new_new_n31293__ = ~new_new_n31291__ & ~new_new_n31292__;
  assign new_new_n31294__ = ys__n602 & ~new_new_n31293__;
  assign ys__n26745 = new_new_n31290__ | new_new_n31294__;
  assign new_new_n31296__ = ~ys__n778 & ys__n26180;
  assign new_new_n31297__ = ys__n26180 & new_new_n16723__;
  assign new_new_n31298__ = ys__n6120 & ~ys__n18173;
  assign new_new_n31299__ = ys__n18173 & ys__n18853;
  assign new_new_n31300__ = ~new_new_n31298__ & ~new_new_n31299__;
  assign new_new_n31301__ = ~new_new_n16723__ & ~new_new_n31300__;
  assign new_new_n31302__ = ~new_new_n31297__ & ~new_new_n31301__;
  assign new_new_n31303__ = ys__n778 & ~new_new_n31302__;
  assign new_new_n31304__ = ~new_new_n31296__ & ~new_new_n31303__;
  assign new_new_n31305__ = ~ys__n602 & ~new_new_n31304__;
  assign new_new_n31306__ = new_new_n16723__ & ~new_new_n31304__;
  assign new_new_n31307__ = ys__n26182 & ~new_new_n16723__;
  assign new_new_n31308__ = ~new_new_n31306__ & ~new_new_n31307__;
  assign new_new_n31309__ = ys__n602 & ~new_new_n31308__;
  assign ys__n26746 = new_new_n31305__ | new_new_n31309__;
  assign new_new_n31311__ = ~ys__n778 & ys__n26182;
  assign new_new_n31312__ = ys__n26182 & new_new_n16723__;
  assign new_new_n31313__ = ys__n6121 & ~ys__n18173;
  assign new_new_n31314__ = ys__n18173 & ys__n18855;
  assign new_new_n31315__ = ~new_new_n31313__ & ~new_new_n31314__;
  assign new_new_n31316__ = ~new_new_n16723__ & ~new_new_n31315__;
  assign new_new_n31317__ = ~new_new_n31312__ & ~new_new_n31316__;
  assign new_new_n31318__ = ys__n778 & ~new_new_n31317__;
  assign new_new_n31319__ = ~new_new_n31311__ & ~new_new_n31318__;
  assign new_new_n31320__ = ~ys__n602 & ~new_new_n31319__;
  assign new_new_n31321__ = new_new_n16723__ & ~new_new_n31319__;
  assign new_new_n31322__ = ys__n26184 & ~new_new_n16723__;
  assign new_new_n31323__ = ~new_new_n31321__ & ~new_new_n31322__;
  assign new_new_n31324__ = ys__n602 & ~new_new_n31323__;
  assign ys__n26747 = new_new_n31320__ | new_new_n31324__;
  assign new_new_n31326__ = ~ys__n778 & ys__n26184;
  assign new_new_n31327__ = ys__n26184 & new_new_n16723__;
  assign new_new_n31328__ = ys__n6123 & ~ys__n18173;
  assign new_new_n31329__ = ys__n18173 & ys__n18857;
  assign new_new_n31330__ = ~new_new_n31328__ & ~new_new_n31329__;
  assign new_new_n31331__ = ~new_new_n16723__ & ~new_new_n31330__;
  assign new_new_n31332__ = ~new_new_n31327__ & ~new_new_n31331__;
  assign new_new_n31333__ = ys__n778 & ~new_new_n31332__;
  assign new_new_n31334__ = ~new_new_n31326__ & ~new_new_n31333__;
  assign new_new_n31335__ = ~ys__n602 & ~new_new_n31334__;
  assign new_new_n31336__ = new_new_n16723__ & ~new_new_n31334__;
  assign new_new_n31337__ = ys__n26186 & ~new_new_n16723__;
  assign new_new_n31338__ = ~new_new_n31336__ & ~new_new_n31337__;
  assign new_new_n31339__ = ys__n602 & ~new_new_n31338__;
  assign ys__n26748 = new_new_n31335__ | new_new_n31339__;
  assign new_new_n31341__ = ~ys__n778 & ys__n26186;
  assign new_new_n31342__ = ys__n26186 & new_new_n16723__;
  assign new_new_n31343__ = ys__n6124 & ~ys__n18173;
  assign new_new_n31344__ = ys__n18173 & ys__n18859;
  assign new_new_n31345__ = ~new_new_n31343__ & ~new_new_n31344__;
  assign new_new_n31346__ = ~new_new_n16723__ & ~new_new_n31345__;
  assign new_new_n31347__ = ~new_new_n31342__ & ~new_new_n31346__;
  assign new_new_n31348__ = ys__n778 & ~new_new_n31347__;
  assign new_new_n31349__ = ~new_new_n31341__ & ~new_new_n31348__;
  assign new_new_n31350__ = ~ys__n602 & ~new_new_n31349__;
  assign new_new_n31351__ = new_new_n16723__ & ~new_new_n31349__;
  assign new_new_n31352__ = ys__n26188 & ~new_new_n16723__;
  assign new_new_n31353__ = ~new_new_n31351__ & ~new_new_n31352__;
  assign new_new_n31354__ = ys__n602 & ~new_new_n31353__;
  assign ys__n26749 = new_new_n31350__ | new_new_n31354__;
  assign new_new_n31356__ = ~ys__n778 & ys__n26188;
  assign new_new_n31357__ = ys__n26188 & new_new_n16723__;
  assign new_new_n31358__ = ys__n6126 & ~ys__n18173;
  assign new_new_n31359__ = ys__n18173 & ys__n18861;
  assign new_new_n31360__ = ~new_new_n31358__ & ~new_new_n31359__;
  assign new_new_n31361__ = ~new_new_n16723__ & ~new_new_n31360__;
  assign new_new_n31362__ = ~new_new_n31357__ & ~new_new_n31361__;
  assign new_new_n31363__ = ys__n778 & ~new_new_n31362__;
  assign new_new_n31364__ = ~new_new_n31356__ & ~new_new_n31363__;
  assign new_new_n31365__ = ~ys__n602 & ~new_new_n31364__;
  assign new_new_n31366__ = new_new_n16723__ & ~new_new_n31364__;
  assign new_new_n31367__ = ys__n26190 & ~new_new_n16723__;
  assign new_new_n31368__ = ~new_new_n31366__ & ~new_new_n31367__;
  assign new_new_n31369__ = ys__n602 & ~new_new_n31368__;
  assign ys__n26750 = new_new_n31365__ | new_new_n31369__;
  assign new_new_n31371__ = ~ys__n778 & ys__n26190;
  assign new_new_n31372__ = ys__n26190 & new_new_n16723__;
  assign new_new_n31373__ = ys__n6127 & ~ys__n18173;
  assign new_new_n31374__ = ys__n18173 & ys__n18863;
  assign new_new_n31375__ = ~new_new_n31373__ & ~new_new_n31374__;
  assign new_new_n31376__ = ~new_new_n16723__ & ~new_new_n31375__;
  assign new_new_n31377__ = ~new_new_n31372__ & ~new_new_n31376__;
  assign new_new_n31378__ = ys__n778 & ~new_new_n31377__;
  assign new_new_n31379__ = ~new_new_n31371__ & ~new_new_n31378__;
  assign new_new_n31380__ = ~ys__n602 & ~new_new_n31379__;
  assign new_new_n31381__ = new_new_n16723__ & ~new_new_n31379__;
  assign new_new_n31382__ = ys__n26192 & ~new_new_n16723__;
  assign new_new_n31383__ = ~new_new_n31381__ & ~new_new_n31382__;
  assign new_new_n31384__ = ys__n602 & ~new_new_n31383__;
  assign ys__n26751 = new_new_n31380__ | new_new_n31384__;
  assign new_new_n31386__ = ~ys__n778 & ys__n26192;
  assign new_new_n31387__ = ys__n26192 & new_new_n16723__;
  assign new_new_n31388__ = ys__n6129 & ~ys__n18173;
  assign new_new_n31389__ = ys__n18173 & ys__n18865;
  assign new_new_n31390__ = ~new_new_n31388__ & ~new_new_n31389__;
  assign new_new_n31391__ = ~new_new_n16723__ & ~new_new_n31390__;
  assign new_new_n31392__ = ~new_new_n31387__ & ~new_new_n31391__;
  assign new_new_n31393__ = ys__n778 & ~new_new_n31392__;
  assign new_new_n31394__ = ~new_new_n31386__ & ~new_new_n31393__;
  assign new_new_n31395__ = ~ys__n602 & ~new_new_n31394__;
  assign new_new_n31396__ = new_new_n16723__ & ~new_new_n31394__;
  assign new_new_n31397__ = ys__n26194 & ~new_new_n16723__;
  assign new_new_n31398__ = ~new_new_n31396__ & ~new_new_n31397__;
  assign new_new_n31399__ = ys__n602 & ~new_new_n31398__;
  assign ys__n26752 = new_new_n31395__ | new_new_n31399__;
  assign new_new_n31401__ = ~ys__n778 & ys__n26194;
  assign new_new_n31402__ = ys__n26194 & new_new_n16723__;
  assign new_new_n31403__ = ys__n6130 & ~ys__n18173;
  assign new_new_n31404__ = ys__n18173 & ys__n18867;
  assign new_new_n31405__ = ~new_new_n31403__ & ~new_new_n31404__;
  assign new_new_n31406__ = ~new_new_n16723__ & ~new_new_n31405__;
  assign new_new_n31407__ = ~new_new_n31402__ & ~new_new_n31406__;
  assign new_new_n31408__ = ys__n778 & ~new_new_n31407__;
  assign new_new_n31409__ = ~new_new_n31401__ & ~new_new_n31408__;
  assign new_new_n31410__ = ~ys__n602 & ~new_new_n31409__;
  assign new_new_n31411__ = new_new_n16723__ & ~new_new_n31409__;
  assign new_new_n31412__ = ys__n26196 & ~new_new_n16723__;
  assign new_new_n31413__ = ~new_new_n31411__ & ~new_new_n31412__;
  assign new_new_n31414__ = ys__n602 & ~new_new_n31413__;
  assign ys__n26753 = new_new_n31410__ | new_new_n31414__;
  assign new_new_n31416__ = ~ys__n778 & ys__n26196;
  assign new_new_n31417__ = ys__n26196 & new_new_n16723__;
  assign new_new_n31418__ = ys__n42 & ~ys__n18173;
  assign new_new_n31419__ = ys__n18173 & ys__n18869;
  assign new_new_n31420__ = ~new_new_n31418__ & ~new_new_n31419__;
  assign new_new_n31421__ = ~new_new_n16723__ & ~new_new_n31420__;
  assign new_new_n31422__ = ~new_new_n31417__ & ~new_new_n31421__;
  assign new_new_n31423__ = ys__n778 & ~new_new_n31422__;
  assign new_new_n31424__ = ~new_new_n31416__ & ~new_new_n31423__;
  assign new_new_n31425__ = ~ys__n602 & ~new_new_n31424__;
  assign new_new_n31426__ = new_new_n16723__ & ~new_new_n31424__;
  assign new_new_n31427__ = ys__n26198 & ~new_new_n16723__;
  assign new_new_n31428__ = ~new_new_n31426__ & ~new_new_n31427__;
  assign new_new_n31429__ = ys__n602 & ~new_new_n31428__;
  assign ys__n26754 = new_new_n31425__ | new_new_n31429__;
  assign new_new_n31431__ = ~ys__n778 & ys__n26198;
  assign new_new_n31432__ = ys__n26198 & new_new_n16723__;
  assign new_new_n31433__ = ys__n40 & ~ys__n18173;
  assign new_new_n31434__ = ys__n18173 & ys__n18871;
  assign new_new_n31435__ = ~new_new_n31433__ & ~new_new_n31434__;
  assign new_new_n31436__ = ~new_new_n16723__ & ~new_new_n31435__;
  assign new_new_n31437__ = ~new_new_n31432__ & ~new_new_n31436__;
  assign new_new_n31438__ = ys__n778 & ~new_new_n31437__;
  assign new_new_n31439__ = ~new_new_n31431__ & ~new_new_n31438__;
  assign new_new_n31440__ = ~ys__n602 & ~new_new_n31439__;
  assign new_new_n31441__ = new_new_n16723__ & ~new_new_n31439__;
  assign new_new_n31442__ = ys__n26200 & ~new_new_n16723__;
  assign new_new_n31443__ = ~new_new_n31441__ & ~new_new_n31442__;
  assign new_new_n31444__ = ys__n602 & ~new_new_n31443__;
  assign ys__n26755 = new_new_n31440__ | new_new_n31444__;
  assign new_new_n31446__ = ~ys__n778 & ys__n26200;
  assign new_new_n31447__ = ys__n26200 & new_new_n16723__;
  assign new_new_n31448__ = ys__n6133 & ~ys__n18173;
  assign new_new_n31449__ = ys__n18173 & ys__n18873;
  assign new_new_n31450__ = ~new_new_n31448__ & ~new_new_n31449__;
  assign new_new_n31451__ = ~new_new_n16723__ & ~new_new_n31450__;
  assign new_new_n31452__ = ~new_new_n31447__ & ~new_new_n31451__;
  assign new_new_n31453__ = ys__n778 & ~new_new_n31452__;
  assign new_new_n31454__ = ~new_new_n31446__ & ~new_new_n31453__;
  assign new_new_n31455__ = ~ys__n602 & ~new_new_n31454__;
  assign new_new_n31456__ = new_new_n16723__ & ~new_new_n31454__;
  assign new_new_n31457__ = ys__n26202 & ~new_new_n16723__;
  assign new_new_n31458__ = ~new_new_n31456__ & ~new_new_n31457__;
  assign new_new_n31459__ = ys__n602 & ~new_new_n31458__;
  assign ys__n26756 = new_new_n31455__ | new_new_n31459__;
  assign new_new_n31461__ = ~ys__n778 & ys__n26202;
  assign new_new_n31462__ = ys__n26202 & new_new_n16723__;
  assign new_new_n31463__ = ys__n6134 & ~ys__n18173;
  assign new_new_n31464__ = ys__n18173 & ys__n18875;
  assign new_new_n31465__ = ~new_new_n31463__ & ~new_new_n31464__;
  assign new_new_n31466__ = ~new_new_n16723__ & ~new_new_n31465__;
  assign new_new_n31467__ = ~new_new_n31462__ & ~new_new_n31466__;
  assign new_new_n31468__ = ys__n778 & ~new_new_n31467__;
  assign new_new_n31469__ = ~new_new_n31461__ & ~new_new_n31468__;
  assign new_new_n31470__ = ~ys__n602 & ~new_new_n31469__;
  assign new_new_n31471__ = new_new_n16723__ & ~new_new_n31469__;
  assign new_new_n31472__ = ys__n26204 & ~new_new_n16723__;
  assign new_new_n31473__ = ~new_new_n31471__ & ~new_new_n31472__;
  assign new_new_n31474__ = ys__n602 & ~new_new_n31473__;
  assign ys__n26757 = new_new_n31470__ | new_new_n31474__;
  assign new_new_n31476__ = ~ys__n778 & ys__n26204;
  assign new_new_n31477__ = ys__n26204 & new_new_n16723__;
  assign new_new_n31478__ = ys__n38 & ~ys__n18173;
  assign new_new_n31479__ = ys__n18173 & ys__n18877;
  assign new_new_n31480__ = ~new_new_n31478__ & ~new_new_n31479__;
  assign new_new_n31481__ = ~new_new_n16723__ & ~new_new_n31480__;
  assign new_new_n31482__ = ~new_new_n31477__ & ~new_new_n31481__;
  assign new_new_n31483__ = ys__n778 & ~new_new_n31482__;
  assign new_new_n31484__ = ~new_new_n31476__ & ~new_new_n31483__;
  assign new_new_n31485__ = ~ys__n602 & ~new_new_n31484__;
  assign new_new_n31486__ = new_new_n16723__ & ~new_new_n31484__;
  assign new_new_n31487__ = ys__n26206 & ~new_new_n16723__;
  assign new_new_n31488__ = ~new_new_n31486__ & ~new_new_n31487__;
  assign new_new_n31489__ = ys__n602 & ~new_new_n31488__;
  assign ys__n26758 = new_new_n31485__ | new_new_n31489__;
  assign new_new_n31491__ = ~ys__n778 & ys__n26206;
  assign new_new_n31492__ = ys__n26206 & new_new_n16723__;
  assign new_new_n31493__ = ys__n36 & ~ys__n18173;
  assign new_new_n31494__ = ys__n18173 & ys__n18879;
  assign new_new_n31495__ = ~new_new_n31493__ & ~new_new_n31494__;
  assign new_new_n31496__ = ~new_new_n16723__ & ~new_new_n31495__;
  assign new_new_n31497__ = ~new_new_n31492__ & ~new_new_n31496__;
  assign new_new_n31498__ = ys__n778 & ~new_new_n31497__;
  assign new_new_n31499__ = ~new_new_n31491__ & ~new_new_n31498__;
  assign new_new_n31500__ = ~ys__n602 & ~new_new_n31499__;
  assign new_new_n31501__ = new_new_n16723__ & ~new_new_n31499__;
  assign new_new_n31502__ = ys__n26208 & ~new_new_n16723__;
  assign new_new_n31503__ = ~new_new_n31501__ & ~new_new_n31502__;
  assign new_new_n31504__ = ys__n602 & ~new_new_n31503__;
  assign ys__n26759 = new_new_n31500__ | new_new_n31504__;
  assign new_new_n31506__ = ~ys__n778 & ys__n26208;
  assign new_new_n31507__ = ys__n26208 & new_new_n16723__;
  assign new_new_n31508__ = ys__n34 & ~ys__n18173;
  assign new_new_n31509__ = ys__n18173 & ys__n18881;
  assign new_new_n31510__ = ~new_new_n31508__ & ~new_new_n31509__;
  assign new_new_n31511__ = ~new_new_n16723__ & ~new_new_n31510__;
  assign new_new_n31512__ = ~new_new_n31507__ & ~new_new_n31511__;
  assign new_new_n31513__ = ys__n778 & ~new_new_n31512__;
  assign new_new_n31514__ = ~new_new_n31506__ & ~new_new_n31513__;
  assign new_new_n31515__ = ~ys__n602 & ~new_new_n31514__;
  assign new_new_n31516__ = new_new_n16723__ & ~new_new_n31514__;
  assign new_new_n31517__ = ys__n26210 & ~new_new_n16723__;
  assign new_new_n31518__ = ~new_new_n31516__ & ~new_new_n31517__;
  assign new_new_n31519__ = ys__n602 & ~new_new_n31518__;
  assign ys__n26760 = new_new_n31515__ | new_new_n31519__;
  assign new_new_n31521__ = ~ys__n778 & ys__n26210;
  assign new_new_n31522__ = ys__n26210 & new_new_n16723__;
  assign new_new_n31523__ = ys__n32 & ~ys__n18173;
  assign new_new_n31524__ = ys__n18173 & ys__n18883;
  assign new_new_n31525__ = ~new_new_n31523__ & ~new_new_n31524__;
  assign new_new_n31526__ = ~new_new_n16723__ & ~new_new_n31525__;
  assign new_new_n31527__ = ~new_new_n31522__ & ~new_new_n31526__;
  assign new_new_n31528__ = ys__n778 & ~new_new_n31527__;
  assign new_new_n31529__ = ~new_new_n31521__ & ~new_new_n31528__;
  assign new_new_n31530__ = ~ys__n602 & ~new_new_n31529__;
  assign new_new_n31531__ = new_new_n16723__ & ~new_new_n31529__;
  assign new_new_n31532__ = ys__n26212 & ~new_new_n16723__;
  assign new_new_n31533__ = ~new_new_n31531__ & ~new_new_n31532__;
  assign new_new_n31534__ = ys__n602 & ~new_new_n31533__;
  assign ys__n26761 = new_new_n31530__ | new_new_n31534__;
  assign new_new_n31536__ = ~ys__n778 & ys__n26212;
  assign new_new_n31537__ = ys__n26212 & new_new_n16723__;
  assign new_new_n31538__ = ys__n30 & ~ys__n18173;
  assign new_new_n31539__ = ys__n18173 & ys__n18885;
  assign new_new_n31540__ = ~new_new_n31538__ & ~new_new_n31539__;
  assign new_new_n31541__ = ~new_new_n16723__ & ~new_new_n31540__;
  assign new_new_n31542__ = ~new_new_n31537__ & ~new_new_n31541__;
  assign new_new_n31543__ = ys__n778 & ~new_new_n31542__;
  assign new_new_n31544__ = ~new_new_n31536__ & ~new_new_n31543__;
  assign new_new_n31545__ = ~ys__n602 & ~new_new_n31544__;
  assign new_new_n31546__ = new_new_n16723__ & ~new_new_n31544__;
  assign new_new_n31547__ = ys__n26214 & ~new_new_n16723__;
  assign new_new_n31548__ = ~new_new_n31546__ & ~new_new_n31547__;
  assign new_new_n31549__ = ys__n602 & ~new_new_n31548__;
  assign ys__n26762 = new_new_n31545__ | new_new_n31549__;
  assign new_new_n31551__ = ~ys__n778 & ys__n26214;
  assign new_new_n31552__ = ys__n26214 & new_new_n16723__;
  assign new_new_n31553__ = ys__n28 & ~ys__n18173;
  assign new_new_n31554__ = ys__n18173 & ys__n18887;
  assign new_new_n31555__ = ~new_new_n31553__ & ~new_new_n31554__;
  assign new_new_n31556__ = ~new_new_n16723__ & ~new_new_n31555__;
  assign new_new_n31557__ = ~new_new_n31552__ & ~new_new_n31556__;
  assign new_new_n31558__ = ys__n778 & ~new_new_n31557__;
  assign new_new_n31559__ = ~new_new_n31551__ & ~new_new_n31558__;
  assign new_new_n31560__ = ~ys__n602 & ~new_new_n31559__;
  assign new_new_n31561__ = new_new_n16723__ & ~new_new_n31559__;
  assign new_new_n31562__ = ys__n26216 & ~new_new_n16723__;
  assign new_new_n31563__ = ~new_new_n31561__ & ~new_new_n31562__;
  assign new_new_n31564__ = ys__n602 & ~new_new_n31563__;
  assign ys__n26763 = new_new_n31560__ | new_new_n31564__;
  assign new_new_n31566__ = ~ys__n778 & ys__n26216;
  assign new_new_n31567__ = ys__n26216 & new_new_n16723__;
  assign new_new_n31568__ = ys__n26 & ~ys__n18173;
  assign new_new_n31569__ = ys__n18173 & ys__n18889;
  assign new_new_n31570__ = ~new_new_n31568__ & ~new_new_n31569__;
  assign new_new_n31571__ = ~new_new_n16723__ & ~new_new_n31570__;
  assign new_new_n31572__ = ~new_new_n31567__ & ~new_new_n31571__;
  assign new_new_n31573__ = ys__n778 & ~new_new_n31572__;
  assign new_new_n31574__ = ~new_new_n31566__ & ~new_new_n31573__;
  assign new_new_n31575__ = ~ys__n602 & ~new_new_n31574__;
  assign new_new_n31576__ = new_new_n16723__ & ~new_new_n31574__;
  assign new_new_n31577__ = ys__n26218 & ~new_new_n16723__;
  assign new_new_n31578__ = ~new_new_n31576__ & ~new_new_n31577__;
  assign new_new_n31579__ = ys__n602 & ~new_new_n31578__;
  assign ys__n26764 = new_new_n31575__ | new_new_n31579__;
  assign new_new_n31581__ = ~ys__n778 & ys__n26218;
  assign new_new_n31582__ = ys__n26218 & new_new_n16723__;
  assign new_new_n31583__ = ys__n24 & ~ys__n18173;
  assign new_new_n31584__ = ys__n18173 & ys__n18891;
  assign new_new_n31585__ = ~new_new_n31583__ & ~new_new_n31584__;
  assign new_new_n31586__ = ~new_new_n16723__ & ~new_new_n31585__;
  assign new_new_n31587__ = ~new_new_n31582__ & ~new_new_n31586__;
  assign new_new_n31588__ = ys__n778 & ~new_new_n31587__;
  assign new_new_n31589__ = ~new_new_n31581__ & ~new_new_n31588__;
  assign new_new_n31590__ = ~ys__n602 & ~new_new_n31589__;
  assign new_new_n31591__ = new_new_n16723__ & ~new_new_n31589__;
  assign new_new_n31592__ = ~new_new_n16723__ & new_new_n30646__;
  assign new_new_n31593__ = ~new_new_n31591__ & ~new_new_n31592__;
  assign new_new_n31594__ = ys__n602 & ~new_new_n31593__;
  assign ys__n26765 = new_new_n31590__ | new_new_n31594__;
  assign ys__n26802 = ys__n18448 & new_new_n12246__;
  assign ys__n26803 = new_new_n12250__ & ys__n26802;
  assign ys__n26804 = ys__n18451 & new_new_n12246__;
  assign ys__n26805 = new_new_n12250__ & ys__n26804;
  assign ys__n26806 = ys__n18454 & new_new_n12246__;
  assign ys__n26807 = new_new_n12250__ & ys__n26806;
  assign ys__n26808 = ys__n18457 & new_new_n12246__;
  assign ys__n26809 = new_new_n12250__ & ys__n26808;
  assign ys__n26810 = ys__n18460 & new_new_n12246__;
  assign ys__n26811 = new_new_n12250__ & ys__n26810;
  assign ys__n26812 = ys__n18463 & new_new_n12246__;
  assign ys__n26813 = new_new_n12250__ & ys__n26812;
  assign ys__n26814 = ys__n18466 & new_new_n12246__;
  assign ys__n26815 = new_new_n12250__ & ys__n26814;
  assign ys__n26816 = ys__n18469 & new_new_n12246__;
  assign ys__n26817 = new_new_n12250__ & ys__n26816;
  assign ys__n26818 = ys__n18472 & new_new_n12246__;
  assign ys__n26819 = new_new_n12250__ & ys__n26818;
  assign ys__n26820 = ys__n18475 & new_new_n12246__;
  assign ys__n26821 = new_new_n12250__ & ys__n26820;
  assign ys__n26822 = ys__n18478 & new_new_n12246__;
  assign ys__n26823 = new_new_n12250__ & ys__n26822;
  assign ys__n26824 = ys__n18481 & new_new_n12246__;
  assign ys__n26825 = new_new_n12250__ & ys__n26824;
  assign ys__n26826 = ys__n18484 & new_new_n12246__;
  assign ys__n26827 = new_new_n12250__ & ys__n26826;
  assign ys__n26828 = ys__n18487 & new_new_n12246__;
  assign ys__n26829 = new_new_n12250__ & ys__n26828;
  assign ys__n26830 = ys__n18490 & new_new_n12246__;
  assign ys__n26831 = new_new_n12250__ & ys__n26830;
  assign ys__n26832 = ys__n18493 & new_new_n12246__;
  assign ys__n26833 = new_new_n12250__ & ys__n26832;
  assign ys__n26834 = ys__n18496 & new_new_n12246__;
  assign ys__n26835 = new_new_n12250__ & ys__n26834;
  assign ys__n26836 = ys__n18499 & new_new_n12246__;
  assign ys__n26837 = new_new_n12250__ & ys__n26836;
  assign ys__n26838 = ys__n18502 & new_new_n12246__;
  assign ys__n26839 = new_new_n12250__ & ys__n26838;
  assign ys__n26840 = ys__n18505 & new_new_n12246__;
  assign ys__n26841 = new_new_n12250__ & ys__n26840;
  assign ys__n26842 = ys__n18508 & new_new_n12246__;
  assign ys__n26843 = new_new_n12250__ & ys__n26842;
  assign ys__n26844 = ys__n18511 & new_new_n12246__;
  assign ys__n26845 = new_new_n12250__ & ys__n26844;
  assign ys__n26846 = ys__n18514 & new_new_n12246__;
  assign ys__n26847 = new_new_n12250__ & ys__n26846;
  assign ys__n26848 = ys__n18517 & new_new_n12246__;
  assign ys__n26849 = new_new_n12250__ & ys__n26848;
  assign ys__n26850 = ys__n18520 & new_new_n12246__;
  assign ys__n26851 = new_new_n12250__ & ys__n26850;
  assign ys__n26852 = ys__n18523 & new_new_n12246__;
  assign ys__n26853 = new_new_n12250__ & ys__n26852;
  assign ys__n26854 = ys__n18526 & new_new_n12246__;
  assign ys__n26855 = new_new_n12250__ & ys__n26854;
  assign ys__n26856 = ys__n18529 & new_new_n12246__;
  assign ys__n26857 = new_new_n12250__ & ys__n26856;
  assign ys__n26858 = ys__n18532 & new_new_n12246__;
  assign ys__n26859 = new_new_n12250__ & ys__n26858;
  assign ys__n26860 = ys__n18535 & new_new_n12246__;
  assign ys__n26861 = new_new_n12250__ & ys__n26860;
  assign ys__n26862 = ys__n18538 & new_new_n12246__;
  assign ys__n26863 = new_new_n12250__ & ys__n26862;
  assign ys__n26864 = ys__n18541 & new_new_n12246__;
  assign ys__n26865 = new_new_n12250__ & ys__n26864;
  assign ys__n26866 = ys__n18448 & new_new_n12245__;
  assign ys__n26867 = new_new_n12250__ & ys__n26866;
  assign ys__n26868 = ys__n18451 & new_new_n12245__;
  assign ys__n26869 = new_new_n12250__ & ys__n26868;
  assign ys__n26870 = ys__n18454 & new_new_n12245__;
  assign ys__n26871 = new_new_n12250__ & ys__n26870;
  assign ys__n26872 = ys__n18457 & new_new_n12245__;
  assign ys__n26873 = new_new_n12250__ & ys__n26872;
  assign ys__n26874 = ys__n18460 & new_new_n12245__;
  assign ys__n26875 = new_new_n12250__ & ys__n26874;
  assign ys__n26876 = ys__n18463 & new_new_n12245__;
  assign ys__n26877 = new_new_n12250__ & ys__n26876;
  assign ys__n26878 = ys__n18466 & new_new_n12245__;
  assign ys__n26879 = new_new_n12250__ & ys__n26878;
  assign ys__n26880 = ys__n18469 & new_new_n12245__;
  assign ys__n26881 = new_new_n12250__ & ys__n26880;
  assign ys__n26882 = ys__n18472 & new_new_n12245__;
  assign ys__n26883 = new_new_n12250__ & ys__n26882;
  assign ys__n26884 = ys__n18475 & new_new_n12245__;
  assign ys__n26885 = new_new_n12250__ & ys__n26884;
  assign ys__n26886 = ys__n18478 & new_new_n12245__;
  assign ys__n26887 = new_new_n12250__ & ys__n26886;
  assign ys__n26888 = ys__n18481 & new_new_n12245__;
  assign ys__n26889 = new_new_n12250__ & ys__n26888;
  assign ys__n26890 = ys__n18484 & new_new_n12245__;
  assign ys__n26891 = new_new_n12250__ & ys__n26890;
  assign ys__n26892 = ys__n18487 & new_new_n12245__;
  assign ys__n26893 = new_new_n12250__ & ys__n26892;
  assign ys__n26894 = ys__n18490 & new_new_n12245__;
  assign ys__n26895 = new_new_n12250__ & ys__n26894;
  assign ys__n26896 = ys__n18493 & new_new_n12245__;
  assign ys__n26897 = new_new_n12250__ & ys__n26896;
  assign ys__n26898 = ys__n18496 & new_new_n12245__;
  assign ys__n26899 = new_new_n12250__ & ys__n26898;
  assign ys__n26900 = ys__n18499 & new_new_n12245__;
  assign ys__n26901 = new_new_n12250__ & ys__n26900;
  assign ys__n26902 = ys__n18502 & new_new_n12245__;
  assign ys__n26903 = new_new_n12250__ & ys__n26902;
  assign ys__n26904 = ys__n18505 & new_new_n12245__;
  assign ys__n26905 = new_new_n12250__ & ys__n26904;
  assign ys__n26906 = ys__n18508 & new_new_n12245__;
  assign ys__n26907 = new_new_n12250__ & ys__n26906;
  assign ys__n26908 = ys__n18511 & new_new_n12245__;
  assign ys__n26909 = new_new_n12250__ & ys__n26908;
  assign ys__n26910 = ys__n18514 & new_new_n12245__;
  assign ys__n26911 = new_new_n12250__ & ys__n26910;
  assign ys__n26912 = ys__n18517 & new_new_n12245__;
  assign ys__n26913 = new_new_n12250__ & ys__n26912;
  assign ys__n26914 = ys__n18520 & new_new_n12245__;
  assign ys__n26915 = new_new_n12250__ & ys__n26914;
  assign ys__n26916 = ys__n18523 & new_new_n12245__;
  assign ys__n26917 = new_new_n12250__ & ys__n26916;
  assign ys__n26918 = ys__n18526 & new_new_n12245__;
  assign ys__n26919 = new_new_n12250__ & ys__n26918;
  assign ys__n26920 = ys__n18529 & new_new_n12245__;
  assign ys__n26921 = new_new_n12250__ & ys__n26920;
  assign ys__n26922 = ys__n18532 & new_new_n12245__;
  assign ys__n26923 = new_new_n12250__ & ys__n26922;
  assign ys__n26924 = ys__n18535 & new_new_n12245__;
  assign ys__n26925 = new_new_n12250__ & ys__n26924;
  assign ys__n26926 = ys__n18538 & new_new_n12245__;
  assign ys__n26927 = new_new_n12250__ & ys__n26926;
  assign ys__n26928 = ys__n18541 & new_new_n12245__;
  assign ys__n26929 = new_new_n12250__ & ys__n26928;
  assign ys__n26930 = ys__n18448 & new_new_n12248__;
  assign ys__n26931 = new_new_n12250__ & ys__n26930;
  assign ys__n26932 = ys__n18451 & new_new_n12248__;
  assign ys__n26933 = new_new_n12250__ & ys__n26932;
  assign ys__n26934 = ys__n18454 & new_new_n12248__;
  assign ys__n26935 = new_new_n12250__ & ys__n26934;
  assign ys__n26936 = ys__n18457 & new_new_n12248__;
  assign ys__n26937 = new_new_n12250__ & ys__n26936;
  assign ys__n26938 = ys__n18460 & new_new_n12248__;
  assign ys__n26939 = new_new_n12250__ & ys__n26938;
  assign ys__n26940 = ys__n18463 & new_new_n12248__;
  assign ys__n26941 = new_new_n12250__ & ys__n26940;
  assign ys__n26942 = ys__n18466 & new_new_n12248__;
  assign ys__n26943 = new_new_n12250__ & ys__n26942;
  assign ys__n26944 = ys__n18469 & new_new_n12248__;
  assign ys__n26945 = new_new_n12250__ & ys__n26944;
  assign ys__n26946 = ys__n18472 & new_new_n12248__;
  assign ys__n26947 = new_new_n12250__ & ys__n26946;
  assign ys__n26948 = ys__n18475 & new_new_n12248__;
  assign ys__n26949 = new_new_n12250__ & ys__n26948;
  assign ys__n26950 = ys__n18478 & new_new_n12248__;
  assign ys__n26951 = new_new_n12250__ & ys__n26950;
  assign ys__n26952 = ys__n18481 & new_new_n12248__;
  assign ys__n26953 = new_new_n12250__ & ys__n26952;
  assign ys__n26954 = ys__n18484 & new_new_n12248__;
  assign ys__n26955 = new_new_n12250__ & ys__n26954;
  assign ys__n26956 = ys__n18487 & new_new_n12248__;
  assign ys__n26957 = new_new_n12250__ & ys__n26956;
  assign ys__n26958 = ys__n18490 & new_new_n12248__;
  assign ys__n26959 = new_new_n12250__ & ys__n26958;
  assign ys__n26960 = ys__n18493 & new_new_n12248__;
  assign ys__n26961 = new_new_n12250__ & ys__n26960;
  assign ys__n26962 = ys__n18496 & new_new_n12248__;
  assign ys__n26963 = new_new_n12250__ & ys__n26962;
  assign ys__n26964 = ys__n18499 & new_new_n12248__;
  assign ys__n26965 = new_new_n12250__ & ys__n26964;
  assign ys__n26966 = ys__n18502 & new_new_n12248__;
  assign ys__n26967 = new_new_n12250__ & ys__n26966;
  assign ys__n26968 = ys__n18505 & new_new_n12248__;
  assign ys__n26969 = new_new_n12250__ & ys__n26968;
  assign ys__n26970 = ys__n18508 & new_new_n12248__;
  assign ys__n26971 = new_new_n12250__ & ys__n26970;
  assign ys__n26972 = ys__n18511 & new_new_n12248__;
  assign ys__n26973 = new_new_n12250__ & ys__n26972;
  assign ys__n26974 = ys__n18514 & new_new_n12248__;
  assign ys__n26975 = new_new_n12250__ & ys__n26974;
  assign ys__n26976 = ys__n18517 & new_new_n12248__;
  assign ys__n26977 = new_new_n12250__ & ys__n26976;
  assign ys__n26978 = ys__n18520 & new_new_n12248__;
  assign ys__n26979 = new_new_n12250__ & ys__n26978;
  assign ys__n26980 = ys__n18523 & new_new_n12248__;
  assign ys__n26981 = new_new_n12250__ & ys__n26980;
  assign ys__n26982 = ys__n18526 & new_new_n12248__;
  assign ys__n26983 = new_new_n12250__ & ys__n26982;
  assign ys__n26984 = ys__n18529 & new_new_n12248__;
  assign ys__n26985 = new_new_n12250__ & ys__n26984;
  assign ys__n26986 = ys__n18532 & new_new_n12248__;
  assign ys__n26987 = new_new_n12250__ & ys__n26986;
  assign ys__n26988 = ys__n18535 & new_new_n12248__;
  assign ys__n26989 = new_new_n12250__ & ys__n26988;
  assign ys__n26990 = ys__n18538 & new_new_n12248__;
  assign ys__n26991 = new_new_n12250__ & ys__n26990;
  assign ys__n26992 = ys__n18541 & new_new_n12248__;
  assign ys__n26993 = new_new_n12250__ & ys__n26992;
  assign ys__n26994 = ys__n18448 & new_new_n12356__;
  assign ys__n26995 = new_new_n12250__ & ys__n26994;
  assign ys__n26996 = ys__n18451 & new_new_n12356__;
  assign ys__n26997 = new_new_n12250__ & ys__n26996;
  assign ys__n26998 = ys__n18454 & new_new_n12356__;
  assign ys__n26999 = new_new_n12250__ & ys__n26998;
  assign ys__n27000 = ys__n18457 & new_new_n12356__;
  assign ys__n27001 = new_new_n12250__ & ys__n27000;
  assign ys__n27002 = ys__n18460 & new_new_n12356__;
  assign ys__n27003 = new_new_n12250__ & ys__n27002;
  assign ys__n27004 = ys__n18463 & new_new_n12356__;
  assign ys__n27005 = new_new_n12250__ & ys__n27004;
  assign ys__n27006 = ys__n18466 & new_new_n12356__;
  assign ys__n27007 = new_new_n12250__ & ys__n27006;
  assign ys__n27008 = ys__n18469 & new_new_n12356__;
  assign ys__n27009 = new_new_n12250__ & ys__n27008;
  assign ys__n27010 = ys__n18472 & new_new_n12356__;
  assign ys__n27011 = new_new_n12250__ & ys__n27010;
  assign ys__n27012 = ys__n18475 & new_new_n12356__;
  assign ys__n27013 = new_new_n12250__ & ys__n27012;
  assign ys__n27014 = ys__n18478 & new_new_n12356__;
  assign ys__n27015 = new_new_n12250__ & ys__n27014;
  assign ys__n27016 = ys__n18481 & new_new_n12356__;
  assign ys__n27017 = new_new_n12250__ & ys__n27016;
  assign ys__n27018 = ys__n18484 & new_new_n12356__;
  assign ys__n27019 = new_new_n12250__ & ys__n27018;
  assign ys__n27020 = ys__n18487 & new_new_n12356__;
  assign ys__n27021 = new_new_n12250__ & ys__n27020;
  assign ys__n27022 = ys__n18490 & new_new_n12356__;
  assign ys__n27023 = new_new_n12250__ & ys__n27022;
  assign ys__n27024 = ys__n18493 & new_new_n12356__;
  assign ys__n27025 = new_new_n12250__ & ys__n27024;
  assign ys__n27026 = ys__n18496 & new_new_n12356__;
  assign ys__n27027 = new_new_n12250__ & ys__n27026;
  assign ys__n27028 = ys__n18499 & new_new_n12356__;
  assign ys__n27029 = new_new_n12250__ & ys__n27028;
  assign ys__n27030 = ys__n18502 & new_new_n12356__;
  assign ys__n27031 = new_new_n12250__ & ys__n27030;
  assign ys__n27032 = ys__n18505 & new_new_n12356__;
  assign ys__n27033 = new_new_n12250__ & ys__n27032;
  assign ys__n27034 = ys__n18508 & new_new_n12356__;
  assign ys__n27035 = new_new_n12250__ & ys__n27034;
  assign ys__n27036 = ys__n18511 & new_new_n12356__;
  assign ys__n27037 = new_new_n12250__ & ys__n27036;
  assign ys__n27038 = ys__n18514 & new_new_n12356__;
  assign ys__n27039 = new_new_n12250__ & ys__n27038;
  assign ys__n27040 = ys__n18517 & new_new_n12356__;
  assign ys__n27041 = new_new_n12250__ & ys__n27040;
  assign ys__n27042 = ys__n18520 & new_new_n12356__;
  assign ys__n27043 = new_new_n12250__ & ys__n27042;
  assign ys__n27044 = ys__n18523 & new_new_n12356__;
  assign ys__n27045 = new_new_n12250__ & ys__n27044;
  assign ys__n27046 = ys__n18526 & new_new_n12356__;
  assign ys__n27047 = new_new_n12250__ & ys__n27046;
  assign ys__n27048 = ys__n18529 & new_new_n12356__;
  assign ys__n27049 = new_new_n12250__ & ys__n27048;
  assign ys__n27050 = ys__n18532 & new_new_n12356__;
  assign ys__n27051 = new_new_n12250__ & ys__n27050;
  assign ys__n27052 = ys__n18535 & new_new_n12356__;
  assign ys__n27053 = new_new_n12250__ & ys__n27052;
  assign ys__n27054 = ys__n18538 & new_new_n12356__;
  assign ys__n27055 = new_new_n12250__ & ys__n27054;
  assign ys__n27056 = ys__n18541 & new_new_n12356__;
  assign ys__n27057 = new_new_n12250__ & ys__n27056;
  assign ys__n27058 = new_new_n12242__ & ys__n26802;
  assign ys__n27059 = new_new_n12242__ & ys__n26804;
  assign ys__n27060 = new_new_n12242__ & ys__n26806;
  assign ys__n27061 = new_new_n12242__ & ys__n26808;
  assign ys__n27062 = new_new_n12242__ & ys__n26810;
  assign ys__n27063 = new_new_n12242__ & ys__n26812;
  assign ys__n27064 = new_new_n12242__ & ys__n26814;
  assign ys__n27065 = new_new_n12242__ & ys__n26816;
  assign ys__n27066 = new_new_n12242__ & ys__n26818;
  assign ys__n27067 = new_new_n12242__ & ys__n26820;
  assign ys__n27068 = new_new_n12242__ & ys__n26822;
  assign ys__n27069 = new_new_n12242__ & ys__n26824;
  assign ys__n27070 = new_new_n12242__ & ys__n26826;
  assign ys__n27071 = new_new_n12242__ & ys__n26828;
  assign ys__n27072 = new_new_n12242__ & ys__n26830;
  assign ys__n27073 = new_new_n12242__ & ys__n26832;
  assign ys__n27074 = new_new_n12242__ & ys__n26834;
  assign ys__n27075 = new_new_n12242__ & ys__n26836;
  assign ys__n27076 = new_new_n12242__ & ys__n26838;
  assign ys__n27077 = new_new_n12242__ & ys__n26840;
  assign ys__n27078 = new_new_n12242__ & ys__n26842;
  assign ys__n27079 = new_new_n12242__ & ys__n26844;
  assign ys__n27080 = new_new_n12242__ & ys__n26846;
  assign ys__n27081 = new_new_n12242__ & ys__n26848;
  assign ys__n27082 = new_new_n12242__ & ys__n26850;
  assign ys__n27083 = new_new_n12242__ & ys__n26852;
  assign ys__n27084 = new_new_n12242__ & ys__n26854;
  assign ys__n27085 = new_new_n12242__ & ys__n26856;
  assign ys__n27086 = new_new_n12242__ & ys__n26858;
  assign ys__n27087 = new_new_n12242__ & ys__n26860;
  assign ys__n27088 = new_new_n12242__ & ys__n26862;
  assign ys__n27089 = new_new_n12242__ & ys__n26864;
  assign ys__n27090 = new_new_n12242__ & ys__n26866;
  assign ys__n27091 = new_new_n12242__ & ys__n26868;
  assign ys__n27092 = new_new_n12242__ & ys__n26870;
  assign ys__n27093 = new_new_n12242__ & ys__n26872;
  assign ys__n27094 = new_new_n12242__ & ys__n26874;
  assign ys__n27095 = new_new_n12242__ & ys__n26876;
  assign ys__n27096 = new_new_n12242__ & ys__n26878;
  assign ys__n27097 = new_new_n12242__ & ys__n26880;
  assign ys__n27098 = new_new_n12242__ & ys__n26882;
  assign ys__n27099 = new_new_n12242__ & ys__n26884;
  assign ys__n27100 = new_new_n12242__ & ys__n26886;
  assign ys__n27101 = new_new_n12242__ & ys__n26888;
  assign ys__n27102 = new_new_n12242__ & ys__n26890;
  assign ys__n27103 = new_new_n12242__ & ys__n26892;
  assign ys__n27104 = new_new_n12242__ & ys__n26894;
  assign ys__n27105 = new_new_n12242__ & ys__n26896;
  assign ys__n27106 = new_new_n12242__ & ys__n26898;
  assign ys__n27107 = new_new_n12242__ & ys__n26900;
  assign ys__n27108 = new_new_n12242__ & ys__n26902;
  assign ys__n27109 = new_new_n12242__ & ys__n26904;
  assign ys__n27110 = new_new_n12242__ & ys__n26906;
  assign ys__n27111 = new_new_n12242__ & ys__n26908;
  assign ys__n27112 = new_new_n12242__ & ys__n26910;
  assign ys__n27113 = new_new_n12242__ & ys__n26912;
  assign ys__n27114 = new_new_n12242__ & ys__n26914;
  assign ys__n27115 = new_new_n12242__ & ys__n26916;
  assign ys__n27116 = new_new_n12242__ & ys__n26918;
  assign ys__n27117 = new_new_n12242__ & ys__n26920;
  assign ys__n27118 = new_new_n12242__ & ys__n26922;
  assign ys__n27119 = new_new_n12242__ & ys__n26924;
  assign ys__n27120 = new_new_n12242__ & ys__n26926;
  assign ys__n27121 = new_new_n12242__ & ys__n26928;
  assign ys__n27122 = new_new_n12242__ & ys__n26930;
  assign ys__n27123 = new_new_n12242__ & ys__n26932;
  assign ys__n27124 = new_new_n12242__ & ys__n26934;
  assign ys__n27125 = new_new_n12242__ & ys__n26936;
  assign ys__n27126 = new_new_n12242__ & ys__n26938;
  assign ys__n27127 = new_new_n12242__ & ys__n26940;
  assign ys__n27128 = new_new_n12242__ & ys__n26942;
  assign ys__n27129 = new_new_n12242__ & ys__n26944;
  assign ys__n27130 = new_new_n12242__ & ys__n26946;
  assign ys__n27131 = new_new_n12242__ & ys__n26948;
  assign ys__n27132 = new_new_n12242__ & ys__n26950;
  assign ys__n27133 = new_new_n12242__ & ys__n26952;
  assign ys__n27134 = new_new_n12242__ & ys__n26954;
  assign ys__n27135 = new_new_n12242__ & ys__n26956;
  assign ys__n27136 = new_new_n12242__ & ys__n26958;
  assign ys__n27137 = new_new_n12242__ & ys__n26960;
  assign ys__n27138 = new_new_n12242__ & ys__n26962;
  assign ys__n27139 = new_new_n12242__ & ys__n26964;
  assign ys__n27140 = new_new_n12242__ & ys__n26966;
  assign ys__n27141 = new_new_n12242__ & ys__n26968;
  assign ys__n27142 = new_new_n12242__ & ys__n26970;
  assign ys__n27143 = new_new_n12242__ & ys__n26972;
  assign ys__n27144 = new_new_n12242__ & ys__n26974;
  assign ys__n27145 = new_new_n12242__ & ys__n26976;
  assign ys__n27146 = new_new_n12242__ & ys__n26978;
  assign ys__n27147 = new_new_n12242__ & ys__n26980;
  assign ys__n27148 = new_new_n12242__ & ys__n26982;
  assign ys__n27149 = new_new_n12242__ & ys__n26984;
  assign ys__n27150 = new_new_n12242__ & ys__n26986;
  assign ys__n27151 = new_new_n12242__ & ys__n26988;
  assign ys__n27152 = new_new_n12242__ & ys__n26990;
  assign ys__n27153 = new_new_n12242__ & ys__n26992;
  assign ys__n27154 = new_new_n12242__ & ys__n26994;
  assign ys__n27155 = new_new_n12242__ & ys__n26996;
  assign ys__n27156 = new_new_n12242__ & ys__n26998;
  assign ys__n27157 = new_new_n12242__ & ys__n27000;
  assign ys__n27158 = new_new_n12242__ & ys__n27002;
  assign ys__n27159 = new_new_n12242__ & ys__n27004;
  assign ys__n27160 = new_new_n12242__ & ys__n27006;
  assign ys__n27161 = new_new_n12242__ & ys__n27008;
  assign ys__n27162 = new_new_n12242__ & ys__n27010;
  assign ys__n27163 = new_new_n12242__ & ys__n27012;
  assign ys__n27164 = new_new_n12242__ & ys__n27014;
  assign ys__n27165 = new_new_n12242__ & ys__n27016;
  assign ys__n27166 = new_new_n12242__ & ys__n27018;
  assign ys__n27167 = new_new_n12242__ & ys__n27020;
  assign ys__n27168 = new_new_n12242__ & ys__n27022;
  assign ys__n27169 = new_new_n12242__ & ys__n27024;
  assign ys__n27170 = new_new_n12242__ & ys__n27026;
  assign ys__n27171 = new_new_n12242__ & ys__n27028;
  assign ys__n27172 = new_new_n12242__ & ys__n27030;
  assign ys__n27173 = new_new_n12242__ & ys__n27032;
  assign ys__n27174 = new_new_n12242__ & ys__n27034;
  assign ys__n27175 = new_new_n12242__ & ys__n27036;
  assign ys__n27176 = new_new_n12242__ & ys__n27038;
  assign ys__n27177 = new_new_n12242__ & ys__n27040;
  assign ys__n27178 = new_new_n12242__ & ys__n27042;
  assign ys__n27179 = new_new_n12242__ & ys__n27044;
  assign ys__n27180 = new_new_n12242__ & ys__n27046;
  assign ys__n27181 = new_new_n12242__ & ys__n27048;
  assign ys__n27182 = new_new_n12242__ & ys__n27050;
  assign ys__n27183 = new_new_n12242__ & ys__n27052;
  assign ys__n27184 = new_new_n12242__ & ys__n27054;
  assign ys__n27185 = new_new_n12242__ & ys__n27056;
  assign ys__n27186 = new_new_n12240__ & ys__n26802;
  assign ys__n27187 = new_new_n12240__ & ys__n26804;
  assign ys__n27188 = new_new_n12240__ & ys__n26806;
  assign ys__n27189 = new_new_n12240__ & ys__n26808;
  assign ys__n27190 = new_new_n12240__ & ys__n26810;
  assign ys__n27191 = new_new_n12240__ & ys__n26812;
  assign ys__n27192 = new_new_n12240__ & ys__n26814;
  assign ys__n27193 = new_new_n12240__ & ys__n26816;
  assign ys__n27194 = new_new_n12240__ & ys__n26818;
  assign ys__n27195 = new_new_n12240__ & ys__n26820;
  assign ys__n27196 = new_new_n12240__ & ys__n26822;
  assign ys__n27197 = new_new_n12240__ & ys__n26824;
  assign ys__n27198 = new_new_n12240__ & ys__n26826;
  assign ys__n27199 = new_new_n12240__ & ys__n26828;
  assign ys__n27200 = new_new_n12240__ & ys__n26830;
  assign ys__n27201 = new_new_n12240__ & ys__n26832;
  assign ys__n27202 = new_new_n12240__ & ys__n26834;
  assign ys__n27203 = new_new_n12240__ & ys__n26836;
  assign ys__n27204 = new_new_n12240__ & ys__n26838;
  assign ys__n27205 = new_new_n12240__ & ys__n26840;
  assign ys__n27206 = new_new_n12240__ & ys__n26842;
  assign ys__n27207 = new_new_n12240__ & ys__n26844;
  assign ys__n27208 = new_new_n12240__ & ys__n26846;
  assign ys__n27209 = new_new_n12240__ & ys__n26848;
  assign ys__n27210 = new_new_n12240__ & ys__n26850;
  assign ys__n27211 = new_new_n12240__ & ys__n26852;
  assign ys__n27212 = new_new_n12240__ & ys__n26854;
  assign ys__n27213 = new_new_n12240__ & ys__n26856;
  assign ys__n27214 = new_new_n12240__ & ys__n26858;
  assign ys__n27215 = new_new_n12240__ & ys__n26860;
  assign ys__n27216 = new_new_n12240__ & ys__n26862;
  assign ys__n27217 = new_new_n12240__ & ys__n26864;
  assign ys__n27218 = new_new_n12240__ & ys__n26866;
  assign ys__n27219 = new_new_n12240__ & ys__n26868;
  assign ys__n27220 = new_new_n12240__ & ys__n26870;
  assign ys__n27221 = new_new_n12240__ & ys__n26872;
  assign ys__n27222 = new_new_n12240__ & ys__n26874;
  assign ys__n27223 = new_new_n12240__ & ys__n26876;
  assign ys__n27224 = new_new_n12240__ & ys__n26878;
  assign ys__n27225 = new_new_n12240__ & ys__n26880;
  assign ys__n27226 = new_new_n12240__ & ys__n26882;
  assign ys__n27227 = new_new_n12240__ & ys__n26884;
  assign ys__n27228 = new_new_n12240__ & ys__n26886;
  assign ys__n27229 = new_new_n12240__ & ys__n26888;
  assign ys__n27230 = new_new_n12240__ & ys__n26890;
  assign ys__n27231 = new_new_n12240__ & ys__n26892;
  assign ys__n27232 = new_new_n12240__ & ys__n26894;
  assign ys__n27233 = new_new_n12240__ & ys__n26896;
  assign ys__n27234 = new_new_n12240__ & ys__n26898;
  assign ys__n27235 = new_new_n12240__ & ys__n26900;
  assign ys__n27236 = new_new_n12240__ & ys__n26902;
  assign ys__n27237 = new_new_n12240__ & ys__n26904;
  assign ys__n27238 = new_new_n12240__ & ys__n26906;
  assign ys__n27239 = new_new_n12240__ & ys__n26908;
  assign ys__n27240 = new_new_n12240__ & ys__n26910;
  assign ys__n27241 = new_new_n12240__ & ys__n26912;
  assign ys__n27242 = new_new_n12240__ & ys__n26914;
  assign ys__n27243 = new_new_n12240__ & ys__n26916;
  assign ys__n27244 = new_new_n12240__ & ys__n26918;
  assign ys__n27245 = new_new_n12240__ & ys__n26920;
  assign ys__n27246 = new_new_n12240__ & ys__n26922;
  assign ys__n27247 = new_new_n12240__ & ys__n26924;
  assign ys__n27248 = new_new_n12240__ & ys__n26926;
  assign ys__n27249 = new_new_n12240__ & ys__n26928;
  assign ys__n27250 = new_new_n12240__ & ys__n26930;
  assign ys__n27251 = new_new_n12240__ & ys__n26932;
  assign ys__n27252 = new_new_n12240__ & ys__n26934;
  assign ys__n27253 = new_new_n12240__ & ys__n26936;
  assign ys__n27254 = new_new_n12240__ & ys__n26938;
  assign ys__n27255 = new_new_n12240__ & ys__n26940;
  assign ys__n27256 = new_new_n12240__ & ys__n26942;
  assign ys__n27257 = new_new_n12240__ & ys__n26944;
  assign ys__n27258 = new_new_n12240__ & ys__n26946;
  assign ys__n27259 = new_new_n12240__ & ys__n26948;
  assign ys__n27260 = new_new_n12240__ & ys__n26950;
  assign ys__n27261 = new_new_n12240__ & ys__n26952;
  assign ys__n27262 = new_new_n12240__ & ys__n26954;
  assign ys__n27263 = new_new_n12240__ & ys__n26956;
  assign ys__n27264 = new_new_n12240__ & ys__n26958;
  assign ys__n27265 = new_new_n12240__ & ys__n26960;
  assign ys__n27266 = new_new_n12240__ & ys__n26962;
  assign ys__n27267 = new_new_n12240__ & ys__n26964;
  assign ys__n27268 = new_new_n12240__ & ys__n26966;
  assign ys__n27269 = new_new_n12240__ & ys__n26968;
  assign ys__n27270 = new_new_n12240__ & ys__n26970;
  assign ys__n27271 = new_new_n12240__ & ys__n26972;
  assign ys__n27272 = new_new_n12240__ & ys__n26974;
  assign ys__n27273 = new_new_n12240__ & ys__n26976;
  assign ys__n27274 = new_new_n12240__ & ys__n26978;
  assign ys__n27275 = new_new_n12240__ & ys__n26980;
  assign ys__n27276 = new_new_n12240__ & ys__n26982;
  assign ys__n27277 = new_new_n12240__ & ys__n26984;
  assign ys__n27278 = new_new_n12240__ & ys__n26986;
  assign ys__n27279 = new_new_n12240__ & ys__n26988;
  assign ys__n27280 = new_new_n12240__ & ys__n26990;
  assign ys__n27281 = new_new_n12240__ & ys__n26992;
  assign ys__n27282 = new_new_n12240__ & ys__n26994;
  assign ys__n27283 = new_new_n12240__ & ys__n26996;
  assign ys__n27284 = new_new_n12240__ & ys__n26998;
  assign ys__n27285 = new_new_n12240__ & ys__n27000;
  assign ys__n27286 = new_new_n12240__ & ys__n27002;
  assign ys__n27287 = new_new_n12240__ & ys__n27004;
  assign ys__n27288 = new_new_n12240__ & ys__n27006;
  assign ys__n27289 = new_new_n12240__ & ys__n27008;
  assign ys__n27290 = new_new_n12240__ & ys__n27010;
  assign ys__n27291 = new_new_n12240__ & ys__n27012;
  assign ys__n27292 = new_new_n12240__ & ys__n27014;
  assign ys__n27293 = new_new_n12240__ & ys__n27016;
  assign ys__n27294 = new_new_n12240__ & ys__n27018;
  assign ys__n27295 = new_new_n12240__ & ys__n27020;
  assign ys__n27296 = new_new_n12240__ & ys__n27022;
  assign ys__n27297 = new_new_n12240__ & ys__n27024;
  assign ys__n27298 = new_new_n12240__ & ys__n27026;
  assign ys__n27299 = new_new_n12240__ & ys__n27028;
  assign ys__n27300 = new_new_n12240__ & ys__n27030;
  assign ys__n27301 = new_new_n12240__ & ys__n27032;
  assign ys__n27302 = new_new_n12240__ & ys__n27034;
  assign ys__n27303 = new_new_n12240__ & ys__n27036;
  assign ys__n27304 = new_new_n12240__ & ys__n27038;
  assign ys__n27305 = new_new_n12240__ & ys__n27040;
  assign ys__n27306 = new_new_n12240__ & ys__n27042;
  assign ys__n27307 = new_new_n12240__ & ys__n27044;
  assign ys__n27308 = new_new_n12240__ & ys__n27046;
  assign ys__n27309 = new_new_n12240__ & ys__n27048;
  assign ys__n27310 = new_new_n12240__ & ys__n27050;
  assign ys__n27311 = new_new_n12240__ & ys__n27052;
  assign ys__n27312 = new_new_n12240__ & ys__n27054;
  assign ys__n27313 = new_new_n12240__ & ys__n27056;
  assign ys__n27314 = new_new_n12241__ & ys__n26804;
  assign ys__n27315 = new_new_n12241__ & ys__n26806;
  assign ys__n27316 = new_new_n12241__ & ys__n26808;
  assign ys__n27317 = new_new_n12241__ & ys__n26810;
  assign ys__n27318 = new_new_n12241__ & ys__n26812;
  assign ys__n27319 = new_new_n12241__ & ys__n26814;
  assign ys__n27320 = new_new_n12241__ & ys__n26816;
  assign ys__n27321 = new_new_n12241__ & ys__n26818;
  assign ys__n27322 = new_new_n12241__ & ys__n26820;
  assign ys__n27323 = new_new_n12241__ & ys__n26822;
  assign ys__n27324 = new_new_n12241__ & ys__n26824;
  assign ys__n27325 = new_new_n12241__ & ys__n26826;
  assign ys__n27326 = new_new_n12241__ & ys__n26828;
  assign ys__n27327 = new_new_n12241__ & ys__n26830;
  assign ys__n27328 = new_new_n12241__ & ys__n26832;
  assign ys__n27329 = new_new_n12241__ & ys__n26834;
  assign ys__n27330 = new_new_n12241__ & ys__n26836;
  assign ys__n27331 = new_new_n12241__ & ys__n26838;
  assign ys__n27332 = new_new_n12241__ & ys__n26840;
  assign ys__n27333 = new_new_n12241__ & ys__n26842;
  assign ys__n27334 = new_new_n12241__ & ys__n26844;
  assign ys__n27335 = new_new_n12241__ & ys__n26846;
  assign ys__n27336 = new_new_n12241__ & ys__n26848;
  assign ys__n27337 = new_new_n12241__ & ys__n26850;
  assign ys__n27338 = new_new_n12241__ & ys__n26852;
  assign ys__n27339 = new_new_n12241__ & ys__n26854;
  assign ys__n27340 = new_new_n12241__ & ys__n26856;
  assign ys__n27341 = new_new_n12241__ & ys__n26858;
  assign ys__n27342 = new_new_n12241__ & ys__n26860;
  assign ys__n27343 = new_new_n12241__ & ys__n26862;
  assign ys__n27344 = new_new_n12241__ & ys__n26864;
  assign ys__n27345 = new_new_n12241__ & ys__n26868;
  assign ys__n27346 = new_new_n12241__ & ys__n26870;
  assign ys__n27347 = new_new_n12241__ & ys__n26872;
  assign ys__n27348 = new_new_n12241__ & ys__n26874;
  assign ys__n27349 = new_new_n12241__ & ys__n26876;
  assign ys__n27350 = new_new_n12241__ & ys__n26878;
  assign ys__n27351 = new_new_n12241__ & ys__n26880;
  assign ys__n27352 = new_new_n12241__ & ys__n26882;
  assign ys__n27353 = new_new_n12241__ & ys__n26884;
  assign ys__n27354 = new_new_n12241__ & ys__n26886;
  assign ys__n27355 = new_new_n12241__ & ys__n26888;
  assign ys__n27356 = new_new_n12241__ & ys__n26890;
  assign ys__n27357 = new_new_n12241__ & ys__n26892;
  assign ys__n27358 = new_new_n12241__ & ys__n26894;
  assign ys__n27359 = new_new_n12241__ & ys__n26896;
  assign ys__n27360 = new_new_n12241__ & ys__n26898;
  assign ys__n27361 = new_new_n12241__ & ys__n26900;
  assign ys__n27362 = new_new_n12241__ & ys__n26902;
  assign ys__n27363 = new_new_n12241__ & ys__n26904;
  assign ys__n27364 = new_new_n12241__ & ys__n26906;
  assign ys__n27365 = new_new_n12241__ & ys__n26908;
  assign ys__n27366 = new_new_n12241__ & ys__n26910;
  assign ys__n27367 = new_new_n12241__ & ys__n26912;
  assign ys__n27368 = new_new_n12241__ & ys__n26914;
  assign ys__n27369 = new_new_n12241__ & ys__n26916;
  assign ys__n27370 = new_new_n12241__ & ys__n26918;
  assign ys__n27371 = new_new_n12241__ & ys__n26920;
  assign ys__n27372 = new_new_n12241__ & ys__n26922;
  assign ys__n27373 = new_new_n12241__ & ys__n26924;
  assign ys__n27374 = new_new_n12241__ & ys__n26926;
  assign ys__n27375 = new_new_n12241__ & ys__n26928;
  assign ys__n27376 = new_new_n12241__ & ys__n26932;
  assign ys__n27377 = new_new_n12241__ & ys__n26934;
  assign ys__n27378 = new_new_n12241__ & ys__n26936;
  assign ys__n27379 = new_new_n12241__ & ys__n26938;
  assign ys__n27380 = new_new_n12241__ & ys__n26940;
  assign ys__n27381 = new_new_n12241__ & ys__n26942;
  assign ys__n27382 = new_new_n12241__ & ys__n26944;
  assign ys__n27383 = new_new_n12241__ & ys__n26946;
  assign ys__n27384 = new_new_n12241__ & ys__n26948;
  assign ys__n27385 = new_new_n12241__ & ys__n26950;
  assign ys__n27386 = new_new_n12241__ & ys__n26952;
  assign ys__n27387 = new_new_n12241__ & ys__n26954;
  assign ys__n27388 = new_new_n12241__ & ys__n26956;
  assign ys__n27389 = new_new_n12241__ & ys__n26958;
  assign ys__n27390 = new_new_n12241__ & ys__n26960;
  assign ys__n27391 = new_new_n12241__ & ys__n26962;
  assign ys__n27392 = new_new_n12241__ & ys__n26964;
  assign ys__n27393 = new_new_n12241__ & ys__n26966;
  assign ys__n27394 = new_new_n12241__ & ys__n26968;
  assign ys__n27395 = new_new_n12241__ & ys__n26970;
  assign ys__n27396 = new_new_n12241__ & ys__n26972;
  assign ys__n27397 = new_new_n12241__ & ys__n26974;
  assign ys__n27398 = new_new_n12241__ & ys__n26976;
  assign ys__n27399 = new_new_n12241__ & ys__n26978;
  assign ys__n27400 = new_new_n12241__ & ys__n26980;
  assign ys__n27401 = new_new_n12241__ & ys__n26982;
  assign ys__n27402 = new_new_n12241__ & ys__n26984;
  assign ys__n27403 = new_new_n12241__ & ys__n26986;
  assign ys__n27404 = new_new_n12241__ & ys__n26988;
  assign ys__n27405 = new_new_n12241__ & ys__n26990;
  assign ys__n27406 = new_new_n12241__ & ys__n26992;
  assign ys__n27407 = new_new_n12241__ & ys__n26996;
  assign ys__n27408 = new_new_n12241__ & ys__n26998;
  assign ys__n27409 = new_new_n12241__ & ys__n27000;
  assign ys__n27410 = new_new_n12241__ & ys__n27002;
  assign ys__n27411 = new_new_n12241__ & ys__n27004;
  assign ys__n27412 = new_new_n12241__ & ys__n27006;
  assign ys__n27413 = new_new_n12241__ & ys__n27008;
  assign ys__n27414 = new_new_n12241__ & ys__n27010;
  assign ys__n27415 = new_new_n12241__ & ys__n27012;
  assign ys__n27416 = new_new_n12241__ & ys__n27014;
  assign ys__n27417 = new_new_n12241__ & ys__n27016;
  assign ys__n27418 = new_new_n12241__ & ys__n27018;
  assign ys__n27419 = new_new_n12241__ & ys__n27020;
  assign ys__n27420 = new_new_n12241__ & ys__n27022;
  assign ys__n27421 = new_new_n12241__ & ys__n27024;
  assign ys__n27422 = new_new_n12241__ & ys__n27026;
  assign ys__n27423 = new_new_n12241__ & ys__n27028;
  assign ys__n27424 = new_new_n12241__ & ys__n27030;
  assign ys__n27425 = new_new_n12241__ & ys__n27032;
  assign ys__n27426 = new_new_n12241__ & ys__n27034;
  assign ys__n27427 = new_new_n12241__ & ys__n27036;
  assign ys__n27428 = new_new_n12241__ & ys__n27038;
  assign ys__n27429 = new_new_n12241__ & ys__n27040;
  assign ys__n27430 = new_new_n12241__ & ys__n27042;
  assign ys__n27431 = new_new_n12241__ & ys__n27044;
  assign ys__n27432 = new_new_n12241__ & ys__n27046;
  assign ys__n27433 = new_new_n12241__ & ys__n27048;
  assign ys__n27434 = new_new_n12241__ & ys__n27050;
  assign ys__n27435 = new_new_n12241__ & ys__n27052;
  assign ys__n27436 = new_new_n12241__ & ys__n27054;
  assign ys__n27437 = new_new_n12241__ & ys__n27056;
  assign new_new_n32232__ = ys__n26766 & ~new_new_n26767__;
  assign new_new_n32233__ = ys__n26766 & ~new_new_n26703__;
  assign new_new_n32234__ = ~new_new_n26705__ & ~new_new_n32233__;
  assign new_new_n32235__ = new_new_n26767__ & ~new_new_n32234__;
  assign new_new_n32236__ = ~new_new_n32232__ & ~new_new_n32235__;
  assign new_new_n32237__ = ys__n6126 & ys__n46936;
  assign new_new_n32238__ = ~ys__n6126 & ~ys__n46936;
  assign new_new_n32239__ = ~ys__n46906 & ~new_new_n32238__;
  assign new_new_n32240__ = ~new_new_n32237__ & new_new_n32239__;
  assign new_new_n32241__ = ys__n6127 & ys__n46937;
  assign new_new_n32242__ = ~ys__n6127 & ~ys__n46937;
  assign new_new_n32243__ = ~ys__n46908 & ~new_new_n32242__;
  assign new_new_n32244__ = ~new_new_n32241__ & new_new_n32243__;
  assign new_new_n32245__ = ~new_new_n32240__ & ~new_new_n32244__;
  assign new_new_n32246__ = ys__n6129 & ys__n46938;
  assign new_new_n32247__ = ~ys__n6129 & ~ys__n46938;
  assign new_new_n32248__ = ~ys__n46910 & ~new_new_n32247__;
  assign new_new_n32249__ = ~new_new_n32246__ & new_new_n32248__;
  assign new_new_n32250__ = ys__n6130 & ys__n46939;
  assign new_new_n32251__ = ~ys__n6130 & ~ys__n46939;
  assign new_new_n32252__ = ~ys__n46912 & ~new_new_n32251__;
  assign new_new_n32253__ = ~new_new_n32250__ & new_new_n32252__;
  assign new_new_n32254__ = ~new_new_n32249__ & ~new_new_n32253__;
  assign new_new_n32255__ = new_new_n32245__ & new_new_n32254__;
  assign new_new_n32256__ = ys__n6120 & ys__n46932;
  assign new_new_n32257__ = ~ys__n6120 & ~ys__n46932;
  assign new_new_n32258__ = ~ys__n46898 & ~new_new_n32257__;
  assign new_new_n32259__ = ~new_new_n32256__ & new_new_n32258__;
  assign new_new_n32260__ = ys__n6121 & ys__n46933;
  assign new_new_n32261__ = ~ys__n6121 & ~ys__n46933;
  assign new_new_n32262__ = ~ys__n46900 & ~new_new_n32261__;
  assign new_new_n32263__ = ~new_new_n32260__ & new_new_n32262__;
  assign new_new_n32264__ = ~new_new_n32259__ & ~new_new_n32263__;
  assign new_new_n32265__ = ys__n6123 & ys__n46934;
  assign new_new_n32266__ = ~ys__n6123 & ~ys__n46934;
  assign new_new_n32267__ = ~ys__n46902 & ~new_new_n32266__;
  assign new_new_n32268__ = ~new_new_n32265__ & new_new_n32267__;
  assign new_new_n32269__ = ys__n6124 & ys__n46935;
  assign new_new_n32270__ = ~ys__n6124 & ~ys__n46935;
  assign new_new_n32271__ = ~ys__n46904 & ~new_new_n32270__;
  assign new_new_n32272__ = ~new_new_n32269__ & new_new_n32271__;
  assign new_new_n32273__ = ~new_new_n32268__ & ~new_new_n32272__;
  assign new_new_n32274__ = new_new_n32264__ & new_new_n32273__;
  assign new_new_n32275__ = new_new_n32255__ & new_new_n32274__;
  assign new_new_n32276__ = ys__n18448 & ys__n46843;
  assign new_new_n32277__ = ~ys__n18448 & ~ys__n46843;
  assign new_new_n32278__ = ~ys__n46780 & ~new_new_n32277__;
  assign new_new_n32279__ = ~new_new_n32276__ & new_new_n32278__;
  assign new_new_n32280__ = ys__n18451 & ys__n46844;
  assign new_new_n32281__ = ~ys__n18451 & ~ys__n46844;
  assign new_new_n32282__ = ~ys__n46782 & ~new_new_n32281__;
  assign new_new_n32283__ = ~new_new_n32280__ & new_new_n32282__;
  assign new_new_n32284__ = ~new_new_n32279__ & ~new_new_n32283__;
  assign new_new_n32285__ = ys__n18454 & ys__n46845;
  assign new_new_n32286__ = ~ys__n18454 & ~ys__n46845;
  assign new_new_n32287__ = ~ys__n46784 & ~new_new_n32286__;
  assign new_new_n32288__ = ~new_new_n32285__ & new_new_n32287__;
  assign new_new_n32289__ = ys__n18457 & ys__n46846;
  assign new_new_n32290__ = ~ys__n18457 & ~ys__n46846;
  assign new_new_n32291__ = ~ys__n46786 & ~new_new_n32290__;
  assign new_new_n32292__ = ~new_new_n32289__ & new_new_n32291__;
  assign new_new_n32293__ = ~new_new_n32288__ & ~new_new_n32292__;
  assign new_new_n32294__ = new_new_n32284__ & new_new_n32293__;
  assign new_new_n32295__ = ys__n42 & ys__n46940;
  assign new_new_n32296__ = ~ys__n42 & ~ys__n46940;
  assign new_new_n32297__ = ~ys__n46914 & ~new_new_n32296__;
  assign new_new_n32298__ = ~new_new_n32295__ & new_new_n32297__;
  assign new_new_n32299__ = ys__n40 & ys__n46941;
  assign new_new_n32300__ = ~ys__n40 & ~ys__n46941;
  assign new_new_n32301__ = ~ys__n46916 & ~new_new_n32300__;
  assign new_new_n32302__ = ~new_new_n32299__ & new_new_n32301__;
  assign new_new_n32303__ = ~new_new_n32298__ & ~new_new_n32302__;
  assign new_new_n32304__ = ys__n6133 & ys__n46942;
  assign new_new_n32305__ = ~ys__n6133 & ~ys__n46942;
  assign new_new_n32306__ = ~ys__n46918 & ~new_new_n32305__;
  assign new_new_n32307__ = ~new_new_n32304__ & new_new_n32306__;
  assign new_new_n32308__ = ys__n6134 & ys__n46943;
  assign new_new_n32309__ = ~ys__n6134 & ~ys__n46943;
  assign new_new_n32310__ = ~ys__n46920 & ~new_new_n32309__;
  assign new_new_n32311__ = ~new_new_n32308__ & new_new_n32310__;
  assign new_new_n32312__ = ~new_new_n32307__ & ~new_new_n32311__;
  assign new_new_n32313__ = new_new_n32303__ & new_new_n32312__;
  assign new_new_n32314__ = new_new_n32294__ & new_new_n32313__;
  assign new_new_n32315__ = new_new_n32275__ & new_new_n32314__;
  assign new_new_n32316__ = ys__n6113 & ys__n46921;
  assign new_new_n32317__ = ~ys__n6113 & ~ys__n46921;
  assign new_new_n32318__ = ~ys__n46876 & ~new_new_n32317__;
  assign new_new_n32319__ = ~new_new_n32316__ & new_new_n32318__;
  assign new_new_n32320__ = ~ys__n38 & ~ys__n46944;
  assign new_new_n32321__ = ys__n38 & ys__n46944;
  assign new_new_n32322__ = ~new_new_n32320__ & ~new_new_n32321__;
  assign new_new_n32323__ = ~ys__n36 & ~ys__n46945;
  assign new_new_n32324__ = ys__n36 & ys__n46945;
  assign new_new_n32325__ = ~new_new_n32323__ & ~new_new_n32324__;
  assign new_new_n32326__ = ~new_new_n32322__ & ~new_new_n32325__;
  assign new_new_n32327__ = ~new_new_n32319__ & new_new_n32326__;
  assign new_new_n32328__ = ys__n172 & ys__n46922;
  assign new_new_n32329__ = ~ys__n172 & ~ys__n46922;
  assign new_new_n32330__ = ~ys__n46878 & ~new_new_n32329__;
  assign new_new_n32331__ = ~new_new_n32328__ & new_new_n32330__;
  assign new_new_n32332__ = ys__n338 & ys__n46923;
  assign new_new_n32333__ = ~ys__n338 & ~ys__n46923;
  assign new_new_n32334__ = ~ys__n46880 & ~new_new_n32333__;
  assign new_new_n32335__ = ~new_new_n32332__ & new_new_n32334__;
  assign new_new_n32336__ = ~new_new_n32331__ & ~new_new_n32335__;
  assign new_new_n32337__ = new_new_n32327__ & new_new_n32336__;
  assign new_new_n32338__ = ~ys__n26 & ~ys__n46950;
  assign new_new_n32339__ = ys__n26 & ys__n46950;
  assign new_new_n32340__ = ~new_new_n32338__ & ~new_new_n32339__;
  assign new_new_n32341__ = ~ys__n24 & ~ys__n46951;
  assign new_new_n32342__ = ys__n24 & ys__n46951;
  assign new_new_n32343__ = ~new_new_n32341__ & ~new_new_n32342__;
  assign new_new_n32344__ = ~new_new_n32340__ & ~new_new_n32343__;
  assign new_new_n32345__ = ~ys__n46230 & ys__n46231;
  assign new_new_n32346__ = ys__n46230 & ~ys__n46231;
  assign new_new_n32347__ = ~new_new_n32345__ & ~new_new_n32346__;
  assign new_new_n32348__ = ys__n18059 & ys__n18065;
  assign new_new_n32349__ = ~ys__n27479 & new_new_n32348__;
  assign new_new_n32350__ = ~new_new_n32347__ & ~new_new_n32349__;
  assign new_new_n32351__ = new_new_n32344__ & new_new_n32350__;
  assign new_new_n32352__ = ~ys__n34 & ~ys__n46946;
  assign new_new_n32353__ = ys__n34 & ys__n46946;
  assign new_new_n32354__ = ~new_new_n32352__ & ~new_new_n32353__;
  assign new_new_n32355__ = ~ys__n32 & ~ys__n46947;
  assign new_new_n32356__ = ys__n32 & ys__n46947;
  assign new_new_n32357__ = ~new_new_n32355__ & ~new_new_n32356__;
  assign new_new_n32358__ = ~new_new_n32354__ & ~new_new_n32357__;
  assign new_new_n32359__ = ~ys__n30 & ~ys__n46948;
  assign new_new_n32360__ = ys__n30 & ys__n46948;
  assign new_new_n32361__ = ~new_new_n32359__ & ~new_new_n32360__;
  assign new_new_n32362__ = ~ys__n28 & ~ys__n46949;
  assign new_new_n32363__ = ys__n28 & ys__n46949;
  assign new_new_n32364__ = ~new_new_n32362__ & ~new_new_n32363__;
  assign new_new_n32365__ = ~new_new_n32361__ & ~new_new_n32364__;
  assign new_new_n32366__ = new_new_n32358__ & new_new_n32365__;
  assign new_new_n32367__ = new_new_n32351__ & new_new_n32366__;
  assign new_new_n32368__ = new_new_n32337__ & new_new_n32367__;
  assign new_new_n32369__ = ys__n340 & ys__n46928;
  assign new_new_n32370__ = ~ys__n340 & ~ys__n46928;
  assign new_new_n32371__ = ~ys__n46890 & ~new_new_n32370__;
  assign new_new_n32372__ = ~new_new_n32369__ & new_new_n32371__;
  assign new_new_n32373__ = ys__n46 & ys__n46929;
  assign new_new_n32374__ = ~ys__n46 & ~ys__n46929;
  assign new_new_n32375__ = ~ys__n46892 & ~new_new_n32374__;
  assign new_new_n32376__ = ~new_new_n32373__ & new_new_n32375__;
  assign new_new_n32377__ = ~new_new_n32372__ & ~new_new_n32376__;
  assign new_new_n32378__ = ys__n6118 & ys__n46930;
  assign new_new_n32379__ = ~ys__n6118 & ~ys__n46930;
  assign new_new_n32380__ = ~ys__n46894 & ~new_new_n32379__;
  assign new_new_n32381__ = ~new_new_n32378__ & new_new_n32380__;
  assign new_new_n32382__ = ys__n6119 & ys__n46931;
  assign new_new_n32383__ = ~ys__n6119 & ~ys__n46931;
  assign new_new_n32384__ = ~ys__n46896 & ~new_new_n32383__;
  assign new_new_n32385__ = ~new_new_n32382__ & new_new_n32384__;
  assign new_new_n32386__ = ~new_new_n32381__ & ~new_new_n32385__;
  assign new_new_n32387__ = new_new_n32377__ & new_new_n32386__;
  assign new_new_n32388__ = ys__n22 & ys__n46924;
  assign new_new_n32389__ = ~ys__n22 & ~ys__n46924;
  assign new_new_n32390__ = ~ys__n46882 & ~new_new_n32389__;
  assign new_new_n32391__ = ~new_new_n32388__ & new_new_n32390__;
  assign new_new_n32392__ = ys__n316 & ys__n46925;
  assign new_new_n32393__ = ~ys__n316 & ~ys__n46925;
  assign new_new_n32394__ = ~ys__n46884 & ~new_new_n32393__;
  assign new_new_n32395__ = ~new_new_n32392__ & new_new_n32394__;
  assign new_new_n32396__ = ~new_new_n32391__ & ~new_new_n32395__;
  assign new_new_n32397__ = ys__n6115 & ys__n46926;
  assign new_new_n32398__ = ~ys__n6115 & ~ys__n46926;
  assign new_new_n32399__ = ~ys__n46886 & ~new_new_n32398__;
  assign new_new_n32400__ = ~new_new_n32397__ & new_new_n32399__;
  assign new_new_n32401__ = ys__n44 & ys__n46927;
  assign new_new_n32402__ = ~ys__n44 & ~ys__n46927;
  assign new_new_n32403__ = ~ys__n46888 & ~new_new_n32402__;
  assign new_new_n32404__ = ~new_new_n32401__ & new_new_n32403__;
  assign new_new_n32405__ = ~new_new_n32400__ & ~new_new_n32404__;
  assign new_new_n32406__ = new_new_n32396__ & new_new_n32405__;
  assign new_new_n32407__ = new_new_n32387__ & new_new_n32406__;
  assign new_new_n32408__ = new_new_n32368__ & new_new_n32407__;
  assign new_new_n32409__ = new_new_n32315__ & new_new_n32408__;
  assign new_new_n32410__ = ys__n18520 & ys__n46867;
  assign new_new_n32411__ = ~ys__n18520 & ~ys__n46867;
  assign new_new_n32412__ = ~ys__n46828 & ~new_new_n32411__;
  assign new_new_n32413__ = ~new_new_n32410__ & new_new_n32412__;
  assign new_new_n32414__ = ys__n18523 & ys__n46868;
  assign new_new_n32415__ = ~ys__n18523 & ~ys__n46868;
  assign new_new_n32416__ = ~ys__n46830 & ~new_new_n32415__;
  assign new_new_n32417__ = ~new_new_n32414__ & new_new_n32416__;
  assign new_new_n32418__ = ~new_new_n32413__ & ~new_new_n32417__;
  assign new_new_n32419__ = ys__n18526 & ys__n46869;
  assign new_new_n32420__ = ~ys__n18526 & ~ys__n46869;
  assign new_new_n32421__ = ~ys__n46832 & ~new_new_n32420__;
  assign new_new_n32422__ = ~new_new_n32419__ & new_new_n32421__;
  assign new_new_n32423__ = ys__n18529 & ys__n46870;
  assign new_new_n32424__ = ~ys__n18529 & ~ys__n46870;
  assign new_new_n32425__ = ~ys__n46834 & ~new_new_n32424__;
  assign new_new_n32426__ = ~new_new_n32423__ & new_new_n32425__;
  assign new_new_n32427__ = ~new_new_n32422__ & ~new_new_n32426__;
  assign new_new_n32428__ = new_new_n32418__ & new_new_n32427__;
  assign new_new_n32429__ = ys__n18508 & ys__n46863;
  assign new_new_n32430__ = ~ys__n18508 & ~ys__n46863;
  assign new_new_n32431__ = ~ys__n46820 & ~new_new_n32430__;
  assign new_new_n32432__ = ~new_new_n32429__ & new_new_n32431__;
  assign new_new_n32433__ = ys__n18511 & ys__n46864;
  assign new_new_n32434__ = ~ys__n18511 & ~ys__n46864;
  assign new_new_n32435__ = ~ys__n46822 & ~new_new_n32434__;
  assign new_new_n32436__ = ~new_new_n32433__ & new_new_n32435__;
  assign new_new_n32437__ = ~new_new_n32432__ & ~new_new_n32436__;
  assign new_new_n32438__ = ys__n18514 & ys__n46865;
  assign new_new_n32439__ = ~ys__n18514 & ~ys__n46865;
  assign new_new_n32440__ = ~ys__n46824 & ~new_new_n32439__;
  assign new_new_n32441__ = ~new_new_n32438__ & new_new_n32440__;
  assign new_new_n32442__ = ys__n18517 & ys__n46866;
  assign new_new_n32443__ = ~ys__n18517 & ~ys__n46866;
  assign new_new_n32444__ = ~ys__n46826 & ~new_new_n32443__;
  assign new_new_n32445__ = ~new_new_n32442__ & new_new_n32444__;
  assign new_new_n32446__ = ~new_new_n32441__ & ~new_new_n32445__;
  assign new_new_n32447__ = new_new_n32437__ & new_new_n32446__;
  assign new_new_n32448__ = new_new_n32428__ & new_new_n32447__;
  assign new_new_n32449__ = ~ys__n18059 & ~ys__n18065;
  assign new_new_n32450__ = ~ys__n18208 & new_new_n32449__;
  assign new_new_n32451__ = ~ys__n18061 & new_new_n32450__;
  assign new_new_n32452__ = ys__n18059 & ~ys__n18065;
  assign new_new_n32453__ = ys__n18208 & new_new_n32452__;
  assign new_new_n32454__ = ~ys__n18067 & new_new_n32453__;
  assign new_new_n32455__ = ~ys__n18208 & new_new_n32452__;
  assign new_new_n32456__ = ~ys__n18063 & new_new_n32455__;
  assign new_new_n32457__ = ~new_new_n32454__ & ~new_new_n32456__;
  assign new_new_n32458__ = ~new_new_n32451__ & new_new_n32457__;
  assign new_new_n32459__ = ys__n18532 & ys__n46871;
  assign new_new_n32460__ = ~ys__n18532 & ~ys__n46871;
  assign new_new_n32461__ = ~ys__n46836 & ~new_new_n32460__;
  assign new_new_n32462__ = ~new_new_n32459__ & new_new_n32461__;
  assign new_new_n32463__ = ys__n18535 & ys__n46872;
  assign new_new_n32464__ = ~ys__n18535 & ~ys__n46872;
  assign new_new_n32465__ = ~ys__n46838 & ~new_new_n32464__;
  assign new_new_n32466__ = ~new_new_n32463__ & new_new_n32465__;
  assign new_new_n32467__ = ~new_new_n32462__ & ~new_new_n32466__;
  assign new_new_n32468__ = ys__n18538 & ys__n46873;
  assign new_new_n32469__ = ~ys__n18538 & ~ys__n46873;
  assign new_new_n32470__ = ~ys__n46840 & ~new_new_n32469__;
  assign new_new_n32471__ = ~new_new_n32468__ & new_new_n32470__;
  assign new_new_n32472__ = ys__n18541 & ys__n46874;
  assign new_new_n32473__ = ~ys__n18541 & ~ys__n46874;
  assign new_new_n32474__ = ~ys__n46842 & ~new_new_n32473__;
  assign new_new_n32475__ = ~new_new_n32472__ & new_new_n32474__;
  assign new_new_n32476__ = ~new_new_n32471__ & ~new_new_n32475__;
  assign new_new_n32477__ = new_new_n32467__ & new_new_n32476__;
  assign new_new_n32478__ = new_new_n32458__ & new_new_n32477__;
  assign new_new_n32479__ = new_new_n32448__ & new_new_n32478__;
  assign new_new_n32480__ = ys__n18472 & ys__n46851;
  assign new_new_n32481__ = ~ys__n18472 & ~ys__n46851;
  assign new_new_n32482__ = ~ys__n46796 & ~new_new_n32481__;
  assign new_new_n32483__ = ~new_new_n32480__ & new_new_n32482__;
  assign new_new_n32484__ = ys__n18475 & ys__n46852;
  assign new_new_n32485__ = ~ys__n18475 & ~ys__n46852;
  assign new_new_n32486__ = ~ys__n46798 & ~new_new_n32485__;
  assign new_new_n32487__ = ~new_new_n32484__ & new_new_n32486__;
  assign new_new_n32488__ = ~new_new_n32483__ & ~new_new_n32487__;
  assign new_new_n32489__ = ys__n18478 & ys__n46853;
  assign new_new_n32490__ = ~ys__n18478 & ~ys__n46853;
  assign new_new_n32491__ = ~ys__n46800 & ~new_new_n32490__;
  assign new_new_n32492__ = ~new_new_n32489__ & new_new_n32491__;
  assign new_new_n32493__ = ys__n18481 & ys__n46854;
  assign new_new_n32494__ = ~ys__n18481 & ~ys__n46854;
  assign new_new_n32495__ = ~ys__n46802 & ~new_new_n32494__;
  assign new_new_n32496__ = ~new_new_n32493__ & new_new_n32495__;
  assign new_new_n32497__ = ~new_new_n32492__ & ~new_new_n32496__;
  assign new_new_n32498__ = new_new_n32488__ & new_new_n32497__;
  assign new_new_n32499__ = ys__n18460 & ys__n46847;
  assign new_new_n32500__ = ~ys__n18460 & ~ys__n46847;
  assign new_new_n32501__ = ~ys__n46788 & ~new_new_n32500__;
  assign new_new_n32502__ = ~new_new_n32499__ & new_new_n32501__;
  assign new_new_n32503__ = ys__n18463 & ys__n46848;
  assign new_new_n32504__ = ~ys__n18463 & ~ys__n46848;
  assign new_new_n32505__ = ~ys__n46790 & ~new_new_n32504__;
  assign new_new_n32506__ = ~new_new_n32503__ & new_new_n32505__;
  assign new_new_n32507__ = ~new_new_n32502__ & ~new_new_n32506__;
  assign new_new_n32508__ = ys__n18466 & ys__n46849;
  assign new_new_n32509__ = ~ys__n18466 & ~ys__n46849;
  assign new_new_n32510__ = ~ys__n46792 & ~new_new_n32509__;
  assign new_new_n32511__ = ~new_new_n32508__ & new_new_n32510__;
  assign new_new_n32512__ = ys__n18469 & ys__n46850;
  assign new_new_n32513__ = ~ys__n18469 & ~ys__n46850;
  assign new_new_n32514__ = ~ys__n46794 & ~new_new_n32513__;
  assign new_new_n32515__ = ~new_new_n32512__ & new_new_n32514__;
  assign new_new_n32516__ = ~new_new_n32511__ & ~new_new_n32515__;
  assign new_new_n32517__ = new_new_n32507__ & new_new_n32516__;
  assign new_new_n32518__ = new_new_n32498__ & new_new_n32517__;
  assign new_new_n32519__ = ys__n18496 & ys__n46859;
  assign new_new_n32520__ = ~ys__n18496 & ~ys__n46859;
  assign new_new_n32521__ = ~ys__n46812 & ~new_new_n32520__;
  assign new_new_n32522__ = ~new_new_n32519__ & new_new_n32521__;
  assign new_new_n32523__ = ys__n18499 & ys__n46860;
  assign new_new_n32524__ = ~ys__n18499 & ~ys__n46860;
  assign new_new_n32525__ = ~ys__n46814 & ~new_new_n32524__;
  assign new_new_n32526__ = ~new_new_n32523__ & new_new_n32525__;
  assign new_new_n32527__ = ~new_new_n32522__ & ~new_new_n32526__;
  assign new_new_n32528__ = ys__n18502 & ys__n46861;
  assign new_new_n32529__ = ~ys__n18502 & ~ys__n46861;
  assign new_new_n32530__ = ~ys__n46816 & ~new_new_n32529__;
  assign new_new_n32531__ = ~new_new_n32528__ & new_new_n32530__;
  assign new_new_n32532__ = ys__n18505 & ys__n46862;
  assign new_new_n32533__ = ~ys__n18505 & ~ys__n46862;
  assign new_new_n32534__ = ~ys__n46818 & ~new_new_n32533__;
  assign new_new_n32535__ = ~new_new_n32532__ & new_new_n32534__;
  assign new_new_n32536__ = ~new_new_n32531__ & ~new_new_n32535__;
  assign new_new_n32537__ = new_new_n32527__ & new_new_n32536__;
  assign new_new_n32538__ = ys__n18484 & ys__n46855;
  assign new_new_n32539__ = ~ys__n18484 & ~ys__n46855;
  assign new_new_n32540__ = ~ys__n46804 & ~new_new_n32539__;
  assign new_new_n32541__ = ~new_new_n32538__ & new_new_n32540__;
  assign new_new_n32542__ = ys__n18487 & ys__n46856;
  assign new_new_n32543__ = ~ys__n18487 & ~ys__n46856;
  assign new_new_n32544__ = ~ys__n46806 & ~new_new_n32543__;
  assign new_new_n32545__ = ~new_new_n32542__ & new_new_n32544__;
  assign new_new_n32546__ = ~new_new_n32541__ & ~new_new_n32545__;
  assign new_new_n32547__ = ys__n18490 & ys__n46857;
  assign new_new_n32548__ = ~ys__n18490 & ~ys__n46857;
  assign new_new_n32549__ = ~ys__n46808 & ~new_new_n32548__;
  assign new_new_n32550__ = ~new_new_n32547__ & new_new_n32549__;
  assign new_new_n32551__ = ys__n18493 & ys__n46858;
  assign new_new_n32552__ = ~ys__n18493 & ~ys__n46858;
  assign new_new_n32553__ = ~ys__n46810 & ~new_new_n32552__;
  assign new_new_n32554__ = ~new_new_n32551__ & new_new_n32553__;
  assign new_new_n32555__ = ~new_new_n32550__ & ~new_new_n32554__;
  assign new_new_n32556__ = new_new_n32546__ & new_new_n32555__;
  assign new_new_n32557__ = new_new_n32537__ & new_new_n32556__;
  assign new_new_n32558__ = new_new_n32518__ & new_new_n32557__;
  assign new_new_n32559__ = new_new_n32479__ & new_new_n32558__;
  assign new_new_n32560__ = new_new_n32409__ & new_new_n32559__;
  assign new_new_n32561__ = ~new_new_n32236__ & ~new_new_n32560__;
  assign new_new_n32562__ = ~ys__n27481 & ~new_new_n32236__;
  assign new_new_n32563__ = ~ys__n27481 & ~new_new_n32562__;
  assign new_new_n32564__ = ~ys__n27485 & ~new_new_n32563__;
  assign new_new_n32565__ = ~ys__n27485 & ~new_new_n32564__;
  assign new_new_n32566__ = new_new_n32560__ & ~new_new_n32565__;
  assign ys__n27484 = new_new_n32561__ | new_new_n32566__;
  assign new_new_n32568__ = ys__n26768 & ~new_new_n26767__;
  assign new_new_n32569__ = ys__n26768 & ~new_new_n26703__;
  assign new_new_n32570__ = ~new_new_n26712__ & ~new_new_n32569__;
  assign new_new_n32571__ = new_new_n26767__ & ~new_new_n32570__;
  assign new_new_n32572__ = ~new_new_n32568__ & ~new_new_n32571__;
  assign new_new_n32573__ = ys__n6126 & ys__n46760;
  assign new_new_n32574__ = ~ys__n6126 & ~ys__n46760;
  assign new_new_n32575__ = ~ys__n46730 & ~new_new_n32574__;
  assign new_new_n32576__ = ~new_new_n32573__ & new_new_n32575__;
  assign new_new_n32577__ = ys__n6127 & ys__n46761;
  assign new_new_n32578__ = ~ys__n6127 & ~ys__n46761;
  assign new_new_n32579__ = ~ys__n46732 & ~new_new_n32578__;
  assign new_new_n32580__ = ~new_new_n32577__ & new_new_n32579__;
  assign new_new_n32581__ = ~new_new_n32576__ & ~new_new_n32580__;
  assign new_new_n32582__ = ys__n6129 & ys__n46762;
  assign new_new_n32583__ = ~ys__n6129 & ~ys__n46762;
  assign new_new_n32584__ = ~ys__n46734 & ~new_new_n32583__;
  assign new_new_n32585__ = ~new_new_n32582__ & new_new_n32584__;
  assign new_new_n32586__ = ys__n6130 & ys__n46763;
  assign new_new_n32587__ = ~ys__n6130 & ~ys__n46763;
  assign new_new_n32588__ = ~ys__n46736 & ~new_new_n32587__;
  assign new_new_n32589__ = ~new_new_n32586__ & new_new_n32588__;
  assign new_new_n32590__ = ~new_new_n32585__ & ~new_new_n32589__;
  assign new_new_n32591__ = new_new_n32581__ & new_new_n32590__;
  assign new_new_n32592__ = ys__n6120 & ys__n46756;
  assign new_new_n32593__ = ~ys__n6120 & ~ys__n46756;
  assign new_new_n32594__ = ~ys__n46722 & ~new_new_n32593__;
  assign new_new_n32595__ = ~new_new_n32592__ & new_new_n32594__;
  assign new_new_n32596__ = ys__n6121 & ys__n46757;
  assign new_new_n32597__ = ~ys__n6121 & ~ys__n46757;
  assign new_new_n32598__ = ~ys__n46724 & ~new_new_n32597__;
  assign new_new_n32599__ = ~new_new_n32596__ & new_new_n32598__;
  assign new_new_n32600__ = ~new_new_n32595__ & ~new_new_n32599__;
  assign new_new_n32601__ = ys__n6123 & ys__n46758;
  assign new_new_n32602__ = ~ys__n6123 & ~ys__n46758;
  assign new_new_n32603__ = ~ys__n46726 & ~new_new_n32602__;
  assign new_new_n32604__ = ~new_new_n32601__ & new_new_n32603__;
  assign new_new_n32605__ = ys__n6124 & ys__n46759;
  assign new_new_n32606__ = ~ys__n6124 & ~ys__n46759;
  assign new_new_n32607__ = ~ys__n46728 & ~new_new_n32606__;
  assign new_new_n32608__ = ~new_new_n32605__ & new_new_n32607__;
  assign new_new_n32609__ = ~new_new_n32604__ & ~new_new_n32608__;
  assign new_new_n32610__ = new_new_n32600__ & new_new_n32609__;
  assign new_new_n32611__ = new_new_n32591__ & new_new_n32610__;
  assign new_new_n32612__ = ys__n18448 & ys__n46667;
  assign new_new_n32613__ = ~ys__n18448 & ~ys__n46667;
  assign new_new_n32614__ = ~ys__n46604 & ~new_new_n32613__;
  assign new_new_n32615__ = ~new_new_n32612__ & new_new_n32614__;
  assign new_new_n32616__ = ys__n18451 & ys__n46668;
  assign new_new_n32617__ = ~ys__n18451 & ~ys__n46668;
  assign new_new_n32618__ = ~ys__n46606 & ~new_new_n32617__;
  assign new_new_n32619__ = ~new_new_n32616__ & new_new_n32618__;
  assign new_new_n32620__ = ~new_new_n32615__ & ~new_new_n32619__;
  assign new_new_n32621__ = ys__n18454 & ys__n46669;
  assign new_new_n32622__ = ~ys__n18454 & ~ys__n46669;
  assign new_new_n32623__ = ~ys__n46608 & ~new_new_n32622__;
  assign new_new_n32624__ = ~new_new_n32621__ & new_new_n32623__;
  assign new_new_n32625__ = ys__n18457 & ys__n46670;
  assign new_new_n32626__ = ~ys__n18457 & ~ys__n46670;
  assign new_new_n32627__ = ~ys__n46610 & ~new_new_n32626__;
  assign new_new_n32628__ = ~new_new_n32625__ & new_new_n32627__;
  assign new_new_n32629__ = ~new_new_n32624__ & ~new_new_n32628__;
  assign new_new_n32630__ = new_new_n32620__ & new_new_n32629__;
  assign new_new_n32631__ = ys__n42 & ys__n46764;
  assign new_new_n32632__ = ~ys__n42 & ~ys__n46764;
  assign new_new_n32633__ = ~ys__n46738 & ~new_new_n32632__;
  assign new_new_n32634__ = ~new_new_n32631__ & new_new_n32633__;
  assign new_new_n32635__ = ys__n40 & ys__n46765;
  assign new_new_n32636__ = ~ys__n40 & ~ys__n46765;
  assign new_new_n32637__ = ~ys__n46740 & ~new_new_n32636__;
  assign new_new_n32638__ = ~new_new_n32635__ & new_new_n32637__;
  assign new_new_n32639__ = ~new_new_n32634__ & ~new_new_n32638__;
  assign new_new_n32640__ = ys__n6133 & ys__n46766;
  assign new_new_n32641__ = ~ys__n6133 & ~ys__n46766;
  assign new_new_n32642__ = ~ys__n46742 & ~new_new_n32641__;
  assign new_new_n32643__ = ~new_new_n32640__ & new_new_n32642__;
  assign new_new_n32644__ = ys__n6134 & ys__n46767;
  assign new_new_n32645__ = ~ys__n6134 & ~ys__n46767;
  assign new_new_n32646__ = ~ys__n46744 & ~new_new_n32645__;
  assign new_new_n32647__ = ~new_new_n32644__ & new_new_n32646__;
  assign new_new_n32648__ = ~new_new_n32643__ & ~new_new_n32647__;
  assign new_new_n32649__ = new_new_n32639__ & new_new_n32648__;
  assign new_new_n32650__ = new_new_n32630__ & new_new_n32649__;
  assign new_new_n32651__ = new_new_n32611__ & new_new_n32650__;
  assign new_new_n32652__ = ys__n6113 & ys__n46745;
  assign new_new_n32653__ = ~ys__n6113 & ~ys__n46745;
  assign new_new_n32654__ = ~ys__n46700 & ~new_new_n32653__;
  assign new_new_n32655__ = ~new_new_n32652__ & new_new_n32654__;
  assign new_new_n32656__ = ~ys__n38 & ~ys__n46768;
  assign new_new_n32657__ = ys__n38 & ys__n46768;
  assign new_new_n32658__ = ~new_new_n32656__ & ~new_new_n32657__;
  assign new_new_n32659__ = ~new_new_n32347__ & ~new_new_n32658__;
  assign new_new_n32660__ = ~new_new_n32655__ & new_new_n32659__;
  assign new_new_n32661__ = ys__n172 & ys__n46746;
  assign new_new_n32662__ = ~ys__n172 & ~ys__n46746;
  assign new_new_n32663__ = ~ys__n46702 & ~new_new_n32662__;
  assign new_new_n32664__ = ~new_new_n32661__ & new_new_n32663__;
  assign new_new_n32665__ = ys__n338 & ys__n46747;
  assign new_new_n32666__ = ~ys__n338 & ~ys__n46747;
  assign new_new_n32667__ = ~ys__n46704 & ~new_new_n32666__;
  assign new_new_n32668__ = ~new_new_n32665__ & new_new_n32667__;
  assign new_new_n32669__ = ~new_new_n32664__ & ~new_new_n32668__;
  assign new_new_n32670__ = new_new_n32660__ & new_new_n32669__;
  assign new_new_n32671__ = ~ys__n28 & ~ys__n46773;
  assign new_new_n32672__ = ys__n28 & ys__n46773;
  assign new_new_n32673__ = ~new_new_n32671__ & ~new_new_n32672__;
  assign new_new_n32674__ = ~ys__n26 & ~ys__n46774;
  assign new_new_n32675__ = ys__n26 & ys__n46774;
  assign new_new_n32676__ = ~new_new_n32674__ & ~new_new_n32675__;
  assign new_new_n32677__ = ~new_new_n32673__ & ~new_new_n32676__;
  assign new_new_n32678__ = ~ys__n24 & ~ys__n46775;
  assign new_new_n32679__ = ys__n24 & ys__n46775;
  assign new_new_n32680__ = ~new_new_n32678__ & ~new_new_n32679__;
  assign new_new_n32681__ = ~ys__n27488 & new_new_n32348__;
  assign new_new_n32682__ = ~new_new_n32680__ & ~new_new_n32681__;
  assign new_new_n32683__ = new_new_n32677__ & new_new_n32682__;
  assign new_new_n32684__ = ~ys__n36 & ~ys__n46769;
  assign new_new_n32685__ = ys__n36 & ys__n46769;
  assign new_new_n32686__ = ~new_new_n32684__ & ~new_new_n32685__;
  assign new_new_n32687__ = ~ys__n34 & ~ys__n46770;
  assign new_new_n32688__ = ys__n34 & ys__n46770;
  assign new_new_n32689__ = ~new_new_n32687__ & ~new_new_n32688__;
  assign new_new_n32690__ = ~new_new_n32686__ & ~new_new_n32689__;
  assign new_new_n32691__ = ~ys__n32 & ~ys__n46771;
  assign new_new_n32692__ = ys__n32 & ys__n46771;
  assign new_new_n32693__ = ~new_new_n32691__ & ~new_new_n32692__;
  assign new_new_n32694__ = ~ys__n30 & ~ys__n46772;
  assign new_new_n32695__ = ys__n30 & ys__n46772;
  assign new_new_n32696__ = ~new_new_n32694__ & ~new_new_n32695__;
  assign new_new_n32697__ = ~new_new_n32693__ & ~new_new_n32696__;
  assign new_new_n32698__ = new_new_n32690__ & new_new_n32697__;
  assign new_new_n32699__ = new_new_n32683__ & new_new_n32698__;
  assign new_new_n32700__ = new_new_n32670__ & new_new_n32699__;
  assign new_new_n32701__ = ys__n340 & ys__n46752;
  assign new_new_n32702__ = ~ys__n340 & ~ys__n46752;
  assign new_new_n32703__ = ~ys__n46714 & ~new_new_n32702__;
  assign new_new_n32704__ = ~new_new_n32701__ & new_new_n32703__;
  assign new_new_n32705__ = ys__n46 & ys__n46753;
  assign new_new_n32706__ = ~ys__n46 & ~ys__n46753;
  assign new_new_n32707__ = ~ys__n46716 & ~new_new_n32706__;
  assign new_new_n32708__ = ~new_new_n32705__ & new_new_n32707__;
  assign new_new_n32709__ = ~new_new_n32704__ & ~new_new_n32708__;
  assign new_new_n32710__ = ys__n6118 & ys__n46754;
  assign new_new_n32711__ = ~ys__n6118 & ~ys__n46754;
  assign new_new_n32712__ = ~ys__n46718 & ~new_new_n32711__;
  assign new_new_n32713__ = ~new_new_n32710__ & new_new_n32712__;
  assign new_new_n32714__ = ys__n6119 & ys__n46755;
  assign new_new_n32715__ = ~ys__n6119 & ~ys__n46755;
  assign new_new_n32716__ = ~ys__n46720 & ~new_new_n32715__;
  assign new_new_n32717__ = ~new_new_n32714__ & new_new_n32716__;
  assign new_new_n32718__ = ~new_new_n32713__ & ~new_new_n32717__;
  assign new_new_n32719__ = new_new_n32709__ & new_new_n32718__;
  assign new_new_n32720__ = ys__n22 & ys__n46748;
  assign new_new_n32721__ = ~ys__n22 & ~ys__n46748;
  assign new_new_n32722__ = ~ys__n46706 & ~new_new_n32721__;
  assign new_new_n32723__ = ~new_new_n32720__ & new_new_n32722__;
  assign new_new_n32724__ = ys__n316 & ys__n46749;
  assign new_new_n32725__ = ~ys__n316 & ~ys__n46749;
  assign new_new_n32726__ = ~ys__n46708 & ~new_new_n32725__;
  assign new_new_n32727__ = ~new_new_n32724__ & new_new_n32726__;
  assign new_new_n32728__ = ~new_new_n32723__ & ~new_new_n32727__;
  assign new_new_n32729__ = ys__n6115 & ys__n46750;
  assign new_new_n32730__ = ~ys__n6115 & ~ys__n46750;
  assign new_new_n32731__ = ~ys__n46710 & ~new_new_n32730__;
  assign new_new_n32732__ = ~new_new_n32729__ & new_new_n32731__;
  assign new_new_n32733__ = ys__n44 & ys__n46751;
  assign new_new_n32734__ = ~ys__n44 & ~ys__n46751;
  assign new_new_n32735__ = ~ys__n46712 & ~new_new_n32734__;
  assign new_new_n32736__ = ~new_new_n32733__ & new_new_n32735__;
  assign new_new_n32737__ = ~new_new_n32732__ & ~new_new_n32736__;
  assign new_new_n32738__ = new_new_n32728__ & new_new_n32737__;
  assign new_new_n32739__ = new_new_n32719__ & new_new_n32738__;
  assign new_new_n32740__ = new_new_n32700__ & new_new_n32739__;
  assign new_new_n32741__ = new_new_n32651__ & new_new_n32740__;
  assign new_new_n32742__ = ys__n18520 & ys__n46691;
  assign new_new_n32743__ = ~ys__n18520 & ~ys__n46691;
  assign new_new_n32744__ = ~ys__n46652 & ~new_new_n32743__;
  assign new_new_n32745__ = ~new_new_n32742__ & new_new_n32744__;
  assign new_new_n32746__ = ys__n18523 & ys__n46692;
  assign new_new_n32747__ = ~ys__n18523 & ~ys__n46692;
  assign new_new_n32748__ = ~ys__n46654 & ~new_new_n32747__;
  assign new_new_n32749__ = ~new_new_n32746__ & new_new_n32748__;
  assign new_new_n32750__ = ~new_new_n32745__ & ~new_new_n32749__;
  assign new_new_n32751__ = ys__n18526 & ys__n46693;
  assign new_new_n32752__ = ~ys__n18526 & ~ys__n46693;
  assign new_new_n32753__ = ~ys__n46656 & ~new_new_n32752__;
  assign new_new_n32754__ = ~new_new_n32751__ & new_new_n32753__;
  assign new_new_n32755__ = ys__n18529 & ys__n46694;
  assign new_new_n32756__ = ~ys__n18529 & ~ys__n46694;
  assign new_new_n32757__ = ~ys__n46658 & ~new_new_n32756__;
  assign new_new_n32758__ = ~new_new_n32755__ & new_new_n32757__;
  assign new_new_n32759__ = ~new_new_n32754__ & ~new_new_n32758__;
  assign new_new_n32760__ = new_new_n32750__ & new_new_n32759__;
  assign new_new_n32761__ = ys__n18508 & ys__n46687;
  assign new_new_n32762__ = ~ys__n18508 & ~ys__n46687;
  assign new_new_n32763__ = ~ys__n46644 & ~new_new_n32762__;
  assign new_new_n32764__ = ~new_new_n32761__ & new_new_n32763__;
  assign new_new_n32765__ = ys__n18511 & ys__n46688;
  assign new_new_n32766__ = ~ys__n18511 & ~ys__n46688;
  assign new_new_n32767__ = ~ys__n46646 & ~new_new_n32766__;
  assign new_new_n32768__ = ~new_new_n32765__ & new_new_n32767__;
  assign new_new_n32769__ = ~new_new_n32764__ & ~new_new_n32768__;
  assign new_new_n32770__ = ys__n18514 & ys__n46689;
  assign new_new_n32771__ = ~ys__n18514 & ~ys__n46689;
  assign new_new_n32772__ = ~ys__n46648 & ~new_new_n32771__;
  assign new_new_n32773__ = ~new_new_n32770__ & new_new_n32772__;
  assign new_new_n32774__ = ys__n18517 & ys__n46690;
  assign new_new_n32775__ = ~ys__n18517 & ~ys__n46690;
  assign new_new_n32776__ = ~ys__n46650 & ~new_new_n32775__;
  assign new_new_n32777__ = ~new_new_n32774__ & new_new_n32776__;
  assign new_new_n32778__ = ~new_new_n32773__ & ~new_new_n32777__;
  assign new_new_n32779__ = new_new_n32769__ & new_new_n32778__;
  assign new_new_n32780__ = new_new_n32760__ & new_new_n32779__;
  assign new_new_n32781__ = ~ys__n18053 & new_new_n32450__;
  assign new_new_n32782__ = ~ys__n18057 & new_new_n32453__;
  assign new_new_n32783__ = ~ys__n18055 & new_new_n32455__;
  assign new_new_n32784__ = ~new_new_n32782__ & ~new_new_n32783__;
  assign new_new_n32785__ = ~new_new_n32781__ & new_new_n32784__;
  assign new_new_n32786__ = ys__n18532 & ys__n46695;
  assign new_new_n32787__ = ~ys__n18532 & ~ys__n46695;
  assign new_new_n32788__ = ~ys__n46660 & ~new_new_n32787__;
  assign new_new_n32789__ = ~new_new_n32786__ & new_new_n32788__;
  assign new_new_n32790__ = ys__n18535 & ys__n46696;
  assign new_new_n32791__ = ~ys__n18535 & ~ys__n46696;
  assign new_new_n32792__ = ~ys__n46662 & ~new_new_n32791__;
  assign new_new_n32793__ = ~new_new_n32790__ & new_new_n32792__;
  assign new_new_n32794__ = ~new_new_n32789__ & ~new_new_n32793__;
  assign new_new_n32795__ = ys__n18538 & ys__n46697;
  assign new_new_n32796__ = ~ys__n18538 & ~ys__n46697;
  assign new_new_n32797__ = ~ys__n46664 & ~new_new_n32796__;
  assign new_new_n32798__ = ~new_new_n32795__ & new_new_n32797__;
  assign new_new_n32799__ = ys__n18541 & ys__n46698;
  assign new_new_n32800__ = ~ys__n18541 & ~ys__n46698;
  assign new_new_n32801__ = ~ys__n46666 & ~new_new_n32800__;
  assign new_new_n32802__ = ~new_new_n32799__ & new_new_n32801__;
  assign new_new_n32803__ = ~new_new_n32798__ & ~new_new_n32802__;
  assign new_new_n32804__ = new_new_n32794__ & new_new_n32803__;
  assign new_new_n32805__ = new_new_n32785__ & new_new_n32804__;
  assign new_new_n32806__ = new_new_n32780__ & new_new_n32805__;
  assign new_new_n32807__ = ys__n18472 & ys__n46675;
  assign new_new_n32808__ = ~ys__n18472 & ~ys__n46675;
  assign new_new_n32809__ = ~ys__n46620 & ~new_new_n32808__;
  assign new_new_n32810__ = ~new_new_n32807__ & new_new_n32809__;
  assign new_new_n32811__ = ys__n18475 & ys__n46676;
  assign new_new_n32812__ = ~ys__n18475 & ~ys__n46676;
  assign new_new_n32813__ = ~ys__n46622 & ~new_new_n32812__;
  assign new_new_n32814__ = ~new_new_n32811__ & new_new_n32813__;
  assign new_new_n32815__ = ~new_new_n32810__ & ~new_new_n32814__;
  assign new_new_n32816__ = ys__n18478 & ys__n46677;
  assign new_new_n32817__ = ~ys__n18478 & ~ys__n46677;
  assign new_new_n32818__ = ~ys__n46624 & ~new_new_n32817__;
  assign new_new_n32819__ = ~new_new_n32816__ & new_new_n32818__;
  assign new_new_n32820__ = ys__n18481 & ys__n46678;
  assign new_new_n32821__ = ~ys__n18481 & ~ys__n46678;
  assign new_new_n32822__ = ~ys__n46626 & ~new_new_n32821__;
  assign new_new_n32823__ = ~new_new_n32820__ & new_new_n32822__;
  assign new_new_n32824__ = ~new_new_n32819__ & ~new_new_n32823__;
  assign new_new_n32825__ = new_new_n32815__ & new_new_n32824__;
  assign new_new_n32826__ = ys__n18460 & ys__n46671;
  assign new_new_n32827__ = ~ys__n18460 & ~ys__n46671;
  assign new_new_n32828__ = ~ys__n46612 & ~new_new_n32827__;
  assign new_new_n32829__ = ~new_new_n32826__ & new_new_n32828__;
  assign new_new_n32830__ = ys__n18463 & ys__n46672;
  assign new_new_n32831__ = ~ys__n18463 & ~ys__n46672;
  assign new_new_n32832__ = ~ys__n46614 & ~new_new_n32831__;
  assign new_new_n32833__ = ~new_new_n32830__ & new_new_n32832__;
  assign new_new_n32834__ = ~new_new_n32829__ & ~new_new_n32833__;
  assign new_new_n32835__ = ys__n18466 & ys__n46673;
  assign new_new_n32836__ = ~ys__n18466 & ~ys__n46673;
  assign new_new_n32837__ = ~ys__n46616 & ~new_new_n32836__;
  assign new_new_n32838__ = ~new_new_n32835__ & new_new_n32837__;
  assign new_new_n32839__ = ys__n18469 & ys__n46674;
  assign new_new_n32840__ = ~ys__n18469 & ~ys__n46674;
  assign new_new_n32841__ = ~ys__n46618 & ~new_new_n32840__;
  assign new_new_n32842__ = ~new_new_n32839__ & new_new_n32841__;
  assign new_new_n32843__ = ~new_new_n32838__ & ~new_new_n32842__;
  assign new_new_n32844__ = new_new_n32834__ & new_new_n32843__;
  assign new_new_n32845__ = new_new_n32825__ & new_new_n32844__;
  assign new_new_n32846__ = ys__n18496 & ys__n46683;
  assign new_new_n32847__ = ~ys__n18496 & ~ys__n46683;
  assign new_new_n32848__ = ~ys__n46636 & ~new_new_n32847__;
  assign new_new_n32849__ = ~new_new_n32846__ & new_new_n32848__;
  assign new_new_n32850__ = ys__n18499 & ys__n46684;
  assign new_new_n32851__ = ~ys__n18499 & ~ys__n46684;
  assign new_new_n32852__ = ~ys__n46638 & ~new_new_n32851__;
  assign new_new_n32853__ = ~new_new_n32850__ & new_new_n32852__;
  assign new_new_n32854__ = ~new_new_n32849__ & ~new_new_n32853__;
  assign new_new_n32855__ = ys__n18502 & ys__n46685;
  assign new_new_n32856__ = ~ys__n18502 & ~ys__n46685;
  assign new_new_n32857__ = ~ys__n46640 & ~new_new_n32856__;
  assign new_new_n32858__ = ~new_new_n32855__ & new_new_n32857__;
  assign new_new_n32859__ = ys__n18505 & ys__n46686;
  assign new_new_n32860__ = ~ys__n18505 & ~ys__n46686;
  assign new_new_n32861__ = ~ys__n46642 & ~new_new_n32860__;
  assign new_new_n32862__ = ~new_new_n32859__ & new_new_n32861__;
  assign new_new_n32863__ = ~new_new_n32858__ & ~new_new_n32862__;
  assign new_new_n32864__ = new_new_n32854__ & new_new_n32863__;
  assign new_new_n32865__ = ys__n18484 & ys__n46679;
  assign new_new_n32866__ = ~ys__n18484 & ~ys__n46679;
  assign new_new_n32867__ = ~ys__n46628 & ~new_new_n32866__;
  assign new_new_n32868__ = ~new_new_n32865__ & new_new_n32867__;
  assign new_new_n32869__ = ys__n18487 & ys__n46680;
  assign new_new_n32870__ = ~ys__n18487 & ~ys__n46680;
  assign new_new_n32871__ = ~ys__n46630 & ~new_new_n32870__;
  assign new_new_n32872__ = ~new_new_n32869__ & new_new_n32871__;
  assign new_new_n32873__ = ~new_new_n32868__ & ~new_new_n32872__;
  assign new_new_n32874__ = ys__n18490 & ys__n46681;
  assign new_new_n32875__ = ~ys__n18490 & ~ys__n46681;
  assign new_new_n32876__ = ~ys__n46632 & ~new_new_n32875__;
  assign new_new_n32877__ = ~new_new_n32874__ & new_new_n32876__;
  assign new_new_n32878__ = ys__n18493 & ys__n46682;
  assign new_new_n32879__ = ~ys__n18493 & ~ys__n46682;
  assign new_new_n32880__ = ~ys__n46634 & ~new_new_n32879__;
  assign new_new_n32881__ = ~new_new_n32878__ & new_new_n32880__;
  assign new_new_n32882__ = ~new_new_n32877__ & ~new_new_n32881__;
  assign new_new_n32883__ = new_new_n32873__ & new_new_n32882__;
  assign new_new_n32884__ = new_new_n32864__ & new_new_n32883__;
  assign new_new_n32885__ = new_new_n32845__ & new_new_n32884__;
  assign new_new_n32886__ = new_new_n32806__ & new_new_n32885__;
  assign new_new_n32887__ = new_new_n32741__ & new_new_n32886__;
  assign new_new_n32888__ = ~new_new_n32572__ & ~new_new_n32887__;
  assign new_new_n32889__ = ~ys__n27496 & ~new_new_n32572__;
  assign new_new_n32890__ = ~ys__n27496 & ~new_new_n32889__;
  assign new_new_n32891__ = ~ys__n27498 & ~new_new_n32890__;
  assign new_new_n32892__ = ~ys__n27498 & ~new_new_n32891__;
  assign new_new_n32893__ = new_new_n32887__ & ~new_new_n32892__;
  assign ys__n27493 = new_new_n32888__ | new_new_n32893__;
  assign new_new_n32895__ = ys__n26770 & ~new_new_n26767__;
  assign new_new_n32896__ = ys__n26770 & ~new_new_n26703__;
  assign new_new_n32897__ = ~new_new_n26719__ & ~new_new_n32896__;
  assign new_new_n32898__ = new_new_n26767__ & ~new_new_n32897__;
  assign new_new_n32899__ = ~new_new_n32895__ & ~new_new_n32898__;
  assign new_new_n32900__ = ys__n6126 & ys__n46584;
  assign new_new_n32901__ = ~ys__n6126 & ~ys__n46584;
  assign new_new_n32902__ = ~ys__n46554 & ~new_new_n32901__;
  assign new_new_n32903__ = ~new_new_n32900__ & new_new_n32902__;
  assign new_new_n32904__ = ys__n6127 & ys__n46585;
  assign new_new_n32905__ = ~ys__n6127 & ~ys__n46585;
  assign new_new_n32906__ = ~ys__n46556 & ~new_new_n32905__;
  assign new_new_n32907__ = ~new_new_n32904__ & new_new_n32906__;
  assign new_new_n32908__ = ~new_new_n32903__ & ~new_new_n32907__;
  assign new_new_n32909__ = ys__n6129 & ys__n46586;
  assign new_new_n32910__ = ~ys__n6129 & ~ys__n46586;
  assign new_new_n32911__ = ~ys__n46558 & ~new_new_n32910__;
  assign new_new_n32912__ = ~new_new_n32909__ & new_new_n32911__;
  assign new_new_n32913__ = ys__n6130 & ys__n46587;
  assign new_new_n32914__ = ~ys__n6130 & ~ys__n46587;
  assign new_new_n32915__ = ~ys__n46560 & ~new_new_n32914__;
  assign new_new_n32916__ = ~new_new_n32913__ & new_new_n32915__;
  assign new_new_n32917__ = ~new_new_n32912__ & ~new_new_n32916__;
  assign new_new_n32918__ = new_new_n32908__ & new_new_n32917__;
  assign new_new_n32919__ = ys__n6120 & ys__n46580;
  assign new_new_n32920__ = ~ys__n6120 & ~ys__n46580;
  assign new_new_n32921__ = ~ys__n46546 & ~new_new_n32920__;
  assign new_new_n32922__ = ~new_new_n32919__ & new_new_n32921__;
  assign new_new_n32923__ = ys__n6121 & ys__n46581;
  assign new_new_n32924__ = ~ys__n6121 & ~ys__n46581;
  assign new_new_n32925__ = ~ys__n46548 & ~new_new_n32924__;
  assign new_new_n32926__ = ~new_new_n32923__ & new_new_n32925__;
  assign new_new_n32927__ = ~new_new_n32922__ & ~new_new_n32926__;
  assign new_new_n32928__ = ys__n6123 & ys__n46582;
  assign new_new_n32929__ = ~ys__n6123 & ~ys__n46582;
  assign new_new_n32930__ = ~ys__n46550 & ~new_new_n32929__;
  assign new_new_n32931__ = ~new_new_n32928__ & new_new_n32930__;
  assign new_new_n32932__ = ys__n6124 & ys__n46583;
  assign new_new_n32933__ = ~ys__n6124 & ~ys__n46583;
  assign new_new_n32934__ = ~ys__n46552 & ~new_new_n32933__;
  assign new_new_n32935__ = ~new_new_n32932__ & new_new_n32934__;
  assign new_new_n32936__ = ~new_new_n32931__ & ~new_new_n32935__;
  assign new_new_n32937__ = new_new_n32927__ & new_new_n32936__;
  assign new_new_n32938__ = new_new_n32918__ & new_new_n32937__;
  assign new_new_n32939__ = ys__n18448 & ys__n46491;
  assign new_new_n32940__ = ~ys__n18448 & ~ys__n46491;
  assign new_new_n32941__ = ~ys__n46428 & ~new_new_n32940__;
  assign new_new_n32942__ = ~new_new_n32939__ & new_new_n32941__;
  assign new_new_n32943__ = ys__n18451 & ys__n46492;
  assign new_new_n32944__ = ~ys__n18451 & ~ys__n46492;
  assign new_new_n32945__ = ~ys__n46430 & ~new_new_n32944__;
  assign new_new_n32946__ = ~new_new_n32943__ & new_new_n32945__;
  assign new_new_n32947__ = ~new_new_n32942__ & ~new_new_n32946__;
  assign new_new_n32948__ = ys__n18454 & ys__n46493;
  assign new_new_n32949__ = ~ys__n18454 & ~ys__n46493;
  assign new_new_n32950__ = ~ys__n46432 & ~new_new_n32949__;
  assign new_new_n32951__ = ~new_new_n32948__ & new_new_n32950__;
  assign new_new_n32952__ = ys__n18457 & ys__n46494;
  assign new_new_n32953__ = ~ys__n18457 & ~ys__n46494;
  assign new_new_n32954__ = ~ys__n46434 & ~new_new_n32953__;
  assign new_new_n32955__ = ~new_new_n32952__ & new_new_n32954__;
  assign new_new_n32956__ = ~new_new_n32951__ & ~new_new_n32955__;
  assign new_new_n32957__ = new_new_n32947__ & new_new_n32956__;
  assign new_new_n32958__ = ys__n42 & ys__n46588;
  assign new_new_n32959__ = ~ys__n42 & ~ys__n46588;
  assign new_new_n32960__ = ~ys__n46562 & ~new_new_n32959__;
  assign new_new_n32961__ = ~new_new_n32958__ & new_new_n32960__;
  assign new_new_n32962__ = ys__n40 & ys__n46589;
  assign new_new_n32963__ = ~ys__n40 & ~ys__n46589;
  assign new_new_n32964__ = ~ys__n46564 & ~new_new_n32963__;
  assign new_new_n32965__ = ~new_new_n32962__ & new_new_n32964__;
  assign new_new_n32966__ = ~new_new_n32961__ & ~new_new_n32965__;
  assign new_new_n32967__ = ys__n6133 & ys__n46590;
  assign new_new_n32968__ = ~ys__n6133 & ~ys__n46590;
  assign new_new_n32969__ = ~ys__n46566 & ~new_new_n32968__;
  assign new_new_n32970__ = ~new_new_n32967__ & new_new_n32969__;
  assign new_new_n32971__ = ys__n6134 & ys__n46591;
  assign new_new_n32972__ = ~ys__n6134 & ~ys__n46591;
  assign new_new_n32973__ = ~ys__n46568 & ~new_new_n32972__;
  assign new_new_n32974__ = ~new_new_n32971__ & new_new_n32973__;
  assign new_new_n32975__ = ~new_new_n32970__ & ~new_new_n32974__;
  assign new_new_n32976__ = new_new_n32966__ & new_new_n32975__;
  assign new_new_n32977__ = new_new_n32957__ & new_new_n32976__;
  assign new_new_n32978__ = new_new_n32938__ & new_new_n32977__;
  assign new_new_n32979__ = ys__n6113 & ys__n46569;
  assign new_new_n32980__ = ~ys__n6113 & ~ys__n46569;
  assign new_new_n32981__ = ~ys__n46524 & ~new_new_n32980__;
  assign new_new_n32982__ = ~new_new_n32979__ & new_new_n32981__;
  assign new_new_n32983__ = ~ys__n38 & ~ys__n46592;
  assign new_new_n32984__ = ys__n38 & ys__n46592;
  assign new_new_n32985__ = ~new_new_n32983__ & ~new_new_n32984__;
  assign new_new_n32986__ = ~new_new_n32347__ & ~new_new_n32985__;
  assign new_new_n32987__ = ~new_new_n32982__ & new_new_n32986__;
  assign new_new_n32988__ = ys__n172 & ys__n46570;
  assign new_new_n32989__ = ~ys__n172 & ~ys__n46570;
  assign new_new_n32990__ = ~ys__n46526 & ~new_new_n32989__;
  assign new_new_n32991__ = ~new_new_n32988__ & new_new_n32990__;
  assign new_new_n32992__ = ys__n338 & ys__n46571;
  assign new_new_n32993__ = ~ys__n338 & ~ys__n46571;
  assign new_new_n32994__ = ~ys__n46528 & ~new_new_n32993__;
  assign new_new_n32995__ = ~new_new_n32992__ & new_new_n32994__;
  assign new_new_n32996__ = ~new_new_n32991__ & ~new_new_n32995__;
  assign new_new_n32997__ = new_new_n32987__ & new_new_n32996__;
  assign new_new_n32998__ = ~ys__n28 & ~ys__n46597;
  assign new_new_n32999__ = ys__n28 & ys__n46597;
  assign new_new_n33000__ = ~new_new_n32998__ & ~new_new_n32999__;
  assign new_new_n33001__ = ~ys__n26 & ~ys__n46598;
  assign new_new_n33002__ = ys__n26 & ys__n46598;
  assign new_new_n33003__ = ~new_new_n33001__ & ~new_new_n33002__;
  assign new_new_n33004__ = ~new_new_n33000__ & ~new_new_n33003__;
  assign new_new_n33005__ = ~ys__n24 & ~ys__n46599;
  assign new_new_n33006__ = ys__n24 & ys__n46599;
  assign new_new_n33007__ = ~new_new_n33005__ & ~new_new_n33006__;
  assign new_new_n33008__ = ~ys__n27499 & new_new_n32348__;
  assign new_new_n33009__ = ~new_new_n33007__ & ~new_new_n33008__;
  assign new_new_n33010__ = new_new_n33004__ & new_new_n33009__;
  assign new_new_n33011__ = ~ys__n36 & ~ys__n46593;
  assign new_new_n33012__ = ys__n36 & ys__n46593;
  assign new_new_n33013__ = ~new_new_n33011__ & ~new_new_n33012__;
  assign new_new_n33014__ = ~ys__n34 & ~ys__n46594;
  assign new_new_n33015__ = ys__n34 & ys__n46594;
  assign new_new_n33016__ = ~new_new_n33014__ & ~new_new_n33015__;
  assign new_new_n33017__ = ~new_new_n33013__ & ~new_new_n33016__;
  assign new_new_n33018__ = ~ys__n32 & ~ys__n46595;
  assign new_new_n33019__ = ys__n32 & ys__n46595;
  assign new_new_n33020__ = ~new_new_n33018__ & ~new_new_n33019__;
  assign new_new_n33021__ = ~ys__n30 & ~ys__n46596;
  assign new_new_n33022__ = ys__n30 & ys__n46596;
  assign new_new_n33023__ = ~new_new_n33021__ & ~new_new_n33022__;
  assign new_new_n33024__ = ~new_new_n33020__ & ~new_new_n33023__;
  assign new_new_n33025__ = new_new_n33017__ & new_new_n33024__;
  assign new_new_n33026__ = new_new_n33010__ & new_new_n33025__;
  assign new_new_n33027__ = new_new_n32997__ & new_new_n33026__;
  assign new_new_n33028__ = ys__n340 & ys__n46576;
  assign new_new_n33029__ = ~ys__n340 & ~ys__n46576;
  assign new_new_n33030__ = ~ys__n46538 & ~new_new_n33029__;
  assign new_new_n33031__ = ~new_new_n33028__ & new_new_n33030__;
  assign new_new_n33032__ = ys__n46 & ys__n46577;
  assign new_new_n33033__ = ~ys__n46 & ~ys__n46577;
  assign new_new_n33034__ = ~ys__n46540 & ~new_new_n33033__;
  assign new_new_n33035__ = ~new_new_n33032__ & new_new_n33034__;
  assign new_new_n33036__ = ~new_new_n33031__ & ~new_new_n33035__;
  assign new_new_n33037__ = ys__n6118 & ys__n46578;
  assign new_new_n33038__ = ~ys__n6118 & ~ys__n46578;
  assign new_new_n33039__ = ~ys__n46542 & ~new_new_n33038__;
  assign new_new_n33040__ = ~new_new_n33037__ & new_new_n33039__;
  assign new_new_n33041__ = ys__n6119 & ys__n46579;
  assign new_new_n33042__ = ~ys__n6119 & ~ys__n46579;
  assign new_new_n33043__ = ~ys__n46544 & ~new_new_n33042__;
  assign new_new_n33044__ = ~new_new_n33041__ & new_new_n33043__;
  assign new_new_n33045__ = ~new_new_n33040__ & ~new_new_n33044__;
  assign new_new_n33046__ = new_new_n33036__ & new_new_n33045__;
  assign new_new_n33047__ = ys__n22 & ys__n46572;
  assign new_new_n33048__ = ~ys__n22 & ~ys__n46572;
  assign new_new_n33049__ = ~ys__n46530 & ~new_new_n33048__;
  assign new_new_n33050__ = ~new_new_n33047__ & new_new_n33049__;
  assign new_new_n33051__ = ys__n316 & ys__n46573;
  assign new_new_n33052__ = ~ys__n316 & ~ys__n46573;
  assign new_new_n33053__ = ~ys__n46532 & ~new_new_n33052__;
  assign new_new_n33054__ = ~new_new_n33051__ & new_new_n33053__;
  assign new_new_n33055__ = ~new_new_n33050__ & ~new_new_n33054__;
  assign new_new_n33056__ = ys__n6115 & ys__n46574;
  assign new_new_n33057__ = ~ys__n6115 & ~ys__n46574;
  assign new_new_n33058__ = ~ys__n46534 & ~new_new_n33057__;
  assign new_new_n33059__ = ~new_new_n33056__ & new_new_n33058__;
  assign new_new_n33060__ = ys__n44 & ys__n46575;
  assign new_new_n33061__ = ~ys__n44 & ~ys__n46575;
  assign new_new_n33062__ = ~ys__n46536 & ~new_new_n33061__;
  assign new_new_n33063__ = ~new_new_n33060__ & new_new_n33062__;
  assign new_new_n33064__ = ~new_new_n33059__ & ~new_new_n33063__;
  assign new_new_n33065__ = new_new_n33055__ & new_new_n33064__;
  assign new_new_n33066__ = new_new_n33046__ & new_new_n33065__;
  assign new_new_n33067__ = new_new_n33027__ & new_new_n33066__;
  assign new_new_n33068__ = new_new_n32978__ & new_new_n33067__;
  assign new_new_n33069__ = ys__n18520 & ys__n46515;
  assign new_new_n33070__ = ~ys__n18520 & ~ys__n46515;
  assign new_new_n33071__ = ~ys__n46476 & ~new_new_n33070__;
  assign new_new_n33072__ = ~new_new_n33069__ & new_new_n33071__;
  assign new_new_n33073__ = ys__n18523 & ys__n46516;
  assign new_new_n33074__ = ~ys__n18523 & ~ys__n46516;
  assign new_new_n33075__ = ~ys__n46478 & ~new_new_n33074__;
  assign new_new_n33076__ = ~new_new_n33073__ & new_new_n33075__;
  assign new_new_n33077__ = ~new_new_n33072__ & ~new_new_n33076__;
  assign new_new_n33078__ = ys__n18526 & ys__n46517;
  assign new_new_n33079__ = ~ys__n18526 & ~ys__n46517;
  assign new_new_n33080__ = ~ys__n46480 & ~new_new_n33079__;
  assign new_new_n33081__ = ~new_new_n33078__ & new_new_n33080__;
  assign new_new_n33082__ = ys__n18529 & ys__n46518;
  assign new_new_n33083__ = ~ys__n18529 & ~ys__n46518;
  assign new_new_n33084__ = ~ys__n46482 & ~new_new_n33083__;
  assign new_new_n33085__ = ~new_new_n33082__ & new_new_n33084__;
  assign new_new_n33086__ = ~new_new_n33081__ & ~new_new_n33085__;
  assign new_new_n33087__ = new_new_n33077__ & new_new_n33086__;
  assign new_new_n33088__ = ys__n18508 & ys__n46511;
  assign new_new_n33089__ = ~ys__n18508 & ~ys__n46511;
  assign new_new_n33090__ = ~ys__n46468 & ~new_new_n33089__;
  assign new_new_n33091__ = ~new_new_n33088__ & new_new_n33090__;
  assign new_new_n33092__ = ys__n18511 & ys__n46512;
  assign new_new_n33093__ = ~ys__n18511 & ~ys__n46512;
  assign new_new_n33094__ = ~ys__n46470 & ~new_new_n33093__;
  assign new_new_n33095__ = ~new_new_n33092__ & new_new_n33094__;
  assign new_new_n33096__ = ~new_new_n33091__ & ~new_new_n33095__;
  assign new_new_n33097__ = ys__n18514 & ys__n46513;
  assign new_new_n33098__ = ~ys__n18514 & ~ys__n46513;
  assign new_new_n33099__ = ~ys__n46472 & ~new_new_n33098__;
  assign new_new_n33100__ = ~new_new_n33097__ & new_new_n33099__;
  assign new_new_n33101__ = ys__n18517 & ys__n46514;
  assign new_new_n33102__ = ~ys__n18517 & ~ys__n46514;
  assign new_new_n33103__ = ~ys__n46474 & ~new_new_n33102__;
  assign new_new_n33104__ = ~new_new_n33101__ & new_new_n33103__;
  assign new_new_n33105__ = ~new_new_n33100__ & ~new_new_n33104__;
  assign new_new_n33106__ = new_new_n33096__ & new_new_n33105__;
  assign new_new_n33107__ = new_new_n33087__ & new_new_n33106__;
  assign new_new_n33108__ = ~ys__n18047 & new_new_n32450__;
  assign new_new_n33109__ = ~ys__n18051 & new_new_n32453__;
  assign new_new_n33110__ = ~ys__n18049 & new_new_n32455__;
  assign new_new_n33111__ = ~new_new_n33109__ & ~new_new_n33110__;
  assign new_new_n33112__ = ~new_new_n33108__ & new_new_n33111__;
  assign new_new_n33113__ = ys__n18532 & ys__n46519;
  assign new_new_n33114__ = ~ys__n18532 & ~ys__n46519;
  assign new_new_n33115__ = ~ys__n46484 & ~new_new_n33114__;
  assign new_new_n33116__ = ~new_new_n33113__ & new_new_n33115__;
  assign new_new_n33117__ = ys__n18535 & ys__n46520;
  assign new_new_n33118__ = ~ys__n18535 & ~ys__n46520;
  assign new_new_n33119__ = ~ys__n46486 & ~new_new_n33118__;
  assign new_new_n33120__ = ~new_new_n33117__ & new_new_n33119__;
  assign new_new_n33121__ = ~new_new_n33116__ & ~new_new_n33120__;
  assign new_new_n33122__ = ys__n18538 & ys__n46521;
  assign new_new_n33123__ = ~ys__n18538 & ~ys__n46521;
  assign new_new_n33124__ = ~ys__n46488 & ~new_new_n33123__;
  assign new_new_n33125__ = ~new_new_n33122__ & new_new_n33124__;
  assign new_new_n33126__ = ys__n18541 & ys__n46522;
  assign new_new_n33127__ = ~ys__n18541 & ~ys__n46522;
  assign new_new_n33128__ = ~ys__n46490 & ~new_new_n33127__;
  assign new_new_n33129__ = ~new_new_n33126__ & new_new_n33128__;
  assign new_new_n33130__ = ~new_new_n33125__ & ~new_new_n33129__;
  assign new_new_n33131__ = new_new_n33121__ & new_new_n33130__;
  assign new_new_n33132__ = new_new_n33112__ & new_new_n33131__;
  assign new_new_n33133__ = new_new_n33107__ & new_new_n33132__;
  assign new_new_n33134__ = ys__n18472 & ys__n46499;
  assign new_new_n33135__ = ~ys__n18472 & ~ys__n46499;
  assign new_new_n33136__ = ~ys__n46444 & ~new_new_n33135__;
  assign new_new_n33137__ = ~new_new_n33134__ & new_new_n33136__;
  assign new_new_n33138__ = ys__n18475 & ys__n46500;
  assign new_new_n33139__ = ~ys__n18475 & ~ys__n46500;
  assign new_new_n33140__ = ~ys__n46446 & ~new_new_n33139__;
  assign new_new_n33141__ = ~new_new_n33138__ & new_new_n33140__;
  assign new_new_n33142__ = ~new_new_n33137__ & ~new_new_n33141__;
  assign new_new_n33143__ = ys__n18478 & ys__n46501;
  assign new_new_n33144__ = ~ys__n18478 & ~ys__n46501;
  assign new_new_n33145__ = ~ys__n46448 & ~new_new_n33144__;
  assign new_new_n33146__ = ~new_new_n33143__ & new_new_n33145__;
  assign new_new_n33147__ = ys__n18481 & ys__n46502;
  assign new_new_n33148__ = ~ys__n18481 & ~ys__n46502;
  assign new_new_n33149__ = ~ys__n46450 & ~new_new_n33148__;
  assign new_new_n33150__ = ~new_new_n33147__ & new_new_n33149__;
  assign new_new_n33151__ = ~new_new_n33146__ & ~new_new_n33150__;
  assign new_new_n33152__ = new_new_n33142__ & new_new_n33151__;
  assign new_new_n33153__ = ys__n18460 & ys__n46495;
  assign new_new_n33154__ = ~ys__n18460 & ~ys__n46495;
  assign new_new_n33155__ = ~ys__n46436 & ~new_new_n33154__;
  assign new_new_n33156__ = ~new_new_n33153__ & new_new_n33155__;
  assign new_new_n33157__ = ys__n18463 & ys__n46496;
  assign new_new_n33158__ = ~ys__n18463 & ~ys__n46496;
  assign new_new_n33159__ = ~ys__n46438 & ~new_new_n33158__;
  assign new_new_n33160__ = ~new_new_n33157__ & new_new_n33159__;
  assign new_new_n33161__ = ~new_new_n33156__ & ~new_new_n33160__;
  assign new_new_n33162__ = ys__n18466 & ys__n46497;
  assign new_new_n33163__ = ~ys__n18466 & ~ys__n46497;
  assign new_new_n33164__ = ~ys__n46440 & ~new_new_n33163__;
  assign new_new_n33165__ = ~new_new_n33162__ & new_new_n33164__;
  assign new_new_n33166__ = ys__n18469 & ys__n46498;
  assign new_new_n33167__ = ~ys__n18469 & ~ys__n46498;
  assign new_new_n33168__ = ~ys__n46442 & ~new_new_n33167__;
  assign new_new_n33169__ = ~new_new_n33166__ & new_new_n33168__;
  assign new_new_n33170__ = ~new_new_n33165__ & ~new_new_n33169__;
  assign new_new_n33171__ = new_new_n33161__ & new_new_n33170__;
  assign new_new_n33172__ = new_new_n33152__ & new_new_n33171__;
  assign new_new_n33173__ = ys__n18496 & ys__n46507;
  assign new_new_n33174__ = ~ys__n18496 & ~ys__n46507;
  assign new_new_n33175__ = ~ys__n46460 & ~new_new_n33174__;
  assign new_new_n33176__ = ~new_new_n33173__ & new_new_n33175__;
  assign new_new_n33177__ = ys__n18499 & ys__n46508;
  assign new_new_n33178__ = ~ys__n18499 & ~ys__n46508;
  assign new_new_n33179__ = ~ys__n46462 & ~new_new_n33178__;
  assign new_new_n33180__ = ~new_new_n33177__ & new_new_n33179__;
  assign new_new_n33181__ = ~new_new_n33176__ & ~new_new_n33180__;
  assign new_new_n33182__ = ys__n18502 & ys__n46509;
  assign new_new_n33183__ = ~ys__n18502 & ~ys__n46509;
  assign new_new_n33184__ = ~ys__n46464 & ~new_new_n33183__;
  assign new_new_n33185__ = ~new_new_n33182__ & new_new_n33184__;
  assign new_new_n33186__ = ys__n18505 & ys__n46510;
  assign new_new_n33187__ = ~ys__n18505 & ~ys__n46510;
  assign new_new_n33188__ = ~ys__n46466 & ~new_new_n33187__;
  assign new_new_n33189__ = ~new_new_n33186__ & new_new_n33188__;
  assign new_new_n33190__ = ~new_new_n33185__ & ~new_new_n33189__;
  assign new_new_n33191__ = new_new_n33181__ & new_new_n33190__;
  assign new_new_n33192__ = ys__n18484 & ys__n46503;
  assign new_new_n33193__ = ~ys__n18484 & ~ys__n46503;
  assign new_new_n33194__ = ~ys__n46452 & ~new_new_n33193__;
  assign new_new_n33195__ = ~new_new_n33192__ & new_new_n33194__;
  assign new_new_n33196__ = ys__n18487 & ys__n46504;
  assign new_new_n33197__ = ~ys__n18487 & ~ys__n46504;
  assign new_new_n33198__ = ~ys__n46454 & ~new_new_n33197__;
  assign new_new_n33199__ = ~new_new_n33196__ & new_new_n33198__;
  assign new_new_n33200__ = ~new_new_n33195__ & ~new_new_n33199__;
  assign new_new_n33201__ = ys__n18490 & ys__n46505;
  assign new_new_n33202__ = ~ys__n18490 & ~ys__n46505;
  assign new_new_n33203__ = ~ys__n46456 & ~new_new_n33202__;
  assign new_new_n33204__ = ~new_new_n33201__ & new_new_n33203__;
  assign new_new_n33205__ = ys__n18493 & ys__n46506;
  assign new_new_n33206__ = ~ys__n18493 & ~ys__n46506;
  assign new_new_n33207__ = ~ys__n46458 & ~new_new_n33206__;
  assign new_new_n33208__ = ~new_new_n33205__ & new_new_n33207__;
  assign new_new_n33209__ = ~new_new_n33204__ & ~new_new_n33208__;
  assign new_new_n33210__ = new_new_n33200__ & new_new_n33209__;
  assign new_new_n33211__ = new_new_n33191__ & new_new_n33210__;
  assign new_new_n33212__ = new_new_n33172__ & new_new_n33211__;
  assign new_new_n33213__ = new_new_n33133__ & new_new_n33212__;
  assign new_new_n33214__ = new_new_n33068__ & new_new_n33213__;
  assign new_new_n33215__ = ~new_new_n32899__ & ~new_new_n33214__;
  assign new_new_n33216__ = ~ys__n27507 & ~new_new_n32899__;
  assign new_new_n33217__ = ~ys__n27507 & ~new_new_n33216__;
  assign new_new_n33218__ = ~ys__n27509 & ~new_new_n33217__;
  assign new_new_n33219__ = ~ys__n27509 & ~new_new_n33218__;
  assign new_new_n33220__ = new_new_n33214__ & ~new_new_n33219__;
  assign ys__n27504 = new_new_n33215__ | new_new_n33220__;
  assign new_new_n33222__ = ys__n27481 & new_new_n32560__;
  assign new_new_n33223__ = ~new_new_n32887__ & new_new_n33222__;
  assign new_new_n33224__ = ~ys__n27496 & new_new_n33222__;
  assign new_new_n33225__ = ~ys__n27496 & ~new_new_n33224__;
  assign new_new_n33226__ = new_new_n32887__ & ~new_new_n33225__;
  assign new_new_n33227__ = ~new_new_n33223__ & ~new_new_n33226__;
  assign new_new_n33228__ = ~new_new_n33214__ & ~new_new_n33227__;
  assign new_new_n33229__ = ~ys__n27507 & ~new_new_n33227__;
  assign new_new_n33230__ = ~ys__n27507 & ~new_new_n33229__;
  assign new_new_n33231__ = new_new_n33214__ & ~new_new_n33230__;
  assign new_new_n33232__ = ~new_new_n33228__ & ~new_new_n33231__;
  assign new_new_n33233__ = ys__n6126 & ys__n46408;
  assign new_new_n33234__ = ~ys__n6126 & ~ys__n46408;
  assign new_new_n33235__ = ~ys__n46378 & ~new_new_n33234__;
  assign new_new_n33236__ = ~new_new_n33233__ & new_new_n33235__;
  assign new_new_n33237__ = ys__n6127 & ys__n46409;
  assign new_new_n33238__ = ~ys__n6127 & ~ys__n46409;
  assign new_new_n33239__ = ~ys__n46380 & ~new_new_n33238__;
  assign new_new_n33240__ = ~new_new_n33237__ & new_new_n33239__;
  assign new_new_n33241__ = ~new_new_n33236__ & ~new_new_n33240__;
  assign new_new_n33242__ = ys__n6129 & ys__n46410;
  assign new_new_n33243__ = ~ys__n6129 & ~ys__n46410;
  assign new_new_n33244__ = ~ys__n46382 & ~new_new_n33243__;
  assign new_new_n33245__ = ~new_new_n33242__ & new_new_n33244__;
  assign new_new_n33246__ = ys__n6130 & ys__n46411;
  assign new_new_n33247__ = ~ys__n6130 & ~ys__n46411;
  assign new_new_n33248__ = ~ys__n46384 & ~new_new_n33247__;
  assign new_new_n33249__ = ~new_new_n33246__ & new_new_n33248__;
  assign new_new_n33250__ = ~new_new_n33245__ & ~new_new_n33249__;
  assign new_new_n33251__ = new_new_n33241__ & new_new_n33250__;
  assign new_new_n33252__ = ys__n6120 & ys__n46404;
  assign new_new_n33253__ = ~ys__n6120 & ~ys__n46404;
  assign new_new_n33254__ = ~ys__n46370 & ~new_new_n33253__;
  assign new_new_n33255__ = ~new_new_n33252__ & new_new_n33254__;
  assign new_new_n33256__ = ys__n6121 & ys__n46405;
  assign new_new_n33257__ = ~ys__n6121 & ~ys__n46405;
  assign new_new_n33258__ = ~ys__n46372 & ~new_new_n33257__;
  assign new_new_n33259__ = ~new_new_n33256__ & new_new_n33258__;
  assign new_new_n33260__ = ~new_new_n33255__ & ~new_new_n33259__;
  assign new_new_n33261__ = ys__n6123 & ys__n46406;
  assign new_new_n33262__ = ~ys__n6123 & ~ys__n46406;
  assign new_new_n33263__ = ~ys__n46374 & ~new_new_n33262__;
  assign new_new_n33264__ = ~new_new_n33261__ & new_new_n33263__;
  assign new_new_n33265__ = ys__n6124 & ys__n46407;
  assign new_new_n33266__ = ~ys__n6124 & ~ys__n46407;
  assign new_new_n33267__ = ~ys__n46376 & ~new_new_n33266__;
  assign new_new_n33268__ = ~new_new_n33265__ & new_new_n33267__;
  assign new_new_n33269__ = ~new_new_n33264__ & ~new_new_n33268__;
  assign new_new_n33270__ = new_new_n33260__ & new_new_n33269__;
  assign new_new_n33271__ = new_new_n33251__ & new_new_n33270__;
  assign new_new_n33272__ = ys__n18448 & ys__n46315;
  assign new_new_n33273__ = ~ys__n18448 & ~ys__n46315;
  assign new_new_n33274__ = ~ys__n46252 & ~new_new_n33273__;
  assign new_new_n33275__ = ~new_new_n33272__ & new_new_n33274__;
  assign new_new_n33276__ = ys__n18451 & ys__n46316;
  assign new_new_n33277__ = ~ys__n18451 & ~ys__n46316;
  assign new_new_n33278__ = ~ys__n46254 & ~new_new_n33277__;
  assign new_new_n33279__ = ~new_new_n33276__ & new_new_n33278__;
  assign new_new_n33280__ = ~new_new_n33275__ & ~new_new_n33279__;
  assign new_new_n33281__ = ys__n18454 & ys__n46317;
  assign new_new_n33282__ = ~ys__n18454 & ~ys__n46317;
  assign new_new_n33283__ = ~ys__n46256 & ~new_new_n33282__;
  assign new_new_n33284__ = ~new_new_n33281__ & new_new_n33283__;
  assign new_new_n33285__ = ys__n18457 & ys__n46318;
  assign new_new_n33286__ = ~ys__n18457 & ~ys__n46318;
  assign new_new_n33287__ = ~ys__n46258 & ~new_new_n33286__;
  assign new_new_n33288__ = ~new_new_n33285__ & new_new_n33287__;
  assign new_new_n33289__ = ~new_new_n33284__ & ~new_new_n33288__;
  assign new_new_n33290__ = new_new_n33280__ & new_new_n33289__;
  assign new_new_n33291__ = ys__n42 & ys__n46412;
  assign new_new_n33292__ = ~ys__n42 & ~ys__n46412;
  assign new_new_n33293__ = ~ys__n46386 & ~new_new_n33292__;
  assign new_new_n33294__ = ~new_new_n33291__ & new_new_n33293__;
  assign new_new_n33295__ = ys__n40 & ys__n46413;
  assign new_new_n33296__ = ~ys__n40 & ~ys__n46413;
  assign new_new_n33297__ = ~ys__n46388 & ~new_new_n33296__;
  assign new_new_n33298__ = ~new_new_n33295__ & new_new_n33297__;
  assign new_new_n33299__ = ~new_new_n33294__ & ~new_new_n33298__;
  assign new_new_n33300__ = ys__n6133 & ys__n46414;
  assign new_new_n33301__ = ~ys__n6133 & ~ys__n46414;
  assign new_new_n33302__ = ~ys__n46390 & ~new_new_n33301__;
  assign new_new_n33303__ = ~new_new_n33300__ & new_new_n33302__;
  assign new_new_n33304__ = ys__n6134 & ys__n46415;
  assign new_new_n33305__ = ~ys__n6134 & ~ys__n46415;
  assign new_new_n33306__ = ~ys__n46392 & ~new_new_n33305__;
  assign new_new_n33307__ = ~new_new_n33304__ & new_new_n33306__;
  assign new_new_n33308__ = ~new_new_n33303__ & ~new_new_n33307__;
  assign new_new_n33309__ = new_new_n33299__ & new_new_n33308__;
  assign new_new_n33310__ = new_new_n33290__ & new_new_n33309__;
  assign new_new_n33311__ = new_new_n33271__ & new_new_n33310__;
  assign new_new_n33312__ = ys__n6113 & ys__n46393;
  assign new_new_n33313__ = ~ys__n6113 & ~ys__n46393;
  assign new_new_n33314__ = ~ys__n46348 & ~new_new_n33313__;
  assign new_new_n33315__ = ~new_new_n33312__ & new_new_n33314__;
  assign new_new_n33316__ = ~ys__n38 & ~ys__n46416;
  assign new_new_n33317__ = ys__n38 & ys__n46416;
  assign new_new_n33318__ = ~new_new_n33316__ & ~new_new_n33317__;
  assign new_new_n33319__ = ~new_new_n32347__ & ~new_new_n33318__;
  assign new_new_n33320__ = ~new_new_n33315__ & new_new_n33319__;
  assign new_new_n33321__ = ys__n172 & ys__n46394;
  assign new_new_n33322__ = ~ys__n172 & ~ys__n46394;
  assign new_new_n33323__ = ~ys__n46350 & ~new_new_n33322__;
  assign new_new_n33324__ = ~new_new_n33321__ & new_new_n33323__;
  assign new_new_n33325__ = ys__n338 & ys__n46395;
  assign new_new_n33326__ = ~ys__n338 & ~ys__n46395;
  assign new_new_n33327__ = ~ys__n46352 & ~new_new_n33326__;
  assign new_new_n33328__ = ~new_new_n33325__ & new_new_n33327__;
  assign new_new_n33329__ = ~new_new_n33324__ & ~new_new_n33328__;
  assign new_new_n33330__ = new_new_n33320__ & new_new_n33329__;
  assign new_new_n33331__ = ~ys__n28 & ~ys__n46421;
  assign new_new_n33332__ = ys__n28 & ys__n46421;
  assign new_new_n33333__ = ~new_new_n33331__ & ~new_new_n33332__;
  assign new_new_n33334__ = ~ys__n26 & ~ys__n46422;
  assign new_new_n33335__ = ys__n26 & ys__n46422;
  assign new_new_n33336__ = ~new_new_n33334__ & ~new_new_n33335__;
  assign new_new_n33337__ = ~new_new_n33333__ & ~new_new_n33336__;
  assign new_new_n33338__ = ~ys__n24 & ~ys__n46423;
  assign new_new_n33339__ = ys__n24 & ys__n46423;
  assign new_new_n33340__ = ~new_new_n33338__ & ~new_new_n33339__;
  assign new_new_n33341__ = ~ys__n27510 & new_new_n32348__;
  assign new_new_n33342__ = ~new_new_n33340__ & ~new_new_n33341__;
  assign new_new_n33343__ = new_new_n33337__ & new_new_n33342__;
  assign new_new_n33344__ = ~ys__n36 & ~ys__n46417;
  assign new_new_n33345__ = ys__n36 & ys__n46417;
  assign new_new_n33346__ = ~new_new_n33344__ & ~new_new_n33345__;
  assign new_new_n33347__ = ~ys__n34 & ~ys__n46418;
  assign new_new_n33348__ = ys__n34 & ys__n46418;
  assign new_new_n33349__ = ~new_new_n33347__ & ~new_new_n33348__;
  assign new_new_n33350__ = ~new_new_n33346__ & ~new_new_n33349__;
  assign new_new_n33351__ = ~ys__n32 & ~ys__n46419;
  assign new_new_n33352__ = ys__n32 & ys__n46419;
  assign new_new_n33353__ = ~new_new_n33351__ & ~new_new_n33352__;
  assign new_new_n33354__ = ~ys__n30 & ~ys__n46420;
  assign new_new_n33355__ = ys__n30 & ys__n46420;
  assign new_new_n33356__ = ~new_new_n33354__ & ~new_new_n33355__;
  assign new_new_n33357__ = ~new_new_n33353__ & ~new_new_n33356__;
  assign new_new_n33358__ = new_new_n33350__ & new_new_n33357__;
  assign new_new_n33359__ = new_new_n33343__ & new_new_n33358__;
  assign new_new_n33360__ = new_new_n33330__ & new_new_n33359__;
  assign new_new_n33361__ = ys__n340 & ys__n46400;
  assign new_new_n33362__ = ~ys__n340 & ~ys__n46400;
  assign new_new_n33363__ = ~ys__n46362 & ~new_new_n33362__;
  assign new_new_n33364__ = ~new_new_n33361__ & new_new_n33363__;
  assign new_new_n33365__ = ys__n46 & ys__n46401;
  assign new_new_n33366__ = ~ys__n46 & ~ys__n46401;
  assign new_new_n33367__ = ~ys__n46364 & ~new_new_n33366__;
  assign new_new_n33368__ = ~new_new_n33365__ & new_new_n33367__;
  assign new_new_n33369__ = ~new_new_n33364__ & ~new_new_n33368__;
  assign new_new_n33370__ = ys__n6118 & ys__n46402;
  assign new_new_n33371__ = ~ys__n6118 & ~ys__n46402;
  assign new_new_n33372__ = ~ys__n46366 & ~new_new_n33371__;
  assign new_new_n33373__ = ~new_new_n33370__ & new_new_n33372__;
  assign new_new_n33374__ = ys__n6119 & ys__n46403;
  assign new_new_n33375__ = ~ys__n6119 & ~ys__n46403;
  assign new_new_n33376__ = ~ys__n46368 & ~new_new_n33375__;
  assign new_new_n33377__ = ~new_new_n33374__ & new_new_n33376__;
  assign new_new_n33378__ = ~new_new_n33373__ & ~new_new_n33377__;
  assign new_new_n33379__ = new_new_n33369__ & new_new_n33378__;
  assign new_new_n33380__ = ys__n22 & ys__n46396;
  assign new_new_n33381__ = ~ys__n22 & ~ys__n46396;
  assign new_new_n33382__ = ~ys__n46354 & ~new_new_n33381__;
  assign new_new_n33383__ = ~new_new_n33380__ & new_new_n33382__;
  assign new_new_n33384__ = ys__n316 & ys__n46397;
  assign new_new_n33385__ = ~ys__n316 & ~ys__n46397;
  assign new_new_n33386__ = ~ys__n46356 & ~new_new_n33385__;
  assign new_new_n33387__ = ~new_new_n33384__ & new_new_n33386__;
  assign new_new_n33388__ = ~new_new_n33383__ & ~new_new_n33387__;
  assign new_new_n33389__ = ys__n6115 & ys__n46398;
  assign new_new_n33390__ = ~ys__n6115 & ~ys__n46398;
  assign new_new_n33391__ = ~ys__n46358 & ~new_new_n33390__;
  assign new_new_n33392__ = ~new_new_n33389__ & new_new_n33391__;
  assign new_new_n33393__ = ys__n44 & ys__n46399;
  assign new_new_n33394__ = ~ys__n44 & ~ys__n46399;
  assign new_new_n33395__ = ~ys__n46360 & ~new_new_n33394__;
  assign new_new_n33396__ = ~new_new_n33393__ & new_new_n33395__;
  assign new_new_n33397__ = ~new_new_n33392__ & ~new_new_n33396__;
  assign new_new_n33398__ = new_new_n33388__ & new_new_n33397__;
  assign new_new_n33399__ = new_new_n33379__ & new_new_n33398__;
  assign new_new_n33400__ = new_new_n33360__ & new_new_n33399__;
  assign new_new_n33401__ = new_new_n33311__ & new_new_n33400__;
  assign new_new_n33402__ = ys__n18520 & ys__n46339;
  assign new_new_n33403__ = ~ys__n18520 & ~ys__n46339;
  assign new_new_n33404__ = ~ys__n46300 & ~new_new_n33403__;
  assign new_new_n33405__ = ~new_new_n33402__ & new_new_n33404__;
  assign new_new_n33406__ = ys__n18523 & ys__n46340;
  assign new_new_n33407__ = ~ys__n18523 & ~ys__n46340;
  assign new_new_n33408__ = ~ys__n46302 & ~new_new_n33407__;
  assign new_new_n33409__ = ~new_new_n33406__ & new_new_n33408__;
  assign new_new_n33410__ = ~new_new_n33405__ & ~new_new_n33409__;
  assign new_new_n33411__ = ys__n18526 & ys__n46341;
  assign new_new_n33412__ = ~ys__n18526 & ~ys__n46341;
  assign new_new_n33413__ = ~ys__n46304 & ~new_new_n33412__;
  assign new_new_n33414__ = ~new_new_n33411__ & new_new_n33413__;
  assign new_new_n33415__ = ys__n18529 & ys__n46342;
  assign new_new_n33416__ = ~ys__n18529 & ~ys__n46342;
  assign new_new_n33417__ = ~ys__n46306 & ~new_new_n33416__;
  assign new_new_n33418__ = ~new_new_n33415__ & new_new_n33417__;
  assign new_new_n33419__ = ~new_new_n33414__ & ~new_new_n33418__;
  assign new_new_n33420__ = new_new_n33410__ & new_new_n33419__;
  assign new_new_n33421__ = ys__n18508 & ys__n46335;
  assign new_new_n33422__ = ~ys__n18508 & ~ys__n46335;
  assign new_new_n33423__ = ~ys__n46292 & ~new_new_n33422__;
  assign new_new_n33424__ = ~new_new_n33421__ & new_new_n33423__;
  assign new_new_n33425__ = ys__n18511 & ys__n46336;
  assign new_new_n33426__ = ~ys__n18511 & ~ys__n46336;
  assign new_new_n33427__ = ~ys__n46294 & ~new_new_n33426__;
  assign new_new_n33428__ = ~new_new_n33425__ & new_new_n33427__;
  assign new_new_n33429__ = ~new_new_n33424__ & ~new_new_n33428__;
  assign new_new_n33430__ = ys__n18514 & ys__n46337;
  assign new_new_n33431__ = ~ys__n18514 & ~ys__n46337;
  assign new_new_n33432__ = ~ys__n46296 & ~new_new_n33431__;
  assign new_new_n33433__ = ~new_new_n33430__ & new_new_n33432__;
  assign new_new_n33434__ = ys__n18517 & ys__n46338;
  assign new_new_n33435__ = ~ys__n18517 & ~ys__n46338;
  assign new_new_n33436__ = ~ys__n46298 & ~new_new_n33435__;
  assign new_new_n33437__ = ~new_new_n33434__ & new_new_n33436__;
  assign new_new_n33438__ = ~new_new_n33433__ & ~new_new_n33437__;
  assign new_new_n33439__ = new_new_n33429__ & new_new_n33438__;
  assign new_new_n33440__ = new_new_n33420__ & new_new_n33439__;
  assign new_new_n33441__ = ~ys__n18041 & new_new_n32450__;
  assign new_new_n33442__ = ~ys__n18045 & new_new_n32453__;
  assign new_new_n33443__ = ~ys__n18043 & new_new_n32455__;
  assign new_new_n33444__ = ~new_new_n33442__ & ~new_new_n33443__;
  assign new_new_n33445__ = ~new_new_n33441__ & new_new_n33444__;
  assign new_new_n33446__ = ys__n18532 & ys__n46343;
  assign new_new_n33447__ = ~ys__n18532 & ~ys__n46343;
  assign new_new_n33448__ = ~ys__n46308 & ~new_new_n33447__;
  assign new_new_n33449__ = ~new_new_n33446__ & new_new_n33448__;
  assign new_new_n33450__ = ys__n18535 & ys__n46344;
  assign new_new_n33451__ = ~ys__n18535 & ~ys__n46344;
  assign new_new_n33452__ = ~ys__n46310 & ~new_new_n33451__;
  assign new_new_n33453__ = ~new_new_n33450__ & new_new_n33452__;
  assign new_new_n33454__ = ~new_new_n33449__ & ~new_new_n33453__;
  assign new_new_n33455__ = ys__n18538 & ys__n46345;
  assign new_new_n33456__ = ~ys__n18538 & ~ys__n46345;
  assign new_new_n33457__ = ~ys__n46312 & ~new_new_n33456__;
  assign new_new_n33458__ = ~new_new_n33455__ & new_new_n33457__;
  assign new_new_n33459__ = ys__n18541 & ys__n46346;
  assign new_new_n33460__ = ~ys__n18541 & ~ys__n46346;
  assign new_new_n33461__ = ~ys__n46314 & ~new_new_n33460__;
  assign new_new_n33462__ = ~new_new_n33459__ & new_new_n33461__;
  assign new_new_n33463__ = ~new_new_n33458__ & ~new_new_n33462__;
  assign new_new_n33464__ = new_new_n33454__ & new_new_n33463__;
  assign new_new_n33465__ = new_new_n33445__ & new_new_n33464__;
  assign new_new_n33466__ = new_new_n33440__ & new_new_n33465__;
  assign new_new_n33467__ = ys__n18472 & ys__n46323;
  assign new_new_n33468__ = ~ys__n18472 & ~ys__n46323;
  assign new_new_n33469__ = ~ys__n46268 & ~new_new_n33468__;
  assign new_new_n33470__ = ~new_new_n33467__ & new_new_n33469__;
  assign new_new_n33471__ = ys__n18475 & ys__n46324;
  assign new_new_n33472__ = ~ys__n18475 & ~ys__n46324;
  assign new_new_n33473__ = ~ys__n46270 & ~new_new_n33472__;
  assign new_new_n33474__ = ~new_new_n33471__ & new_new_n33473__;
  assign new_new_n33475__ = ~new_new_n33470__ & ~new_new_n33474__;
  assign new_new_n33476__ = ys__n18478 & ys__n46325;
  assign new_new_n33477__ = ~ys__n18478 & ~ys__n46325;
  assign new_new_n33478__ = ~ys__n46272 & ~new_new_n33477__;
  assign new_new_n33479__ = ~new_new_n33476__ & new_new_n33478__;
  assign new_new_n33480__ = ys__n18481 & ys__n46326;
  assign new_new_n33481__ = ~ys__n18481 & ~ys__n46326;
  assign new_new_n33482__ = ~ys__n46274 & ~new_new_n33481__;
  assign new_new_n33483__ = ~new_new_n33480__ & new_new_n33482__;
  assign new_new_n33484__ = ~new_new_n33479__ & ~new_new_n33483__;
  assign new_new_n33485__ = new_new_n33475__ & new_new_n33484__;
  assign new_new_n33486__ = ys__n18460 & ys__n46319;
  assign new_new_n33487__ = ~ys__n18460 & ~ys__n46319;
  assign new_new_n33488__ = ~ys__n46260 & ~new_new_n33487__;
  assign new_new_n33489__ = ~new_new_n33486__ & new_new_n33488__;
  assign new_new_n33490__ = ys__n18463 & ys__n46320;
  assign new_new_n33491__ = ~ys__n18463 & ~ys__n46320;
  assign new_new_n33492__ = ~ys__n46262 & ~new_new_n33491__;
  assign new_new_n33493__ = ~new_new_n33490__ & new_new_n33492__;
  assign new_new_n33494__ = ~new_new_n33489__ & ~new_new_n33493__;
  assign new_new_n33495__ = ys__n18466 & ys__n46321;
  assign new_new_n33496__ = ~ys__n18466 & ~ys__n46321;
  assign new_new_n33497__ = ~ys__n46264 & ~new_new_n33496__;
  assign new_new_n33498__ = ~new_new_n33495__ & new_new_n33497__;
  assign new_new_n33499__ = ys__n18469 & ys__n46322;
  assign new_new_n33500__ = ~ys__n18469 & ~ys__n46322;
  assign new_new_n33501__ = ~ys__n46266 & ~new_new_n33500__;
  assign new_new_n33502__ = ~new_new_n33499__ & new_new_n33501__;
  assign new_new_n33503__ = ~new_new_n33498__ & ~new_new_n33502__;
  assign new_new_n33504__ = new_new_n33494__ & new_new_n33503__;
  assign new_new_n33505__ = new_new_n33485__ & new_new_n33504__;
  assign new_new_n33506__ = ys__n18496 & ys__n46331;
  assign new_new_n33507__ = ~ys__n18496 & ~ys__n46331;
  assign new_new_n33508__ = ~ys__n46284 & ~new_new_n33507__;
  assign new_new_n33509__ = ~new_new_n33506__ & new_new_n33508__;
  assign new_new_n33510__ = ys__n18499 & ys__n46332;
  assign new_new_n33511__ = ~ys__n18499 & ~ys__n46332;
  assign new_new_n33512__ = ~ys__n46286 & ~new_new_n33511__;
  assign new_new_n33513__ = ~new_new_n33510__ & new_new_n33512__;
  assign new_new_n33514__ = ~new_new_n33509__ & ~new_new_n33513__;
  assign new_new_n33515__ = ys__n18502 & ys__n46333;
  assign new_new_n33516__ = ~ys__n18502 & ~ys__n46333;
  assign new_new_n33517__ = ~ys__n46288 & ~new_new_n33516__;
  assign new_new_n33518__ = ~new_new_n33515__ & new_new_n33517__;
  assign new_new_n33519__ = ys__n18505 & ys__n46334;
  assign new_new_n33520__ = ~ys__n18505 & ~ys__n46334;
  assign new_new_n33521__ = ~ys__n46290 & ~new_new_n33520__;
  assign new_new_n33522__ = ~new_new_n33519__ & new_new_n33521__;
  assign new_new_n33523__ = ~new_new_n33518__ & ~new_new_n33522__;
  assign new_new_n33524__ = new_new_n33514__ & new_new_n33523__;
  assign new_new_n33525__ = ys__n18484 & ys__n46327;
  assign new_new_n33526__ = ~ys__n18484 & ~ys__n46327;
  assign new_new_n33527__ = ~ys__n46276 & ~new_new_n33526__;
  assign new_new_n33528__ = ~new_new_n33525__ & new_new_n33527__;
  assign new_new_n33529__ = ys__n18487 & ys__n46328;
  assign new_new_n33530__ = ~ys__n18487 & ~ys__n46328;
  assign new_new_n33531__ = ~ys__n46278 & ~new_new_n33530__;
  assign new_new_n33532__ = ~new_new_n33529__ & new_new_n33531__;
  assign new_new_n33533__ = ~new_new_n33528__ & ~new_new_n33532__;
  assign new_new_n33534__ = ys__n18490 & ys__n46329;
  assign new_new_n33535__ = ~ys__n18490 & ~ys__n46329;
  assign new_new_n33536__ = ~ys__n46280 & ~new_new_n33535__;
  assign new_new_n33537__ = ~new_new_n33534__ & new_new_n33536__;
  assign new_new_n33538__ = ys__n18493 & ys__n46330;
  assign new_new_n33539__ = ~ys__n18493 & ~ys__n46330;
  assign new_new_n33540__ = ~ys__n46282 & ~new_new_n33539__;
  assign new_new_n33541__ = ~new_new_n33538__ & new_new_n33540__;
  assign new_new_n33542__ = ~new_new_n33537__ & ~new_new_n33541__;
  assign new_new_n33543__ = new_new_n33533__ & new_new_n33542__;
  assign new_new_n33544__ = new_new_n33524__ & new_new_n33543__;
  assign new_new_n33545__ = new_new_n33505__ & new_new_n33544__;
  assign new_new_n33546__ = new_new_n33466__ & new_new_n33545__;
  assign new_new_n33547__ = new_new_n33401__ & new_new_n33546__;
  assign new_new_n33548__ = ~new_new_n33232__ & ~new_new_n33547__;
  assign new_new_n33549__ = ~ys__n27518 & ~new_new_n33232__;
  assign new_new_n33550__ = ~ys__n27518 & ~new_new_n33549__;
  assign new_new_n33551__ = new_new_n33547__ & ~new_new_n33550__;
  assign ys__n27513 = new_new_n33548__ | new_new_n33551__;
  assign new_new_n33553__ = ys__n26772 & ~new_new_n26767__;
  assign new_new_n33554__ = ys__n26772 & ~new_new_n26703__;
  assign new_new_n33555__ = ~new_new_n26726__ & ~new_new_n33554__;
  assign new_new_n33556__ = new_new_n26767__ & ~new_new_n33555__;
  assign new_new_n33557__ = ~new_new_n33553__ & ~new_new_n33556__;
  assign new_new_n33558__ = ~new_new_n33547__ & ~new_new_n33557__;
  assign new_new_n33559__ = ~ys__n27518 & ~new_new_n33557__;
  assign new_new_n33560__ = ~ys__n27518 & ~new_new_n33559__;
  assign new_new_n33561__ = ~ys__n27520 & ~new_new_n33560__;
  assign new_new_n33562__ = ~ys__n27520 & ~new_new_n33561__;
  assign new_new_n33563__ = new_new_n33547__ & ~new_new_n33562__;
  assign ys__n27515 = new_new_n33558__ | new_new_n33563__;
  assign new_new_n33565__ = ys__n27485 & new_new_n32560__;
  assign new_new_n33566__ = ~new_new_n32887__ & new_new_n33565__;
  assign new_new_n33567__ = ~ys__n27498 & new_new_n33565__;
  assign new_new_n33568__ = ~ys__n27498 & ~new_new_n33567__;
  assign new_new_n33569__ = new_new_n32887__ & ~new_new_n33568__;
  assign new_new_n33570__ = ~new_new_n33566__ & ~new_new_n33569__;
  assign new_new_n33571__ = ~new_new_n33214__ & ~new_new_n33570__;
  assign new_new_n33572__ = ~ys__n27509 & ~new_new_n33570__;
  assign new_new_n33573__ = ~ys__n27509 & ~new_new_n33572__;
  assign new_new_n33574__ = new_new_n33214__ & ~new_new_n33573__;
  assign new_new_n33575__ = ~new_new_n33571__ & ~new_new_n33574__;
  assign new_new_n33576__ = ~new_new_n33547__ & ~new_new_n33575__;
  assign new_new_n33577__ = ~ys__n27520 & ~new_new_n33575__;
  assign new_new_n33578__ = ~ys__n27520 & ~new_new_n33577__;
  assign new_new_n33579__ = new_new_n33547__ & ~new_new_n33578__;
  assign ys__n27517 = new_new_n33576__ | new_new_n33579__;
  assign new_new_n33581__ = ys__n874 & ys__n18214;
  assign new_new_n33582__ = ys__n874 & ys__n18218;
  assign new_new_n33583__ = new_new_n33581__ & ~new_new_n33582__;
  assign new_new_n33584__ = ys__n18217 & new_new_n33581__;
  assign new_new_n33585__ = new_new_n33582__ & new_new_n33584__;
  assign ys__n27550 = new_new_n33583__ | new_new_n33585__;
  assign new_new_n33587__ = ~ys__n18217 & ~new_new_n33582__;
  assign new_new_n33588__ = ys__n18217 & new_new_n33582__;
  assign ys__n27551 = new_new_n33587__ | new_new_n33588__;
  assign new_new_n33590__ = ~ys__n18393 & ys__n27737;
  assign new_new_n33591__ = ys__n828 & ys__n18393;
  assign ys__n27598 = new_new_n33590__ | new_new_n33591__;
  assign new_new_n33593__ = ~ys__n18317 & new_new_n12094__;
  assign new_new_n33594__ = ys__n18317 & new_new_n12099__;
  assign new_new_n33595__ = ~new_new_n33593__ & ~new_new_n33594__;
  assign new_new_n33596__ = ys__n18065 & ~new_new_n33595__;
  assign new_new_n33597__ = ys__n27607 & ~new_new_n33596__;
  assign new_new_n33598__ = ys__n27608 & new_new_n33596__;
  assign ys__n27610 = new_new_n33597__ | new_new_n33598__;
  assign new_new_n33600__ = ys__n27611 & ~new_new_n33596__;
  assign new_new_n33601__ = ys__n27612 & new_new_n33596__;
  assign ys__n27613 = new_new_n33600__ | new_new_n33601__;
  assign new_new_n33603__ = ys__n27614 & ~new_new_n33596__;
  assign new_new_n33604__ = ys__n27615 & new_new_n33596__;
  assign ys__n27616 = new_new_n33603__ | new_new_n33604__;
  assign new_new_n33606__ = ys__n27617 & ~new_new_n33596__;
  assign new_new_n33607__ = ys__n27618 & new_new_n33596__;
  assign ys__n27619 = new_new_n33606__ | new_new_n33607__;
  assign new_new_n33609__ = ys__n27620 & ~new_new_n33596__;
  assign new_new_n33610__ = ys__n27621 & new_new_n33596__;
  assign ys__n27622 = new_new_n33609__ | new_new_n33610__;
  assign new_new_n33612__ = ys__n27623 & ~new_new_n33596__;
  assign new_new_n33613__ = ys__n27624 & new_new_n33596__;
  assign ys__n27625 = new_new_n33612__ | new_new_n33613__;
  assign new_new_n33615__ = ys__n27626 & ~new_new_n33596__;
  assign new_new_n33616__ = ys__n27627 & new_new_n33596__;
  assign ys__n27628 = new_new_n33615__ | new_new_n33616__;
  assign new_new_n33618__ = ys__n27629 & ~new_new_n33596__;
  assign new_new_n33619__ = ys__n27630 & new_new_n33596__;
  assign ys__n27631 = new_new_n33618__ | new_new_n33619__;
  assign new_new_n33621__ = ys__n27632 & ~new_new_n33596__;
  assign new_new_n33622__ = ys__n27633 & new_new_n33596__;
  assign ys__n27634 = new_new_n33621__ | new_new_n33622__;
  assign new_new_n33624__ = ys__n27635 & ~new_new_n33596__;
  assign new_new_n33625__ = ys__n27636 & new_new_n33596__;
  assign ys__n27637 = new_new_n33624__ | new_new_n33625__;
  assign new_new_n33627__ = ys__n27638 & ~new_new_n33596__;
  assign new_new_n33628__ = ys__n27639 & new_new_n33596__;
  assign ys__n27640 = new_new_n33627__ | new_new_n33628__;
  assign new_new_n33630__ = ys__n27641 & ~new_new_n33596__;
  assign new_new_n33631__ = ys__n27642 & new_new_n33596__;
  assign ys__n27643 = new_new_n33630__ | new_new_n33631__;
  assign new_new_n33633__ = ys__n27644 & ~new_new_n33596__;
  assign new_new_n33634__ = ys__n27645 & new_new_n33596__;
  assign ys__n27646 = new_new_n33633__ | new_new_n33634__;
  assign new_new_n33636__ = ys__n27647 & ~new_new_n33596__;
  assign new_new_n33637__ = ys__n27648 & new_new_n33596__;
  assign ys__n27649 = new_new_n33636__ | new_new_n33637__;
  assign new_new_n33639__ = ys__n27650 & ~new_new_n33596__;
  assign new_new_n33640__ = ys__n27651 & new_new_n33596__;
  assign ys__n27652 = new_new_n33639__ | new_new_n33640__;
  assign new_new_n33642__ = ys__n27653 & ~new_new_n33596__;
  assign new_new_n33643__ = ys__n27654 & new_new_n33596__;
  assign ys__n27655 = new_new_n33642__ | new_new_n33643__;
  assign new_new_n33645__ = ys__n27656 & ~new_new_n33596__;
  assign new_new_n33646__ = ys__n27657 & new_new_n33596__;
  assign ys__n27658 = new_new_n33645__ | new_new_n33646__;
  assign new_new_n33648__ = ys__n27659 & ~new_new_n33596__;
  assign new_new_n33649__ = ys__n27660 & new_new_n33596__;
  assign ys__n27661 = new_new_n33648__ | new_new_n33649__;
  assign new_new_n33651__ = ys__n27662 & ~new_new_n33596__;
  assign new_new_n33652__ = ys__n27663 & new_new_n33596__;
  assign ys__n27664 = new_new_n33651__ | new_new_n33652__;
  assign new_new_n33654__ = ys__n27665 & ~new_new_n33596__;
  assign new_new_n33655__ = ys__n27666 & new_new_n33596__;
  assign ys__n27667 = new_new_n33654__ | new_new_n33655__;
  assign new_new_n33657__ = ys__n27668 & ~new_new_n33596__;
  assign new_new_n33658__ = ys__n27669 & new_new_n33596__;
  assign ys__n27670 = new_new_n33657__ | new_new_n33658__;
  assign new_new_n33660__ = ys__n27671 & ~new_new_n33596__;
  assign new_new_n33661__ = ys__n27672 & new_new_n33596__;
  assign ys__n27673 = new_new_n33660__ | new_new_n33661__;
  assign new_new_n33663__ = ys__n27674 & ~new_new_n33596__;
  assign new_new_n33664__ = ys__n27675 & new_new_n33596__;
  assign ys__n27676 = new_new_n33663__ | new_new_n33664__;
  assign new_new_n33666__ = ys__n27677 & ~new_new_n33596__;
  assign new_new_n33667__ = ys__n27678 & new_new_n33596__;
  assign ys__n27679 = new_new_n33666__ | new_new_n33667__;
  assign new_new_n33669__ = ys__n27680 & ~new_new_n33596__;
  assign new_new_n33670__ = ys__n27681 & new_new_n33596__;
  assign ys__n27682 = new_new_n33669__ | new_new_n33670__;
  assign new_new_n33672__ = ys__n27683 & ~new_new_n33596__;
  assign new_new_n33673__ = ys__n27684 & new_new_n33596__;
  assign ys__n27685 = new_new_n33672__ | new_new_n33673__;
  assign new_new_n33675__ = ys__n27686 & ~new_new_n33596__;
  assign new_new_n33676__ = ys__n27687 & new_new_n33596__;
  assign ys__n27688 = new_new_n33675__ | new_new_n33676__;
  assign new_new_n33678__ = ys__n27689 & ~new_new_n33596__;
  assign new_new_n33679__ = ys__n27690 & new_new_n33596__;
  assign ys__n27691 = new_new_n33678__ | new_new_n33679__;
  assign new_new_n33681__ = ys__n27692 & ~new_new_n33596__;
  assign new_new_n33682__ = ys__n27693 & new_new_n33596__;
  assign ys__n27694 = new_new_n33681__ | new_new_n33682__;
  assign new_new_n33684__ = ys__n27695 & ~new_new_n33596__;
  assign new_new_n33685__ = ys__n27696 & new_new_n33596__;
  assign ys__n27697 = new_new_n33684__ | new_new_n33685__;
  assign new_new_n33687__ = ys__n27698 & ~new_new_n33596__;
  assign new_new_n33688__ = ys__n27699 & new_new_n33596__;
  assign ys__n27700 = new_new_n33687__ | new_new_n33688__;
  assign new_new_n33690__ = ys__n27701 & ~new_new_n33596__;
  assign new_new_n33691__ = ys__n27702 & new_new_n33596__;
  assign ys__n27703 = new_new_n33690__ | new_new_n33691__;
  assign new_new_n33693__ = ~ys__n18065 & ~new_new_n33595__;
  assign new_new_n33694__ = ys__n27607 & ~new_new_n33693__;
  assign new_new_n33695__ = ys__n27608 & new_new_n33693__;
  assign ys__n27705 = new_new_n33694__ | new_new_n33695__;
  assign new_new_n33697__ = ys__n27611 & ~new_new_n33693__;
  assign new_new_n33698__ = ys__n27612 & new_new_n33693__;
  assign ys__n27706 = new_new_n33697__ | new_new_n33698__;
  assign new_new_n33700__ = ys__n27614 & ~new_new_n33693__;
  assign new_new_n33701__ = ys__n27615 & new_new_n33693__;
  assign ys__n27707 = new_new_n33700__ | new_new_n33701__;
  assign new_new_n33703__ = ys__n27617 & ~new_new_n33693__;
  assign new_new_n33704__ = ys__n27618 & new_new_n33693__;
  assign ys__n27708 = new_new_n33703__ | new_new_n33704__;
  assign new_new_n33706__ = ys__n27620 & ~new_new_n33693__;
  assign new_new_n33707__ = ys__n27621 & new_new_n33693__;
  assign ys__n27709 = new_new_n33706__ | new_new_n33707__;
  assign new_new_n33709__ = ys__n27623 & ~new_new_n33693__;
  assign new_new_n33710__ = ys__n27624 & new_new_n33693__;
  assign ys__n27710 = new_new_n33709__ | new_new_n33710__;
  assign new_new_n33712__ = ys__n27626 & ~new_new_n33693__;
  assign new_new_n33713__ = ys__n27627 & new_new_n33693__;
  assign ys__n27711 = new_new_n33712__ | new_new_n33713__;
  assign new_new_n33715__ = ys__n27629 & ~new_new_n33693__;
  assign new_new_n33716__ = ys__n27630 & new_new_n33693__;
  assign ys__n27712 = new_new_n33715__ | new_new_n33716__;
  assign new_new_n33718__ = ys__n27632 & ~new_new_n33693__;
  assign new_new_n33719__ = ys__n27633 & new_new_n33693__;
  assign ys__n27713 = new_new_n33718__ | new_new_n33719__;
  assign new_new_n33721__ = ys__n27635 & ~new_new_n33693__;
  assign new_new_n33722__ = ys__n27636 & new_new_n33693__;
  assign ys__n27714 = new_new_n33721__ | new_new_n33722__;
  assign new_new_n33724__ = ys__n27638 & ~new_new_n33693__;
  assign new_new_n33725__ = ys__n27639 & new_new_n33693__;
  assign ys__n27715 = new_new_n33724__ | new_new_n33725__;
  assign new_new_n33727__ = ys__n27641 & ~new_new_n33693__;
  assign new_new_n33728__ = ys__n27642 & new_new_n33693__;
  assign ys__n27716 = new_new_n33727__ | new_new_n33728__;
  assign new_new_n33730__ = ys__n27644 & ~new_new_n33693__;
  assign new_new_n33731__ = ys__n27645 & new_new_n33693__;
  assign ys__n27717 = new_new_n33730__ | new_new_n33731__;
  assign new_new_n33733__ = ys__n27647 & ~new_new_n33693__;
  assign new_new_n33734__ = ys__n27648 & new_new_n33693__;
  assign ys__n27718 = new_new_n33733__ | new_new_n33734__;
  assign new_new_n33736__ = ys__n27650 & ~new_new_n33693__;
  assign new_new_n33737__ = ys__n27651 & new_new_n33693__;
  assign ys__n27719 = new_new_n33736__ | new_new_n33737__;
  assign new_new_n33739__ = ys__n27653 & ~new_new_n33693__;
  assign new_new_n33740__ = ys__n27654 & new_new_n33693__;
  assign ys__n27720 = new_new_n33739__ | new_new_n33740__;
  assign new_new_n33742__ = ys__n27656 & ~new_new_n33693__;
  assign new_new_n33743__ = ys__n27657 & new_new_n33693__;
  assign ys__n27721 = new_new_n33742__ | new_new_n33743__;
  assign new_new_n33745__ = ys__n27659 & ~new_new_n33693__;
  assign new_new_n33746__ = ys__n27660 & new_new_n33693__;
  assign ys__n27722 = new_new_n33745__ | new_new_n33746__;
  assign new_new_n33748__ = ys__n27662 & ~new_new_n33693__;
  assign new_new_n33749__ = ys__n27663 & new_new_n33693__;
  assign ys__n27723 = new_new_n33748__ | new_new_n33749__;
  assign new_new_n33751__ = ys__n27665 & ~new_new_n33693__;
  assign new_new_n33752__ = ys__n27666 & new_new_n33693__;
  assign ys__n27724 = new_new_n33751__ | new_new_n33752__;
  assign new_new_n33754__ = ys__n27668 & ~new_new_n33693__;
  assign new_new_n33755__ = ys__n27669 & new_new_n33693__;
  assign ys__n27725 = new_new_n33754__ | new_new_n33755__;
  assign new_new_n33757__ = ys__n27671 & ~new_new_n33693__;
  assign new_new_n33758__ = ys__n27672 & new_new_n33693__;
  assign ys__n27726 = new_new_n33757__ | new_new_n33758__;
  assign new_new_n33760__ = ys__n27674 & ~new_new_n33693__;
  assign new_new_n33761__ = ys__n27675 & new_new_n33693__;
  assign ys__n27727 = new_new_n33760__ | new_new_n33761__;
  assign new_new_n33763__ = ys__n27677 & ~new_new_n33693__;
  assign new_new_n33764__ = ys__n27678 & new_new_n33693__;
  assign ys__n27728 = new_new_n33763__ | new_new_n33764__;
  assign new_new_n33766__ = ys__n27680 & ~new_new_n33693__;
  assign new_new_n33767__ = ys__n27681 & new_new_n33693__;
  assign ys__n27729 = new_new_n33766__ | new_new_n33767__;
  assign new_new_n33769__ = ys__n27683 & ~new_new_n33693__;
  assign new_new_n33770__ = ys__n27684 & new_new_n33693__;
  assign ys__n27730 = new_new_n33769__ | new_new_n33770__;
  assign new_new_n33772__ = ys__n27686 & ~new_new_n33693__;
  assign new_new_n33773__ = ys__n27687 & new_new_n33693__;
  assign ys__n27731 = new_new_n33772__ | new_new_n33773__;
  assign new_new_n33775__ = ys__n27689 & ~new_new_n33693__;
  assign new_new_n33776__ = ys__n27690 & new_new_n33693__;
  assign ys__n27732 = new_new_n33775__ | new_new_n33776__;
  assign new_new_n33778__ = ys__n27692 & ~new_new_n33693__;
  assign new_new_n33779__ = ys__n27693 & new_new_n33693__;
  assign ys__n27733 = new_new_n33778__ | new_new_n33779__;
  assign new_new_n33781__ = ys__n27695 & ~new_new_n33693__;
  assign new_new_n33782__ = ys__n27696 & new_new_n33693__;
  assign ys__n27734 = new_new_n33781__ | new_new_n33782__;
  assign new_new_n33784__ = ys__n27698 & ~new_new_n33693__;
  assign new_new_n33785__ = ys__n27699 & new_new_n33693__;
  assign ys__n27735 = new_new_n33784__ | new_new_n33785__;
  assign new_new_n33787__ = ys__n27701 & ~new_new_n33693__;
  assign new_new_n33788__ = ys__n27702 & new_new_n33693__;
  assign ys__n27736 = new_new_n33787__ | new_new_n33788__;
  assign ys__n27739 = ~ys__n35065 & ~new_new_n11141__;
  assign new_new_n33791__ = ~ys__n18393 & ys__n27739;
  assign new_new_n33792__ = ys__n18393 & ys__n27740;
  assign ys__n27741 = new_new_n33791__ | new_new_n33792__;
  assign ys__n28258 = ~ys__n1535 & ys__n28243;
  assign ys__n28276 = ys__n1535 & ys__n28243;
  assign new_new_n33796__ = ys__n240 & ~ys__n1535;
  assign new_new_n33797__ = ~ys__n1535 & ~new_new_n33796__;
  assign ys__n28328 = ys__n28243 & ~new_new_n33797__;
  assign new_new_n33799__ = ys__n238 & ~ys__n1535;
  assign new_new_n33800__ = ~ys__n1535 & ~new_new_n33799__;
  assign ys__n28330 = ys__n28243 & ~new_new_n33800__;
  assign new_new_n33802__ = ys__n242 & ~ys__n1535;
  assign new_new_n33803__ = ~ys__n1535 & ~new_new_n33802__;
  assign ys__n28332 = ys__n28243 & ~new_new_n33803__;
  assign new_new_n33805__ = ~ys__n238 & ~ys__n242;
  assign new_new_n33806__ = ~ys__n1535 & new_new_n33805__;
  assign new_new_n33807__ = ~ys__n1535 & ~new_new_n33806__;
  assign ys__n28336 = ys__n28243 & ~new_new_n33807__;
  assign new_new_n33809__ = ys__n758 & ~ys__n760;
  assign new_new_n33810__ = ~ys__n762 & ~ys__n764;
  assign new_new_n33811__ = new_new_n33809__ & new_new_n33810__;
  assign new_new_n33812__ = ~ys__n766 & ys__n38198;
  assign new_new_n33813__ = new_new_n33811__ & new_new_n33812__;
  assign ys__n28343 = ~ys__n4566 & new_new_n33813__;
  assign new_new_n33815__ = ~ys__n758 & ys__n760;
  assign new_new_n33816__ = new_new_n33810__ & new_new_n33815__;
  assign new_new_n33817__ = new_new_n33812__ & new_new_n33816__;
  assign ys__n28345 = ~ys__n4566 & new_new_n33817__;
  assign new_new_n33819__ = ys__n758 & ys__n760;
  assign new_new_n33820__ = new_new_n33810__ & new_new_n33819__;
  assign new_new_n33821__ = new_new_n33812__ & new_new_n33820__;
  assign ys__n28347 = ~ys__n4566 & new_new_n33821__;
  assign new_new_n33823__ = ~ys__n758 & ~ys__n760;
  assign new_new_n33824__ = ys__n762 & ~ys__n764;
  assign new_new_n33825__ = new_new_n33823__ & new_new_n33824__;
  assign new_new_n33826__ = new_new_n33812__ & new_new_n33825__;
  assign ys__n28349 = ~ys__n4566 & new_new_n33826__;
  assign new_new_n33828__ = new_new_n33809__ & new_new_n33824__;
  assign new_new_n33829__ = new_new_n33812__ & new_new_n33828__;
  assign ys__n28351 = ~ys__n4566 & new_new_n33829__;
  assign new_new_n33831__ = new_new_n33815__ & new_new_n33824__;
  assign new_new_n33832__ = new_new_n33812__ & new_new_n33831__;
  assign ys__n28353 = ~ys__n4566 & new_new_n33832__;
  assign new_new_n33834__ = new_new_n33819__ & new_new_n33824__;
  assign new_new_n33835__ = new_new_n33812__ & new_new_n33834__;
  assign ys__n28355 = ~ys__n4566 & new_new_n33835__;
  assign new_new_n33837__ = ~ys__n762 & ys__n764;
  assign new_new_n33838__ = new_new_n33823__ & new_new_n33837__;
  assign new_new_n33839__ = new_new_n33812__ & new_new_n33838__;
  assign ys__n28357 = ~ys__n4566 & new_new_n33839__;
  assign new_new_n33841__ = new_new_n33809__ & new_new_n33837__;
  assign new_new_n33842__ = new_new_n33812__ & new_new_n33841__;
  assign ys__n28359 = ~ys__n4566 & new_new_n33842__;
  assign new_new_n33844__ = new_new_n33815__ & new_new_n33837__;
  assign new_new_n33845__ = new_new_n33812__ & new_new_n33844__;
  assign ys__n28361 = ~ys__n4566 & new_new_n33845__;
  assign new_new_n33847__ = new_new_n33819__ & new_new_n33837__;
  assign new_new_n33848__ = new_new_n33812__ & new_new_n33847__;
  assign ys__n28363 = ~ys__n4566 & new_new_n33848__;
  assign new_new_n33850__ = ys__n762 & ys__n764;
  assign new_new_n33851__ = new_new_n33823__ & new_new_n33850__;
  assign new_new_n33852__ = new_new_n33812__ & new_new_n33851__;
  assign ys__n28365 = ~ys__n4566 & new_new_n33852__;
  assign new_new_n33854__ = new_new_n33809__ & new_new_n33850__;
  assign new_new_n33855__ = new_new_n33812__ & new_new_n33854__;
  assign ys__n28367 = ~ys__n4566 & new_new_n33855__;
  assign new_new_n33857__ = new_new_n33815__ & new_new_n33850__;
  assign new_new_n33858__ = new_new_n33812__ & new_new_n33857__;
  assign ys__n28369 = ~ys__n4566 & new_new_n33858__;
  assign new_new_n33860__ = new_new_n33819__ & new_new_n33850__;
  assign new_new_n33861__ = new_new_n33812__ & new_new_n33860__;
  assign ys__n28371 = ~ys__n4566 & new_new_n33861__;
  assign new_new_n33863__ = ys__n766 & ys__n38198;
  assign new_new_n33864__ = new_new_n33810__ & new_new_n33863__;
  assign new_new_n33865__ = new_new_n33823__ & new_new_n33864__;
  assign ys__n28373 = ~ys__n4566 & new_new_n33865__;
  assign new_new_n33867__ = new_new_n33811__ & new_new_n33863__;
  assign ys__n28375 = ~ys__n4566 & new_new_n33867__;
  assign new_new_n33869__ = new_new_n33816__ & new_new_n33863__;
  assign ys__n28377 = ~ys__n4566 & new_new_n33869__;
  assign new_new_n33871__ = new_new_n33820__ & new_new_n33863__;
  assign ys__n28379 = ~ys__n4566 & new_new_n33871__;
  assign new_new_n33873__ = new_new_n33825__ & new_new_n33863__;
  assign ys__n28381 = ~ys__n4566 & new_new_n33873__;
  assign new_new_n33875__ = new_new_n33828__ & new_new_n33863__;
  assign ys__n28383 = ~ys__n4566 & new_new_n33875__;
  assign new_new_n33877__ = new_new_n33831__ & new_new_n33863__;
  assign ys__n28385 = ~ys__n4566 & new_new_n33877__;
  assign new_new_n33879__ = new_new_n33834__ & new_new_n33863__;
  assign ys__n28387 = ~ys__n4566 & new_new_n33879__;
  assign new_new_n33881__ = new_new_n33838__ & new_new_n33863__;
  assign ys__n28389 = ~ys__n4566 & new_new_n33881__;
  assign new_new_n33883__ = new_new_n33841__ & new_new_n33863__;
  assign ys__n28391 = ~ys__n4566 & new_new_n33883__;
  assign new_new_n33885__ = new_new_n33844__ & new_new_n33863__;
  assign ys__n28393 = ~ys__n4566 & new_new_n33885__;
  assign new_new_n33887__ = new_new_n33847__ & new_new_n33863__;
  assign ys__n28395 = ~ys__n4566 & new_new_n33887__;
  assign new_new_n33889__ = new_new_n33851__ & new_new_n33863__;
  assign ys__n28397 = ~ys__n4566 & new_new_n33889__;
  assign new_new_n33891__ = new_new_n33854__ & new_new_n33863__;
  assign ys__n28399 = ~ys__n4566 & new_new_n33891__;
  assign new_new_n33893__ = new_new_n33857__ & new_new_n33863__;
  assign ys__n28401 = ~ys__n4566 & new_new_n33893__;
  assign new_new_n33895__ = new_new_n33860__ & new_new_n33863__;
  assign ys__n28403 = ~ys__n4566 & new_new_n33895__;
  assign new_new_n33897__ = ~new_new_n13884__ & new_new_n13910__;
  assign new_new_n33898__ = new_new_n13884__ & new_new_n13917__;
  assign ys__n28406 = new_new_n33897__ | new_new_n33898__;
  assign new_new_n33900__ = ~ys__n738 & new_new_n13887__;
  assign new_new_n33901__ = new_new_n13902__ & new_new_n33900__;
  assign new_new_n33902__ = ~new_new_n13899__ & ~new_new_n33901__;
  assign new_new_n33903__ = ~new_new_n13884__ & new_new_n33902__;
  assign new_new_n33904__ = new_new_n13884__ & ~new_new_n13899__;
  assign ys__n28409 = new_new_n33903__ | new_new_n33904__;
  assign new_new_n33906__ = ys__n935 & ~ys__n478;
  assign new_new_n33907__ = ~ys__n232 & ~ys__n935;
  assign new_new_n33908__ = ~ys__n478 & new_new_n33907__;
  assign new_new_n33909__ = ~new_new_n33906__ & ~new_new_n33908__;
  assign new_new_n33910__ = ys__n38427 & ~new_new_n33909__;
  assign new_new_n33911__ = ys__n232 & ~ys__n935;
  assign new_new_n33912__ = ~ys__n478 & new_new_n33911__;
  assign new_new_n33913__ = ys__n47755 & new_new_n33912__;
  assign new_new_n33914__ = ~new_new_n33910__ & ~new_new_n33913__;
  assign new_new_n33915__ = ~ys__n478 & ~new_new_n33912__;
  assign new_new_n33916__ = new_new_n33909__ & new_new_n33915__;
  assign new_new_n33917__ = ~new_new_n12635__ & ~new_new_n33916__;
  assign new_new_n33918__ = ~new_new_n33914__ & new_new_n33917__;
  assign new_new_n33919__ = ys__n28462 & new_new_n12635__;
  assign ys__n28410 = new_new_n33918__ | new_new_n33919__;
  assign new_new_n33921__ = ~ys__n4454 & ys__n4455;
  assign new_new_n33922__ = ys__n22885 & new_new_n33921__;
  assign new_new_n33923__ = ys__n4454 & ys__n22822;
  assign new_new_n33924__ = ~new_new_n33922__ & ~new_new_n33923__;
  assign new_new_n33925__ = ~ys__n4452 & ~new_new_n33924__;
  assign new_new_n33926__ = ys__n4452 & ys__n22779;
  assign new_new_n33927__ = ~new_new_n33925__ & ~new_new_n33926__;
  assign new_new_n33928__ = ~ys__n4457 & ~new_new_n33927__;
  assign new_new_n33929__ = ys__n4457 & ys__n22715;
  assign new_new_n33930__ = ~new_new_n33928__ & ~new_new_n33929__;
  assign new_new_n33931__ = ~ys__n4451 & ~new_new_n33930__;
  assign new_new_n33932__ = ys__n4451 & ys__n22675;
  assign new_new_n33933__ = ~new_new_n33931__ & ~new_new_n33932__;
  assign new_new_n33934__ = ~ys__n4449 & ~ys__n4458;
  assign new_new_n33935__ = ~new_new_n33933__ & new_new_n33934__;
  assign new_new_n33936__ = ys__n4458 & ys__n22564;
  assign new_new_n33937__ = ~new_new_n33935__ & ~new_new_n33936__;
  assign new_new_n33938__ = ~ys__n4460 & ~ys__n4461;
  assign new_new_n33939__ = ~new_new_n33937__ & new_new_n33938__;
  assign new_new_n33940__ = ~ys__n4460 & ~new_new_n33939__;
  assign new_new_n33941__ = ~ys__n4448 & ~new_new_n33940__;
  assign new_new_n33942__ = ys__n4448 & ys__n28410;
  assign ys__n28411 = new_new_n33941__ | new_new_n33942__;
  assign new_new_n33944__ = ys__n38315 & ~new_new_n33909__;
  assign new_new_n33945__ = ys__n47756 & new_new_n33912__;
  assign new_new_n33946__ = ~new_new_n33944__ & ~new_new_n33945__;
  assign new_new_n33947__ = new_new_n33917__ & ~new_new_n33946__;
  assign new_new_n33948__ = ys__n28464 & new_new_n12635__;
  assign ys__n28412 = new_new_n33947__ | new_new_n33948__;
  assign new_new_n33950__ = ys__n22886 & new_new_n33921__;
  assign new_new_n33951__ = ys__n4454 & ys__n22824;
  assign new_new_n33952__ = ~new_new_n33950__ & ~new_new_n33951__;
  assign new_new_n33953__ = ~ys__n4452 & ~new_new_n33952__;
  assign new_new_n33954__ = ys__n4452 & ys__n22781;
  assign new_new_n33955__ = ~new_new_n33953__ & ~new_new_n33954__;
  assign new_new_n33956__ = ~ys__n4457 & ~new_new_n33955__;
  assign new_new_n33957__ = ys__n4457 & ys__n22717;
  assign new_new_n33958__ = ~new_new_n33956__ & ~new_new_n33957__;
  assign new_new_n33959__ = ~ys__n4451 & ~new_new_n33958__;
  assign new_new_n33960__ = ys__n4451 & ys__n22677;
  assign new_new_n33961__ = ~new_new_n33959__ & ~new_new_n33960__;
  assign new_new_n33962__ = new_new_n33934__ & ~new_new_n33961__;
  assign new_new_n33963__ = ys__n4458 & ys__n22566;
  assign new_new_n33964__ = ~new_new_n33962__ & ~new_new_n33963__;
  assign new_new_n33965__ = ~ys__n4448 & ~ys__n4460;
  assign new_new_n33966__ = ~ys__n4461 & new_new_n33965__;
  assign new_new_n33967__ = ~new_new_n33964__ & new_new_n33966__;
  assign new_new_n33968__ = ys__n4448 & ys__n28412;
  assign ys__n28413 = new_new_n33967__ | new_new_n33968__;
  assign new_new_n33970__ = ys__n47755 & ~new_new_n33909__;
  assign new_new_n33971__ = ys__n47757 & new_new_n33912__;
  assign new_new_n33972__ = ys__n38427 & ys__n478;
  assign new_new_n33973__ = ~new_new_n33971__ & ~new_new_n33972__;
  assign new_new_n33974__ = ~new_new_n33970__ & new_new_n33973__;
  assign new_new_n33975__ = new_new_n33917__ & ~new_new_n33974__;
  assign new_new_n33976__ = ys__n28466 & new_new_n12635__;
  assign ys__n28414 = new_new_n33975__ | new_new_n33976__;
  assign new_new_n33978__ = ys__n22887 & new_new_n33921__;
  assign new_new_n33979__ = ys__n4454 & ys__n22826;
  assign new_new_n33980__ = ~new_new_n33978__ & ~new_new_n33979__;
  assign new_new_n33981__ = ~ys__n4452 & ~new_new_n33980__;
  assign new_new_n33982__ = ys__n4452 & ys__n22783;
  assign new_new_n33983__ = ~new_new_n33981__ & ~new_new_n33982__;
  assign new_new_n33984__ = ~ys__n4457 & ~new_new_n33983__;
  assign new_new_n33985__ = ys__n4457 & ys__n22719;
  assign new_new_n33986__ = ~new_new_n33984__ & ~new_new_n33985__;
  assign new_new_n33987__ = ~ys__n4451 & ~new_new_n33986__;
  assign new_new_n33988__ = ys__n4451 & ys__n22679;
  assign new_new_n33989__ = ~new_new_n33987__ & ~new_new_n33988__;
  assign new_new_n33990__ = ~ys__n4449 & ~new_new_n33989__;
  assign new_new_n33991__ = ys__n4449 & ys__n22630;
  assign new_new_n33992__ = ~new_new_n33990__ & ~new_new_n33991__;
  assign new_new_n33993__ = ~ys__n4458 & ~new_new_n33992__;
  assign new_new_n33994__ = ys__n4458 & ys__n22568;
  assign new_new_n33995__ = ~new_new_n33993__ & ~new_new_n33994__;
  assign new_new_n33996__ = new_new_n33966__ & ~new_new_n33995__;
  assign new_new_n33997__ = ys__n4448 & ys__n28414;
  assign ys__n28415 = new_new_n33996__ | new_new_n33997__;
  assign new_new_n33999__ = ys__n47756 & ~new_new_n33909__;
  assign new_new_n34000__ = ys__n47758 & new_new_n33912__;
  assign new_new_n34001__ = ys__n38315 & ys__n478;
  assign new_new_n34002__ = ~new_new_n34000__ & ~new_new_n34001__;
  assign new_new_n34003__ = ~new_new_n33999__ & new_new_n34002__;
  assign new_new_n34004__ = new_new_n33917__ & ~new_new_n34003__;
  assign new_new_n34005__ = ys__n28468 & new_new_n12635__;
  assign ys__n28416 = new_new_n34004__ | new_new_n34005__;
  assign new_new_n34007__ = ys__n22888 & new_new_n33921__;
  assign new_new_n34008__ = ys__n4454 & ys__n22828;
  assign new_new_n34009__ = ~new_new_n34007__ & ~new_new_n34008__;
  assign new_new_n34010__ = ~ys__n4452 & ~new_new_n34009__;
  assign new_new_n34011__ = ys__n4452 & ys__n22785;
  assign new_new_n34012__ = ~new_new_n34010__ & ~new_new_n34011__;
  assign new_new_n34013__ = ~ys__n4457 & ~new_new_n34012__;
  assign new_new_n34014__ = ys__n4457 & ys__n22721;
  assign new_new_n34015__ = ~new_new_n34013__ & ~new_new_n34014__;
  assign new_new_n34016__ = ~ys__n4451 & ~new_new_n34015__;
  assign new_new_n34017__ = ys__n4451 & ys__n22681;
  assign new_new_n34018__ = ~new_new_n34016__ & ~new_new_n34017__;
  assign new_new_n34019__ = ~ys__n4449 & ~new_new_n34018__;
  assign new_new_n34020__ = ys__n4449 & ys__n22632;
  assign new_new_n34021__ = ~new_new_n34019__ & ~new_new_n34020__;
  assign new_new_n34022__ = ~ys__n4458 & ~new_new_n34021__;
  assign new_new_n34023__ = ys__n4458 & ys__n22570;
  assign new_new_n34024__ = ~new_new_n34022__ & ~new_new_n34023__;
  assign new_new_n34025__ = ~ys__n4461 & ~new_new_n34024__;
  assign new_new_n34026__ = ~ys__n4461 & ~new_new_n34025__;
  assign new_new_n34027__ = new_new_n33965__ & ~new_new_n34026__;
  assign new_new_n34028__ = ys__n4448 & ys__n28416;
  assign ys__n28417 = new_new_n34027__ | new_new_n34028__;
  assign new_new_n34030__ = ys__n47757 & ~new_new_n33909__;
  assign new_new_n34031__ = ys__n47755 & ys__n478;
  assign new_new_n34032__ = ~new_new_n33971__ & ~new_new_n34031__;
  assign new_new_n34033__ = ~new_new_n34030__ & new_new_n34032__;
  assign new_new_n34034__ = new_new_n33917__ & ~new_new_n34033__;
  assign new_new_n34035__ = ys__n28470 & new_new_n12635__;
  assign ys__n28418 = new_new_n34034__ | new_new_n34035__;
  assign new_new_n34037__ = ys__n22889 & new_new_n33921__;
  assign new_new_n34038__ = ys__n4454 & ys__n22830;
  assign new_new_n34039__ = ~new_new_n34037__ & ~new_new_n34038__;
  assign new_new_n34040__ = ~ys__n4452 & ~new_new_n34039__;
  assign new_new_n34041__ = ys__n4452 & ys__n22787;
  assign new_new_n34042__ = ~new_new_n34040__ & ~new_new_n34041__;
  assign new_new_n34043__ = ~ys__n4457 & ~new_new_n34042__;
  assign new_new_n34044__ = ys__n4457 & ys__n22723;
  assign new_new_n34045__ = ~new_new_n34043__ & ~new_new_n34044__;
  assign new_new_n34046__ = ~ys__n4451 & ~new_new_n34045__;
  assign new_new_n34047__ = ys__n4451 & ys__n22683;
  assign new_new_n34048__ = ~new_new_n34046__ & ~new_new_n34047__;
  assign new_new_n34049__ = ~ys__n4449 & ~new_new_n34048__;
  assign new_new_n34050__ = ys__n4449 & ys__n22634;
  assign new_new_n34051__ = ~new_new_n34049__ & ~new_new_n34050__;
  assign new_new_n34052__ = ~ys__n4458 & ~new_new_n34051__;
  assign new_new_n34053__ = ys__n4458 & ys__n22572;
  assign new_new_n34054__ = ~new_new_n34052__ & ~new_new_n34053__;
  assign new_new_n34055__ = new_new_n33966__ & ~new_new_n34054__;
  assign new_new_n34056__ = ys__n4448 & ys__n28418;
  assign ys__n28419 = new_new_n34055__ | new_new_n34056__;
  assign new_new_n34058__ = ys__n47758 & ~new_new_n33909__;
  assign new_new_n34059__ = ys__n47756 & ys__n478;
  assign new_new_n34060__ = ~new_new_n34000__ & ~new_new_n34059__;
  assign new_new_n34061__ = ~new_new_n34058__ & new_new_n34060__;
  assign new_new_n34062__ = new_new_n33917__ & ~new_new_n34061__;
  assign new_new_n34063__ = ys__n28472 & new_new_n12635__;
  assign ys__n28420 = new_new_n34062__ | new_new_n34063__;
  assign new_new_n34065__ = ys__n22890 & new_new_n33921__;
  assign new_new_n34066__ = ys__n4454 & ys__n22832;
  assign new_new_n34067__ = ~new_new_n34065__ & ~new_new_n34066__;
  assign new_new_n34068__ = ~ys__n4452 & ~new_new_n34067__;
  assign new_new_n34069__ = ys__n4452 & ys__n22789;
  assign new_new_n34070__ = ~new_new_n34068__ & ~new_new_n34069__;
  assign new_new_n34071__ = ~ys__n4457 & ~new_new_n34070__;
  assign new_new_n34072__ = ys__n4457 & ys__n22725;
  assign new_new_n34073__ = ~new_new_n34071__ & ~new_new_n34072__;
  assign new_new_n34074__ = ~ys__n4451 & ~new_new_n34073__;
  assign new_new_n34075__ = ys__n4451 & ys__n22685;
  assign new_new_n34076__ = ~new_new_n34074__ & ~new_new_n34075__;
  assign new_new_n34077__ = ~ys__n4449 & ~new_new_n34076__;
  assign new_new_n34078__ = ys__n4449 & ys__n22636;
  assign new_new_n34079__ = ~new_new_n34077__ & ~new_new_n34078__;
  assign new_new_n34080__ = ~ys__n4458 & ~new_new_n34079__;
  assign new_new_n34081__ = ys__n4458 & ys__n22574;
  assign new_new_n34082__ = ~new_new_n34080__ & ~new_new_n34081__;
  assign new_new_n34083__ = new_new_n33966__ & ~new_new_n34082__;
  assign new_new_n34084__ = ys__n4448 & ys__n28420;
  assign ys__n28421 = new_new_n34083__ | new_new_n34084__;
  assign new_new_n34086__ = ys__n22891 & new_new_n33921__;
  assign new_new_n34087__ = ys__n4454 & ys__n22834;
  assign new_new_n34088__ = ~new_new_n34086__ & ~new_new_n34087__;
  assign new_new_n34089__ = ~ys__n4452 & ~ys__n4457;
  assign new_new_n34090__ = ~new_new_n34088__ & new_new_n34089__;
  assign new_new_n34091__ = ys__n4457 & ys__n22727;
  assign new_new_n34092__ = ~new_new_n34090__ & ~new_new_n34091__;
  assign new_new_n34093__ = ~ys__n4451 & ~new_new_n34092__;
  assign new_new_n34094__ = ys__n4451 & ys__n22687;
  assign new_new_n34095__ = ~new_new_n34093__ & ~new_new_n34094__;
  assign new_new_n34096__ = new_new_n33934__ & ~new_new_n34095__;
  assign new_new_n34097__ = ys__n4458 & ys__n22576;
  assign new_new_n34098__ = ~new_new_n34096__ & ~new_new_n34097__;
  assign ys__n28422 = new_new_n33966__ & ~new_new_n34098__;
  assign new_new_n34100__ = ys__n22892 & new_new_n33921__;
  assign new_new_n34101__ = ys__n4454 & ys__n22836;
  assign new_new_n34102__ = ~new_new_n34100__ & ~new_new_n34101__;
  assign new_new_n34103__ = ~ys__n4452 & ~new_new_n34102__;
  assign new_new_n34104__ = ys__n4452 & ys__n22792;
  assign new_new_n34105__ = ~new_new_n34103__ & ~new_new_n34104__;
  assign new_new_n34106__ = ~ys__n4457 & ~new_new_n34105__;
  assign new_new_n34107__ = ys__n4457 & ys__n22729;
  assign new_new_n34108__ = ~new_new_n34106__ & ~new_new_n34107__;
  assign new_new_n34109__ = ~ys__n4451 & ~new_new_n34108__;
  assign new_new_n34110__ = ys__n4451 & ys__n22689;
  assign new_new_n34111__ = ~new_new_n34109__ & ~new_new_n34110__;
  assign new_new_n34112__ = new_new_n33934__ & ~new_new_n34111__;
  assign new_new_n34113__ = ys__n4458 & ys__n22578;
  assign new_new_n34114__ = ~new_new_n34112__ & ~new_new_n34113__;
  assign new_new_n34115__ = ~ys__n4461 & ~new_new_n34114__;
  assign new_new_n34116__ = ~ys__n4461 & ~new_new_n34115__;
  assign ys__n28423 = new_new_n33965__ & ~new_new_n34116__;
  assign new_new_n34118__ = ys__n22893 & new_new_n33921__;
  assign new_new_n34119__ = ys__n4454 & ys__n22838;
  assign new_new_n34120__ = ~new_new_n34118__ & ~new_new_n34119__;
  assign new_new_n34121__ = ~ys__n4452 & ~new_new_n34120__;
  assign new_new_n34122__ = ys__n4452 & ys__n22794;
  assign new_new_n34123__ = ~new_new_n34121__ & ~new_new_n34122__;
  assign new_new_n34124__ = ~ys__n4457 & ~new_new_n34123__;
  assign new_new_n34125__ = ys__n4457 & ys__n22731;
  assign new_new_n34126__ = ~new_new_n34124__ & ~new_new_n34125__;
  assign new_new_n34127__ = ~ys__n4449 & ~ys__n4451;
  assign new_new_n34128__ = ~new_new_n34126__ & new_new_n34127__;
  assign new_new_n34129__ = ys__n4449 & ys__n22640;
  assign new_new_n34130__ = ~new_new_n34128__ & ~new_new_n34129__;
  assign new_new_n34131__ = ~ys__n4458 & ~new_new_n34130__;
  assign new_new_n34132__ = ys__n4458 & ys__n22580;
  assign new_new_n34133__ = ~new_new_n34131__ & ~new_new_n34132__;
  assign new_new_n34134__ = ~ys__n4461 & ~new_new_n34133__;
  assign new_new_n34135__ = ~ys__n4461 & ~new_new_n34134__;
  assign new_new_n34136__ = ~ys__n4460 & ~new_new_n34135__;
  assign new_new_n34137__ = ~ys__n4460 & ~new_new_n34136__;
  assign new_new_n34138__ = ~ys__n4448 & ~new_new_n34137__;
  assign new_new_n34139__ = ys__n4448 & ys__n28424;
  assign ys__n28425 = new_new_n34138__ | new_new_n34139__;
  assign new_new_n34141__ = ys__n22894 & new_new_n33921__;
  assign new_new_n34142__ = ys__n4454 & ys__n22840;
  assign new_new_n34143__ = ~new_new_n34141__ & ~new_new_n34142__;
  assign new_new_n34144__ = new_new_n34089__ & ~new_new_n34143__;
  assign new_new_n34145__ = ys__n4457 & ys__n22733;
  assign new_new_n34146__ = ~new_new_n34144__ & ~new_new_n34145__;
  assign new_new_n34147__ = new_new_n34127__ & ~new_new_n34146__;
  assign new_new_n34148__ = ys__n4449 & ys__n22642;
  assign new_new_n34149__ = ~new_new_n34147__ & ~new_new_n34148__;
  assign new_new_n34150__ = ~ys__n4458 & ~new_new_n34149__;
  assign new_new_n34151__ = ys__n4458 & ys__n22582;
  assign new_new_n34152__ = ~new_new_n34150__ & ~new_new_n34151__;
  assign new_new_n34153__ = new_new_n33966__ & ~new_new_n34152__;
  assign new_new_n34154__ = ys__n4448 & ys__n28426;
  assign ys__n28427 = new_new_n34153__ | new_new_n34154__;
  assign new_new_n34156__ = ys__n22895 & new_new_n33921__;
  assign new_new_n34157__ = ys__n4454 & ys__n22842;
  assign new_new_n34158__ = ~new_new_n34156__ & ~new_new_n34157__;
  assign new_new_n34159__ = new_new_n34089__ & ~new_new_n34158__;
  assign new_new_n34160__ = ys__n4457 & ys__n22735;
  assign new_new_n34161__ = ~new_new_n34159__ & ~new_new_n34160__;
  assign new_new_n34162__ = new_new_n34127__ & ~new_new_n34161__;
  assign new_new_n34163__ = ys__n4449 & ys__n22644;
  assign new_new_n34164__ = ~new_new_n34162__ & ~new_new_n34163__;
  assign new_new_n34165__ = ~ys__n4458 & ~new_new_n34164__;
  assign new_new_n34166__ = ys__n4458 & ys__n22584;
  assign new_new_n34167__ = ~new_new_n34165__ & ~new_new_n34166__;
  assign new_new_n34168__ = new_new_n33966__ & ~new_new_n34167__;
  assign new_new_n34169__ = ys__n4448 & ys__n28428;
  assign ys__n28429 = new_new_n34168__ | new_new_n34169__;
  assign new_new_n34171__ = ys__n22896 & new_new_n33921__;
  assign new_new_n34172__ = ys__n4454 & ys__n22844;
  assign new_new_n34173__ = ~new_new_n34171__ & ~new_new_n34172__;
  assign new_new_n34174__ = new_new_n34089__ & ~new_new_n34173__;
  assign new_new_n34175__ = ys__n4457 & ys__n22737;
  assign new_new_n34176__ = ~new_new_n34174__ & ~new_new_n34175__;
  assign new_new_n34177__ = new_new_n34127__ & ~new_new_n34176__;
  assign new_new_n34178__ = ys__n4449 & ys__n22646;
  assign new_new_n34179__ = ~new_new_n34177__ & ~new_new_n34178__;
  assign new_new_n34180__ = ~ys__n4458 & ~new_new_n34179__;
  assign new_new_n34181__ = ys__n4458 & ys__n22586;
  assign new_new_n34182__ = ~new_new_n34180__ & ~new_new_n34181__;
  assign new_new_n34183__ = new_new_n33966__ & ~new_new_n34182__;
  assign new_new_n34184__ = ys__n4448 & ys__n28430;
  assign ys__n28431 = new_new_n34183__ | new_new_n34184__;
  assign new_new_n34186__ = ys__n22897 & new_new_n33921__;
  assign new_new_n34187__ = ys__n4454 & ys__n22846;
  assign new_new_n34188__ = ~new_new_n34186__ & ~new_new_n34187__;
  assign new_new_n34189__ = ~ys__n4452 & ~new_new_n34188__;
  assign new_new_n34190__ = ys__n4452 & ys__n22799;
  assign new_new_n34191__ = ~new_new_n34189__ & ~new_new_n34190__;
  assign new_new_n34192__ = ~ys__n4457 & ~new_new_n34191__;
  assign new_new_n34193__ = ys__n4457 & ys__n22739;
  assign new_new_n34194__ = ~new_new_n34192__ & ~new_new_n34193__;
  assign new_new_n34195__ = new_new_n34127__ & ~new_new_n34194__;
  assign new_new_n34196__ = ys__n4449 & ys__n22648;
  assign new_new_n34197__ = ~new_new_n34195__ & ~new_new_n34196__;
  assign new_new_n34198__ = ~ys__n4458 & ~new_new_n34197__;
  assign new_new_n34199__ = ys__n4458 & ys__n22588;
  assign new_new_n34200__ = ~new_new_n34198__ & ~new_new_n34199__;
  assign new_new_n34201__ = new_new_n33966__ & ~new_new_n34200__;
  assign new_new_n34202__ = ys__n4448 & ys__n28432;
  assign ys__n28433 = new_new_n34201__ | new_new_n34202__;
  assign new_new_n34204__ = ys__n22898 & new_new_n33921__;
  assign new_new_n34205__ = ys__n4454 & ys__n22848;
  assign new_new_n34206__ = ~new_new_n34204__ & ~new_new_n34205__;
  assign new_new_n34207__ = new_new_n34089__ & ~new_new_n34206__;
  assign new_new_n34208__ = ys__n4457 & ys__n22741;
  assign new_new_n34209__ = ~new_new_n34207__ & ~new_new_n34208__;
  assign new_new_n34210__ = new_new_n34127__ & ~new_new_n34209__;
  assign new_new_n34211__ = ys__n4449 & ys__n22650;
  assign new_new_n34212__ = ~new_new_n34210__ & ~new_new_n34211__;
  assign new_new_n34213__ = ~ys__n4458 & ~new_new_n34212__;
  assign new_new_n34214__ = ys__n4458 & ys__n22590;
  assign new_new_n34215__ = ~new_new_n34213__ & ~new_new_n34214__;
  assign new_new_n34216__ = new_new_n33966__ & ~new_new_n34215__;
  assign new_new_n34217__ = ys__n4448 & ys__n28434;
  assign ys__n28435 = new_new_n34216__ | new_new_n34217__;
  assign new_new_n34219__ = ys__n22899 & new_new_n33921__;
  assign new_new_n34220__ = ys__n4454 & ys__n22850;
  assign new_new_n34221__ = ~new_new_n34219__ & ~new_new_n34220__;
  assign new_new_n34222__ = new_new_n34089__ & ~new_new_n34221__;
  assign new_new_n34223__ = ys__n4457 & ys__n22743;
  assign new_new_n34224__ = ~new_new_n34222__ & ~new_new_n34223__;
  assign new_new_n34225__ = new_new_n34127__ & ~new_new_n34224__;
  assign new_new_n34226__ = ys__n4449 & ys__n22652;
  assign new_new_n34227__ = ~new_new_n34225__ & ~new_new_n34226__;
  assign new_new_n34228__ = ~ys__n4458 & ~new_new_n34227__;
  assign new_new_n34229__ = ys__n4458 & ys__n22592;
  assign new_new_n34230__ = ~new_new_n34228__ & ~new_new_n34229__;
  assign new_new_n34231__ = new_new_n33938__ & ~new_new_n34230__;
  assign new_new_n34232__ = ~ys__n4460 & ~new_new_n34231__;
  assign new_new_n34233__ = ~ys__n4448 & ~new_new_n34232__;
  assign new_new_n34234__ = ys__n4448 & ys__n28436;
  assign ys__n28437 = new_new_n34233__ | new_new_n34234__;
  assign new_new_n34236__ = ys__n22900 & new_new_n33921__;
  assign new_new_n34237__ = ys__n4454 & ys__n22852;
  assign new_new_n34238__ = ~new_new_n34236__ & ~new_new_n34237__;
  assign new_new_n34239__ = new_new_n34089__ & ~new_new_n34238__;
  assign new_new_n34240__ = ys__n4457 & ys__n22745;
  assign new_new_n34241__ = ~new_new_n34239__ & ~new_new_n34240__;
  assign new_new_n34242__ = new_new_n34127__ & ~new_new_n34241__;
  assign new_new_n34243__ = ys__n4449 & ys__n22654;
  assign new_new_n34244__ = ~new_new_n34242__ & ~new_new_n34243__;
  assign new_new_n34245__ = ~ys__n4458 & ~new_new_n34244__;
  assign new_new_n34246__ = ys__n4458 & ys__n22594;
  assign new_new_n34247__ = ~new_new_n34245__ & ~new_new_n34246__;
  assign new_new_n34248__ = new_new_n33938__ & ~new_new_n34247__;
  assign new_new_n34249__ = ~ys__n4460 & ~new_new_n34248__;
  assign new_new_n34250__ = ~ys__n4448 & ~new_new_n34249__;
  assign new_new_n34251__ = ys__n4448 & ys__n28438;
  assign ys__n28439 = new_new_n34250__ | new_new_n34251__;
  assign new_new_n34253__ = ys__n22901 & new_new_n33921__;
  assign new_new_n34254__ = ys__n4454 & ys__n22854;
  assign new_new_n34255__ = ~new_new_n34253__ & ~new_new_n34254__;
  assign new_new_n34256__ = new_new_n34089__ & ~new_new_n34255__;
  assign new_new_n34257__ = ys__n4457 & ys__n22747;
  assign new_new_n34258__ = ~new_new_n34256__ & ~new_new_n34257__;
  assign new_new_n34259__ = ~ys__n4458 & new_new_n34127__;
  assign new_new_n34260__ = ~new_new_n34258__ & new_new_n34259__;
  assign new_new_n34261__ = ys__n4458 & ys__n22596;
  assign new_new_n34262__ = ~new_new_n34260__ & ~new_new_n34261__;
  assign new_new_n34263__ = ~ys__n4461 & ~new_new_n34262__;
  assign new_new_n34264__ = ~ys__n4461 & ~new_new_n34263__;
  assign ys__n28440 = new_new_n33965__ & ~new_new_n34264__;
  assign new_new_n34266__ = ys__n22902 & new_new_n33921__;
  assign new_new_n34267__ = ys__n4454 & ys__n22856;
  assign new_new_n34268__ = ~new_new_n34266__ & ~new_new_n34267__;
  assign new_new_n34269__ = new_new_n34089__ & ~new_new_n34268__;
  assign new_new_n34270__ = ys__n4457 & ys__n22749;
  assign new_new_n34271__ = ~new_new_n34269__ & ~new_new_n34270__;
  assign new_new_n34272__ = new_new_n34259__ & ~new_new_n34271__;
  assign new_new_n34273__ = ys__n4458 & ys__n22598;
  assign new_new_n34274__ = ~new_new_n34272__ & ~new_new_n34273__;
  assign ys__n28441 = new_new_n33966__ & ~new_new_n34274__;
  assign new_new_n34276__ = ys__n22903 & new_new_n33921__;
  assign new_new_n34277__ = ys__n4454 & ys__n22858;
  assign new_new_n34278__ = ~new_new_n34276__ & ~new_new_n34277__;
  assign new_new_n34279__ = new_new_n34089__ & ~new_new_n34278__;
  assign new_new_n34280__ = ys__n4457 & ys__n22751;
  assign new_new_n34281__ = ~new_new_n34279__ & ~new_new_n34280__;
  assign new_new_n34282__ = new_new_n34259__ & ~new_new_n34281__;
  assign new_new_n34283__ = ys__n4458 & ys__n22600;
  assign new_new_n34284__ = ~new_new_n34282__ & ~new_new_n34283__;
  assign new_new_n34285__ = ~ys__n4461 & ~new_new_n34284__;
  assign new_new_n34286__ = ~ys__n4461 & ~new_new_n34285__;
  assign ys__n28442 = new_new_n33965__ & ~new_new_n34286__;
  assign new_new_n34288__ = ys__n22904 & new_new_n33921__;
  assign new_new_n34289__ = ys__n4454 & ys__n22860;
  assign new_new_n34290__ = ~new_new_n34288__ & ~new_new_n34289__;
  assign new_new_n34291__ = new_new_n34089__ & ~new_new_n34290__;
  assign new_new_n34292__ = ys__n4457 & ys__n22753;
  assign new_new_n34293__ = ~new_new_n34291__ & ~new_new_n34292__;
  assign new_new_n34294__ = new_new_n34259__ & ~new_new_n34293__;
  assign new_new_n34295__ = ys__n4458 & ys__n22602;
  assign new_new_n34296__ = ~new_new_n34294__ & ~new_new_n34295__;
  assign new_new_n34297__ = ~ys__n4461 & ~new_new_n34296__;
  assign new_new_n34298__ = ~ys__n4461 & ~new_new_n34297__;
  assign ys__n28443 = new_new_n33965__ & ~new_new_n34298__;
  assign new_new_n34300__ = ys__n22905 & new_new_n33921__;
  assign new_new_n34301__ = ys__n4454 & ys__n22862;
  assign new_new_n34302__ = ~new_new_n34300__ & ~new_new_n34301__;
  assign new_new_n34303__ = new_new_n34089__ & ~new_new_n34302__;
  assign new_new_n34304__ = ys__n4457 & ys__n22755;
  assign new_new_n34305__ = ~new_new_n34303__ & ~new_new_n34304__;
  assign new_new_n34306__ = new_new_n34259__ & ~new_new_n34305__;
  assign new_new_n34307__ = ys__n4458 & ys__n22604;
  assign new_new_n34308__ = ~new_new_n34306__ & ~new_new_n34307__;
  assign ys__n28444 = new_new_n33966__ & ~new_new_n34308__;
  assign new_new_n34310__ = ys__n22906 & new_new_n33921__;
  assign new_new_n34311__ = ys__n4454 & ys__n22864;
  assign new_new_n34312__ = ~new_new_n34310__ & ~new_new_n34311__;
  assign new_new_n34313__ = new_new_n34089__ & ~new_new_n34312__;
  assign new_new_n34314__ = ys__n4457 & ys__n22757;
  assign new_new_n34315__ = ~new_new_n34313__ & ~new_new_n34314__;
  assign new_new_n34316__ = new_new_n34259__ & ~new_new_n34315__;
  assign new_new_n34317__ = ys__n4458 & ys__n22606;
  assign new_new_n34318__ = ~new_new_n34316__ & ~new_new_n34317__;
  assign ys__n28445 = new_new_n33966__ & ~new_new_n34318__;
  assign new_new_n34320__ = ys__n22907 & new_new_n33921__;
  assign new_new_n34321__ = ys__n4454 & ys__n22866;
  assign new_new_n34322__ = ~new_new_n34320__ & ~new_new_n34321__;
  assign new_new_n34323__ = new_new_n34089__ & ~new_new_n34322__;
  assign new_new_n34324__ = ys__n4457 & ys__n22759;
  assign new_new_n34325__ = ~new_new_n34323__ & ~new_new_n34324__;
  assign new_new_n34326__ = new_new_n34259__ & ~new_new_n34325__;
  assign new_new_n34327__ = ys__n4458 & ys__n22608;
  assign new_new_n34328__ = ~new_new_n34326__ & ~new_new_n34327__;
  assign new_new_n34329__ = ~ys__n4461 & ~new_new_n34328__;
  assign new_new_n34330__ = ~ys__n4461 & ~new_new_n34329__;
  assign new_new_n34331__ = new_new_n33965__ & ~new_new_n34330__;
  assign new_new_n34332__ = ys__n4448 & ys__n28446;
  assign ys__n28447 = new_new_n34331__ | new_new_n34332__;
  assign new_new_n34334__ = ys__n22908 & new_new_n33921__;
  assign new_new_n34335__ = ys__n4454 & ys__n22868;
  assign new_new_n34336__ = ~new_new_n34334__ & ~new_new_n34335__;
  assign new_new_n34337__ = new_new_n34089__ & ~new_new_n34336__;
  assign new_new_n34338__ = ys__n4457 & ys__n22761;
  assign new_new_n34339__ = ~new_new_n34337__ & ~new_new_n34338__;
  assign new_new_n34340__ = new_new_n34259__ & ~new_new_n34339__;
  assign new_new_n34341__ = ys__n4458 & ys__n22610;
  assign new_new_n34342__ = ~new_new_n34340__ & ~new_new_n34341__;
  assign ys__n28448 = new_new_n33966__ & ~new_new_n34342__;
  assign new_new_n34344__ = ys__n22909 & new_new_n33921__;
  assign new_new_n34345__ = ys__n4454 & ys__n22870;
  assign new_new_n34346__ = ~new_new_n34344__ & ~new_new_n34345__;
  assign new_new_n34347__ = new_new_n34089__ & ~new_new_n34346__;
  assign new_new_n34348__ = ys__n4457 & ys__n22763;
  assign new_new_n34349__ = ~new_new_n34347__ & ~new_new_n34348__;
  assign new_new_n34350__ = new_new_n34259__ & ~new_new_n34349__;
  assign new_new_n34351__ = ys__n4458 & ys__n22612;
  assign new_new_n34352__ = ~new_new_n34350__ & ~new_new_n34351__;
  assign ys__n28449 = new_new_n33966__ & ~new_new_n34352__;
  assign new_new_n34354__ = ys__n22910 & new_new_n33921__;
  assign new_new_n34355__ = ys__n4454 & ys__n22872;
  assign new_new_n34356__ = ~new_new_n34354__ & ~new_new_n34355__;
  assign new_new_n34357__ = new_new_n34089__ & ~new_new_n34356__;
  assign new_new_n34358__ = ys__n4457 & ys__n22765;
  assign new_new_n34359__ = ~new_new_n34357__ & ~new_new_n34358__;
  assign new_new_n34360__ = new_new_n34259__ & ~new_new_n34359__;
  assign new_new_n34361__ = ys__n4458 & ys__n22614;
  assign new_new_n34362__ = ~new_new_n34360__ & ~new_new_n34361__;
  assign ys__n28450 = new_new_n33966__ & ~new_new_n34362__;
  assign new_new_n34364__ = ys__n22911 & new_new_n33921__;
  assign new_new_n34365__ = ys__n4454 & ys__n22874;
  assign new_new_n34366__ = ~new_new_n34364__ & ~new_new_n34365__;
  assign new_new_n34367__ = new_new_n34089__ & ~new_new_n34366__;
  assign new_new_n34368__ = ys__n4457 & ys__n22767;
  assign new_new_n34369__ = ~new_new_n34367__ & ~new_new_n34368__;
  assign new_new_n34370__ = new_new_n34259__ & ~new_new_n34369__;
  assign new_new_n34371__ = ys__n4458 & ys__n22616;
  assign new_new_n34372__ = ~new_new_n34370__ & ~new_new_n34371__;
  assign ys__n28451 = new_new_n33966__ & ~new_new_n34372__;
  assign new_new_n34374__ = ys__n22912 & new_new_n33921__;
  assign new_new_n34375__ = ys__n4454 & ys__n22876;
  assign new_new_n34376__ = ~new_new_n34374__ & ~new_new_n34375__;
  assign new_new_n34377__ = new_new_n34089__ & ~new_new_n34376__;
  assign new_new_n34378__ = ys__n4457 & ys__n22769;
  assign new_new_n34379__ = ~new_new_n34377__ & ~new_new_n34378__;
  assign new_new_n34380__ = new_new_n34259__ & ~new_new_n34379__;
  assign new_new_n34381__ = ys__n4458 & ys__n22618;
  assign new_new_n34382__ = ~new_new_n34380__ & ~new_new_n34381__;
  assign ys__n28452 = new_new_n33966__ & ~new_new_n34382__;
  assign new_new_n34384__ = ys__n22913 & new_new_n33921__;
  assign new_new_n34385__ = ys__n4454 & ys__n22878;
  assign new_new_n34386__ = ~new_new_n34384__ & ~new_new_n34385__;
  assign new_new_n34387__ = new_new_n34089__ & ~new_new_n34386__;
  assign new_new_n34388__ = ys__n4457 & ys__n22771;
  assign new_new_n34389__ = ~new_new_n34387__ & ~new_new_n34388__;
  assign new_new_n34390__ = new_new_n34127__ & ~new_new_n34389__;
  assign new_new_n34391__ = ys__n4449 & ys__n22668;
  assign new_new_n34392__ = ~new_new_n34390__ & ~new_new_n34391__;
  assign new_new_n34393__ = ~ys__n4458 & ~new_new_n34392__;
  assign new_new_n34394__ = ys__n4458 & ys__n22620;
  assign new_new_n34395__ = ~new_new_n34393__ & ~new_new_n34394__;
  assign new_new_n34396__ = new_new_n33966__ & ~new_new_n34395__;
  assign new_new_n34397__ = ys__n4448 & ys__n28453;
  assign ys__n28454 = new_new_n34396__ | new_new_n34397__;
  assign new_new_n34399__ = ys__n22914 & new_new_n33921__;
  assign new_new_n34400__ = ys__n4454 & ys__n22880;
  assign new_new_n34401__ = ~new_new_n34399__ & ~new_new_n34400__;
  assign new_new_n34402__ = new_new_n34089__ & ~new_new_n34401__;
  assign new_new_n34403__ = ys__n4457 & ys__n22773;
  assign new_new_n34404__ = ~new_new_n34402__ & ~new_new_n34403__;
  assign new_new_n34405__ = new_new_n34127__ & ~new_new_n34404__;
  assign new_new_n34406__ = ys__n4449 & ys__n22670;
  assign new_new_n34407__ = ~new_new_n34405__ & ~new_new_n34406__;
  assign new_new_n34408__ = ~ys__n4458 & ~new_new_n34407__;
  assign new_new_n34409__ = ys__n4458 & ys__n22622;
  assign new_new_n34410__ = ~new_new_n34408__ & ~new_new_n34409__;
  assign new_new_n34411__ = ~ys__n4461 & ~new_new_n34410__;
  assign new_new_n34412__ = ~ys__n4461 & ~new_new_n34411__;
  assign new_new_n34413__ = new_new_n33965__ & ~new_new_n34412__;
  assign new_new_n34414__ = ys__n4448 & ys__n28455;
  assign ys__n28456 = new_new_n34413__ | new_new_n34414__;
  assign new_new_n34416__ = ys__n22915 & new_new_n33921__;
  assign new_new_n34417__ = ys__n4454 & ys__n22882;
  assign new_new_n34418__ = ~new_new_n34416__ & ~new_new_n34417__;
  assign new_new_n34419__ = ~ys__n4452 & ~new_new_n34418__;
  assign new_new_n34420__ = ys__n4452 & ys__n22818;
  assign new_new_n34421__ = ~new_new_n34419__ & ~new_new_n34420__;
  assign new_new_n34422__ = ~ys__n4457 & ~new_new_n34421__;
  assign new_new_n34423__ = ys__n4457 & ys__n22775;
  assign new_new_n34424__ = ~new_new_n34422__ & ~new_new_n34423__;
  assign new_new_n34425__ = new_new_n34259__ & ~new_new_n34424__;
  assign new_new_n34426__ = ys__n4458 & ys__n22624;
  assign new_new_n34427__ = ~new_new_n34425__ & ~new_new_n34426__;
  assign new_new_n34428__ = new_new_n33966__ & ~new_new_n34427__;
  assign new_new_n34429__ = ys__n4448 & ys__n28457;
  assign ys__n28458 = new_new_n34428__ | new_new_n34429__;
  assign new_new_n34431__ = ys__n22916 & new_new_n33921__;
  assign new_new_n34432__ = ys__n4454 & ys__n22884;
  assign new_new_n34433__ = ~new_new_n34431__ & ~new_new_n34432__;
  assign new_new_n34434__ = ~ys__n4452 & ~new_new_n34433__;
  assign new_new_n34435__ = ys__n4452 & ys__n22820;
  assign new_new_n34436__ = ~new_new_n34434__ & ~new_new_n34435__;
  assign new_new_n34437__ = ~ys__n4457 & ~new_new_n34436__;
  assign new_new_n34438__ = ys__n4457 & ys__n22777;
  assign new_new_n34439__ = ~new_new_n34437__ & ~new_new_n34438__;
  assign new_new_n34440__ = new_new_n34127__ & ~new_new_n34439__;
  assign new_new_n34441__ = ys__n4449 & ys__n22673;
  assign new_new_n34442__ = ~new_new_n34440__ & ~new_new_n34441__;
  assign new_new_n34443__ = ~ys__n4458 & ~new_new_n34442__;
  assign new_new_n34444__ = ys__n4458 & ys__n22626;
  assign new_new_n34445__ = ~new_new_n34443__ & ~new_new_n34444__;
  assign new_new_n34446__ = new_new_n33966__ & ~new_new_n34445__;
  assign new_new_n34447__ = ys__n4448 & ys__n28459;
  assign ys__n28460 = new_new_n34446__ | new_new_n34447__;
  assign new_new_n34449__ = ~ys__n24256 & ~ys__n24260;
  assign new_new_n34450__ = ~ys__n28412 & ~new_new_n34449__;
  assign new_new_n34451__ = ys__n20053 & new_new_n34450__;
  assign new_new_n34452__ = ~ys__n33375 & ys__n18218;
  assign new_new_n34453__ = ~ys__n20053 & ~new_new_n34452__;
  assign new_new_n34454__ = ys__n28412 & ~new_new_n34449__;
  assign new_new_n34455__ = ~new_new_n34453__ & new_new_n34454__;
  assign ys__n28475 = new_new_n34451__ | new_new_n34455__;
  assign new_new_n34457__ = ~ys__n28243 & ys__n23483;
  assign new_new_n34458__ = ys__n22464 & ys__n28243;
  assign ys__n28476 = new_new_n34457__ | new_new_n34458__;
  assign new_new_n34460__ = ~ys__n28243 & ys__n23485;
  assign new_new_n34461__ = ys__n23548 & ys__n28243;
  assign ys__n28477 = new_new_n34460__ | new_new_n34461__;
  assign new_new_n34463__ = ~ys__n28243 & ys__n23487;
  assign new_new_n34464__ = ys__n23550 & ys__n28243;
  assign ys__n28478 = new_new_n34463__ | new_new_n34464__;
  assign new_new_n34466__ = ~ys__n28243 & ys__n23489;
  assign new_new_n34467__ = ys__n23552 & ys__n28243;
  assign ys__n28479 = new_new_n34466__ | new_new_n34467__;
  assign new_new_n34469__ = ~ys__n28243 & ys__n23491;
  assign new_new_n34470__ = ys__n23554 & ys__n28243;
  assign ys__n28480 = new_new_n34469__ | new_new_n34470__;
  assign new_new_n34472__ = ~ys__n28243 & ys__n23493;
  assign new_new_n34473__ = ys__n23556 & ys__n28243;
  assign ys__n28481 = new_new_n34472__ | new_new_n34473__;
  assign new_new_n34475__ = ~ys__n28243 & ys__n23495;
  assign new_new_n34476__ = ys__n23558 & ys__n28243;
  assign ys__n28482 = new_new_n34475__ | new_new_n34476__;
  assign new_new_n34478__ = ~ys__n28243 & ys__n23497;
  assign new_new_n34479__ = ys__n23560 & ys__n28243;
  assign ys__n28483 = new_new_n34478__ | new_new_n34479__;
  assign new_new_n34481__ = ~ys__n28243 & ys__n23499;
  assign new_new_n34482__ = ys__n23562 & ys__n28243;
  assign ys__n28484 = new_new_n34481__ | new_new_n34482__;
  assign new_new_n34484__ = ~ys__n28243 & ys__n23501;
  assign new_new_n34485__ = ys__n23564 & ys__n28243;
  assign ys__n28485 = new_new_n34484__ | new_new_n34485__;
  assign new_new_n34487__ = ~ys__n28243 & ys__n23503;
  assign new_new_n34488__ = ys__n23566 & ys__n28243;
  assign ys__n28486 = new_new_n34487__ | new_new_n34488__;
  assign new_new_n34490__ = ~ys__n28243 & ys__n23505;
  assign new_new_n34491__ = ys__n23568 & ys__n28243;
  assign ys__n28487 = new_new_n34490__ | new_new_n34491__;
  assign new_new_n34493__ = ~ys__n28243 & ys__n23507;
  assign new_new_n34494__ = ys__n23570 & ys__n28243;
  assign ys__n28488 = new_new_n34493__ | new_new_n34494__;
  assign new_new_n34496__ = ~ys__n28243 & ys__n23509;
  assign new_new_n34497__ = ys__n23572 & ys__n28243;
  assign ys__n28489 = new_new_n34496__ | new_new_n34497__;
  assign new_new_n34499__ = ~ys__n28243 & ys__n23511;
  assign new_new_n34500__ = ys__n23574 & ys__n28243;
  assign ys__n28490 = new_new_n34499__ | new_new_n34500__;
  assign new_new_n34502__ = ~ys__n28243 & ys__n23513;
  assign new_new_n34503__ = ys__n420 & ys__n28243;
  assign ys__n28491 = new_new_n34502__ | new_new_n34503__;
  assign new_new_n34505__ = ~ys__n28243 & ys__n23515;
  assign new_new_n34506__ = ys__n442 & ys__n28243;
  assign ys__n28492 = new_new_n34505__ | new_new_n34506__;
  assign new_new_n34508__ = ~ys__n28243 & ys__n23517;
  assign new_new_n34509__ = ys__n440 & ys__n28243;
  assign ys__n28493 = new_new_n34508__ | new_new_n34509__;
  assign new_new_n34511__ = ~ys__n28243 & ys__n23519;
  assign new_new_n34512__ = ys__n444 & ys__n28243;
  assign ys__n28494 = new_new_n34511__ | new_new_n34512__;
  assign new_new_n34514__ = ~ys__n28243 & ys__n23521;
  assign new_new_n34515__ = ys__n438 & ys__n28243;
  assign ys__n28495 = new_new_n34514__ | new_new_n34515__;
  assign new_new_n34517__ = ~ys__n28243 & ys__n23523;
  assign new_new_n34518__ = ys__n446 & ys__n28243;
  assign ys__n28496 = new_new_n34517__ | new_new_n34518__;
  assign new_new_n34520__ = ~ys__n28243 & ys__n23525;
  assign new_new_n34521__ = ys__n434 & ys__n28243;
  assign ys__n28497 = new_new_n34520__ | new_new_n34521__;
  assign new_new_n34523__ = ~ys__n28243 & ys__n23527;
  assign new_new_n34524__ = ys__n436 & ys__n28243;
  assign ys__n28498 = new_new_n34523__ | new_new_n34524__;
  assign new_new_n34526__ = ~ys__n28243 & ys__n23529;
  assign new_new_n34527__ = ys__n432 & ys__n28243;
  assign ys__n28499 = new_new_n34526__ | new_new_n34527__;
  assign new_new_n34529__ = ~ys__n28243 & ys__n23531;
  assign new_new_n34530__ = ys__n448 & ys__n28243;
  assign ys__n28500 = new_new_n34529__ | new_new_n34530__;
  assign new_new_n34532__ = ~ys__n28243 & ys__n23533;
  assign new_new_n34533__ = ys__n428 & ys__n28243;
  assign ys__n28501 = new_new_n34532__ | new_new_n34533__;
  assign new_new_n34535__ = ~ys__n28243 & ys__n23535;
  assign new_new_n34536__ = ys__n430 & ys__n28243;
  assign ys__n28502 = new_new_n34535__ | new_new_n34536__;
  assign new_new_n34538__ = ~ys__n28243 & ys__n23537;
  assign new_new_n34539__ = ys__n426 & ys__n28243;
  assign ys__n28503 = new_new_n34538__ | new_new_n34539__;
  assign new_new_n34541__ = ~ys__n28243 & ys__n23539;
  assign new_new_n34542__ = ys__n450 & ys__n28243;
  assign ys__n28504 = new_new_n34541__ | new_new_n34542__;
  assign new_new_n34544__ = ~ys__n28243 & ys__n23541;
  assign new_new_n34545__ = ys__n424 & ys__n28243;
  assign ys__n28505 = new_new_n34544__ | new_new_n34545__;
  assign new_new_n34547__ = ~ys__n28243 & ys__n23543;
  assign new_new_n34548__ = ys__n422 & ys__n28243;
  assign ys__n28506 = new_new_n34547__ | new_new_n34548__;
  assign new_new_n34550__ = ys__n47661 & new_new_n11634__;
  assign new_new_n34551__ = ys__n22822 & new_new_n11175__;
  assign new_new_n34552__ = ~new_new_n11180__ & new_new_n34551__;
  assign new_new_n34553__ = ~new_new_n11186__ & new_new_n34552__;
  assign new_new_n34554__ = ys__n23480 & new_new_n11186__;
  assign new_new_n34555__ = ~new_new_n34553__ & ~new_new_n34554__;
  assign new_new_n34556__ = ~new_new_n11270__ & ~new_new_n34555__;
  assign new_new_n34557__ = ys__n23480 & new_new_n11270__;
  assign new_new_n34558__ = ~new_new_n34556__ & ~new_new_n34557__;
  assign new_new_n34559__ = new_new_n11324__ & ~new_new_n11343__;
  assign new_new_n34560__ = ~new_new_n34558__ & new_new_n34559__;
  assign new_new_n34561__ = ys__n23480 & new_new_n11343__;
  assign new_new_n34562__ = ~new_new_n34560__ & ~new_new_n34561__;
  assign new_new_n34563__ = new_new_n11629__ & ~new_new_n34562__;
  assign new_new_n34564__ = ~new_new_n34550__ & ~new_new_n34563__;
  assign new_new_n34565__ = new_new_n11640__ & ~new_new_n34564__;
  assign new_new_n34566__ = ys__n47661 & new_new_n11644__;
  assign new_new_n34567__ = new_new_n11642__ & ~new_new_n34562__;
  assign new_new_n34568__ = ~new_new_n34566__ & ~new_new_n34567__;
  assign new_new_n34569__ = new_new_n11650__ & ~new_new_n34568__;
  assign ys__n28510 = new_new_n34565__ | new_new_n34569__;
  assign new_new_n34571__ = ys__n47662 & new_new_n11634__;
  assign new_new_n34572__ = ys__n22824 & ~new_new_n11180__;
  assign new_new_n34573__ = new_new_n11175__ & new_new_n34572__;
  assign new_new_n34574__ = ~new_new_n16277__ & ~new_new_n34573__;
  assign new_new_n34575__ = ~new_new_n11186__ & ~new_new_n34574__;
  assign new_new_n34576__ = ys__n22464 & new_new_n11186__;
  assign new_new_n34577__ = ~new_new_n34575__ & ~new_new_n34576__;
  assign new_new_n34578__ = ~new_new_n11270__ & ~new_new_n34577__;
  assign new_new_n34579__ = new_new_n11270__ & ys__n23483;
  assign new_new_n34580__ = ~new_new_n34578__ & ~new_new_n34579__;
  assign new_new_n34581__ = new_new_n34559__ & ~new_new_n34580__;
  assign new_new_n34582__ = ~ys__n22464 & new_new_n11389__;
  assign new_new_n34583__ = ys__n22464 & ~new_new_n11389__;
  assign new_new_n34584__ = ~new_new_n34582__ & ~new_new_n34583__;
  assign new_new_n34585__ = new_new_n11343__ & ~new_new_n34584__;
  assign new_new_n34586__ = ~new_new_n34581__ & ~new_new_n34585__;
  assign new_new_n34587__ = new_new_n11629__ & ~new_new_n34586__;
  assign new_new_n34588__ = ~new_new_n34571__ & ~new_new_n34587__;
  assign new_new_n34589__ = new_new_n11640__ & ~new_new_n34588__;
  assign new_new_n34590__ = ys__n47662 & new_new_n11644__;
  assign new_new_n34591__ = new_new_n11642__ & ~new_new_n34586__;
  assign new_new_n34592__ = ~new_new_n34590__ & ~new_new_n34591__;
  assign new_new_n34593__ = new_new_n11650__ & ~new_new_n34592__;
  assign ys__n28513 = new_new_n34589__ | new_new_n34593__;
  assign new_new_n34595__ = ys__n47664 & new_new_n11634__;
  assign new_new_n34596__ = ys__n22828 & ~new_new_n11180__;
  assign new_new_n34597__ = new_new_n11175__ & new_new_n34596__;
  assign new_new_n34598__ = ~new_new_n16289__ & ~new_new_n34597__;
  assign new_new_n34599__ = ~new_new_n11186__ & ~new_new_n34598__;
  assign new_new_n34600__ = ys__n23550 & new_new_n11186__;
  assign new_new_n34601__ = ~new_new_n34599__ & ~new_new_n34600__;
  assign new_new_n34602__ = ~new_new_n11270__ & ~new_new_n34601__;
  assign new_new_n34603__ = new_new_n11270__ & ys__n23487;
  assign new_new_n34604__ = ~new_new_n34602__ & ~new_new_n34603__;
  assign new_new_n34605__ = new_new_n11324__ & ~new_new_n34604__;
  assign new_new_n34606__ = ys__n526 & ~new_new_n11324__;
  assign new_new_n34607__ = ~new_new_n34605__ & ~new_new_n34606__;
  assign new_new_n34608__ = ~new_new_n11343__ & ~new_new_n34607__;
  assign new_new_n34609__ = ~new_new_n11372__ & new_new_n11390__;
  assign new_new_n34610__ = ~new_new_n11394__ & ~new_new_n34609__;
  assign new_new_n34611__ = new_new_n11383__ & ~new_new_n34610__;
  assign new_new_n34612__ = ~new_new_n11383__ & new_new_n34610__;
  assign new_new_n34613__ = ~new_new_n34611__ & ~new_new_n34612__;
  assign new_new_n34614__ = new_new_n11343__ & ~new_new_n34613__;
  assign new_new_n34615__ = ~new_new_n34608__ & ~new_new_n34614__;
  assign new_new_n34616__ = new_new_n11629__ & ~new_new_n34615__;
  assign new_new_n34617__ = ~new_new_n34595__ & ~new_new_n34616__;
  assign new_new_n34618__ = new_new_n11640__ & ~new_new_n34617__;
  assign new_new_n34619__ = ys__n47664 & new_new_n11644__;
  assign new_new_n34620__ = new_new_n11642__ & ~new_new_n34615__;
  assign new_new_n34621__ = ~new_new_n34619__ & ~new_new_n34620__;
  assign new_new_n34622__ = new_new_n11650__ & ~new_new_n34621__;
  assign ys__n28518 = new_new_n34618__ | new_new_n34622__;
  assign new_new_n34624__ = ys__n47671 & new_new_n11634__;
  assign new_new_n34625__ = ys__n22842 & ~new_new_n11180__;
  assign new_new_n34626__ = new_new_n11175__ & new_new_n34625__;
  assign new_new_n34627__ = ~new_new_n16331__ & ~new_new_n34626__;
  assign new_new_n34628__ = ~new_new_n11186__ & ~new_new_n34627__;
  assign new_new_n34629__ = ys__n23564 & new_new_n11186__;
  assign new_new_n34630__ = ~new_new_n34628__ & ~new_new_n34629__;
  assign new_new_n34631__ = ~new_new_n11270__ & ~new_new_n34630__;
  assign new_new_n34632__ = new_new_n11270__ & ys__n23501;
  assign new_new_n34633__ = ~new_new_n34631__ & ~new_new_n34632__;
  assign new_new_n34634__ = new_new_n11324__ & ~new_new_n34633__;
  assign new_new_n34635__ = ys__n518 & ~new_new_n11324__;
  assign new_new_n34636__ = ~new_new_n34634__ & ~new_new_n34635__;
  assign new_new_n34637__ = ~new_new_n11343__ & ~new_new_n34636__;
  assign new_new_n34638__ = ~new_new_n11456__ & new_new_n11536__;
  assign new_new_n34639__ = new_new_n11543__ & ~new_new_n34638__;
  assign new_new_n34640__ = new_new_n11514__ & ~new_new_n34639__;
  assign new_new_n34641__ = ~new_new_n11514__ & new_new_n34639__;
  assign new_new_n34642__ = ~new_new_n34640__ & ~new_new_n34641__;
  assign new_new_n34643__ = new_new_n11343__ & ~new_new_n34642__;
  assign new_new_n34644__ = ~new_new_n34637__ & ~new_new_n34643__;
  assign new_new_n34645__ = new_new_n11629__ & ~new_new_n34644__;
  assign new_new_n34646__ = ~new_new_n34624__ & ~new_new_n34645__;
  assign new_new_n34647__ = new_new_n11640__ & ~new_new_n34646__;
  assign new_new_n34648__ = ys__n47671 & new_new_n11644__;
  assign new_new_n34649__ = new_new_n11642__ & ~new_new_n34644__;
  assign new_new_n34650__ = ~new_new_n34648__ & ~new_new_n34649__;
  assign new_new_n34651__ = new_new_n11650__ & ~new_new_n34650__;
  assign ys__n28533 = new_new_n34647__ | new_new_n34651__;
  assign new_new_n34653__ = ys__n47672 & new_new_n11634__;
  assign new_new_n34654__ = ys__n22844 & ~new_new_n11180__;
  assign new_new_n34655__ = new_new_n11175__ & new_new_n34654__;
  assign new_new_n34656__ = ~new_new_n16337__ & ~new_new_n34655__;
  assign new_new_n34657__ = ~new_new_n11186__ & ~new_new_n34656__;
  assign new_new_n34658__ = ys__n23566 & new_new_n11186__;
  assign new_new_n34659__ = ~new_new_n34657__ & ~new_new_n34658__;
  assign new_new_n34660__ = ~new_new_n11270__ & ~new_new_n34659__;
  assign new_new_n34661__ = new_new_n11270__ & ys__n23503;
  assign new_new_n34662__ = ~new_new_n34660__ & ~new_new_n34661__;
  assign new_new_n34663__ = new_new_n11324__ & ~new_new_n34662__;
  assign new_new_n34664__ = ys__n548 & ~new_new_n11324__;
  assign new_new_n34665__ = ~new_new_n34663__ & ~new_new_n34664__;
  assign new_new_n34666__ = ~new_new_n11343__ & ~new_new_n34665__;
  assign new_new_n34667__ = ~new_new_n11514__ & ~new_new_n34639__;
  assign new_new_n34668__ = ~new_new_n11546__ & ~new_new_n34667__;
  assign new_new_n34669__ = new_new_n11504__ & ~new_new_n34668__;
  assign new_new_n34670__ = ~new_new_n11504__ & new_new_n34668__;
  assign new_new_n34671__ = ~new_new_n34669__ & ~new_new_n34670__;
  assign new_new_n34672__ = new_new_n11343__ & ~new_new_n34671__;
  assign new_new_n34673__ = ~new_new_n34666__ & ~new_new_n34672__;
  assign new_new_n34674__ = new_new_n11629__ & ~new_new_n34673__;
  assign new_new_n34675__ = ~new_new_n34653__ & ~new_new_n34674__;
  assign new_new_n34676__ = new_new_n11640__ & ~new_new_n34675__;
  assign new_new_n34677__ = ys__n47672 & new_new_n11644__;
  assign new_new_n34678__ = new_new_n11642__ & ~new_new_n34673__;
  assign new_new_n34679__ = ~new_new_n34677__ & ~new_new_n34678__;
  assign new_new_n34680__ = new_new_n11650__ & ~new_new_n34679__;
  assign ys__n28536 = new_new_n34676__ | new_new_n34680__;
  assign new_new_n34682__ = ys__n47673 & new_new_n11634__;
  assign new_new_n34683__ = ys__n22846 & ~new_new_n11180__;
  assign new_new_n34684__ = new_new_n11175__ & new_new_n34683__;
  assign new_new_n34685__ = ~new_new_n16343__ & ~new_new_n34684__;
  assign new_new_n34686__ = ~new_new_n11186__ & ~new_new_n34685__;
  assign new_new_n34687__ = ys__n23568 & new_new_n11186__;
  assign new_new_n34688__ = ~new_new_n34686__ & ~new_new_n34687__;
  assign new_new_n34689__ = ~new_new_n11270__ & ~new_new_n34688__;
  assign new_new_n34690__ = new_new_n11270__ & ys__n23505;
  assign new_new_n34691__ = ~new_new_n34689__ & ~new_new_n34690__;
  assign new_new_n34692__ = new_new_n11324__ & ~new_new_n34691__;
  assign new_new_n34693__ = ys__n550 & ~new_new_n11324__;
  assign new_new_n34694__ = ~new_new_n34692__ & ~new_new_n34693__;
  assign new_new_n34695__ = ~new_new_n11343__ & ~new_new_n34694__;
  assign new_new_n34696__ = ~new_new_n11456__ & new_new_n11537__;
  assign new_new_n34697__ = new_new_n11549__ & ~new_new_n34696__;
  assign new_new_n34698__ = new_new_n11493__ & ~new_new_n34697__;
  assign new_new_n34699__ = ~new_new_n11493__ & new_new_n34697__;
  assign new_new_n34700__ = ~new_new_n34698__ & ~new_new_n34699__;
  assign new_new_n34701__ = new_new_n11343__ & ~new_new_n34700__;
  assign new_new_n34702__ = ~new_new_n34695__ & ~new_new_n34701__;
  assign new_new_n34703__ = new_new_n11629__ & ~new_new_n34702__;
  assign new_new_n34704__ = ~new_new_n34682__ & ~new_new_n34703__;
  assign new_new_n34705__ = new_new_n11640__ & ~new_new_n34704__;
  assign new_new_n34706__ = ys__n47673 & new_new_n11644__;
  assign new_new_n34707__ = new_new_n11642__ & ~new_new_n34702__;
  assign new_new_n34708__ = ~new_new_n34706__ & ~new_new_n34707__;
  assign new_new_n34709__ = new_new_n11650__ & ~new_new_n34708__;
  assign ys__n28539 = new_new_n34705__ | new_new_n34709__;
  assign new_new_n34711__ = ys__n47674 & new_new_n11634__;
  assign new_new_n34712__ = ys__n22848 & ~new_new_n11180__;
  assign new_new_n34713__ = new_new_n11175__ & new_new_n34712__;
  assign new_new_n34714__ = ~new_new_n16349__ & ~new_new_n34713__;
  assign new_new_n34715__ = ~new_new_n11186__ & ~new_new_n34714__;
  assign new_new_n34716__ = ys__n23570 & new_new_n11186__;
  assign new_new_n34717__ = ~new_new_n34715__ & ~new_new_n34716__;
  assign new_new_n34718__ = ~new_new_n11270__ & ~new_new_n34717__;
  assign new_new_n34719__ = new_new_n11270__ & ys__n23507;
  assign new_new_n34720__ = ~new_new_n34718__ & ~new_new_n34719__;
  assign new_new_n34721__ = new_new_n11324__ & ~new_new_n34720__;
  assign new_new_n34722__ = ys__n640 & ~new_new_n11324__;
  assign new_new_n34723__ = ~new_new_n34721__ & ~new_new_n34722__;
  assign new_new_n34724__ = ~new_new_n11343__ & ~new_new_n34723__;
  assign new_new_n34725__ = ~new_new_n11493__ & ~new_new_n34697__;
  assign new_new_n34726__ = ~new_new_n11552__ & ~new_new_n34725__;
  assign new_new_n34727__ = new_new_n11484__ & ~new_new_n34726__;
  assign new_new_n34728__ = ~new_new_n11484__ & new_new_n34726__;
  assign new_new_n34729__ = ~new_new_n34727__ & ~new_new_n34728__;
  assign new_new_n34730__ = new_new_n11343__ & ~new_new_n34729__;
  assign new_new_n34731__ = ~new_new_n34724__ & ~new_new_n34730__;
  assign new_new_n34732__ = new_new_n11629__ & ~new_new_n34731__;
  assign new_new_n34733__ = ~new_new_n34711__ & ~new_new_n34732__;
  assign new_new_n34734__ = new_new_n11640__ & ~new_new_n34733__;
  assign new_new_n34735__ = ys__n47674 & new_new_n11644__;
  assign new_new_n34736__ = new_new_n11642__ & ~new_new_n34731__;
  assign new_new_n34737__ = ~new_new_n34735__ & ~new_new_n34736__;
  assign new_new_n34738__ = new_new_n11650__ & ~new_new_n34737__;
  assign ys__n28542 = new_new_n34734__ | new_new_n34738__;
  assign new_new_n34740__ = ys__n47675 & new_new_n11634__;
  assign new_new_n34741__ = ys__n22850 & ~new_new_n11180__;
  assign new_new_n34742__ = new_new_n11175__ & new_new_n34741__;
  assign new_new_n34743__ = ~new_new_n16355__ & ~new_new_n34742__;
  assign new_new_n34744__ = ~new_new_n11186__ & ~new_new_n34743__;
  assign new_new_n34745__ = ys__n23572 & new_new_n11186__;
  assign new_new_n34746__ = ~new_new_n34744__ & ~new_new_n34745__;
  assign new_new_n34747__ = ~new_new_n11270__ & ~new_new_n34746__;
  assign new_new_n34748__ = new_new_n11270__ & ys__n23509;
  assign new_new_n34749__ = ~new_new_n34747__ & ~new_new_n34748__;
  assign new_new_n34750__ = new_new_n11324__ & ~new_new_n34749__;
  assign new_new_n34751__ = ys__n638 & ~new_new_n11324__;
  assign new_new_n34752__ = ~new_new_n34750__ & ~new_new_n34751__;
  assign new_new_n34753__ = ~new_new_n11343__ & ~new_new_n34752__;
  assign new_new_n34754__ = new_new_n11494__ & ~new_new_n34697__;
  assign new_new_n34755__ = new_new_n11554__ & ~new_new_n34754__;
  assign new_new_n34756__ = new_new_n11474__ & ~new_new_n34755__;
  assign new_new_n34757__ = ~new_new_n11474__ & new_new_n34755__;
  assign new_new_n34758__ = ~new_new_n34756__ & ~new_new_n34757__;
  assign new_new_n34759__ = new_new_n11343__ & ~new_new_n34758__;
  assign new_new_n34760__ = ~new_new_n34753__ & ~new_new_n34759__;
  assign new_new_n34761__ = new_new_n11629__ & ~new_new_n34760__;
  assign new_new_n34762__ = ~new_new_n34740__ & ~new_new_n34761__;
  assign new_new_n34763__ = new_new_n11640__ & ~new_new_n34762__;
  assign new_new_n34764__ = ys__n47675 & new_new_n11644__;
  assign new_new_n34765__ = new_new_n11642__ & ~new_new_n34760__;
  assign new_new_n34766__ = ~new_new_n34764__ & ~new_new_n34765__;
  assign new_new_n34767__ = new_new_n11650__ & ~new_new_n34766__;
  assign ys__n28545 = new_new_n34763__ | new_new_n34767__;
  assign new_new_n34769__ = ys__n47676 & new_new_n11634__;
  assign new_new_n34770__ = ys__n22852 & ~new_new_n11180__;
  assign new_new_n34771__ = new_new_n11175__ & new_new_n34770__;
  assign new_new_n34772__ = ~new_new_n16361__ & ~new_new_n34771__;
  assign new_new_n34773__ = ~new_new_n11186__ & ~new_new_n34772__;
  assign new_new_n34774__ = ys__n23574 & new_new_n11186__;
  assign new_new_n34775__ = ~new_new_n34773__ & ~new_new_n34774__;
  assign new_new_n34776__ = ~new_new_n11270__ & ~new_new_n34775__;
  assign new_new_n34777__ = new_new_n11270__ & ys__n23511;
  assign new_new_n34778__ = ~new_new_n34776__ & ~new_new_n34777__;
  assign new_new_n34779__ = new_new_n11324__ & ~new_new_n34778__;
  assign new_new_n34780__ = ys__n636 & ~new_new_n11324__;
  assign new_new_n34781__ = ~new_new_n34779__ & ~new_new_n34780__;
  assign new_new_n34782__ = ~new_new_n11343__ & ~new_new_n34781__;
  assign new_new_n34783__ = ~new_new_n11474__ & ~new_new_n34755__;
  assign new_new_n34784__ = ~new_new_n11557__ & ~new_new_n34783__;
  assign new_new_n34785__ = new_new_n11465__ & ~new_new_n34784__;
  assign new_new_n34786__ = ~new_new_n11465__ & new_new_n34784__;
  assign new_new_n34787__ = ~new_new_n34785__ & ~new_new_n34786__;
  assign new_new_n34788__ = new_new_n11343__ & ~new_new_n34787__;
  assign new_new_n34789__ = ~new_new_n34782__ & ~new_new_n34788__;
  assign new_new_n34790__ = new_new_n11629__ & ~new_new_n34789__;
  assign new_new_n34791__ = ~new_new_n34769__ & ~new_new_n34790__;
  assign new_new_n34792__ = new_new_n11640__ & ~new_new_n34791__;
  assign new_new_n34793__ = ys__n47676 & new_new_n11644__;
  assign new_new_n34794__ = new_new_n11642__ & ~new_new_n34789__;
  assign new_new_n34795__ = ~new_new_n34793__ & ~new_new_n34794__;
  assign new_new_n34796__ = new_new_n11650__ & ~new_new_n34795__;
  assign ys__n28548 = new_new_n34792__ | new_new_n34796__;
  assign new_new_n34798__ = ys__n47677 & new_new_n11634__;
  assign new_new_n34799__ = ys__n22854 & ~new_new_n11180__;
  assign new_new_n34800__ = new_new_n11175__ & new_new_n34799__;
  assign new_new_n34801__ = ~new_new_n16367__ & ~new_new_n34800__;
  assign new_new_n34802__ = ~new_new_n11186__ & ~new_new_n34801__;
  assign new_new_n34803__ = ys__n420 & new_new_n11186__;
  assign new_new_n34804__ = ~new_new_n34802__ & ~new_new_n34803__;
  assign new_new_n34805__ = ~new_new_n11270__ & ~new_new_n34804__;
  assign new_new_n34806__ = new_new_n11270__ & ys__n23513;
  assign new_new_n34807__ = ~new_new_n34805__ & ~new_new_n34806__;
  assign new_new_n34808__ = new_new_n11324__ & ~new_new_n34807__;
  assign new_new_n34809__ = ys__n634 & ~new_new_n11324__;
  assign new_new_n34810__ = ~new_new_n34808__ & ~new_new_n34809__;
  assign new_new_n34811__ = ~new_new_n11343__ & ~new_new_n34810__;
  assign new_new_n34812__ = new_new_n11361__ & ~new_new_n11562__;
  assign new_new_n34813__ = ~new_new_n11361__ & new_new_n11562__;
  assign new_new_n34814__ = ~new_new_n34812__ & ~new_new_n34813__;
  assign new_new_n34815__ = new_new_n11343__ & ~new_new_n34814__;
  assign new_new_n34816__ = ~new_new_n34811__ & ~new_new_n34815__;
  assign new_new_n34817__ = new_new_n11629__ & ~new_new_n34816__;
  assign new_new_n34818__ = ~new_new_n34798__ & ~new_new_n34817__;
  assign new_new_n34819__ = new_new_n11640__ & ~new_new_n34818__;
  assign new_new_n34820__ = ys__n47677 & new_new_n11644__;
  assign new_new_n34821__ = new_new_n11642__ & ~new_new_n34816__;
  assign new_new_n34822__ = ~new_new_n34820__ & ~new_new_n34821__;
  assign new_new_n34823__ = new_new_n11650__ & ~new_new_n34822__;
  assign ys__n28551 = new_new_n34819__ | new_new_n34823__;
  assign new_new_n34825__ = ys__n47678 & new_new_n11634__;
  assign new_new_n34826__ = ys__n22856 & ~new_new_n11180__;
  assign new_new_n34827__ = new_new_n11175__ & new_new_n34826__;
  assign new_new_n34828__ = ~new_new_n16373__ & ~new_new_n34827__;
  assign new_new_n34829__ = ~new_new_n11186__ & ~new_new_n34828__;
  assign new_new_n34830__ = ys__n442 & new_new_n11186__;
  assign new_new_n34831__ = ~new_new_n34829__ & ~new_new_n34830__;
  assign new_new_n34832__ = ~new_new_n11270__ & ~new_new_n34831__;
  assign new_new_n34833__ = new_new_n11270__ & ys__n23515;
  assign new_new_n34834__ = ~new_new_n34832__ & ~new_new_n34833__;
  assign new_new_n34835__ = new_new_n11324__ & ~new_new_n34834__;
  assign new_new_n34836__ = ys__n642 & ~new_new_n11324__;
  assign new_new_n34837__ = ~new_new_n34835__ & ~new_new_n34836__;
  assign new_new_n34838__ = ~new_new_n11343__ & ~new_new_n34837__;
  assign new_new_n34839__ = ys__n442 & ~new_new_n11569__;
  assign new_new_n34840__ = ~ys__n442 & new_new_n11603__;
  assign new_new_n34841__ = ~ys__n442 & new_new_n11619__;
  assign new_new_n34842__ = ~new_new_n34840__ & ~new_new_n34841__;
  assign new_new_n34843__ = ~new_new_n34839__ & new_new_n34842__;
  assign new_new_n34844__ = new_new_n11625__ & ~new_new_n34843__;
  assign new_new_n34845__ = ~new_new_n34838__ & ~new_new_n34844__;
  assign new_new_n34846__ = new_new_n11629__ & ~new_new_n34845__;
  assign new_new_n34847__ = ~new_new_n34825__ & ~new_new_n34846__;
  assign new_new_n34848__ = new_new_n11640__ & ~new_new_n34847__;
  assign new_new_n34849__ = ys__n47678 & new_new_n11644__;
  assign new_new_n34850__ = new_new_n11642__ & ~new_new_n34845__;
  assign new_new_n34851__ = ~new_new_n34849__ & ~new_new_n34850__;
  assign new_new_n34852__ = new_new_n11650__ & ~new_new_n34851__;
  assign ys__n28554 = new_new_n34848__ | new_new_n34852__;
  assign new_new_n34854__ = ys__n47679 & new_new_n11634__;
  assign new_new_n34855__ = ys__n22858 & ~new_new_n11180__;
  assign new_new_n34856__ = new_new_n11175__ & new_new_n34855__;
  assign new_new_n34857__ = ~new_new_n16379__ & ~new_new_n34856__;
  assign new_new_n34858__ = ~new_new_n11186__ & ~new_new_n34857__;
  assign new_new_n34859__ = ys__n440 & new_new_n11186__;
  assign new_new_n34860__ = ~new_new_n34858__ & ~new_new_n34859__;
  assign new_new_n34861__ = ~new_new_n11270__ & ~new_new_n34860__;
  assign new_new_n34862__ = new_new_n11270__ & ys__n23517;
  assign new_new_n34863__ = ~new_new_n34861__ & ~new_new_n34862__;
  assign new_new_n34864__ = new_new_n11324__ & ~new_new_n34863__;
  assign new_new_n34865__ = ys__n514 & ~ys__n28243;
  assign new_new_n34866__ = ys__n28243 & ys__n28632;
  assign new_new_n34867__ = ~new_new_n34865__ & ~new_new_n34866__;
  assign new_new_n34868__ = ~new_new_n11324__ & ~new_new_n34867__;
  assign new_new_n34869__ = ~new_new_n34864__ & ~new_new_n34868__;
  assign new_new_n34870__ = ~new_new_n11343__ & ~new_new_n34869__;
  assign new_new_n34871__ = ys__n440 & ~new_new_n11569__;
  assign new_new_n34872__ = ~ys__n440 & ~ys__n442;
  assign new_new_n34873__ = ~new_new_n11608__ & ~new_new_n34872__;
  assign new_new_n34874__ = new_new_n11603__ & ~new_new_n34873__;
  assign new_new_n34875__ = ys__n440 & ~ys__n442;
  assign new_new_n34876__ = ~new_new_n11571__ & ~new_new_n34875__;
  assign new_new_n34877__ = new_new_n11619__ & ~new_new_n34876__;
  assign new_new_n34878__ = ~new_new_n34874__ & ~new_new_n34877__;
  assign new_new_n34879__ = ~new_new_n34871__ & new_new_n34878__;
  assign new_new_n34880__ = new_new_n11625__ & ~new_new_n34879__;
  assign new_new_n34881__ = ~new_new_n34870__ & ~new_new_n34880__;
  assign new_new_n34882__ = new_new_n11629__ & ~new_new_n34881__;
  assign new_new_n34883__ = ~new_new_n34854__ & ~new_new_n34882__;
  assign new_new_n34884__ = new_new_n11640__ & ~new_new_n34883__;
  assign new_new_n34885__ = ys__n47679 & new_new_n11644__;
  assign new_new_n34886__ = new_new_n11642__ & ~new_new_n34881__;
  assign new_new_n34887__ = ~new_new_n34885__ & ~new_new_n34886__;
  assign new_new_n34888__ = new_new_n11650__ & ~new_new_n34887__;
  assign ys__n28557 = new_new_n34884__ | new_new_n34888__;
  assign new_new_n34890__ = ys__n47680 & new_new_n11634__;
  assign new_new_n34891__ = ys__n22860 & ~new_new_n11180__;
  assign new_new_n34892__ = new_new_n11175__ & new_new_n34891__;
  assign new_new_n34893__ = ~new_new_n16385__ & ~new_new_n34892__;
  assign new_new_n34894__ = ~new_new_n11186__ & ~new_new_n34893__;
  assign new_new_n34895__ = ys__n444 & new_new_n11186__;
  assign new_new_n34896__ = ~new_new_n34894__ & ~new_new_n34895__;
  assign new_new_n34897__ = ~new_new_n11270__ & ~new_new_n34896__;
  assign new_new_n34898__ = new_new_n11270__ & ys__n23519;
  assign new_new_n34899__ = ~new_new_n34897__ & ~new_new_n34898__;
  assign new_new_n34900__ = new_new_n11324__ & ~new_new_n34899__;
  assign new_new_n34901__ = ys__n2024 & ~ys__n28243;
  assign new_new_n34902__ = ys__n28243 & ys__n28633;
  assign new_new_n34903__ = ~new_new_n34901__ & ~new_new_n34902__;
  assign new_new_n34904__ = ~new_new_n11324__ & ~new_new_n34903__;
  assign new_new_n34905__ = ~new_new_n34900__ & ~new_new_n34904__;
  assign new_new_n34906__ = ~new_new_n11343__ & ~new_new_n34905__;
  assign new_new_n34907__ = ys__n444 & ~new_new_n11569__;
  assign new_new_n34908__ = ys__n444 & ~new_new_n11572__;
  assign new_new_n34909__ = ~ys__n444 & new_new_n11572__;
  assign new_new_n34910__ = ~new_new_n34908__ & ~new_new_n34909__;
  assign new_new_n34911__ = new_new_n11603__ & ~new_new_n34910__;
  assign new_new_n34912__ = ~ys__n444 & new_new_n11608__;
  assign new_new_n34913__ = ys__n444 & ~new_new_n11608__;
  assign new_new_n34914__ = ~new_new_n34912__ & ~new_new_n34913__;
  assign new_new_n34915__ = new_new_n11619__ & ~new_new_n34914__;
  assign new_new_n34916__ = ~new_new_n34911__ & ~new_new_n34915__;
  assign new_new_n34917__ = ~new_new_n34907__ & new_new_n34916__;
  assign new_new_n34918__ = new_new_n11625__ & ~new_new_n34917__;
  assign new_new_n34919__ = ~new_new_n34906__ & ~new_new_n34918__;
  assign new_new_n34920__ = new_new_n11629__ & ~new_new_n34919__;
  assign new_new_n34921__ = ~new_new_n34890__ & ~new_new_n34920__;
  assign new_new_n34922__ = new_new_n11640__ & ~new_new_n34921__;
  assign new_new_n34923__ = ys__n47680 & new_new_n11644__;
  assign new_new_n34924__ = new_new_n11642__ & ~new_new_n34919__;
  assign new_new_n34925__ = ~new_new_n34923__ & ~new_new_n34924__;
  assign new_new_n34926__ = new_new_n11650__ & ~new_new_n34925__;
  assign ys__n28560 = new_new_n34922__ | new_new_n34926__;
  assign new_new_n34928__ = ys__n47681 & new_new_n11634__;
  assign new_new_n34929__ = ys__n22862 & ~new_new_n11180__;
  assign new_new_n34930__ = new_new_n11175__ & new_new_n34929__;
  assign new_new_n34931__ = ~new_new_n16391__ & ~new_new_n34930__;
  assign new_new_n34932__ = ~new_new_n11186__ & ~new_new_n34931__;
  assign new_new_n34933__ = ys__n438 & new_new_n11186__;
  assign new_new_n34934__ = ~new_new_n34932__ & ~new_new_n34933__;
  assign new_new_n34935__ = ~new_new_n11270__ & ~new_new_n34934__;
  assign new_new_n34936__ = new_new_n11270__ & ys__n23521;
  assign new_new_n34937__ = ~new_new_n34935__ & ~new_new_n34936__;
  assign new_new_n34938__ = new_new_n11324__ & ~new_new_n34937__;
  assign new_new_n34939__ = ys__n4478 & ~ys__n28243;
  assign new_new_n34940__ = ys__n28243 & ys__n28634;
  assign new_new_n34941__ = ~new_new_n34939__ & ~new_new_n34940__;
  assign new_new_n34942__ = ~new_new_n11324__ & ~new_new_n34941__;
  assign new_new_n34943__ = ~new_new_n34938__ & ~new_new_n34942__;
  assign new_new_n34944__ = ~new_new_n11343__ & ~new_new_n34943__;
  assign new_new_n34945__ = ys__n438 & ~new_new_n11569__;
  assign new_new_n34946__ = ~ys__n444 & ~new_new_n11572__;
  assign new_new_n34947__ = ~ys__n444 & ~new_new_n34946__;
  assign new_new_n34948__ = ys__n438 & ~new_new_n34947__;
  assign new_new_n34949__ = ~ys__n438 & new_new_n34947__;
  assign new_new_n34950__ = ~new_new_n34948__ & ~new_new_n34949__;
  assign new_new_n34951__ = new_new_n11603__ & ~new_new_n34950__;
  assign new_new_n34952__ = ys__n444 & new_new_n11608__;
  assign new_new_n34953__ = ~ys__n438 & new_new_n34952__;
  assign new_new_n34954__ = ys__n438 & ~new_new_n34952__;
  assign new_new_n34955__ = ~new_new_n34953__ & ~new_new_n34954__;
  assign new_new_n34956__ = new_new_n11619__ & ~new_new_n34955__;
  assign new_new_n34957__ = ~new_new_n34951__ & ~new_new_n34956__;
  assign new_new_n34958__ = ~new_new_n34945__ & new_new_n34957__;
  assign new_new_n34959__ = new_new_n11625__ & ~new_new_n34958__;
  assign new_new_n34960__ = ~new_new_n34944__ & ~new_new_n34959__;
  assign new_new_n34961__ = new_new_n11629__ & ~new_new_n34960__;
  assign new_new_n34962__ = ~new_new_n34928__ & ~new_new_n34961__;
  assign new_new_n34963__ = new_new_n11640__ & ~new_new_n34962__;
  assign new_new_n34964__ = ys__n47681 & new_new_n11644__;
  assign new_new_n34965__ = new_new_n11642__ & ~new_new_n34960__;
  assign new_new_n34966__ = ~new_new_n34964__ & ~new_new_n34965__;
  assign new_new_n34967__ = new_new_n11650__ & ~new_new_n34966__;
  assign ys__n28563 = new_new_n34963__ | new_new_n34967__;
  assign new_new_n34969__ = ys__n22864 & new_new_n11175__;
  assign new_new_n34970__ = ~new_new_n15981__ & ~new_new_n34969__;
  assign new_new_n34971__ = ~new_new_n11180__ & ~new_new_n34970__;
  assign new_new_n34972__ = ~new_new_n16397__ & ~new_new_n34971__;
  assign new_new_n34973__ = ~new_new_n11186__ & ~new_new_n34972__;
  assign new_new_n34974__ = ys__n446 & new_new_n11186__;
  assign new_new_n34975__ = ~new_new_n34973__ & ~new_new_n34974__;
  assign new_new_n34976__ = ~new_new_n11270__ & ~new_new_n34975__;
  assign new_new_n34977__ = new_new_n11270__ & ys__n23523;
  assign new_new_n34978__ = ~new_new_n34976__ & ~new_new_n34977__;
  assign new_new_n34979__ = new_new_n11324__ & ~new_new_n34978__;
  assign new_new_n34980__ = ys__n4480 & ~ys__n28243;
  assign new_new_n34981__ = ys__n28243 & ys__n28635;
  assign new_new_n34982__ = ~new_new_n34980__ & ~new_new_n34981__;
  assign new_new_n34983__ = ~new_new_n11324__ & ~new_new_n34982__;
  assign new_new_n34984__ = ~new_new_n34979__ & ~new_new_n34983__;
  assign new_new_n34985__ = ~new_new_n11343__ & ~new_new_n34984__;
  assign new_new_n34986__ = ys__n446 & ~new_new_n11569__;
  assign new_new_n34987__ = ys__n446 & ~new_new_n11577__;
  assign new_new_n34988__ = ~ys__n446 & new_new_n11577__;
  assign new_new_n34989__ = ~new_new_n34987__ & ~new_new_n34988__;
  assign new_new_n34990__ = new_new_n11603__ & ~new_new_n34989__;
  assign new_new_n34991__ = ~ys__n446 & new_new_n11610__;
  assign new_new_n34992__ = ys__n446 & ~new_new_n11610__;
  assign new_new_n34993__ = ~new_new_n34991__ & ~new_new_n34992__;
  assign new_new_n34994__ = new_new_n11619__ & ~new_new_n34993__;
  assign new_new_n34995__ = ~new_new_n34990__ & ~new_new_n34994__;
  assign new_new_n34996__ = ~new_new_n34986__ & new_new_n34995__;
  assign new_new_n34997__ = new_new_n11625__ & ~new_new_n34996__;
  assign new_new_n34998__ = ~new_new_n34985__ & ~new_new_n34997__;
  assign new_new_n34999__ = new_new_n11629__ & ~new_new_n34998__;
  assign new_new_n35000__ = ys__n47682 & new_new_n11634__;
  assign new_new_n35001__ = ~new_new_n16021__ & ~new_new_n35000__;
  assign new_new_n35002__ = ~new_new_n34999__ & new_new_n35001__;
  assign new_new_n35003__ = new_new_n11640__ & ~new_new_n35002__;
  assign new_new_n35004__ = new_new_n11642__ & ~new_new_n34998__;
  assign new_new_n35005__ = ys__n47682 & new_new_n11644__;
  assign new_new_n35006__ = ~new_new_n16021__ & ~new_new_n35005__;
  assign new_new_n35007__ = ~new_new_n35004__ & new_new_n35006__;
  assign new_new_n35008__ = new_new_n11650__ & ~new_new_n35007__;
  assign ys__n28566 = new_new_n35003__ | new_new_n35008__;
  assign new_new_n35010__ = ~ys__n23627 & ~ys__n23629;
  assign new_new_n35011__ = ~new_new_n11175__ & new_new_n35010__;
  assign new_new_n35012__ = ys__n22866 & new_new_n11175__;
  assign new_new_n35013__ = ~new_new_n35011__ & ~new_new_n35012__;
  assign new_new_n35014__ = ~new_new_n11180__ & ~new_new_n35013__;
  assign new_new_n35015__ = ~new_new_n16403__ & ~new_new_n35014__;
  assign new_new_n35016__ = ~new_new_n11186__ & ~new_new_n35015__;
  assign new_new_n35017__ = ys__n434 & new_new_n11186__;
  assign new_new_n35018__ = ~new_new_n35016__ & ~new_new_n35017__;
  assign new_new_n35019__ = ~new_new_n11270__ & ~new_new_n35018__;
  assign new_new_n35020__ = new_new_n11270__ & ys__n23525;
  assign new_new_n35021__ = ~new_new_n35019__ & ~new_new_n35020__;
  assign new_new_n35022__ = new_new_n11324__ & ~new_new_n35021__;
  assign new_new_n35023__ = ys__n516 & ~ys__n28243;
  assign new_new_n35024__ = ys__n28243 & ys__n28636;
  assign new_new_n35025__ = ~new_new_n35023__ & ~new_new_n35024__;
  assign new_new_n35026__ = ~new_new_n11324__ & ~new_new_n35025__;
  assign new_new_n35027__ = ~new_new_n35022__ & ~new_new_n35026__;
  assign new_new_n35028__ = ~new_new_n11343__ & ~new_new_n35027__;
  assign new_new_n35029__ = ys__n434 & ~new_new_n11569__;
  assign new_new_n35030__ = ~ys__n446 & ~new_new_n11577__;
  assign new_new_n35031__ = ~ys__n446 & ~new_new_n35030__;
  assign new_new_n35032__ = ys__n434 & ~new_new_n35031__;
  assign new_new_n35033__ = ~ys__n434 & new_new_n35031__;
  assign new_new_n35034__ = ~new_new_n35032__ & ~new_new_n35033__;
  assign new_new_n35035__ = new_new_n11603__ & ~new_new_n35034__;
  assign new_new_n35036__ = ys__n446 & new_new_n11610__;
  assign new_new_n35037__ = ~ys__n434 & new_new_n35036__;
  assign new_new_n35038__ = ys__n434 & ~new_new_n35036__;
  assign new_new_n35039__ = ~new_new_n35037__ & ~new_new_n35038__;
  assign new_new_n35040__ = new_new_n11619__ & ~new_new_n35039__;
  assign new_new_n35041__ = ~new_new_n35035__ & ~new_new_n35040__;
  assign new_new_n35042__ = ~new_new_n35029__ & new_new_n35041__;
  assign new_new_n35043__ = new_new_n11625__ & ~new_new_n35042__;
  assign new_new_n35044__ = ~new_new_n35028__ & ~new_new_n35043__;
  assign new_new_n35045__ = new_new_n11629__ & ~new_new_n35044__;
  assign new_new_n35046__ = ys__n935 & ~ys__n23629;
  assign new_new_n35047__ = ~new_new_n11631__ & ~new_new_n35046__;
  assign new_new_n35048__ = new_new_n11628__ & ~new_new_n35047__;
  assign new_new_n35049__ = ys__n47683 & new_new_n11634__;
  assign new_new_n35050__ = ~new_new_n35048__ & ~new_new_n35049__;
  assign new_new_n35051__ = ~new_new_n35045__ & new_new_n35050__;
  assign new_new_n35052__ = new_new_n11640__ & ~new_new_n35051__;
  assign new_new_n35053__ = new_new_n11642__ & ~new_new_n35044__;
  assign new_new_n35054__ = ys__n47683 & new_new_n11644__;
  assign new_new_n35055__ = ~new_new_n35048__ & ~new_new_n35054__;
  assign new_new_n35056__ = ~new_new_n35053__ & new_new_n35055__;
  assign new_new_n35057__ = new_new_n11650__ & ~new_new_n35056__;
  assign ys__n28569 = new_new_n35052__ | new_new_n35057__;
  assign new_new_n35059__ = ys__n22868 & new_new_n11175__;
  assign new_new_n35060__ = ~new_new_n35011__ & ~new_new_n35059__;
  assign new_new_n35061__ = ~new_new_n11180__ & ~new_new_n35060__;
  assign new_new_n35062__ = ~new_new_n16409__ & ~new_new_n35061__;
  assign new_new_n35063__ = ~new_new_n11186__ & ~new_new_n35062__;
  assign new_new_n35064__ = ys__n436 & new_new_n11186__;
  assign new_new_n35065__ = ~new_new_n35063__ & ~new_new_n35064__;
  assign new_new_n35066__ = ~new_new_n11270__ & ~new_new_n35065__;
  assign new_new_n35067__ = new_new_n11270__ & ys__n23527;
  assign new_new_n35068__ = ~new_new_n35066__ & ~new_new_n35067__;
  assign new_new_n35069__ = new_new_n11324__ & ~new_new_n35068__;
  assign new_new_n35070__ = ys__n4494 & ~ys__n28243;
  assign new_new_n35071__ = ys__n28243 & ys__n28637;
  assign new_new_n35072__ = ~new_new_n35070__ & ~new_new_n35071__;
  assign new_new_n35073__ = ~new_new_n11324__ & ~new_new_n35072__;
  assign new_new_n35074__ = ~new_new_n35069__ & ~new_new_n35073__;
  assign new_new_n35075__ = ~new_new_n11343__ & ~new_new_n35074__;
  assign new_new_n35076__ = ys__n436 & ~new_new_n11569__;
  assign new_new_n35077__ = ~new_new_n11577__ & new_new_n11579__;
  assign new_new_n35078__ = new_new_n11583__ & ~new_new_n35077__;
  assign new_new_n35079__ = ys__n436 & ~new_new_n35078__;
  assign new_new_n35080__ = ~ys__n436 & new_new_n35078__;
  assign new_new_n35081__ = ~new_new_n35079__ & ~new_new_n35080__;
  assign new_new_n35082__ = new_new_n11603__ & ~new_new_n35081__;
  assign new_new_n35083__ = new_new_n11610__ & new_new_n11611__;
  assign new_new_n35084__ = ~ys__n436 & new_new_n35083__;
  assign new_new_n35085__ = ys__n436 & ~new_new_n35083__;
  assign new_new_n35086__ = ~new_new_n35084__ & ~new_new_n35085__;
  assign new_new_n35087__ = new_new_n11619__ & ~new_new_n35086__;
  assign new_new_n35088__ = ~new_new_n35082__ & ~new_new_n35087__;
  assign new_new_n35089__ = ~new_new_n35076__ & new_new_n35088__;
  assign new_new_n35090__ = new_new_n11625__ & ~new_new_n35089__;
  assign new_new_n35091__ = ~new_new_n35075__ & ~new_new_n35090__;
  assign new_new_n35092__ = new_new_n11629__ & ~new_new_n35091__;
  assign new_new_n35093__ = ys__n47684 & new_new_n11634__;
  assign new_new_n35094__ = ~new_new_n35048__ & ~new_new_n35093__;
  assign new_new_n35095__ = ~new_new_n35092__ & new_new_n35094__;
  assign new_new_n35096__ = new_new_n11640__ & ~new_new_n35095__;
  assign new_new_n35097__ = new_new_n11642__ & ~new_new_n35091__;
  assign new_new_n35098__ = ys__n47684 & new_new_n11644__;
  assign new_new_n35099__ = ~new_new_n35048__ & ~new_new_n35098__;
  assign new_new_n35100__ = ~new_new_n35097__ & new_new_n35099__;
  assign new_new_n35101__ = new_new_n11650__ & ~new_new_n35100__;
  assign ys__n28572 = new_new_n35096__ | new_new_n35101__;
  assign new_new_n35103__ = ys__n22870 & new_new_n11175__;
  assign new_new_n35104__ = ~new_new_n11176__ & ~new_new_n35103__;
  assign new_new_n35105__ = ~new_new_n11180__ & ~new_new_n35104__;
  assign new_new_n35106__ = ~new_new_n16415__ & ~new_new_n35105__;
  assign new_new_n35107__ = ~new_new_n11186__ & ~new_new_n35106__;
  assign new_new_n35108__ = ys__n432 & new_new_n11186__;
  assign new_new_n35109__ = ~new_new_n35107__ & ~new_new_n35108__;
  assign new_new_n35110__ = ~new_new_n11270__ & ~new_new_n35109__;
  assign new_new_n35111__ = new_new_n11270__ & ys__n23529;
  assign new_new_n35112__ = ~new_new_n35110__ & ~new_new_n35111__;
  assign new_new_n35113__ = new_new_n11324__ & ~new_new_n35112__;
  assign new_new_n35114__ = ys__n4496 & ~ys__n28243;
  assign new_new_n35115__ = ys__n28243 & ys__n28638;
  assign new_new_n35116__ = ~new_new_n35114__ & ~new_new_n35115__;
  assign new_new_n35117__ = ~new_new_n11324__ & ~new_new_n35116__;
  assign new_new_n35118__ = ~new_new_n35113__ & ~new_new_n35117__;
  assign new_new_n35119__ = ~new_new_n11343__ & ~new_new_n35118__;
  assign new_new_n35120__ = ys__n432 & ~new_new_n11569__;
  assign new_new_n35121__ = ~ys__n436 & ~new_new_n35078__;
  assign new_new_n35122__ = ~ys__n436 & ~new_new_n35121__;
  assign new_new_n35123__ = ys__n432 & ~new_new_n35122__;
  assign new_new_n35124__ = ~ys__n432 & new_new_n35122__;
  assign new_new_n35125__ = ~new_new_n35123__ & ~new_new_n35124__;
  assign new_new_n35126__ = new_new_n11603__ & ~new_new_n35125__;
  assign new_new_n35127__ = ys__n436 & new_new_n35083__;
  assign new_new_n35128__ = ~ys__n432 & new_new_n35127__;
  assign new_new_n35129__ = ys__n432 & ~new_new_n35127__;
  assign new_new_n35130__ = ~new_new_n35128__ & ~new_new_n35129__;
  assign new_new_n35131__ = new_new_n11619__ & ~new_new_n35130__;
  assign new_new_n35132__ = ~new_new_n35126__ & ~new_new_n35131__;
  assign new_new_n35133__ = ~new_new_n35120__ & new_new_n35132__;
  assign new_new_n35134__ = new_new_n11625__ & ~new_new_n35133__;
  assign new_new_n35135__ = ~new_new_n35119__ & ~new_new_n35134__;
  assign new_new_n35136__ = new_new_n11629__ & ~new_new_n35135__;
  assign new_new_n35137__ = ys__n47685 & new_new_n11634__;
  assign new_new_n35138__ = ~new_new_n11633__ & ~new_new_n35137__;
  assign new_new_n35139__ = ~new_new_n35136__ & new_new_n35138__;
  assign new_new_n35140__ = new_new_n11640__ & ~new_new_n35139__;
  assign new_new_n35141__ = new_new_n11642__ & ~new_new_n35135__;
  assign new_new_n35142__ = ys__n47685 & new_new_n11644__;
  assign new_new_n35143__ = ~new_new_n11633__ & ~new_new_n35142__;
  assign new_new_n35144__ = ~new_new_n35141__ & new_new_n35143__;
  assign new_new_n35145__ = new_new_n11650__ & ~new_new_n35144__;
  assign ys__n28575 = new_new_n35140__ | new_new_n35145__;
  assign new_new_n35147__ = ys__n22872 & new_new_n11175__;
  assign new_new_n35148__ = ~new_new_n11176__ & ~new_new_n35147__;
  assign new_new_n35149__ = ~new_new_n11180__ & ~new_new_n35148__;
  assign new_new_n35150__ = ~new_new_n16421__ & ~new_new_n35149__;
  assign new_new_n35151__ = ~new_new_n11186__ & ~new_new_n35150__;
  assign new_new_n35152__ = ys__n448 & new_new_n11186__;
  assign new_new_n35153__ = ~new_new_n35151__ & ~new_new_n35152__;
  assign new_new_n35154__ = ~new_new_n11270__ & ~new_new_n35153__;
  assign new_new_n35155__ = new_new_n11270__ & ys__n23531;
  assign new_new_n35156__ = ~new_new_n35154__ & ~new_new_n35155__;
  assign new_new_n35157__ = new_new_n11324__ & ~new_new_n35156__;
  assign new_new_n35158__ = ys__n632 & ~ys__n28243;
  assign new_new_n35159__ = ys__n28243 & ys__n28639;
  assign new_new_n35160__ = ~new_new_n35158__ & ~new_new_n35159__;
  assign new_new_n35161__ = ~new_new_n11324__ & ~new_new_n35160__;
  assign new_new_n35162__ = ~new_new_n35157__ & ~new_new_n35161__;
  assign new_new_n35163__ = ~new_new_n11343__ & ~new_new_n35162__;
  assign new_new_n35164__ = ys__n448 & ~new_new_n11569__;
  assign new_new_n35165__ = ys__n448 & ~new_new_n11588__;
  assign new_new_n35166__ = ~ys__n448 & new_new_n11588__;
  assign new_new_n35167__ = ~new_new_n35165__ & ~new_new_n35166__;
  assign new_new_n35168__ = new_new_n11603__ & ~new_new_n35167__;
  assign new_new_n35169__ = ~ys__n448 & new_new_n11614__;
  assign new_new_n35170__ = ys__n448 & ~new_new_n11614__;
  assign new_new_n35171__ = ~new_new_n35169__ & ~new_new_n35170__;
  assign new_new_n35172__ = new_new_n11619__ & ~new_new_n35171__;
  assign new_new_n35173__ = ~new_new_n35168__ & ~new_new_n35172__;
  assign new_new_n35174__ = ~new_new_n35164__ & new_new_n35173__;
  assign new_new_n35175__ = new_new_n11625__ & ~new_new_n35174__;
  assign new_new_n35176__ = ~new_new_n35163__ & ~new_new_n35175__;
  assign new_new_n35177__ = new_new_n11629__ & ~new_new_n35176__;
  assign new_new_n35178__ = ys__n47686 & new_new_n11634__;
  assign new_new_n35179__ = ~new_new_n11633__ & ~new_new_n35178__;
  assign new_new_n35180__ = ~new_new_n35177__ & new_new_n35179__;
  assign new_new_n35181__ = new_new_n11640__ & ~new_new_n35180__;
  assign new_new_n35182__ = new_new_n11642__ & ~new_new_n35176__;
  assign new_new_n35183__ = ys__n47686 & new_new_n11644__;
  assign new_new_n35184__ = ~new_new_n11633__ & ~new_new_n35183__;
  assign new_new_n35185__ = ~new_new_n35182__ & new_new_n35184__;
  assign new_new_n35186__ = new_new_n11650__ & ~new_new_n35185__;
  assign ys__n28578 = new_new_n35181__ | new_new_n35186__;
  assign new_new_n35188__ = ys__n22874 & new_new_n11175__;
  assign new_new_n35189__ = ~new_new_n11176__ & ~new_new_n35188__;
  assign new_new_n35190__ = ~new_new_n11180__ & ~new_new_n35189__;
  assign new_new_n35191__ = ~new_new_n16427__ & ~new_new_n35190__;
  assign new_new_n35192__ = ~new_new_n11186__ & ~new_new_n35191__;
  assign new_new_n35193__ = ys__n428 & new_new_n11186__;
  assign new_new_n35194__ = ~new_new_n35192__ & ~new_new_n35193__;
  assign new_new_n35195__ = ~new_new_n11270__ & ~new_new_n35194__;
  assign new_new_n35196__ = new_new_n11270__ & ys__n23533;
  assign new_new_n35197__ = ~new_new_n35195__ & ~new_new_n35196__;
  assign new_new_n35198__ = new_new_n11324__ & ~new_new_n35197__;
  assign new_new_n35199__ = ys__n512 & ~ys__n28243;
  assign new_new_n35200__ = ys__n28243 & ys__n28640;
  assign new_new_n35201__ = ~new_new_n35199__ & ~new_new_n35200__;
  assign new_new_n35202__ = ~new_new_n11324__ & ~new_new_n35201__;
  assign new_new_n35203__ = ~new_new_n35198__ & ~new_new_n35202__;
  assign new_new_n35204__ = ~new_new_n11343__ & ~new_new_n35203__;
  assign new_new_n35205__ = ys__n428 & ~new_new_n11569__;
  assign new_new_n35206__ = ~ys__n448 & ~new_new_n11588__;
  assign new_new_n35207__ = ~ys__n448 & ~new_new_n35206__;
  assign new_new_n35208__ = ys__n428 & ~new_new_n35207__;
  assign new_new_n35209__ = ~ys__n428 & new_new_n35207__;
  assign new_new_n35210__ = ~new_new_n35208__ & ~new_new_n35209__;
  assign new_new_n35211__ = new_new_n11603__ & ~new_new_n35210__;
  assign new_new_n35212__ = ys__n448 & new_new_n11614__;
  assign new_new_n35213__ = ~ys__n428 & new_new_n35212__;
  assign new_new_n35214__ = ys__n428 & ~new_new_n35212__;
  assign new_new_n35215__ = ~new_new_n35213__ & ~new_new_n35214__;
  assign new_new_n35216__ = new_new_n11619__ & ~new_new_n35215__;
  assign new_new_n35217__ = ~new_new_n35211__ & ~new_new_n35216__;
  assign new_new_n35218__ = ~new_new_n35205__ & new_new_n35217__;
  assign new_new_n35219__ = new_new_n11625__ & ~new_new_n35218__;
  assign new_new_n35220__ = ~new_new_n35204__ & ~new_new_n35219__;
  assign new_new_n35221__ = new_new_n11629__ & ~new_new_n35220__;
  assign new_new_n35222__ = ys__n47687 & new_new_n11634__;
  assign new_new_n35223__ = ~new_new_n11633__ & ~new_new_n35222__;
  assign new_new_n35224__ = ~new_new_n35221__ & new_new_n35223__;
  assign new_new_n35225__ = new_new_n11640__ & ~new_new_n35224__;
  assign new_new_n35226__ = new_new_n11642__ & ~new_new_n35220__;
  assign new_new_n35227__ = ys__n47687 & new_new_n11644__;
  assign new_new_n35228__ = ~new_new_n11633__ & ~new_new_n35227__;
  assign new_new_n35229__ = ~new_new_n35226__ & new_new_n35228__;
  assign new_new_n35230__ = new_new_n11650__ & ~new_new_n35229__;
  assign ys__n28581 = new_new_n35225__ | new_new_n35230__;
  assign new_new_n35232__ = ys__n22876 & new_new_n11175__;
  assign new_new_n35233__ = ~new_new_n11176__ & ~new_new_n35232__;
  assign new_new_n35234__ = ~new_new_n11180__ & ~new_new_n35233__;
  assign new_new_n35235__ = ~new_new_n16433__ & ~new_new_n35234__;
  assign new_new_n35236__ = ~new_new_n11186__ & ~new_new_n35235__;
  assign new_new_n35237__ = ys__n430 & new_new_n11186__;
  assign new_new_n35238__ = ~new_new_n35236__ & ~new_new_n35237__;
  assign new_new_n35239__ = ~new_new_n11270__ & ~new_new_n35238__;
  assign new_new_n35240__ = new_new_n11270__ & ys__n23535;
  assign new_new_n35241__ = ~new_new_n35239__ & ~new_new_n35240__;
  assign new_new_n35242__ = new_new_n11324__ & ~new_new_n35241__;
  assign new_new_n35243__ = ys__n520 & ~ys__n28243;
  assign new_new_n35244__ = ys__n28243 & ys__n28641;
  assign new_new_n35245__ = ~new_new_n35243__ & ~new_new_n35244__;
  assign new_new_n35246__ = ~new_new_n11324__ & ~new_new_n35245__;
  assign new_new_n35247__ = ~new_new_n35242__ & ~new_new_n35246__;
  assign new_new_n35248__ = ~new_new_n11343__ & ~new_new_n35247__;
  assign new_new_n35249__ = ys__n430 & ~new_new_n11569__;
  assign new_new_n35250__ = ~new_new_n11588__ & new_new_n11590__;
  assign new_new_n35251__ = new_new_n11594__ & ~new_new_n35250__;
  assign new_new_n35252__ = ys__n430 & ~new_new_n35251__;
  assign new_new_n35253__ = ~ys__n430 & new_new_n35251__;
  assign new_new_n35254__ = ~new_new_n35252__ & ~new_new_n35253__;
  assign new_new_n35255__ = new_new_n11603__ & ~new_new_n35254__;
  assign new_new_n35256__ = new_new_n11605__ & new_new_n11614__;
  assign new_new_n35257__ = ~ys__n430 & new_new_n35256__;
  assign new_new_n35258__ = ys__n430 & ~new_new_n35256__;
  assign new_new_n35259__ = ~new_new_n35257__ & ~new_new_n35258__;
  assign new_new_n35260__ = new_new_n11619__ & ~new_new_n35259__;
  assign new_new_n35261__ = ~new_new_n35255__ & ~new_new_n35260__;
  assign new_new_n35262__ = ~new_new_n35249__ & new_new_n35261__;
  assign new_new_n35263__ = new_new_n11625__ & ~new_new_n35262__;
  assign new_new_n35264__ = ~new_new_n35248__ & ~new_new_n35263__;
  assign new_new_n35265__ = new_new_n11629__ & ~new_new_n35264__;
  assign new_new_n35266__ = ys__n47688 & new_new_n11634__;
  assign new_new_n35267__ = ~new_new_n11633__ & ~new_new_n35266__;
  assign new_new_n35268__ = ~new_new_n35265__ & new_new_n35267__;
  assign new_new_n35269__ = new_new_n11640__ & ~new_new_n35268__;
  assign new_new_n35270__ = new_new_n11642__ & ~new_new_n35264__;
  assign new_new_n35271__ = ys__n47688 & new_new_n11644__;
  assign new_new_n35272__ = ~new_new_n11633__ & ~new_new_n35271__;
  assign new_new_n35273__ = ~new_new_n35270__ & new_new_n35272__;
  assign new_new_n35274__ = new_new_n11650__ & ~new_new_n35273__;
  assign ys__n28584 = new_new_n35269__ | new_new_n35274__;
  assign new_new_n35276__ = ys__n22878 & new_new_n11175__;
  assign new_new_n35277__ = ~new_new_n11176__ & ~new_new_n35276__;
  assign new_new_n35278__ = ~new_new_n11180__ & ~new_new_n35277__;
  assign new_new_n35279__ = ~new_new_n16439__ & ~new_new_n35278__;
  assign new_new_n35280__ = ~new_new_n11186__ & ~new_new_n35279__;
  assign new_new_n35281__ = ys__n426 & new_new_n11186__;
  assign new_new_n35282__ = ~new_new_n35280__ & ~new_new_n35281__;
  assign new_new_n35283__ = ~new_new_n11270__ & ~new_new_n35282__;
  assign new_new_n35284__ = new_new_n11270__ & ys__n23537;
  assign new_new_n35285__ = ~new_new_n35283__ & ~new_new_n35284__;
  assign new_new_n35286__ = new_new_n11324__ & ~new_new_n35285__;
  assign new_new_n35287__ = ys__n426 & ~new_new_n11324__;
  assign new_new_n35288__ = ~new_new_n35286__ & ~new_new_n35287__;
  assign new_new_n35289__ = ~new_new_n11343__ & ~new_new_n35288__;
  assign new_new_n35290__ = ys__n426 & ~new_new_n11569__;
  assign new_new_n35291__ = ~ys__n430 & ~new_new_n35251__;
  assign new_new_n35292__ = ~ys__n430 & ~new_new_n35291__;
  assign new_new_n35293__ = ys__n426 & ~new_new_n35292__;
  assign new_new_n35294__ = ~ys__n426 & new_new_n35292__;
  assign new_new_n35295__ = ~new_new_n35293__ & ~new_new_n35294__;
  assign new_new_n35296__ = new_new_n11603__ & ~new_new_n35295__;
  assign new_new_n35297__ = ys__n430 & new_new_n35256__;
  assign new_new_n35298__ = ~ys__n426 & new_new_n35297__;
  assign new_new_n35299__ = ys__n426 & ~new_new_n35297__;
  assign new_new_n35300__ = ~new_new_n35298__ & ~new_new_n35299__;
  assign new_new_n35301__ = new_new_n11619__ & ~new_new_n35300__;
  assign new_new_n35302__ = ~new_new_n35296__ & ~new_new_n35301__;
  assign new_new_n35303__ = ~new_new_n35290__ & new_new_n35302__;
  assign new_new_n35304__ = new_new_n11625__ & ~new_new_n35303__;
  assign new_new_n35305__ = ~new_new_n35289__ & ~new_new_n35304__;
  assign new_new_n35306__ = new_new_n11629__ & ~new_new_n35305__;
  assign new_new_n35307__ = ys__n47689 & new_new_n11634__;
  assign new_new_n35308__ = ~new_new_n11633__ & ~new_new_n35307__;
  assign new_new_n35309__ = ~new_new_n35306__ & new_new_n35308__;
  assign new_new_n35310__ = new_new_n11640__ & ~new_new_n35309__;
  assign new_new_n35311__ = new_new_n11642__ & ~new_new_n35305__;
  assign new_new_n35312__ = ys__n47689 & new_new_n11644__;
  assign new_new_n35313__ = ~new_new_n11633__ & ~new_new_n35312__;
  assign new_new_n35314__ = ~new_new_n35311__ & new_new_n35313__;
  assign new_new_n35315__ = new_new_n11650__ & ~new_new_n35314__;
  assign ys__n28587 = new_new_n35310__ | new_new_n35315__;
  assign ys__n28661 = ys__n532 & ~ys__n28243;
  assign ys__n28662 = ys__n746 & ~ys__n28243;
  assign new_new_n35319__ = ~ys__n860 & new_new_n10986__;
  assign new_new_n35320__ = ~ys__n204 & new_new_n35319__;
  assign new_new_n35321__ = ~ys__n182 & ys__n192;
  assign new_new_n35322__ = new_new_n35320__ & new_new_n35321__;
  assign new_new_n35323__ = ys__n182 & ~ys__n184;
  assign new_new_n35324__ = ys__n204 & new_new_n35319__;
  assign new_new_n35325__ = new_new_n35323__ & new_new_n35324__;
  assign new_new_n35326__ = ~ys__n182 & ys__n204;
  assign new_new_n35327__ = new_new_n35319__ & new_new_n35326__;
  assign new_new_n35328__ = new_new_n35319__ & ~new_new_n35327__;
  assign new_new_n35329__ = ~new_new_n35325__ & new_new_n35328__;
  assign new_new_n35330__ = ~new_new_n35322__ & new_new_n35329__;
  assign new_new_n35331__ = ys__n182 & ys__n192;
  assign new_new_n35332__ = new_new_n35320__ & new_new_n35331__;
  assign new_new_n35333__ = ys__n182 & ys__n184;
  assign new_new_n35334__ = new_new_n35324__ & new_new_n35333__;
  assign new_new_n35335__ = ~ys__n192 & ~ys__n204;
  assign new_new_n35336__ = new_new_n35319__ & new_new_n35335__;
  assign new_new_n35337__ = ~new_new_n35334__ & ~new_new_n35336__;
  assign new_new_n35338__ = ~new_new_n35332__ & new_new_n35337__;
  assign new_new_n35339__ = new_new_n35330__ & new_new_n35338__;
  assign new_new_n35340__ = ys__n190 & new_new_n35333__;
  assign new_new_n35341__ = ys__n190 & new_new_n35323__;
  assign new_new_n35342__ = ~new_new_n35340__ & ~new_new_n35341__;
  assign new_new_n35343__ = ~ys__n182 & ys__n184;
  assign new_new_n35344__ = ys__n190 & new_new_n35343__;
  assign new_new_n35345__ = ~ys__n182 & ~ys__n184;
  assign new_new_n35346__ = ~ys__n190 & new_new_n35345__;
  assign new_new_n35347__ = ~new_new_n35344__ & ~new_new_n35346__;
  assign new_new_n35348__ = new_new_n35342__ & new_new_n35347__;
  assign new_new_n35349__ = ~new_new_n35323__ & ~new_new_n35333__;
  assign new_new_n35350__ = ~new_new_n35343__ & ~new_new_n35345__;
  assign new_new_n35351__ = new_new_n35349__ & new_new_n35350__;
  assign new_new_n35352__ = ~new_new_n35348__ & ~new_new_n35351__;
  assign new_new_n35353__ = ~new_new_n35330__ & new_new_n35352__;
  assign new_new_n35354__ = ~new_new_n35339__ & new_new_n35353__;
  assign new_new_n35355__ = ys__n4566 & new_new_n12582__;
  assign new_new_n35356__ = new_new_n35354__ & new_new_n35355__;
  assign new_new_n35357__ = ~new_new_n11005__ & new_new_n12579__;
  assign new_new_n35358__ = new_new_n35354__ & new_new_n35357__;
  assign new_new_n35359__ = ys__n186 & ~ys__n202;
  assign new_new_n35360__ = new_new_n35343__ & new_new_n35359__;
  assign new_new_n35361__ = ~ys__n38453 & new_new_n35360__;
  assign new_new_n35362__ = ~ys__n186 & ~ys__n202;
  assign new_new_n35363__ = new_new_n35343__ & new_new_n35362__;
  assign new_new_n35364__ = ~ys__n38453 & new_new_n35363__;
  assign new_new_n35365__ = ~new_new_n35361__ & ~new_new_n35364__;
  assign new_new_n35366__ = new_new_n35323__ & new_new_n35359__;
  assign new_new_n35367__ = ~ys__n38453 & new_new_n35366__;
  assign new_new_n35368__ = ~ys__n186 & ys__n202;
  assign new_new_n35369__ = new_new_n35323__ & new_new_n35368__;
  assign new_new_n35370__ = ~ys__n38453 & new_new_n35369__;
  assign new_new_n35371__ = ~new_new_n35367__ & ~new_new_n35370__;
  assign new_new_n35372__ = new_new_n35365__ & new_new_n35371__;
  assign new_new_n35373__ = ys__n38453 & new_new_n35368__;
  assign new_new_n35374__ = ys__n186 & ys__n202;
  assign new_new_n35375__ = new_new_n35333__ & new_new_n35374__;
  assign new_new_n35376__ = ~ys__n38453 & new_new_n35375__;
  assign new_new_n35377__ = ~new_new_n35373__ & ~new_new_n35376__;
  assign new_new_n35378__ = new_new_n35333__ & new_new_n35362__;
  assign new_new_n35379__ = ~ys__n38453 & new_new_n35378__;
  assign new_new_n35380__ = new_new_n35333__ & new_new_n35368__;
  assign new_new_n35381__ = ~ys__n38453 & new_new_n35380__;
  assign new_new_n35382__ = ~new_new_n35379__ & ~new_new_n35381__;
  assign new_new_n35383__ = new_new_n35377__ & new_new_n35382__;
  assign new_new_n35384__ = new_new_n35372__ & new_new_n35383__;
  assign new_new_n35385__ = new_new_n35333__ & new_new_n35359__;
  assign new_new_n35386__ = ~ys__n38453 & new_new_n35385__;
  assign new_new_n35387__ = ys__n38453 & new_new_n35362__;
  assign new_new_n35388__ = new_new_n35345__ & new_new_n35368__;
  assign new_new_n35389__ = ~ys__n38453 & new_new_n35388__;
  assign new_new_n35390__ = ~new_new_n35387__ & ~new_new_n35389__;
  assign new_new_n35391__ = ~new_new_n35386__ & new_new_n35390__;
  assign new_new_n35392__ = new_new_n35345__ & new_new_n35362__;
  assign new_new_n35393__ = ~ys__n38453 & new_new_n35392__;
  assign new_new_n35394__ = new_new_n35343__ & new_new_n35368__;
  assign new_new_n35395__ = ~ys__n38453 & new_new_n35394__;
  assign new_new_n35396__ = ~new_new_n35393__ & ~new_new_n35395__;
  assign new_new_n35397__ = new_new_n35323__ & new_new_n35374__;
  assign new_new_n35398__ = ~ys__n38453 & new_new_n35397__;
  assign new_new_n35399__ = new_new_n35396__ & ~new_new_n35398__;
  assign new_new_n35400__ = new_new_n35391__ & new_new_n35399__;
  assign new_new_n35401__ = new_new_n35323__ & new_new_n35362__;
  assign new_new_n35402__ = ~ys__n38453 & new_new_n35401__;
  assign new_new_n35403__ = new_new_n35345__ & new_new_n35359__;
  assign new_new_n35404__ = ~ys__n38453 & new_new_n35403__;
  assign new_new_n35405__ = new_new_n35343__ & new_new_n35374__;
  assign new_new_n35406__ = ~ys__n38453 & new_new_n35405__;
  assign new_new_n35407__ = ~new_new_n35404__ & ~new_new_n35406__;
  assign new_new_n35408__ = ~new_new_n35402__ & new_new_n35407__;
  assign new_new_n35409__ = ys__n38453 & new_new_n35359__;
  assign new_new_n35410__ = new_new_n35345__ & new_new_n35374__;
  assign new_new_n35411__ = ~ys__n38453 & new_new_n35410__;
  assign new_new_n35412__ = ~new_new_n35409__ & ~new_new_n35411__;
  assign new_new_n35413__ = ys__n38453 & new_new_n35374__;
  assign new_new_n35414__ = new_new_n35412__ & ~new_new_n35413__;
  assign new_new_n35415__ = new_new_n35408__ & new_new_n35414__;
  assign new_new_n35416__ = new_new_n35400__ & new_new_n35415__;
  assign new_new_n35417__ = new_new_n35384__ & new_new_n35416__;
  assign new_new_n35418__ = ~new_new_n35379__ & new_new_n35391__;
  assign new_new_n35419__ = ~new_new_n35367__ & ~new_new_n35402__;
  assign new_new_n35420__ = new_new_n35365__ & new_new_n35419__;
  assign new_new_n35421__ = new_new_n35412__ & new_new_n35420__;
  assign new_new_n35422__ = new_new_n35418__ & new_new_n35421__;
  assign new_new_n35423__ = new_new_n11005__ & ~new_new_n35422__;
  assign new_new_n35424__ = ~new_new_n35417__ & new_new_n35423__;
  assign new_new_n35425__ = ~new_new_n35358__ & ~new_new_n35424__;
  assign new_new_n35426__ = ~new_new_n11005__ & ~new_new_n35357__;
  assign new_new_n35427__ = ~ys__n4566 & ~new_new_n35426__;
  assign new_new_n35428__ = ~new_new_n35425__ & new_new_n35427__;
  assign new_new_n35429__ = ~new_new_n35356__ & ~new_new_n35428__;
  assign new_new_n35430__ = ~ys__n738 & ~new_new_n35429__;
  assign new_new_n35431__ = ys__n738 & new_new_n12579__;
  assign new_new_n35432__ = new_new_n35354__ & new_new_n35431__;
  assign ys__n28781 = new_new_n35430__ | new_new_n35432__;
  assign new_new_n35434__ = ys__n190 & ys__n192;
  assign new_new_n35435__ = ~new_new_n10987__ & ~new_new_n35434__;
  assign new_new_n35436__ = new_new_n35345__ & ~new_new_n35435__;
  assign new_new_n35437__ = ~ys__n192 & new_new_n35343__;
  assign new_new_n35438__ = ys__n192 & new_new_n35333__;
  assign new_new_n35439__ = ys__n192 & new_new_n35323__;
  assign new_new_n35440__ = ~new_new_n35438__ & ~new_new_n35439__;
  assign new_new_n35441__ = ~new_new_n35437__ & new_new_n35440__;
  assign new_new_n35442__ = ~new_new_n35436__ & new_new_n35441__;
  assign new_new_n35443__ = ~new_new_n35351__ & ~new_new_n35442__;
  assign new_new_n35444__ = ~new_new_n35330__ & new_new_n35443__;
  assign new_new_n35445__ = ~new_new_n35339__ & new_new_n35444__;
  assign new_new_n35446__ = new_new_n35355__ & new_new_n35445__;
  assign new_new_n35447__ = new_new_n35357__ & new_new_n35445__;
  assign new_new_n35448__ = ~new_new_n35367__ & new_new_n35412__;
  assign new_new_n35449__ = new_new_n35396__ & new_new_n35448__;
  assign new_new_n35450__ = new_new_n35408__ & new_new_n35449__;
  assign new_new_n35451__ = new_new_n35418__ & new_new_n35450__;
  assign new_new_n35452__ = new_new_n11005__ & ~new_new_n35417__;
  assign new_new_n35453__ = ~new_new_n35451__ & new_new_n35452__;
  assign new_new_n35454__ = ~new_new_n35447__ & ~new_new_n35453__;
  assign new_new_n35455__ = new_new_n35427__ & ~new_new_n35454__;
  assign new_new_n35456__ = ~new_new_n35446__ & ~new_new_n35455__;
  assign new_new_n35457__ = ~ys__n738 & ~new_new_n35456__;
  assign new_new_n35458__ = new_new_n35431__ & new_new_n35445__;
  assign ys__n28782 = new_new_n35457__ | new_new_n35458__;
  assign new_new_n35460__ = ys__n190 & ~ys__n192;
  assign new_new_n35461__ = ~ys__n192 & ~new_new_n35460__;
  assign new_new_n35462__ = ys__n204 & ~new_new_n35461__;
  assign new_new_n35463__ = ~ys__n204 & new_new_n35461__;
  assign new_new_n35464__ = ~new_new_n35462__ & ~new_new_n35463__;
  assign new_new_n35465__ = new_new_n35345__ & ~new_new_n35464__;
  assign new_new_n35466__ = ys__n192 & ys__n204;
  assign new_new_n35467__ = ~new_new_n35335__ & ~new_new_n35466__;
  assign new_new_n35468__ = new_new_n35343__ & ~new_new_n35467__;
  assign new_new_n35469__ = ys__n204 & new_new_n35333__;
  assign new_new_n35470__ = ~ys__n204 & new_new_n35323__;
  assign new_new_n35471__ = ~new_new_n35469__ & ~new_new_n35470__;
  assign new_new_n35472__ = ~new_new_n35468__ & new_new_n35471__;
  assign new_new_n35473__ = ~new_new_n35465__ & new_new_n35472__;
  assign new_new_n35474__ = ~new_new_n35330__ & ~new_new_n35351__;
  assign new_new_n35475__ = ~new_new_n35473__ & new_new_n35474__;
  assign new_new_n35476__ = ~new_new_n35339__ & new_new_n35475__;
  assign new_new_n35477__ = new_new_n35355__ & new_new_n35476__;
  assign new_new_n35478__ = new_new_n35357__ & new_new_n35476__;
  assign new_new_n35479__ = new_new_n35365__ & ~new_new_n35370__;
  assign new_new_n35480__ = new_new_n35407__ & new_new_n35412__;
  assign new_new_n35481__ = new_new_n35479__ & new_new_n35480__;
  assign new_new_n35482__ = new_new_n35399__ & new_new_n35481__;
  assign new_new_n35483__ = new_new_n35418__ & new_new_n35482__;
  assign new_new_n35484__ = new_new_n35452__ & ~new_new_n35483__;
  assign new_new_n35485__ = ~new_new_n35478__ & ~new_new_n35484__;
  assign new_new_n35486__ = new_new_n35427__ & ~new_new_n35485__;
  assign new_new_n35487__ = ~new_new_n35477__ & ~new_new_n35486__;
  assign new_new_n35488__ = ~ys__n738 & ~new_new_n35487__;
  assign new_new_n35489__ = new_new_n35431__ & new_new_n35476__;
  assign ys__n28783 = new_new_n35488__ | new_new_n35489__;
  assign new_new_n35491__ = ~ys__n204 & ~new_new_n35461__;
  assign new_new_n35492__ = ~ys__n204 & ~new_new_n35491__;
  assign new_new_n35493__ = ys__n860 & ~new_new_n35492__;
  assign new_new_n35494__ = ~ys__n860 & new_new_n35492__;
  assign new_new_n35495__ = ~new_new_n35493__ & ~new_new_n35494__;
  assign new_new_n35496__ = new_new_n35345__ & ~new_new_n35495__;
  assign new_new_n35497__ = ys__n192 & ~ys__n204;
  assign new_new_n35498__ = ~ys__n204 & ~new_new_n35497__;
  assign new_new_n35499__ = ys__n860 & ~new_new_n35498__;
  assign new_new_n35500__ = ~ys__n860 & new_new_n35498__;
  assign new_new_n35501__ = ~new_new_n35499__ & ~new_new_n35500__;
  assign new_new_n35502__ = new_new_n35343__ & ~new_new_n35501__;
  assign new_new_n35503__ = ~ys__n860 & new_new_n35333__;
  assign new_new_n35504__ = ys__n204 & ys__n860;
  assign new_new_n35505__ = ~new_new_n10988__ & ~new_new_n35504__;
  assign new_new_n35506__ = new_new_n35323__ & ~new_new_n35505__;
  assign new_new_n35507__ = ~new_new_n35503__ & ~new_new_n35506__;
  assign new_new_n35508__ = ~new_new_n35502__ & new_new_n35507__;
  assign new_new_n35509__ = ~new_new_n35496__ & new_new_n35508__;
  assign new_new_n35510__ = ~new_new_n35339__ & new_new_n35474__;
  assign new_new_n35511__ = ~new_new_n35509__ & new_new_n35510__;
  assign new_new_n35512__ = new_new_n35355__ & new_new_n35511__;
  assign new_new_n35513__ = new_new_n35357__ & new_new_n35511__;
  assign new_new_n35514__ = ~new_new_n35370__ & new_new_n35396__;
  assign new_new_n35515__ = ~new_new_n35364__ & ~new_new_n35402__;
  assign new_new_n35516__ = ~new_new_n35381__ & ~new_new_n35413__;
  assign new_new_n35517__ = new_new_n35515__ & new_new_n35516__;
  assign new_new_n35518__ = new_new_n35391__ & new_new_n35517__;
  assign new_new_n35519__ = new_new_n35514__ & new_new_n35518__;
  assign new_new_n35520__ = new_new_n11005__ & ~new_new_n35519__;
  assign new_new_n35521__ = ~new_new_n35417__ & new_new_n35520__;
  assign new_new_n35522__ = ~new_new_n35513__ & ~new_new_n35521__;
  assign new_new_n35523__ = new_new_n35427__ & ~new_new_n35522__;
  assign new_new_n35524__ = ~new_new_n35512__ & ~new_new_n35523__;
  assign new_new_n35525__ = ~ys__n738 & ~new_new_n35524__;
  assign new_new_n35526__ = new_new_n35431__ & new_new_n35511__;
  assign ys__n28784 = new_new_n35525__ | new_new_n35526__;
  assign new_new_n35528__ = ys__n204 & ~ys__n860;
  assign new_new_n35529__ = ~ys__n860 & ~new_new_n35528__;
  assign new_new_n35530__ = new_new_n10988__ & ~new_new_n35461__;
  assign new_new_n35531__ = new_new_n35529__ & ~new_new_n35530__;
  assign new_new_n35532__ = ys__n208 & ~new_new_n35531__;
  assign new_new_n35533__ = ~ys__n208 & new_new_n35531__;
  assign new_new_n35534__ = ~new_new_n35532__ & ~new_new_n35533__;
  assign new_new_n35535__ = new_new_n35345__ & ~new_new_n35534__;
  assign new_new_n35536__ = ys__n192 & new_new_n10988__;
  assign new_new_n35537__ = new_new_n35529__ & ~new_new_n35536__;
  assign new_new_n35538__ = ys__n208 & ~new_new_n35537__;
  assign new_new_n35539__ = ~ys__n208 & new_new_n35537__;
  assign new_new_n35540__ = ~new_new_n35538__ & ~new_new_n35539__;
  assign new_new_n35541__ = new_new_n35343__ & ~new_new_n35540__;
  assign new_new_n35542__ = ~ys__n204 & ys__n860;
  assign new_new_n35543__ = ~new_new_n35504__ & ~new_new_n35542__;
  assign new_new_n35544__ = ys__n208 & ~new_new_n35543__;
  assign new_new_n35545__ = ~ys__n208 & new_new_n35543__;
  assign new_new_n35546__ = ~new_new_n35544__ & ~new_new_n35545__;
  assign new_new_n35547__ = new_new_n35333__ & ~new_new_n35546__;
  assign new_new_n35548__ = ys__n208 & ~new_new_n35529__;
  assign new_new_n35549__ = ~ys__n208 & new_new_n35529__;
  assign new_new_n35550__ = ~new_new_n35548__ & ~new_new_n35549__;
  assign new_new_n35551__ = new_new_n35323__ & ~new_new_n35550__;
  assign new_new_n35552__ = ~new_new_n35547__ & ~new_new_n35551__;
  assign new_new_n35553__ = ~new_new_n35541__ & new_new_n35552__;
  assign new_new_n35554__ = ~new_new_n35535__ & new_new_n35553__;
  assign new_new_n35555__ = new_new_n35510__ & ~new_new_n35554__;
  assign new_new_n35556__ = new_new_n35355__ & new_new_n35555__;
  assign new_new_n35557__ = new_new_n35357__ & new_new_n35555__;
  assign new_new_n35558__ = new_new_n35382__ & new_new_n35515__;
  assign new_new_n35559__ = new_new_n35391__ & new_new_n35558__;
  assign new_new_n35560__ = new_new_n35514__ & new_new_n35559__;
  assign new_new_n35561__ = new_new_n11005__ & ~new_new_n35560__;
  assign new_new_n35562__ = ~new_new_n35417__ & new_new_n35561__;
  assign new_new_n35563__ = ~new_new_n35557__ & ~new_new_n35562__;
  assign new_new_n35564__ = new_new_n35427__ & ~new_new_n35563__;
  assign new_new_n35565__ = ~new_new_n35556__ & ~new_new_n35564__;
  assign new_new_n35566__ = ~ys__n738 & ~new_new_n35565__;
  assign new_new_n35567__ = new_new_n35431__ & new_new_n35555__;
  assign ys__n28785 = new_new_n35566__ | new_new_n35567__;
  assign new_new_n35569__ = ~ys__n208 & ~new_new_n35531__;
  assign new_new_n35570__ = ~ys__n208 & ~new_new_n35569__;
  assign new_new_n35571__ = ys__n206 & ~new_new_n35570__;
  assign new_new_n35572__ = ~ys__n206 & new_new_n35570__;
  assign new_new_n35573__ = ~new_new_n35571__ & ~new_new_n35572__;
  assign new_new_n35574__ = new_new_n35345__ & ~new_new_n35573__;
  assign new_new_n35575__ = ~ys__n208 & ~new_new_n35537__;
  assign new_new_n35576__ = ~ys__n208 & ~new_new_n35575__;
  assign new_new_n35577__ = ys__n206 & ~new_new_n35576__;
  assign new_new_n35578__ = ~ys__n206 & new_new_n35576__;
  assign new_new_n35579__ = ~new_new_n35577__ & ~new_new_n35578__;
  assign new_new_n35580__ = new_new_n35343__ & ~new_new_n35579__;
  assign new_new_n35581__ = ~ys__n208 & ~new_new_n35543__;
  assign new_new_n35582__ = ~ys__n208 & ~new_new_n35581__;
  assign new_new_n35583__ = ys__n206 & ~new_new_n35582__;
  assign new_new_n35584__ = ~ys__n206 & new_new_n35582__;
  assign new_new_n35585__ = ~new_new_n35583__ & ~new_new_n35584__;
  assign new_new_n35586__ = new_new_n35333__ & ~new_new_n35585__;
  assign new_new_n35587__ = ~ys__n208 & ~new_new_n35529__;
  assign new_new_n35588__ = ~ys__n208 & ~new_new_n35587__;
  assign new_new_n35589__ = ys__n206 & ~new_new_n35588__;
  assign new_new_n35590__ = ~ys__n206 & new_new_n35588__;
  assign new_new_n35591__ = ~new_new_n35589__ & ~new_new_n35590__;
  assign new_new_n35592__ = new_new_n35323__ & ~new_new_n35591__;
  assign new_new_n35593__ = ~new_new_n35586__ & ~new_new_n35592__;
  assign new_new_n35594__ = ~new_new_n35580__ & new_new_n35593__;
  assign new_new_n35595__ = ~new_new_n35574__ & new_new_n35594__;
  assign new_new_n35596__ = new_new_n35510__ & ~new_new_n35595__;
  assign new_new_n35597__ = new_new_n35355__ & new_new_n35596__;
  assign new_new_n35598__ = new_new_n35357__ & new_new_n35596__;
  assign new_new_n35599__ = ~new_new_n35361__ & ~new_new_n35367__;
  assign new_new_n35600__ = ~new_new_n35398__ & new_new_n35599__;
  assign new_new_n35601__ = new_new_n35377__ & new_new_n35407__;
  assign new_new_n35602__ = new_new_n35600__ & new_new_n35601__;
  assign new_new_n35603__ = new_new_n35414__ & new_new_n35602__;
  assign new_new_n35604__ = new_new_n11005__ & ~new_new_n35603__;
  assign new_new_n35605__ = ~new_new_n35417__ & new_new_n35604__;
  assign new_new_n35606__ = ~new_new_n35598__ & ~new_new_n35605__;
  assign new_new_n35607__ = new_new_n35427__ & ~new_new_n35606__;
  assign new_new_n35608__ = ~new_new_n35597__ & ~new_new_n35607__;
  assign new_new_n35609__ = ~ys__n738 & ~new_new_n35608__;
  assign new_new_n35610__ = new_new_n35431__ & new_new_n35596__;
  assign ys__n28786 = new_new_n35609__ | new_new_n35610__;
  assign new_new_n35612__ = ys__n47185 & ~new_new_n12582__;
  assign new_new_n35613__ = ys__n46962 & new_new_n35333__;
  assign new_new_n35614__ = ys__n46958 & new_new_n35323__;
  assign new_new_n35615__ = ~new_new_n35613__ & ~new_new_n35614__;
  assign new_new_n35616__ = ys__n46956 & new_new_n35343__;
  assign new_new_n35617__ = ys__n47184 & new_new_n35345__;
  assign new_new_n35618__ = ~new_new_n35616__ & ~new_new_n35617__;
  assign new_new_n35619__ = new_new_n35615__ & new_new_n35618__;
  assign new_new_n35620__ = ~new_new_n35351__ & ~new_new_n35619__;
  assign new_new_n35621__ = new_new_n12582__ & new_new_n35620__;
  assign new_new_n35622__ = ~new_new_n35612__ & ~new_new_n35621__;
  assign new_new_n35623__ = ys__n4566 & ~new_new_n35622__;
  assign new_new_n35624__ = new_new_n10993__ & ~new_new_n11004__;
  assign new_new_n35625__ = ys__n202 & new_new_n35624__;
  assign new_new_n35626__ = ys__n23339 & new_new_n35625__;
  assign new_new_n35627__ = ~ys__n202 & new_new_n35624__;
  assign new_new_n35628__ = ys__n22464 & new_new_n35627__;
  assign new_new_n35629__ = ~new_new_n35626__ & ~new_new_n35628__;
  assign new_new_n35630__ = ys__n202 & ~new_new_n35624__;
  assign new_new_n35631__ = ys__n28243 & new_new_n35630__;
  assign new_new_n35632__ = ~ys__n202 & ~new_new_n35624__;
  assign new_new_n35633__ = ys__n47106 & new_new_n35632__;
  assign new_new_n35634__ = ~new_new_n35631__ & ~new_new_n35633__;
  assign new_new_n35635__ = new_new_n35629__ & new_new_n35634__;
  assign new_new_n35636__ = ~new_new_n35625__ & ~new_new_n35627__;
  assign new_new_n35637__ = ~new_new_n35630__ & ~new_new_n35632__;
  assign new_new_n35638__ = new_new_n35636__ & new_new_n35637__;
  assign new_new_n35639__ = new_new_n11005__ & ~new_new_n35638__;
  assign new_new_n35640__ = ~new_new_n35635__ & new_new_n35639__;
  assign new_new_n35641__ = ys__n47185 & new_new_n12580__;
  assign new_new_n35642__ = new_new_n35357__ & new_new_n35620__;
  assign new_new_n35643__ = ~new_new_n35641__ & ~new_new_n35642__;
  assign new_new_n35644__ = ~new_new_n35640__ & new_new_n35643__;
  assign new_new_n35645__ = ~new_new_n12580__ & new_new_n35426__;
  assign new_new_n35646__ = ~ys__n4566 & ~new_new_n35645__;
  assign new_new_n35647__ = ~new_new_n35644__ & new_new_n35646__;
  assign new_new_n35648__ = ~new_new_n35623__ & ~new_new_n35647__;
  assign new_new_n35649__ = ~ys__n738 & ~new_new_n35648__;
  assign new_new_n35650__ = ys__n47185 & ~new_new_n12579__;
  assign new_new_n35651__ = new_new_n12579__ & new_new_n35620__;
  assign new_new_n35652__ = ~new_new_n35650__ & ~new_new_n35651__;
  assign new_new_n35653__ = ys__n738 & ~new_new_n35652__;
  assign ys__n28787 = new_new_n35649__ | new_new_n35653__;
  assign new_new_n35655__ = ys__n47184 & ~new_new_n12582__;
  assign new_new_n35656__ = ys__n46963 & new_new_n35333__;
  assign new_new_n35657__ = ys__n46959 & new_new_n35323__;
  assign new_new_n35658__ = ~new_new_n35656__ & ~new_new_n35657__;
  assign new_new_n35659__ = ys__n46957 & new_new_n35343__;
  assign new_new_n35660__ = ys__n46956 & new_new_n35345__;
  assign new_new_n35661__ = ~new_new_n35659__ & ~new_new_n35660__;
  assign new_new_n35662__ = new_new_n35658__ & new_new_n35661__;
  assign new_new_n35663__ = ~new_new_n35351__ & ~new_new_n35662__;
  assign new_new_n35664__ = new_new_n12582__ & new_new_n35663__;
  assign new_new_n35665__ = ~new_new_n35655__ & ~new_new_n35664__;
  assign new_new_n35666__ = ys__n4566 & ~new_new_n35665__;
  assign new_new_n35667__ = ys__n22464 & new_new_n35625__;
  assign new_new_n35668__ = ys__n23548 & new_new_n35627__;
  assign new_new_n35669__ = ~new_new_n35667__ & ~new_new_n35668__;
  assign new_new_n35670__ = ys__n47106 & new_new_n35630__;
  assign new_new_n35671__ = ys__n23111 & new_new_n35632__;
  assign new_new_n35672__ = ~new_new_n35670__ & ~new_new_n35671__;
  assign new_new_n35673__ = new_new_n35669__ & new_new_n35672__;
  assign new_new_n35674__ = new_new_n35639__ & ~new_new_n35673__;
  assign new_new_n35675__ = ys__n47184 & new_new_n12580__;
  assign new_new_n35676__ = new_new_n35357__ & new_new_n35663__;
  assign new_new_n35677__ = ~new_new_n35675__ & ~new_new_n35676__;
  assign new_new_n35678__ = ~new_new_n35674__ & new_new_n35677__;
  assign new_new_n35679__ = new_new_n35646__ & ~new_new_n35678__;
  assign new_new_n35680__ = ~new_new_n35666__ & ~new_new_n35679__;
  assign new_new_n35681__ = ~ys__n738 & ~new_new_n35680__;
  assign new_new_n35682__ = ys__n47184 & ~new_new_n12579__;
  assign new_new_n35683__ = new_new_n12579__ & new_new_n35663__;
  assign new_new_n35684__ = ~new_new_n35682__ & ~new_new_n35683__;
  assign new_new_n35685__ = ys__n738 & ~new_new_n35684__;
  assign ys__n28788 = new_new_n35681__ | new_new_n35685__;
  assign new_new_n35687__ = ys__n46956 & ~new_new_n12582__;
  assign new_new_n35688__ = ys__n46964 & new_new_n35333__;
  assign new_new_n35689__ = ys__n46960 & new_new_n35323__;
  assign new_new_n35690__ = ~new_new_n35688__ & ~new_new_n35689__;
  assign new_new_n35691__ = ys__n46958 & new_new_n35343__;
  assign new_new_n35692__ = ys__n46957 & new_new_n35345__;
  assign new_new_n35693__ = ~new_new_n35691__ & ~new_new_n35692__;
  assign new_new_n35694__ = new_new_n35690__ & new_new_n35693__;
  assign new_new_n35695__ = ~new_new_n35351__ & ~new_new_n35694__;
  assign new_new_n35696__ = new_new_n12582__ & new_new_n35695__;
  assign new_new_n35697__ = ~new_new_n35687__ & ~new_new_n35696__;
  assign new_new_n35698__ = ys__n4566 & ~new_new_n35697__;
  assign new_new_n35699__ = ys__n23548 & new_new_n35625__;
  assign new_new_n35700__ = ys__n23550 & new_new_n35627__;
  assign new_new_n35701__ = ~new_new_n35699__ & ~new_new_n35700__;
  assign new_new_n35702__ = ys__n23111 & new_new_n35630__;
  assign new_new_n35703__ = ys__n23114 & new_new_n35632__;
  assign new_new_n35704__ = ~new_new_n35702__ & ~new_new_n35703__;
  assign new_new_n35705__ = new_new_n35701__ & new_new_n35704__;
  assign new_new_n35706__ = new_new_n35639__ & ~new_new_n35705__;
  assign new_new_n35707__ = ys__n46956 & new_new_n12580__;
  assign new_new_n35708__ = new_new_n35357__ & new_new_n35695__;
  assign new_new_n35709__ = ~new_new_n35707__ & ~new_new_n35708__;
  assign new_new_n35710__ = ~new_new_n35706__ & new_new_n35709__;
  assign new_new_n35711__ = new_new_n35646__ & ~new_new_n35710__;
  assign new_new_n35712__ = ~new_new_n35698__ & ~new_new_n35711__;
  assign new_new_n35713__ = ~ys__n738 & ~new_new_n35712__;
  assign new_new_n35714__ = ys__n46956 & ~new_new_n12579__;
  assign new_new_n35715__ = new_new_n12579__ & new_new_n35695__;
  assign new_new_n35716__ = ~new_new_n35714__ & ~new_new_n35715__;
  assign new_new_n35717__ = ys__n738 & ~new_new_n35716__;
  assign ys__n28789 = new_new_n35713__ | new_new_n35717__;
  assign new_new_n35719__ = ys__n46957 & ~new_new_n12582__;
  assign new_new_n35720__ = ys__n46965 & new_new_n35333__;
  assign new_new_n35721__ = ys__n46961 & new_new_n35323__;
  assign new_new_n35722__ = ~new_new_n35720__ & ~new_new_n35721__;
  assign new_new_n35723__ = ys__n46959 & new_new_n35343__;
  assign new_new_n35724__ = ys__n46958 & new_new_n35345__;
  assign new_new_n35725__ = ~new_new_n35723__ & ~new_new_n35724__;
  assign new_new_n35726__ = new_new_n35722__ & new_new_n35725__;
  assign new_new_n35727__ = ~new_new_n35351__ & ~new_new_n35726__;
  assign new_new_n35728__ = new_new_n12582__ & new_new_n35727__;
  assign new_new_n35729__ = ~new_new_n35719__ & ~new_new_n35728__;
  assign new_new_n35730__ = ys__n4566 & ~new_new_n35729__;
  assign new_new_n35731__ = ys__n23550 & new_new_n35625__;
  assign new_new_n35732__ = ys__n23552 & new_new_n35627__;
  assign new_new_n35733__ = ~new_new_n35731__ & ~new_new_n35732__;
  assign new_new_n35734__ = ys__n23114 & new_new_n35630__;
  assign new_new_n35735__ = ys__n23117 & new_new_n35632__;
  assign new_new_n35736__ = ~new_new_n35734__ & ~new_new_n35735__;
  assign new_new_n35737__ = new_new_n35733__ & new_new_n35736__;
  assign new_new_n35738__ = new_new_n35639__ & ~new_new_n35737__;
  assign new_new_n35739__ = ys__n46957 & new_new_n12580__;
  assign new_new_n35740__ = new_new_n35357__ & new_new_n35727__;
  assign new_new_n35741__ = ~new_new_n35739__ & ~new_new_n35740__;
  assign new_new_n35742__ = ~new_new_n35738__ & new_new_n35741__;
  assign new_new_n35743__ = new_new_n35646__ & ~new_new_n35742__;
  assign new_new_n35744__ = ~new_new_n35730__ & ~new_new_n35743__;
  assign new_new_n35745__ = ~ys__n738 & ~new_new_n35744__;
  assign new_new_n35746__ = ys__n46957 & ~new_new_n12579__;
  assign new_new_n35747__ = new_new_n12579__ & new_new_n35727__;
  assign new_new_n35748__ = ~new_new_n35746__ & ~new_new_n35747__;
  assign new_new_n35749__ = ys__n738 & ~new_new_n35748__;
  assign ys__n28790 = new_new_n35745__ | new_new_n35749__;
  assign new_new_n35751__ = ys__n46958 & ~new_new_n12582__;
  assign new_new_n35752__ = ys__n46966 & new_new_n35333__;
  assign new_new_n35753__ = ys__n46962 & new_new_n35323__;
  assign new_new_n35754__ = ~new_new_n35752__ & ~new_new_n35753__;
  assign new_new_n35755__ = ys__n46960 & new_new_n35343__;
  assign new_new_n35756__ = ys__n46959 & new_new_n35345__;
  assign new_new_n35757__ = ~new_new_n35755__ & ~new_new_n35756__;
  assign new_new_n35758__ = new_new_n35754__ & new_new_n35757__;
  assign new_new_n35759__ = ~new_new_n35351__ & ~new_new_n35758__;
  assign new_new_n35760__ = new_new_n12582__ & new_new_n35759__;
  assign new_new_n35761__ = ~new_new_n35751__ & ~new_new_n35760__;
  assign new_new_n35762__ = ys__n4566 & ~new_new_n35761__;
  assign new_new_n35763__ = ys__n23552 & new_new_n35625__;
  assign new_new_n35764__ = ys__n23554 & new_new_n35627__;
  assign new_new_n35765__ = ~new_new_n35763__ & ~new_new_n35764__;
  assign new_new_n35766__ = ys__n23117 & new_new_n35630__;
  assign new_new_n35767__ = ys__n23120 & new_new_n35632__;
  assign new_new_n35768__ = ~new_new_n35766__ & ~new_new_n35767__;
  assign new_new_n35769__ = new_new_n35765__ & new_new_n35768__;
  assign new_new_n35770__ = new_new_n35639__ & ~new_new_n35769__;
  assign new_new_n35771__ = ys__n46958 & new_new_n12580__;
  assign new_new_n35772__ = new_new_n35357__ & new_new_n35759__;
  assign new_new_n35773__ = ~new_new_n35771__ & ~new_new_n35772__;
  assign new_new_n35774__ = ~new_new_n35770__ & new_new_n35773__;
  assign new_new_n35775__ = new_new_n35646__ & ~new_new_n35774__;
  assign new_new_n35776__ = ~new_new_n35762__ & ~new_new_n35775__;
  assign new_new_n35777__ = ~ys__n738 & ~new_new_n35776__;
  assign new_new_n35778__ = ys__n46958 & ~new_new_n12579__;
  assign new_new_n35779__ = new_new_n12579__ & new_new_n35759__;
  assign new_new_n35780__ = ~new_new_n35778__ & ~new_new_n35779__;
  assign new_new_n35781__ = ys__n738 & ~new_new_n35780__;
  assign ys__n28791 = new_new_n35777__ | new_new_n35781__;
  assign new_new_n35783__ = ys__n46959 & ~new_new_n12582__;
  assign new_new_n35784__ = ys__n46967 & new_new_n35333__;
  assign new_new_n35785__ = ys__n46963 & new_new_n35323__;
  assign new_new_n35786__ = ~new_new_n35784__ & ~new_new_n35785__;
  assign new_new_n35787__ = ys__n46961 & new_new_n35343__;
  assign new_new_n35788__ = ys__n46960 & new_new_n35345__;
  assign new_new_n35789__ = ~new_new_n35787__ & ~new_new_n35788__;
  assign new_new_n35790__ = new_new_n35786__ & new_new_n35789__;
  assign new_new_n35791__ = ~new_new_n35351__ & ~new_new_n35790__;
  assign new_new_n35792__ = new_new_n12582__ & new_new_n35791__;
  assign new_new_n35793__ = ~new_new_n35783__ & ~new_new_n35792__;
  assign new_new_n35794__ = ys__n4566 & ~new_new_n35793__;
  assign new_new_n35795__ = ys__n23554 & new_new_n35625__;
  assign new_new_n35796__ = ys__n23556 & new_new_n35627__;
  assign new_new_n35797__ = ~new_new_n35795__ & ~new_new_n35796__;
  assign new_new_n35798__ = ys__n23120 & new_new_n35630__;
  assign new_new_n35799__ = ys__n23123 & new_new_n35632__;
  assign new_new_n35800__ = ~new_new_n35798__ & ~new_new_n35799__;
  assign new_new_n35801__ = new_new_n35797__ & new_new_n35800__;
  assign new_new_n35802__ = new_new_n35639__ & ~new_new_n35801__;
  assign new_new_n35803__ = ys__n46959 & new_new_n12580__;
  assign new_new_n35804__ = new_new_n35357__ & new_new_n35791__;
  assign new_new_n35805__ = ~new_new_n35803__ & ~new_new_n35804__;
  assign new_new_n35806__ = ~new_new_n35802__ & new_new_n35805__;
  assign new_new_n35807__ = new_new_n35646__ & ~new_new_n35806__;
  assign new_new_n35808__ = ~new_new_n35794__ & ~new_new_n35807__;
  assign new_new_n35809__ = ~ys__n738 & ~new_new_n35808__;
  assign new_new_n35810__ = ys__n46959 & ~new_new_n12579__;
  assign new_new_n35811__ = new_new_n12579__ & new_new_n35791__;
  assign new_new_n35812__ = ~new_new_n35810__ & ~new_new_n35811__;
  assign new_new_n35813__ = ys__n738 & ~new_new_n35812__;
  assign ys__n28792 = new_new_n35809__ | new_new_n35813__;
  assign new_new_n35815__ = ys__n46960 & ~new_new_n12582__;
  assign new_new_n35816__ = ys__n46968 & new_new_n35333__;
  assign new_new_n35817__ = ys__n46964 & new_new_n35323__;
  assign new_new_n35818__ = ~new_new_n35816__ & ~new_new_n35817__;
  assign new_new_n35819__ = ys__n46962 & new_new_n35343__;
  assign new_new_n35820__ = ys__n46961 & new_new_n35345__;
  assign new_new_n35821__ = ~new_new_n35819__ & ~new_new_n35820__;
  assign new_new_n35822__ = new_new_n35818__ & new_new_n35821__;
  assign new_new_n35823__ = ~new_new_n35351__ & ~new_new_n35822__;
  assign new_new_n35824__ = new_new_n12582__ & new_new_n35823__;
  assign new_new_n35825__ = ~new_new_n35815__ & ~new_new_n35824__;
  assign new_new_n35826__ = ys__n4566 & ~new_new_n35825__;
  assign new_new_n35827__ = ys__n23556 & new_new_n35625__;
  assign new_new_n35828__ = ys__n23558 & new_new_n35627__;
  assign new_new_n35829__ = ~new_new_n35827__ & ~new_new_n35828__;
  assign new_new_n35830__ = ys__n23123 & new_new_n35630__;
  assign new_new_n35831__ = ys__n23126 & new_new_n35632__;
  assign new_new_n35832__ = ~new_new_n35830__ & ~new_new_n35831__;
  assign new_new_n35833__ = new_new_n35829__ & new_new_n35832__;
  assign new_new_n35834__ = new_new_n35639__ & ~new_new_n35833__;
  assign new_new_n35835__ = ys__n46960 & new_new_n12580__;
  assign new_new_n35836__ = new_new_n35357__ & new_new_n35823__;
  assign new_new_n35837__ = ~new_new_n35835__ & ~new_new_n35836__;
  assign new_new_n35838__ = ~new_new_n35834__ & new_new_n35837__;
  assign new_new_n35839__ = new_new_n35646__ & ~new_new_n35838__;
  assign new_new_n35840__ = ~new_new_n35826__ & ~new_new_n35839__;
  assign new_new_n35841__ = ~ys__n738 & ~new_new_n35840__;
  assign new_new_n35842__ = ys__n46960 & ~new_new_n12579__;
  assign new_new_n35843__ = new_new_n12579__ & new_new_n35823__;
  assign new_new_n35844__ = ~new_new_n35842__ & ~new_new_n35843__;
  assign new_new_n35845__ = ys__n738 & ~new_new_n35844__;
  assign ys__n28793 = new_new_n35841__ | new_new_n35845__;
  assign new_new_n35847__ = ys__n46961 & ~new_new_n12582__;
  assign new_new_n35848__ = ys__n46969 & new_new_n35333__;
  assign new_new_n35849__ = ys__n46965 & new_new_n35323__;
  assign new_new_n35850__ = ~new_new_n35848__ & ~new_new_n35849__;
  assign new_new_n35851__ = ys__n46963 & new_new_n35343__;
  assign new_new_n35852__ = ys__n46962 & new_new_n35345__;
  assign new_new_n35853__ = ~new_new_n35851__ & ~new_new_n35852__;
  assign new_new_n35854__ = new_new_n35850__ & new_new_n35853__;
  assign new_new_n35855__ = ~new_new_n35351__ & ~new_new_n35854__;
  assign new_new_n35856__ = new_new_n12582__ & new_new_n35855__;
  assign new_new_n35857__ = ~new_new_n35847__ & ~new_new_n35856__;
  assign new_new_n35858__ = ys__n4566 & ~new_new_n35857__;
  assign new_new_n35859__ = ys__n23558 & new_new_n35625__;
  assign new_new_n35860__ = ys__n23560 & new_new_n35627__;
  assign new_new_n35861__ = ~new_new_n35859__ & ~new_new_n35860__;
  assign new_new_n35862__ = ys__n23126 & new_new_n35630__;
  assign new_new_n35863__ = ys__n23129 & new_new_n35632__;
  assign new_new_n35864__ = ~new_new_n35862__ & ~new_new_n35863__;
  assign new_new_n35865__ = new_new_n35861__ & new_new_n35864__;
  assign new_new_n35866__ = new_new_n35639__ & ~new_new_n35865__;
  assign new_new_n35867__ = ys__n46961 & new_new_n12580__;
  assign new_new_n35868__ = new_new_n35357__ & new_new_n35855__;
  assign new_new_n35869__ = ~new_new_n35867__ & ~new_new_n35868__;
  assign new_new_n35870__ = ~new_new_n35866__ & new_new_n35869__;
  assign new_new_n35871__ = new_new_n35646__ & ~new_new_n35870__;
  assign new_new_n35872__ = ~new_new_n35858__ & ~new_new_n35871__;
  assign new_new_n35873__ = ~ys__n738 & ~new_new_n35872__;
  assign new_new_n35874__ = ys__n46961 & ~new_new_n12579__;
  assign new_new_n35875__ = new_new_n12579__ & new_new_n35855__;
  assign new_new_n35876__ = ~new_new_n35874__ & ~new_new_n35875__;
  assign new_new_n35877__ = ys__n738 & ~new_new_n35876__;
  assign ys__n28794 = new_new_n35873__ | new_new_n35877__;
  assign new_new_n35879__ = ys__n46970 & new_new_n35333__;
  assign new_new_n35880__ = ys__n46966 & new_new_n35323__;
  assign new_new_n35881__ = ~new_new_n35879__ & ~new_new_n35880__;
  assign new_new_n35882__ = ys__n46964 & new_new_n35343__;
  assign new_new_n35883__ = ys__n46963 & new_new_n35345__;
  assign new_new_n35884__ = ~new_new_n35882__ & ~new_new_n35883__;
  assign new_new_n35885__ = new_new_n35881__ & new_new_n35884__;
  assign new_new_n35886__ = ~new_new_n35351__ & ~new_new_n35885__;
  assign new_new_n35887__ = new_new_n35355__ & new_new_n35886__;
  assign new_new_n35888__ = new_new_n35357__ & new_new_n35886__;
  assign new_new_n35889__ = ys__n23560 & new_new_n35625__;
  assign new_new_n35890__ = ys__n23562 & new_new_n35627__;
  assign new_new_n35891__ = ~new_new_n35889__ & ~new_new_n35890__;
  assign new_new_n35892__ = ys__n23129 & new_new_n35630__;
  assign new_new_n35893__ = ys__n23132 & new_new_n35632__;
  assign new_new_n35894__ = ~new_new_n35892__ & ~new_new_n35893__;
  assign new_new_n35895__ = new_new_n35891__ & new_new_n35894__;
  assign new_new_n35896__ = new_new_n35639__ & ~new_new_n35895__;
  assign new_new_n35897__ = ~new_new_n35888__ & ~new_new_n35896__;
  assign new_new_n35898__ = new_new_n35646__ & ~new_new_n35897__;
  assign new_new_n35899__ = ~new_new_n35887__ & ~new_new_n35898__;
  assign new_new_n35900__ = ~ys__n738 & ~new_new_n35899__;
  assign new_new_n35901__ = new_new_n35431__ & new_new_n35886__;
  assign ys__n28796 = new_new_n35900__ | new_new_n35901__;
  assign new_new_n35903__ = ys__n46971 & new_new_n35333__;
  assign new_new_n35904__ = ys__n46967 & new_new_n35323__;
  assign new_new_n35905__ = ~new_new_n35903__ & ~new_new_n35904__;
  assign new_new_n35906__ = ys__n46965 & new_new_n35343__;
  assign new_new_n35907__ = ys__n46964 & new_new_n35345__;
  assign new_new_n35908__ = ~new_new_n35906__ & ~new_new_n35907__;
  assign new_new_n35909__ = new_new_n35905__ & new_new_n35908__;
  assign new_new_n35910__ = ~new_new_n35351__ & ~new_new_n35909__;
  assign new_new_n35911__ = new_new_n35355__ & new_new_n35910__;
  assign new_new_n35912__ = new_new_n35357__ & new_new_n35910__;
  assign new_new_n35913__ = ys__n23562 & new_new_n35625__;
  assign new_new_n35914__ = ys__n23564 & new_new_n35627__;
  assign new_new_n35915__ = ~new_new_n35913__ & ~new_new_n35914__;
  assign new_new_n35916__ = ys__n23132 & new_new_n35630__;
  assign new_new_n35917__ = ys__n23135 & new_new_n35632__;
  assign new_new_n35918__ = ~new_new_n35916__ & ~new_new_n35917__;
  assign new_new_n35919__ = new_new_n35915__ & new_new_n35918__;
  assign new_new_n35920__ = new_new_n35639__ & ~new_new_n35919__;
  assign new_new_n35921__ = ~new_new_n35912__ & ~new_new_n35920__;
  assign new_new_n35922__ = new_new_n35646__ & ~new_new_n35921__;
  assign new_new_n35923__ = ~new_new_n35911__ & ~new_new_n35922__;
  assign new_new_n35924__ = ~ys__n738 & ~new_new_n35923__;
  assign new_new_n35925__ = new_new_n35431__ & new_new_n35910__;
  assign ys__n28798 = new_new_n35924__ | new_new_n35925__;
  assign new_new_n35927__ = ys__n46972 & new_new_n35333__;
  assign new_new_n35928__ = ys__n46968 & new_new_n35323__;
  assign new_new_n35929__ = ~new_new_n35927__ & ~new_new_n35928__;
  assign new_new_n35930__ = ys__n46966 & new_new_n35343__;
  assign new_new_n35931__ = ys__n46965 & new_new_n35345__;
  assign new_new_n35932__ = ~new_new_n35930__ & ~new_new_n35931__;
  assign new_new_n35933__ = new_new_n35929__ & new_new_n35932__;
  assign new_new_n35934__ = ~new_new_n35351__ & ~new_new_n35933__;
  assign new_new_n35935__ = new_new_n35355__ & new_new_n35934__;
  assign new_new_n35936__ = new_new_n35357__ & new_new_n35934__;
  assign new_new_n35937__ = ys__n23564 & new_new_n35625__;
  assign new_new_n35938__ = ys__n23566 & new_new_n35627__;
  assign new_new_n35939__ = ~new_new_n35937__ & ~new_new_n35938__;
  assign new_new_n35940__ = ys__n23135 & new_new_n35630__;
  assign new_new_n35941__ = ys__n23138 & new_new_n35632__;
  assign new_new_n35942__ = ~new_new_n35940__ & ~new_new_n35941__;
  assign new_new_n35943__ = new_new_n35939__ & new_new_n35942__;
  assign new_new_n35944__ = new_new_n35639__ & ~new_new_n35943__;
  assign new_new_n35945__ = ~new_new_n35936__ & ~new_new_n35944__;
  assign new_new_n35946__ = new_new_n35646__ & ~new_new_n35945__;
  assign new_new_n35947__ = ~new_new_n35935__ & ~new_new_n35946__;
  assign new_new_n35948__ = ~ys__n738 & ~new_new_n35947__;
  assign new_new_n35949__ = new_new_n35431__ & new_new_n35934__;
  assign ys__n28800 = new_new_n35948__ | new_new_n35949__;
  assign new_new_n35951__ = ys__n46973 & new_new_n35333__;
  assign new_new_n35952__ = ys__n46969 & new_new_n35323__;
  assign new_new_n35953__ = ~new_new_n35951__ & ~new_new_n35952__;
  assign new_new_n35954__ = ys__n46967 & new_new_n35343__;
  assign new_new_n35955__ = ys__n46966 & new_new_n35345__;
  assign new_new_n35956__ = ~new_new_n35954__ & ~new_new_n35955__;
  assign new_new_n35957__ = new_new_n35953__ & new_new_n35956__;
  assign new_new_n35958__ = ~new_new_n35351__ & ~new_new_n35957__;
  assign new_new_n35959__ = new_new_n35355__ & new_new_n35958__;
  assign new_new_n35960__ = new_new_n35357__ & new_new_n35958__;
  assign new_new_n35961__ = ys__n23566 & new_new_n35625__;
  assign new_new_n35962__ = ys__n23568 & new_new_n35627__;
  assign new_new_n35963__ = ~new_new_n35961__ & ~new_new_n35962__;
  assign new_new_n35964__ = ys__n23138 & new_new_n35630__;
  assign new_new_n35965__ = ys__n23141 & new_new_n35632__;
  assign new_new_n35966__ = ~new_new_n35964__ & ~new_new_n35965__;
  assign new_new_n35967__ = new_new_n35963__ & new_new_n35966__;
  assign new_new_n35968__ = new_new_n35639__ & ~new_new_n35967__;
  assign new_new_n35969__ = ~new_new_n35960__ & ~new_new_n35968__;
  assign new_new_n35970__ = new_new_n35646__ & ~new_new_n35969__;
  assign new_new_n35971__ = ~new_new_n35959__ & ~new_new_n35970__;
  assign new_new_n35972__ = ~ys__n738 & ~new_new_n35971__;
  assign new_new_n35973__ = new_new_n35431__ & new_new_n35958__;
  assign ys__n28802 = new_new_n35972__ | new_new_n35973__;
  assign new_new_n35975__ = ys__n46974 & new_new_n35333__;
  assign new_new_n35976__ = ys__n46970 & new_new_n35323__;
  assign new_new_n35977__ = ~new_new_n35975__ & ~new_new_n35976__;
  assign new_new_n35978__ = ys__n46968 & new_new_n35343__;
  assign new_new_n35979__ = ys__n46967 & new_new_n35345__;
  assign new_new_n35980__ = ~new_new_n35978__ & ~new_new_n35979__;
  assign new_new_n35981__ = new_new_n35977__ & new_new_n35980__;
  assign new_new_n35982__ = ~new_new_n35351__ & ~new_new_n35981__;
  assign new_new_n35983__ = new_new_n35355__ & new_new_n35982__;
  assign new_new_n35984__ = new_new_n35357__ & new_new_n35982__;
  assign new_new_n35985__ = ys__n23568 & new_new_n35625__;
  assign new_new_n35986__ = ys__n23570 & new_new_n35627__;
  assign new_new_n35987__ = ~new_new_n35985__ & ~new_new_n35986__;
  assign new_new_n35988__ = ys__n23141 & new_new_n35630__;
  assign new_new_n35989__ = ys__n23144 & new_new_n35632__;
  assign new_new_n35990__ = ~new_new_n35988__ & ~new_new_n35989__;
  assign new_new_n35991__ = new_new_n35987__ & new_new_n35990__;
  assign new_new_n35992__ = new_new_n35639__ & ~new_new_n35991__;
  assign new_new_n35993__ = ~new_new_n35984__ & ~new_new_n35992__;
  assign new_new_n35994__ = new_new_n35646__ & ~new_new_n35993__;
  assign new_new_n35995__ = ~new_new_n35983__ & ~new_new_n35994__;
  assign new_new_n35996__ = ~ys__n738 & ~new_new_n35995__;
  assign new_new_n35997__ = new_new_n35431__ & new_new_n35982__;
  assign ys__n28804 = new_new_n35996__ | new_new_n35997__;
  assign new_new_n35999__ = ys__n46975 & new_new_n35333__;
  assign new_new_n36000__ = ys__n46971 & new_new_n35323__;
  assign new_new_n36001__ = ~new_new_n35999__ & ~new_new_n36000__;
  assign new_new_n36002__ = ys__n46969 & new_new_n35343__;
  assign new_new_n36003__ = ys__n46968 & new_new_n35345__;
  assign new_new_n36004__ = ~new_new_n36002__ & ~new_new_n36003__;
  assign new_new_n36005__ = new_new_n36001__ & new_new_n36004__;
  assign new_new_n36006__ = ~new_new_n35351__ & ~new_new_n36005__;
  assign new_new_n36007__ = new_new_n35355__ & new_new_n36006__;
  assign new_new_n36008__ = new_new_n35357__ & new_new_n36006__;
  assign new_new_n36009__ = ys__n23570 & new_new_n35625__;
  assign new_new_n36010__ = ys__n23572 & new_new_n35627__;
  assign new_new_n36011__ = ~new_new_n36009__ & ~new_new_n36010__;
  assign new_new_n36012__ = ys__n23144 & new_new_n35630__;
  assign new_new_n36013__ = ys__n23147 & new_new_n35632__;
  assign new_new_n36014__ = ~new_new_n36012__ & ~new_new_n36013__;
  assign new_new_n36015__ = new_new_n36011__ & new_new_n36014__;
  assign new_new_n36016__ = new_new_n35639__ & ~new_new_n36015__;
  assign new_new_n36017__ = ~new_new_n36008__ & ~new_new_n36016__;
  assign new_new_n36018__ = new_new_n35646__ & ~new_new_n36017__;
  assign new_new_n36019__ = ~new_new_n36007__ & ~new_new_n36018__;
  assign new_new_n36020__ = ~ys__n738 & ~new_new_n36019__;
  assign new_new_n36021__ = new_new_n35431__ & new_new_n36006__;
  assign ys__n28806 = new_new_n36020__ | new_new_n36021__;
  assign new_new_n36023__ = ys__n46976 & new_new_n35333__;
  assign new_new_n36024__ = ys__n46972 & new_new_n35323__;
  assign new_new_n36025__ = ~new_new_n36023__ & ~new_new_n36024__;
  assign new_new_n36026__ = ys__n46970 & new_new_n35343__;
  assign new_new_n36027__ = ys__n46969 & new_new_n35345__;
  assign new_new_n36028__ = ~new_new_n36026__ & ~new_new_n36027__;
  assign new_new_n36029__ = new_new_n36025__ & new_new_n36028__;
  assign new_new_n36030__ = ~new_new_n35351__ & ~new_new_n36029__;
  assign new_new_n36031__ = new_new_n35355__ & new_new_n36030__;
  assign new_new_n36032__ = new_new_n35357__ & new_new_n36030__;
  assign new_new_n36033__ = ys__n23572 & new_new_n35625__;
  assign new_new_n36034__ = ys__n23574 & new_new_n35627__;
  assign new_new_n36035__ = ~new_new_n36033__ & ~new_new_n36034__;
  assign new_new_n36036__ = ys__n23147 & new_new_n35630__;
  assign new_new_n36037__ = ys__n23150 & new_new_n35632__;
  assign new_new_n36038__ = ~new_new_n36036__ & ~new_new_n36037__;
  assign new_new_n36039__ = new_new_n36035__ & new_new_n36038__;
  assign new_new_n36040__ = new_new_n35639__ & ~new_new_n36039__;
  assign new_new_n36041__ = ~new_new_n36032__ & ~new_new_n36040__;
  assign new_new_n36042__ = new_new_n35646__ & ~new_new_n36041__;
  assign new_new_n36043__ = ~new_new_n36031__ & ~new_new_n36042__;
  assign new_new_n36044__ = ~ys__n738 & ~new_new_n36043__;
  assign new_new_n36045__ = new_new_n35431__ & new_new_n36030__;
  assign ys__n28808 = new_new_n36044__ | new_new_n36045__;
  assign new_new_n36047__ = ys__n46977 & new_new_n35333__;
  assign new_new_n36048__ = ys__n46973 & new_new_n35323__;
  assign new_new_n36049__ = ~new_new_n36047__ & ~new_new_n36048__;
  assign new_new_n36050__ = ys__n46971 & new_new_n35343__;
  assign new_new_n36051__ = ys__n46970 & new_new_n35345__;
  assign new_new_n36052__ = ~new_new_n36050__ & ~new_new_n36051__;
  assign new_new_n36053__ = new_new_n36049__ & new_new_n36052__;
  assign new_new_n36054__ = ~new_new_n35351__ & ~new_new_n36053__;
  assign new_new_n36055__ = new_new_n35355__ & new_new_n36054__;
  assign new_new_n36056__ = new_new_n35357__ & new_new_n36054__;
  assign new_new_n36057__ = ys__n23574 & new_new_n35625__;
  assign new_new_n36058__ = ys__n420 & new_new_n35627__;
  assign new_new_n36059__ = ~new_new_n36057__ & ~new_new_n36058__;
  assign new_new_n36060__ = ys__n23150 & new_new_n35630__;
  assign new_new_n36061__ = ys__n23153 & new_new_n35632__;
  assign new_new_n36062__ = ~new_new_n36060__ & ~new_new_n36061__;
  assign new_new_n36063__ = new_new_n36059__ & new_new_n36062__;
  assign new_new_n36064__ = new_new_n35639__ & ~new_new_n36063__;
  assign new_new_n36065__ = ~new_new_n36056__ & ~new_new_n36064__;
  assign new_new_n36066__ = new_new_n35646__ & ~new_new_n36065__;
  assign new_new_n36067__ = ~new_new_n36055__ & ~new_new_n36066__;
  assign new_new_n36068__ = ~ys__n738 & ~new_new_n36067__;
  assign new_new_n36069__ = new_new_n35431__ & new_new_n36054__;
  assign ys__n28810 = new_new_n36068__ | new_new_n36069__;
  assign new_new_n36071__ = ys__n46978 & new_new_n35333__;
  assign new_new_n36072__ = ys__n46974 & new_new_n35323__;
  assign new_new_n36073__ = ~new_new_n36071__ & ~new_new_n36072__;
  assign new_new_n36074__ = ys__n46972 & new_new_n35343__;
  assign new_new_n36075__ = ys__n46971 & new_new_n35345__;
  assign new_new_n36076__ = ~new_new_n36074__ & ~new_new_n36075__;
  assign new_new_n36077__ = new_new_n36073__ & new_new_n36076__;
  assign new_new_n36078__ = ~new_new_n35351__ & ~new_new_n36077__;
  assign new_new_n36079__ = new_new_n35355__ & new_new_n36078__;
  assign new_new_n36080__ = new_new_n35357__ & new_new_n36078__;
  assign new_new_n36081__ = ys__n420 & new_new_n35625__;
  assign new_new_n36082__ = ys__n442 & new_new_n35627__;
  assign new_new_n36083__ = ~new_new_n36081__ & ~new_new_n36082__;
  assign new_new_n36084__ = ys__n23153 & new_new_n35630__;
  assign new_new_n36085__ = ys__n23156 & new_new_n35632__;
  assign new_new_n36086__ = ~new_new_n36084__ & ~new_new_n36085__;
  assign new_new_n36087__ = new_new_n36083__ & new_new_n36086__;
  assign new_new_n36088__ = new_new_n35639__ & ~new_new_n36087__;
  assign new_new_n36089__ = ~new_new_n36080__ & ~new_new_n36088__;
  assign new_new_n36090__ = new_new_n35646__ & ~new_new_n36089__;
  assign new_new_n36091__ = ~new_new_n36079__ & ~new_new_n36090__;
  assign new_new_n36092__ = ~ys__n738 & ~new_new_n36091__;
  assign new_new_n36093__ = new_new_n35431__ & new_new_n36078__;
  assign ys__n28812 = new_new_n36092__ | new_new_n36093__;
  assign new_new_n36095__ = ys__n46979 & new_new_n35333__;
  assign new_new_n36096__ = ys__n46975 & new_new_n35323__;
  assign new_new_n36097__ = ~new_new_n36095__ & ~new_new_n36096__;
  assign new_new_n36098__ = ys__n46973 & new_new_n35343__;
  assign new_new_n36099__ = ys__n46972 & new_new_n35345__;
  assign new_new_n36100__ = ~new_new_n36098__ & ~new_new_n36099__;
  assign new_new_n36101__ = new_new_n36097__ & new_new_n36100__;
  assign new_new_n36102__ = ~new_new_n35351__ & ~new_new_n36101__;
  assign new_new_n36103__ = new_new_n35355__ & new_new_n36102__;
  assign new_new_n36104__ = new_new_n35357__ & new_new_n36102__;
  assign new_new_n36105__ = ys__n442 & new_new_n35625__;
  assign new_new_n36106__ = ys__n440 & new_new_n35627__;
  assign new_new_n36107__ = ~new_new_n36105__ & ~new_new_n36106__;
  assign new_new_n36108__ = ys__n23156 & new_new_n35630__;
  assign new_new_n36109__ = ys__n23159 & new_new_n35632__;
  assign new_new_n36110__ = ~new_new_n36108__ & ~new_new_n36109__;
  assign new_new_n36111__ = new_new_n36107__ & new_new_n36110__;
  assign new_new_n36112__ = new_new_n35639__ & ~new_new_n36111__;
  assign new_new_n36113__ = ~new_new_n36104__ & ~new_new_n36112__;
  assign new_new_n36114__ = new_new_n35646__ & ~new_new_n36113__;
  assign new_new_n36115__ = ~new_new_n36103__ & ~new_new_n36114__;
  assign new_new_n36116__ = ~ys__n738 & ~new_new_n36115__;
  assign new_new_n36117__ = new_new_n35431__ & new_new_n36102__;
  assign ys__n28814 = new_new_n36116__ | new_new_n36117__;
  assign new_new_n36119__ = ys__n46980 & new_new_n35333__;
  assign new_new_n36120__ = ys__n46976 & new_new_n35323__;
  assign new_new_n36121__ = ~new_new_n36119__ & ~new_new_n36120__;
  assign new_new_n36122__ = ys__n46974 & new_new_n35343__;
  assign new_new_n36123__ = ys__n46973 & new_new_n35345__;
  assign new_new_n36124__ = ~new_new_n36122__ & ~new_new_n36123__;
  assign new_new_n36125__ = new_new_n36121__ & new_new_n36124__;
  assign new_new_n36126__ = ~new_new_n35351__ & ~new_new_n36125__;
  assign new_new_n36127__ = new_new_n35355__ & new_new_n36126__;
  assign new_new_n36128__ = new_new_n35357__ & new_new_n36126__;
  assign new_new_n36129__ = ys__n440 & new_new_n35625__;
  assign new_new_n36130__ = ys__n444 & new_new_n35627__;
  assign new_new_n36131__ = ~new_new_n36129__ & ~new_new_n36130__;
  assign new_new_n36132__ = ys__n23159 & new_new_n35630__;
  assign new_new_n36133__ = ys__n23162 & new_new_n35632__;
  assign new_new_n36134__ = ~new_new_n36132__ & ~new_new_n36133__;
  assign new_new_n36135__ = new_new_n36131__ & new_new_n36134__;
  assign new_new_n36136__ = new_new_n35639__ & ~new_new_n36135__;
  assign new_new_n36137__ = ~new_new_n36128__ & ~new_new_n36136__;
  assign new_new_n36138__ = new_new_n35646__ & ~new_new_n36137__;
  assign new_new_n36139__ = ~new_new_n36127__ & ~new_new_n36138__;
  assign new_new_n36140__ = ~ys__n738 & ~new_new_n36139__;
  assign new_new_n36141__ = new_new_n35431__ & new_new_n36126__;
  assign ys__n28816 = new_new_n36140__ | new_new_n36141__;
  assign new_new_n36143__ = ys__n46981 & new_new_n35333__;
  assign new_new_n36144__ = ys__n46977 & new_new_n35323__;
  assign new_new_n36145__ = ~new_new_n36143__ & ~new_new_n36144__;
  assign new_new_n36146__ = ys__n46975 & new_new_n35343__;
  assign new_new_n36147__ = ys__n46974 & new_new_n35345__;
  assign new_new_n36148__ = ~new_new_n36146__ & ~new_new_n36147__;
  assign new_new_n36149__ = new_new_n36145__ & new_new_n36148__;
  assign new_new_n36150__ = ~new_new_n35351__ & ~new_new_n36149__;
  assign new_new_n36151__ = new_new_n35355__ & new_new_n36150__;
  assign new_new_n36152__ = new_new_n35357__ & new_new_n36150__;
  assign new_new_n36153__ = ys__n444 & new_new_n35625__;
  assign new_new_n36154__ = ys__n438 & new_new_n35627__;
  assign new_new_n36155__ = ~new_new_n36153__ & ~new_new_n36154__;
  assign new_new_n36156__ = ys__n23162 & new_new_n35630__;
  assign new_new_n36157__ = ys__n23165 & new_new_n35632__;
  assign new_new_n36158__ = ~new_new_n36156__ & ~new_new_n36157__;
  assign new_new_n36159__ = new_new_n36155__ & new_new_n36158__;
  assign new_new_n36160__ = new_new_n35639__ & ~new_new_n36159__;
  assign new_new_n36161__ = ~new_new_n36152__ & ~new_new_n36160__;
  assign new_new_n36162__ = new_new_n35646__ & ~new_new_n36161__;
  assign new_new_n36163__ = ~new_new_n36151__ & ~new_new_n36162__;
  assign new_new_n36164__ = ~ys__n738 & ~new_new_n36163__;
  assign new_new_n36165__ = new_new_n35431__ & new_new_n36150__;
  assign ys__n28818 = new_new_n36164__ | new_new_n36165__;
  assign new_new_n36167__ = ys__n46982 & new_new_n35333__;
  assign new_new_n36168__ = ys__n46978 & new_new_n35323__;
  assign new_new_n36169__ = ~new_new_n36167__ & ~new_new_n36168__;
  assign new_new_n36170__ = ys__n46976 & new_new_n35343__;
  assign new_new_n36171__ = ys__n46975 & new_new_n35345__;
  assign new_new_n36172__ = ~new_new_n36170__ & ~new_new_n36171__;
  assign new_new_n36173__ = new_new_n36169__ & new_new_n36172__;
  assign new_new_n36174__ = ~new_new_n35351__ & ~new_new_n36173__;
  assign new_new_n36175__ = new_new_n35355__ & new_new_n36174__;
  assign new_new_n36176__ = new_new_n35357__ & new_new_n36174__;
  assign new_new_n36177__ = ys__n438 & new_new_n35625__;
  assign new_new_n36178__ = ys__n446 & new_new_n35627__;
  assign new_new_n36179__ = ~new_new_n36177__ & ~new_new_n36178__;
  assign new_new_n36180__ = ys__n23165 & new_new_n35630__;
  assign new_new_n36181__ = ys__n23168 & new_new_n35632__;
  assign new_new_n36182__ = ~new_new_n36180__ & ~new_new_n36181__;
  assign new_new_n36183__ = new_new_n36179__ & new_new_n36182__;
  assign new_new_n36184__ = new_new_n35639__ & ~new_new_n36183__;
  assign new_new_n36185__ = ~new_new_n36176__ & ~new_new_n36184__;
  assign new_new_n36186__ = new_new_n35646__ & ~new_new_n36185__;
  assign new_new_n36187__ = ~new_new_n36175__ & ~new_new_n36186__;
  assign new_new_n36188__ = ~ys__n738 & ~new_new_n36187__;
  assign new_new_n36189__ = new_new_n35431__ & new_new_n36174__;
  assign ys__n28820 = new_new_n36188__ | new_new_n36189__;
  assign new_new_n36191__ = ys__n46983 & new_new_n35333__;
  assign new_new_n36192__ = ys__n46979 & new_new_n35323__;
  assign new_new_n36193__ = ~new_new_n36191__ & ~new_new_n36192__;
  assign new_new_n36194__ = ys__n46977 & new_new_n35343__;
  assign new_new_n36195__ = ys__n46976 & new_new_n35345__;
  assign new_new_n36196__ = ~new_new_n36194__ & ~new_new_n36195__;
  assign new_new_n36197__ = new_new_n36193__ & new_new_n36196__;
  assign new_new_n36198__ = ~new_new_n35351__ & ~new_new_n36197__;
  assign new_new_n36199__ = new_new_n35355__ & new_new_n36198__;
  assign new_new_n36200__ = new_new_n35357__ & new_new_n36198__;
  assign new_new_n36201__ = ys__n446 & new_new_n35625__;
  assign new_new_n36202__ = ys__n434 & new_new_n35627__;
  assign new_new_n36203__ = ~new_new_n36201__ & ~new_new_n36202__;
  assign new_new_n36204__ = ys__n23168 & new_new_n35630__;
  assign new_new_n36205__ = ys__n23171 & new_new_n35632__;
  assign new_new_n36206__ = ~new_new_n36204__ & ~new_new_n36205__;
  assign new_new_n36207__ = new_new_n36203__ & new_new_n36206__;
  assign new_new_n36208__ = new_new_n35639__ & ~new_new_n36207__;
  assign new_new_n36209__ = ~new_new_n36200__ & ~new_new_n36208__;
  assign new_new_n36210__ = new_new_n35646__ & ~new_new_n36209__;
  assign new_new_n36211__ = ~new_new_n36199__ & ~new_new_n36210__;
  assign new_new_n36212__ = ~ys__n738 & ~new_new_n36211__;
  assign new_new_n36213__ = new_new_n35431__ & new_new_n36198__;
  assign ys__n28822 = new_new_n36212__ | new_new_n36213__;
  assign new_new_n36215__ = ys__n46984 & new_new_n35333__;
  assign new_new_n36216__ = ys__n46980 & new_new_n35323__;
  assign new_new_n36217__ = ~new_new_n36215__ & ~new_new_n36216__;
  assign new_new_n36218__ = ys__n46978 & new_new_n35343__;
  assign new_new_n36219__ = ys__n46977 & new_new_n35345__;
  assign new_new_n36220__ = ~new_new_n36218__ & ~new_new_n36219__;
  assign new_new_n36221__ = new_new_n36217__ & new_new_n36220__;
  assign new_new_n36222__ = ~new_new_n35351__ & ~new_new_n36221__;
  assign new_new_n36223__ = new_new_n35355__ & new_new_n36222__;
  assign new_new_n36224__ = new_new_n35357__ & new_new_n36222__;
  assign new_new_n36225__ = ys__n434 & new_new_n35625__;
  assign new_new_n36226__ = ys__n436 & new_new_n35627__;
  assign new_new_n36227__ = ~new_new_n36225__ & ~new_new_n36226__;
  assign new_new_n36228__ = ys__n23171 & new_new_n35630__;
  assign new_new_n36229__ = ys__n23174 & new_new_n35632__;
  assign new_new_n36230__ = ~new_new_n36228__ & ~new_new_n36229__;
  assign new_new_n36231__ = new_new_n36227__ & new_new_n36230__;
  assign new_new_n36232__ = new_new_n35639__ & ~new_new_n36231__;
  assign new_new_n36233__ = ~new_new_n36224__ & ~new_new_n36232__;
  assign new_new_n36234__ = new_new_n35646__ & ~new_new_n36233__;
  assign new_new_n36235__ = ~new_new_n36223__ & ~new_new_n36234__;
  assign new_new_n36236__ = ~ys__n738 & ~new_new_n36235__;
  assign new_new_n36237__ = new_new_n35431__ & new_new_n36222__;
  assign ys__n28824 = new_new_n36236__ | new_new_n36237__;
  assign new_new_n36239__ = ys__n46985 & new_new_n35333__;
  assign new_new_n36240__ = ys__n46981 & new_new_n35323__;
  assign new_new_n36241__ = ~new_new_n36239__ & ~new_new_n36240__;
  assign new_new_n36242__ = ys__n46979 & new_new_n35343__;
  assign new_new_n36243__ = ys__n46978 & new_new_n35345__;
  assign new_new_n36244__ = ~new_new_n36242__ & ~new_new_n36243__;
  assign new_new_n36245__ = new_new_n36241__ & new_new_n36244__;
  assign new_new_n36246__ = ~new_new_n35351__ & ~new_new_n36245__;
  assign new_new_n36247__ = new_new_n35355__ & new_new_n36246__;
  assign new_new_n36248__ = new_new_n35357__ & new_new_n36246__;
  assign new_new_n36249__ = ys__n436 & new_new_n35625__;
  assign new_new_n36250__ = ys__n432 & new_new_n35627__;
  assign new_new_n36251__ = ~new_new_n36249__ & ~new_new_n36250__;
  assign new_new_n36252__ = ys__n23174 & new_new_n35630__;
  assign new_new_n36253__ = ys__n23177 & new_new_n35632__;
  assign new_new_n36254__ = ~new_new_n36252__ & ~new_new_n36253__;
  assign new_new_n36255__ = new_new_n36251__ & new_new_n36254__;
  assign new_new_n36256__ = new_new_n35639__ & ~new_new_n36255__;
  assign new_new_n36257__ = ~new_new_n36248__ & ~new_new_n36256__;
  assign new_new_n36258__ = new_new_n35646__ & ~new_new_n36257__;
  assign new_new_n36259__ = ~new_new_n36247__ & ~new_new_n36258__;
  assign new_new_n36260__ = ~ys__n738 & ~new_new_n36259__;
  assign new_new_n36261__ = new_new_n35431__ & new_new_n36246__;
  assign ys__n28826 = new_new_n36260__ | new_new_n36261__;
  assign new_new_n36263__ = ys__n46986 & new_new_n35333__;
  assign new_new_n36264__ = ys__n46982 & new_new_n35323__;
  assign new_new_n36265__ = ~new_new_n36263__ & ~new_new_n36264__;
  assign new_new_n36266__ = ys__n46980 & new_new_n35343__;
  assign new_new_n36267__ = ys__n46979 & new_new_n35345__;
  assign new_new_n36268__ = ~new_new_n36266__ & ~new_new_n36267__;
  assign new_new_n36269__ = new_new_n36265__ & new_new_n36268__;
  assign new_new_n36270__ = ~new_new_n35351__ & ~new_new_n36269__;
  assign new_new_n36271__ = new_new_n35355__ & new_new_n36270__;
  assign new_new_n36272__ = new_new_n35357__ & new_new_n36270__;
  assign new_new_n36273__ = ys__n432 & new_new_n35625__;
  assign new_new_n36274__ = ys__n448 & new_new_n35627__;
  assign new_new_n36275__ = ~new_new_n36273__ & ~new_new_n36274__;
  assign new_new_n36276__ = ys__n23177 & new_new_n35630__;
  assign new_new_n36277__ = ys__n23180 & new_new_n35632__;
  assign new_new_n36278__ = ~new_new_n36276__ & ~new_new_n36277__;
  assign new_new_n36279__ = new_new_n36275__ & new_new_n36278__;
  assign new_new_n36280__ = new_new_n35639__ & ~new_new_n36279__;
  assign new_new_n36281__ = ~new_new_n36272__ & ~new_new_n36280__;
  assign new_new_n36282__ = new_new_n35646__ & ~new_new_n36281__;
  assign new_new_n36283__ = ~new_new_n36271__ & ~new_new_n36282__;
  assign new_new_n36284__ = ~ys__n738 & ~new_new_n36283__;
  assign new_new_n36285__ = new_new_n35431__ & new_new_n36270__;
  assign ys__n28828 = new_new_n36284__ | new_new_n36285__;
  assign new_new_n36287__ = ys__n46987 & new_new_n35333__;
  assign new_new_n36288__ = ys__n46983 & new_new_n35323__;
  assign new_new_n36289__ = ~new_new_n36287__ & ~new_new_n36288__;
  assign new_new_n36290__ = ys__n46981 & new_new_n35343__;
  assign new_new_n36291__ = ys__n46980 & new_new_n35345__;
  assign new_new_n36292__ = ~new_new_n36290__ & ~new_new_n36291__;
  assign new_new_n36293__ = new_new_n36289__ & new_new_n36292__;
  assign new_new_n36294__ = ~new_new_n35351__ & ~new_new_n36293__;
  assign new_new_n36295__ = new_new_n35355__ & new_new_n36294__;
  assign new_new_n36296__ = new_new_n35357__ & new_new_n36294__;
  assign new_new_n36297__ = ys__n448 & new_new_n35625__;
  assign new_new_n36298__ = ys__n428 & new_new_n35627__;
  assign new_new_n36299__ = ~new_new_n36297__ & ~new_new_n36298__;
  assign new_new_n36300__ = ys__n23180 & new_new_n35630__;
  assign new_new_n36301__ = ys__n23183 & new_new_n35632__;
  assign new_new_n36302__ = ~new_new_n36300__ & ~new_new_n36301__;
  assign new_new_n36303__ = new_new_n36299__ & new_new_n36302__;
  assign new_new_n36304__ = new_new_n35639__ & ~new_new_n36303__;
  assign new_new_n36305__ = ~new_new_n36296__ & ~new_new_n36304__;
  assign new_new_n36306__ = new_new_n35646__ & ~new_new_n36305__;
  assign new_new_n36307__ = ~new_new_n36295__ & ~new_new_n36306__;
  assign new_new_n36308__ = ~ys__n738 & ~new_new_n36307__;
  assign new_new_n36309__ = new_new_n35431__ & new_new_n36294__;
  assign ys__n28830 = new_new_n36308__ | new_new_n36309__;
  assign new_new_n36311__ = ys__n46988 & new_new_n35333__;
  assign new_new_n36312__ = ys__n46984 & new_new_n35323__;
  assign new_new_n36313__ = ~new_new_n36311__ & ~new_new_n36312__;
  assign new_new_n36314__ = ys__n46982 & new_new_n35343__;
  assign new_new_n36315__ = ys__n46981 & new_new_n35345__;
  assign new_new_n36316__ = ~new_new_n36314__ & ~new_new_n36315__;
  assign new_new_n36317__ = new_new_n36313__ & new_new_n36316__;
  assign new_new_n36318__ = ~new_new_n35351__ & ~new_new_n36317__;
  assign new_new_n36319__ = new_new_n35355__ & new_new_n36318__;
  assign new_new_n36320__ = new_new_n35357__ & new_new_n36318__;
  assign new_new_n36321__ = ys__n428 & new_new_n35625__;
  assign new_new_n36322__ = ys__n430 & new_new_n35627__;
  assign new_new_n36323__ = ~new_new_n36321__ & ~new_new_n36322__;
  assign new_new_n36324__ = ys__n23183 & new_new_n35630__;
  assign new_new_n36325__ = ys__n23186 & new_new_n35632__;
  assign new_new_n36326__ = ~new_new_n36324__ & ~new_new_n36325__;
  assign new_new_n36327__ = new_new_n36323__ & new_new_n36326__;
  assign new_new_n36328__ = new_new_n35639__ & ~new_new_n36327__;
  assign new_new_n36329__ = ~new_new_n36320__ & ~new_new_n36328__;
  assign new_new_n36330__ = new_new_n35646__ & ~new_new_n36329__;
  assign new_new_n36331__ = ~new_new_n36319__ & ~new_new_n36330__;
  assign new_new_n36332__ = ~ys__n738 & ~new_new_n36331__;
  assign new_new_n36333__ = new_new_n35431__ & new_new_n36318__;
  assign ys__n28832 = new_new_n36332__ | new_new_n36333__;
  assign new_new_n36335__ = ys__n46989 & new_new_n35333__;
  assign new_new_n36336__ = ys__n46985 & new_new_n35323__;
  assign new_new_n36337__ = ~new_new_n36335__ & ~new_new_n36336__;
  assign new_new_n36338__ = ys__n46983 & new_new_n35343__;
  assign new_new_n36339__ = ys__n46982 & new_new_n35345__;
  assign new_new_n36340__ = ~new_new_n36338__ & ~new_new_n36339__;
  assign new_new_n36341__ = new_new_n36337__ & new_new_n36340__;
  assign new_new_n36342__ = ~new_new_n35351__ & ~new_new_n36341__;
  assign new_new_n36343__ = new_new_n35355__ & new_new_n36342__;
  assign new_new_n36344__ = new_new_n35357__ & new_new_n36342__;
  assign new_new_n36345__ = ys__n430 & new_new_n35625__;
  assign new_new_n36346__ = ys__n426 & new_new_n35627__;
  assign new_new_n36347__ = ~new_new_n36345__ & ~new_new_n36346__;
  assign new_new_n36348__ = ys__n23186 & new_new_n35630__;
  assign new_new_n36349__ = ys__n23189 & new_new_n35632__;
  assign new_new_n36350__ = ~new_new_n36348__ & ~new_new_n36349__;
  assign new_new_n36351__ = new_new_n36347__ & new_new_n36350__;
  assign new_new_n36352__ = new_new_n35639__ & ~new_new_n36351__;
  assign new_new_n36353__ = ~new_new_n36344__ & ~new_new_n36352__;
  assign new_new_n36354__ = new_new_n35646__ & ~new_new_n36353__;
  assign new_new_n36355__ = ~new_new_n36343__ & ~new_new_n36354__;
  assign new_new_n36356__ = ~ys__n738 & ~new_new_n36355__;
  assign new_new_n36357__ = new_new_n35431__ & new_new_n36342__;
  assign ys__n28834 = new_new_n36356__ | new_new_n36357__;
  assign new_new_n36359__ = ys__n46990 & new_new_n35333__;
  assign new_new_n36360__ = ys__n46986 & new_new_n35323__;
  assign new_new_n36361__ = ~new_new_n36359__ & ~new_new_n36360__;
  assign new_new_n36362__ = ys__n46984 & new_new_n35343__;
  assign new_new_n36363__ = ys__n46983 & new_new_n35345__;
  assign new_new_n36364__ = ~new_new_n36362__ & ~new_new_n36363__;
  assign new_new_n36365__ = new_new_n36361__ & new_new_n36364__;
  assign new_new_n36366__ = ~new_new_n35351__ & ~new_new_n36365__;
  assign new_new_n36367__ = new_new_n35355__ & new_new_n36366__;
  assign new_new_n36368__ = new_new_n35357__ & new_new_n36366__;
  assign new_new_n36369__ = ys__n426 & new_new_n35625__;
  assign new_new_n36370__ = ys__n450 & new_new_n35627__;
  assign new_new_n36371__ = ~new_new_n36369__ & ~new_new_n36370__;
  assign new_new_n36372__ = ys__n23189 & new_new_n35630__;
  assign new_new_n36373__ = ys__n23192 & new_new_n35632__;
  assign new_new_n36374__ = ~new_new_n36372__ & ~new_new_n36373__;
  assign new_new_n36375__ = new_new_n36371__ & new_new_n36374__;
  assign new_new_n36376__ = new_new_n35639__ & ~new_new_n36375__;
  assign new_new_n36377__ = ~new_new_n36368__ & ~new_new_n36376__;
  assign new_new_n36378__ = new_new_n35646__ & ~new_new_n36377__;
  assign new_new_n36379__ = ~new_new_n36367__ & ~new_new_n36378__;
  assign new_new_n36380__ = ~ys__n738 & ~new_new_n36379__;
  assign new_new_n36381__ = new_new_n35431__ & new_new_n36366__;
  assign ys__n28836 = new_new_n36380__ | new_new_n36381__;
  assign new_new_n36383__ = ys__n46991 & new_new_n35333__;
  assign new_new_n36384__ = ys__n46987 & new_new_n35323__;
  assign new_new_n36385__ = ~new_new_n36383__ & ~new_new_n36384__;
  assign new_new_n36386__ = ys__n46985 & new_new_n35343__;
  assign new_new_n36387__ = ys__n46984 & new_new_n35345__;
  assign new_new_n36388__ = ~new_new_n36386__ & ~new_new_n36387__;
  assign new_new_n36389__ = new_new_n36385__ & new_new_n36388__;
  assign new_new_n36390__ = ~new_new_n35351__ & ~new_new_n36389__;
  assign new_new_n36391__ = new_new_n35355__ & new_new_n36390__;
  assign new_new_n36392__ = new_new_n35357__ & new_new_n36390__;
  assign new_new_n36393__ = ys__n450 & new_new_n35625__;
  assign new_new_n36394__ = ys__n424 & new_new_n35627__;
  assign new_new_n36395__ = ~new_new_n36393__ & ~new_new_n36394__;
  assign new_new_n36396__ = ys__n23192 & new_new_n35630__;
  assign new_new_n36397__ = ys__n23195 & new_new_n35632__;
  assign new_new_n36398__ = ~new_new_n36396__ & ~new_new_n36397__;
  assign new_new_n36399__ = new_new_n36395__ & new_new_n36398__;
  assign new_new_n36400__ = new_new_n35639__ & ~new_new_n36399__;
  assign new_new_n36401__ = ~new_new_n36392__ & ~new_new_n36400__;
  assign new_new_n36402__ = new_new_n35646__ & ~new_new_n36401__;
  assign new_new_n36403__ = ~new_new_n36391__ & ~new_new_n36402__;
  assign new_new_n36404__ = ~ys__n738 & ~new_new_n36403__;
  assign new_new_n36405__ = new_new_n35431__ & new_new_n36390__;
  assign ys__n28838 = new_new_n36404__ | new_new_n36405__;
  assign new_new_n36407__ = ys__n46992 & new_new_n35333__;
  assign new_new_n36408__ = ys__n46988 & new_new_n35323__;
  assign new_new_n36409__ = ~new_new_n36407__ & ~new_new_n36408__;
  assign new_new_n36410__ = ys__n46986 & new_new_n35343__;
  assign new_new_n36411__ = ys__n46985 & new_new_n35345__;
  assign new_new_n36412__ = ~new_new_n36410__ & ~new_new_n36411__;
  assign new_new_n36413__ = new_new_n36409__ & new_new_n36412__;
  assign new_new_n36414__ = ~new_new_n35351__ & ~new_new_n36413__;
  assign new_new_n36415__ = new_new_n35355__ & new_new_n36414__;
  assign new_new_n36416__ = new_new_n35357__ & new_new_n36414__;
  assign new_new_n36417__ = ys__n424 & new_new_n35625__;
  assign new_new_n36418__ = ys__n422 & new_new_n35627__;
  assign new_new_n36419__ = ~new_new_n36417__ & ~new_new_n36418__;
  assign new_new_n36420__ = ys__n23195 & new_new_n35630__;
  assign new_new_n36421__ = ys__n23198 & new_new_n35632__;
  assign new_new_n36422__ = ~new_new_n36420__ & ~new_new_n36421__;
  assign new_new_n36423__ = new_new_n36419__ & new_new_n36422__;
  assign new_new_n36424__ = new_new_n35639__ & ~new_new_n36423__;
  assign new_new_n36425__ = ~new_new_n36416__ & ~new_new_n36424__;
  assign new_new_n36426__ = new_new_n35646__ & ~new_new_n36425__;
  assign new_new_n36427__ = ~new_new_n36415__ & ~new_new_n36426__;
  assign new_new_n36428__ = ~ys__n738 & ~new_new_n36427__;
  assign new_new_n36429__ = new_new_n35431__ & new_new_n36414__;
  assign ys__n28840 = new_new_n36428__ | new_new_n36429__;
  assign new_new_n36431__ = ys__n46993 & new_new_n35333__;
  assign new_new_n36432__ = ys__n46989 & new_new_n35323__;
  assign new_new_n36433__ = ~new_new_n36431__ & ~new_new_n36432__;
  assign new_new_n36434__ = ys__n46987 & new_new_n35343__;
  assign new_new_n36435__ = ys__n46986 & new_new_n35345__;
  assign new_new_n36436__ = ~new_new_n36434__ & ~new_new_n36435__;
  assign new_new_n36437__ = new_new_n36433__ & new_new_n36436__;
  assign new_new_n36438__ = ~new_new_n35351__ & ~new_new_n36437__;
  assign new_new_n36439__ = new_new_n35355__ & new_new_n36438__;
  assign new_new_n36440__ = new_new_n35357__ & new_new_n36438__;
  assign new_new_n36441__ = ys__n422 & new_new_n35625__;
  assign new_new_n36442__ = ys__n23198 & new_new_n35630__;
  assign new_new_n36443__ = ~new_new_n36441__ & ~new_new_n36442__;
  assign new_new_n36444__ = new_new_n35639__ & ~new_new_n36443__;
  assign new_new_n36445__ = ~new_new_n36440__ & ~new_new_n36444__;
  assign new_new_n36446__ = new_new_n35646__ & ~new_new_n36445__;
  assign new_new_n36447__ = ~new_new_n36439__ & ~new_new_n36446__;
  assign new_new_n36448__ = ~ys__n738 & ~new_new_n36447__;
  assign new_new_n36449__ = new_new_n35431__ & new_new_n36438__;
  assign ys__n28842 = new_new_n36448__ | new_new_n36449__;
  assign new_new_n36451__ = ys__n46987 & new_new_n35345__;
  assign new_new_n36452__ = ys__n46990 & new_new_n35323__;
  assign new_new_n36453__ = ys__n46988 & new_new_n35343__;
  assign new_new_n36454__ = ~new_new_n36452__ & ~new_new_n36453__;
  assign new_new_n36455__ = ~new_new_n36451__ & new_new_n36454__;
  assign new_new_n36456__ = ~new_new_n35351__ & ~new_new_n36455__;
  assign new_new_n36457__ = new_new_n35355__ & new_new_n36456__;
  assign new_new_n36458__ = ~ys__n4566 & new_new_n36456__;
  assign new_new_n36459__ = new_new_n35357__ & new_new_n36458__;
  assign new_new_n36460__ = ~new_new_n35645__ & new_new_n36459__;
  assign new_new_n36461__ = ~new_new_n36457__ & ~new_new_n36460__;
  assign new_new_n36462__ = ~ys__n738 & ~new_new_n36461__;
  assign new_new_n36463__ = new_new_n35431__ & new_new_n36456__;
  assign ys__n28844 = new_new_n36462__ | new_new_n36463__;
  assign new_new_n36465__ = ys__n46988 & new_new_n35345__;
  assign new_new_n36466__ = ys__n46991 & new_new_n35323__;
  assign new_new_n36467__ = ys__n46989 & new_new_n35343__;
  assign new_new_n36468__ = ~new_new_n36466__ & ~new_new_n36467__;
  assign new_new_n36469__ = ~new_new_n36465__ & new_new_n36468__;
  assign new_new_n36470__ = ~new_new_n35351__ & ~new_new_n36469__;
  assign new_new_n36471__ = new_new_n35355__ & new_new_n36470__;
  assign new_new_n36472__ = ~ys__n4566 & new_new_n36470__;
  assign new_new_n36473__ = new_new_n35357__ & new_new_n36472__;
  assign new_new_n36474__ = ~new_new_n35645__ & new_new_n36473__;
  assign new_new_n36475__ = ~new_new_n36471__ & ~new_new_n36474__;
  assign new_new_n36476__ = ~ys__n738 & ~new_new_n36475__;
  assign new_new_n36477__ = new_new_n35431__ & new_new_n36470__;
  assign ys__n28846 = new_new_n36476__ | new_new_n36477__;
  assign new_new_n36479__ = ys__n46989 & new_new_n35345__;
  assign new_new_n36480__ = ys__n46992 & new_new_n35323__;
  assign new_new_n36481__ = ys__n46990 & new_new_n35343__;
  assign new_new_n36482__ = ~new_new_n36480__ & ~new_new_n36481__;
  assign new_new_n36483__ = ~new_new_n36479__ & new_new_n36482__;
  assign new_new_n36484__ = ~new_new_n35351__ & ~new_new_n36483__;
  assign new_new_n36485__ = new_new_n35355__ & new_new_n36484__;
  assign new_new_n36486__ = ~ys__n4566 & new_new_n36484__;
  assign new_new_n36487__ = new_new_n35357__ & new_new_n36486__;
  assign new_new_n36488__ = ~new_new_n35645__ & new_new_n36487__;
  assign new_new_n36489__ = ~new_new_n36485__ & ~new_new_n36488__;
  assign new_new_n36490__ = ~ys__n738 & ~new_new_n36489__;
  assign new_new_n36491__ = new_new_n35431__ & new_new_n36484__;
  assign ys__n28848 = new_new_n36490__ | new_new_n36491__;
  assign new_new_n36493__ = ys__n46990 & new_new_n35345__;
  assign new_new_n36494__ = ys__n46993 & new_new_n35323__;
  assign new_new_n36495__ = ys__n46991 & new_new_n35343__;
  assign new_new_n36496__ = ~new_new_n36494__ & ~new_new_n36495__;
  assign new_new_n36497__ = ~new_new_n36493__ & new_new_n36496__;
  assign new_new_n36498__ = ~new_new_n35351__ & ~new_new_n36497__;
  assign new_new_n36499__ = new_new_n35355__ & new_new_n36498__;
  assign new_new_n36500__ = ~ys__n4566 & new_new_n36498__;
  assign new_new_n36501__ = new_new_n35357__ & new_new_n36500__;
  assign new_new_n36502__ = ~new_new_n35645__ & new_new_n36501__;
  assign new_new_n36503__ = ~new_new_n36499__ & ~new_new_n36502__;
  assign new_new_n36504__ = ~ys__n738 & ~new_new_n36503__;
  assign new_new_n36505__ = new_new_n35431__ & new_new_n36498__;
  assign ys__n28850 = new_new_n36504__ | new_new_n36505__;
  assign new_new_n36507__ = ys__n46992 & new_new_n35343__;
  assign new_new_n36508__ = ys__n46991 & new_new_n35345__;
  assign new_new_n36509__ = ~new_new_n36507__ & ~new_new_n36508__;
  assign new_new_n36510__ = ~new_new_n35351__ & ~new_new_n36509__;
  assign new_new_n36511__ = ys__n4566 & new_new_n36510__;
  assign new_new_n36512__ = new_new_n12582__ & new_new_n36511__;
  assign new_new_n36513__ = ~ys__n4566 & new_new_n36510__;
  assign new_new_n36514__ = new_new_n35357__ & new_new_n36513__;
  assign new_new_n36515__ = ~new_new_n35645__ & new_new_n36514__;
  assign new_new_n36516__ = ~new_new_n36512__ & ~new_new_n36515__;
  assign new_new_n36517__ = ~ys__n738 & ~new_new_n36516__;
  assign new_new_n36518__ = new_new_n35431__ & new_new_n36510__;
  assign ys__n28852 = new_new_n36517__ | new_new_n36518__;
  assign new_new_n36520__ = ys__n46993 & new_new_n35343__;
  assign new_new_n36521__ = ys__n46992 & new_new_n35345__;
  assign new_new_n36522__ = ~new_new_n36520__ & ~new_new_n36521__;
  assign new_new_n36523__ = ~new_new_n35351__ & ~new_new_n36522__;
  assign new_new_n36524__ = ys__n4566 & new_new_n36523__;
  assign new_new_n36525__ = new_new_n12582__ & new_new_n36524__;
  assign new_new_n36526__ = ~ys__n4566 & new_new_n36523__;
  assign new_new_n36527__ = new_new_n35357__ & new_new_n36526__;
  assign new_new_n36528__ = ~new_new_n35645__ & new_new_n36527__;
  assign new_new_n36529__ = ~new_new_n36525__ & ~new_new_n36528__;
  assign new_new_n36530__ = ~ys__n738 & ~new_new_n36529__;
  assign new_new_n36531__ = new_new_n35431__ & new_new_n36523__;
  assign ys__n28854 = new_new_n36530__ | new_new_n36531__;
  assign new_new_n36533__ = ys__n46993 & new_new_n35345__;
  assign new_new_n36534__ = ~new_new_n35351__ & new_new_n36533__;
  assign new_new_n36535__ = ys__n4566 & new_new_n36534__;
  assign new_new_n36536__ = new_new_n12582__ & new_new_n36535__;
  assign new_new_n36537__ = ~ys__n4566 & new_new_n36534__;
  assign new_new_n36538__ = new_new_n35357__ & new_new_n36537__;
  assign new_new_n36539__ = ~new_new_n35645__ & new_new_n36538__;
  assign new_new_n36540__ = ~new_new_n36536__ & ~new_new_n36539__;
  assign new_new_n36541__ = ~ys__n738 & ~new_new_n36540__;
  assign new_new_n36542__ = new_new_n35431__ & new_new_n36534__;
  assign ys__n28856 = new_new_n36541__ | new_new_n36542__;
  assign new_new_n36544__ = ~ys__n4625 & ~ys__n38494;
  assign new_new_n36545__ = new_new_n12225__ & new_new_n36544__;
  assign new_new_n36546__ = ~new_new_n23122__ & new_new_n36545__;
  assign new_new_n36547__ = ~new_new_n23114__ & ~new_new_n23442__;
  assign new_new_n36548__ = ~new_new_n23443__ & ~new_new_n36547__;
  assign new_new_n36549__ = ~new_new_n36545__ & ~new_new_n36548__;
  assign new_new_n36550__ = ~new_new_n36546__ & ~new_new_n36549__;
  assign new_new_n36551__ = new_new_n12210__ & ~new_new_n36550__;
  assign new_new_n36552__ = ~ys__n740 & ~new_new_n12210__;
  assign new_new_n36553__ = ~new_new_n36550__ & new_new_n36552__;
  assign ys__n29022 = new_new_n36551__ | new_new_n36553__;
  assign new_new_n36555__ = ~new_new_n23141__ & new_new_n36545__;
  assign new_new_n36556__ = ys__n30014 & ~new_new_n23415__;
  assign new_new_n36557__ = ys__n30046 & new_new_n23415__;
  assign new_new_n36558__ = ~new_new_n36556__ & ~new_new_n36557__;
  assign new_new_n36559__ = ~new_new_n23419__ & ~new_new_n36558__;
  assign new_new_n36560__ = ys__n30030 & ~new_new_n23415__;
  assign new_new_n36561__ = ys__n30062 & new_new_n23415__;
  assign new_new_n36562__ = ~new_new_n36560__ & ~new_new_n36561__;
  assign new_new_n36563__ = new_new_n23419__ & ~new_new_n36562__;
  assign new_new_n36564__ = ~new_new_n36559__ & ~new_new_n36563__;
  assign new_new_n36565__ = ~new_new_n23427__ & ~new_new_n36564__;
  assign new_new_n36566__ = ys__n30014 & new_new_n23427__;
  assign new_new_n36567__ = ~new_new_n36565__ & ~new_new_n36566__;
  assign new_new_n36568__ = ~new_new_n23431__ & ~new_new_n36567__;
  assign new_new_n36569__ = new_new_n23442__ & new_new_n36568__;
  assign new_new_n36570__ = new_new_n23133__ & ~new_new_n23442__;
  assign new_new_n36571__ = ~new_new_n36569__ & ~new_new_n36570__;
  assign new_new_n36572__ = ~new_new_n36545__ & ~new_new_n36571__;
  assign new_new_n36573__ = ~new_new_n36555__ & ~new_new_n36572__;
  assign new_new_n36574__ = new_new_n12210__ & ~new_new_n36573__;
  assign new_new_n36575__ = new_new_n36552__ & ~new_new_n36573__;
  assign ys__n29025 = new_new_n36574__ | new_new_n36575__;
  assign new_new_n36577__ = ~new_new_n23160__ & new_new_n36545__;
  assign new_new_n36578__ = ys__n30016 & ~new_new_n23415__;
  assign new_new_n36579__ = ys__n30048 & new_new_n23415__;
  assign new_new_n36580__ = ~new_new_n36578__ & ~new_new_n36579__;
  assign new_new_n36581__ = ~new_new_n23419__ & ~new_new_n36580__;
  assign new_new_n36582__ = ys__n30032 & ~new_new_n23415__;
  assign new_new_n36583__ = ys__n30064 & new_new_n23415__;
  assign new_new_n36584__ = ~new_new_n36582__ & ~new_new_n36583__;
  assign new_new_n36585__ = new_new_n23419__ & ~new_new_n36584__;
  assign new_new_n36586__ = ~new_new_n36581__ & ~new_new_n36585__;
  assign new_new_n36587__ = ~new_new_n23427__ & ~new_new_n36586__;
  assign new_new_n36588__ = ys__n30016 & new_new_n23427__;
  assign new_new_n36589__ = ~new_new_n36587__ & ~new_new_n36588__;
  assign new_new_n36590__ = ~new_new_n23431__ & ~new_new_n36589__;
  assign new_new_n36591__ = new_new_n23442__ & new_new_n36590__;
  assign new_new_n36592__ = new_new_n23152__ & ~new_new_n23442__;
  assign new_new_n36593__ = ~new_new_n36591__ & ~new_new_n36592__;
  assign new_new_n36594__ = ~new_new_n36545__ & ~new_new_n36593__;
  assign new_new_n36595__ = ~new_new_n36577__ & ~new_new_n36594__;
  assign new_new_n36596__ = new_new_n12210__ & ~new_new_n36595__;
  assign new_new_n36597__ = new_new_n36552__ & ~new_new_n36595__;
  assign ys__n29028 = new_new_n36596__ | new_new_n36597__;
  assign new_new_n36599__ = ~new_new_n23179__ & new_new_n36545__;
  assign new_new_n36600__ = ys__n30018 & ~new_new_n23415__;
  assign new_new_n36601__ = ys__n30050 & new_new_n23415__;
  assign new_new_n36602__ = ~new_new_n36600__ & ~new_new_n36601__;
  assign new_new_n36603__ = ~new_new_n23419__ & ~new_new_n36602__;
  assign new_new_n36604__ = ys__n30034 & ~new_new_n23415__;
  assign new_new_n36605__ = ys__n30066 & new_new_n23415__;
  assign new_new_n36606__ = ~new_new_n36604__ & ~new_new_n36605__;
  assign new_new_n36607__ = new_new_n23419__ & ~new_new_n36606__;
  assign new_new_n36608__ = ~new_new_n36603__ & ~new_new_n36607__;
  assign new_new_n36609__ = ~new_new_n23427__ & ~new_new_n36608__;
  assign new_new_n36610__ = ys__n30018 & new_new_n23427__;
  assign new_new_n36611__ = ~new_new_n36609__ & ~new_new_n36610__;
  assign new_new_n36612__ = ~new_new_n23431__ & ~new_new_n36611__;
  assign new_new_n36613__ = new_new_n23442__ & new_new_n36612__;
  assign new_new_n36614__ = new_new_n23171__ & ~new_new_n23442__;
  assign new_new_n36615__ = ~new_new_n36613__ & ~new_new_n36614__;
  assign new_new_n36616__ = ~new_new_n36545__ & ~new_new_n36615__;
  assign new_new_n36617__ = ~new_new_n36599__ & ~new_new_n36616__;
  assign new_new_n36618__ = new_new_n12210__ & ~new_new_n36617__;
  assign new_new_n36619__ = new_new_n36552__ & ~new_new_n36617__;
  assign ys__n29031 = new_new_n36618__ | new_new_n36619__;
  assign new_new_n36621__ = ~new_new_n23198__ & new_new_n36545__;
  assign new_new_n36622__ = ys__n30020 & ~new_new_n23415__;
  assign new_new_n36623__ = ys__n30052 & new_new_n23415__;
  assign new_new_n36624__ = ~new_new_n36622__ & ~new_new_n36623__;
  assign new_new_n36625__ = ~new_new_n23419__ & ~new_new_n36624__;
  assign new_new_n36626__ = ys__n30036 & ~new_new_n23415__;
  assign new_new_n36627__ = ys__n30068 & new_new_n23415__;
  assign new_new_n36628__ = ~new_new_n36626__ & ~new_new_n36627__;
  assign new_new_n36629__ = new_new_n23419__ & ~new_new_n36628__;
  assign new_new_n36630__ = ~new_new_n36625__ & ~new_new_n36629__;
  assign new_new_n36631__ = ~new_new_n23427__ & ~new_new_n36630__;
  assign new_new_n36632__ = ys__n30020 & new_new_n23427__;
  assign new_new_n36633__ = ~new_new_n36631__ & ~new_new_n36632__;
  assign new_new_n36634__ = ~new_new_n23431__ & ~new_new_n36633__;
  assign new_new_n36635__ = new_new_n23442__ & new_new_n36634__;
  assign new_new_n36636__ = new_new_n23190__ & ~new_new_n23442__;
  assign new_new_n36637__ = ~new_new_n36635__ & ~new_new_n36636__;
  assign new_new_n36638__ = ~new_new_n36545__ & ~new_new_n36637__;
  assign new_new_n36639__ = ~new_new_n36621__ & ~new_new_n36638__;
  assign new_new_n36640__ = new_new_n12210__ & ~new_new_n36639__;
  assign new_new_n36641__ = new_new_n36552__ & ~new_new_n36639__;
  assign ys__n29034 = new_new_n36640__ | new_new_n36641__;
  assign new_new_n36643__ = ~new_new_n23217__ & new_new_n36545__;
  assign new_new_n36644__ = ys__n30022 & ~new_new_n23415__;
  assign new_new_n36645__ = ys__n30054 & new_new_n23415__;
  assign new_new_n36646__ = ~new_new_n36644__ & ~new_new_n36645__;
  assign new_new_n36647__ = ~new_new_n23419__ & ~new_new_n36646__;
  assign new_new_n36648__ = ys__n30038 & ~new_new_n23415__;
  assign new_new_n36649__ = ys__n30070 & new_new_n23415__;
  assign new_new_n36650__ = ~new_new_n36648__ & ~new_new_n36649__;
  assign new_new_n36651__ = new_new_n23419__ & ~new_new_n36650__;
  assign new_new_n36652__ = ~new_new_n36647__ & ~new_new_n36651__;
  assign new_new_n36653__ = ~new_new_n23427__ & ~new_new_n36652__;
  assign new_new_n36654__ = ys__n30022 & new_new_n23427__;
  assign new_new_n36655__ = ~new_new_n36653__ & ~new_new_n36654__;
  assign new_new_n36656__ = ~new_new_n23431__ & ~new_new_n36655__;
  assign new_new_n36657__ = new_new_n23442__ & new_new_n36656__;
  assign new_new_n36658__ = new_new_n23209__ & ~new_new_n23442__;
  assign new_new_n36659__ = ~new_new_n36657__ & ~new_new_n36658__;
  assign new_new_n36660__ = ~new_new_n36545__ & ~new_new_n36659__;
  assign new_new_n36661__ = ~new_new_n36643__ & ~new_new_n36660__;
  assign new_new_n36662__ = new_new_n12210__ & ~new_new_n36661__;
  assign new_new_n36663__ = new_new_n36552__ & ~new_new_n36661__;
  assign ys__n29037 = new_new_n36662__ | new_new_n36663__;
  assign new_new_n36665__ = ~new_new_n23236__ & new_new_n36545__;
  assign new_new_n36666__ = ys__n30024 & ~new_new_n23415__;
  assign new_new_n36667__ = ys__n30056 & new_new_n23415__;
  assign new_new_n36668__ = ~new_new_n36666__ & ~new_new_n36667__;
  assign new_new_n36669__ = ~new_new_n23419__ & ~new_new_n36668__;
  assign new_new_n36670__ = ys__n30040 & ~new_new_n23415__;
  assign new_new_n36671__ = ys__n30072 & new_new_n23415__;
  assign new_new_n36672__ = ~new_new_n36670__ & ~new_new_n36671__;
  assign new_new_n36673__ = new_new_n23419__ & ~new_new_n36672__;
  assign new_new_n36674__ = ~new_new_n36669__ & ~new_new_n36673__;
  assign new_new_n36675__ = ~new_new_n23427__ & ~new_new_n36674__;
  assign new_new_n36676__ = ys__n30024 & new_new_n23427__;
  assign new_new_n36677__ = ~new_new_n36675__ & ~new_new_n36676__;
  assign new_new_n36678__ = ~new_new_n23431__ & ~new_new_n36677__;
  assign new_new_n36679__ = new_new_n23442__ & new_new_n36678__;
  assign new_new_n36680__ = new_new_n23228__ & ~new_new_n23442__;
  assign new_new_n36681__ = ~new_new_n36679__ & ~new_new_n36680__;
  assign new_new_n36682__ = ~new_new_n36545__ & ~new_new_n36681__;
  assign new_new_n36683__ = ~new_new_n36665__ & ~new_new_n36682__;
  assign new_new_n36684__ = new_new_n12210__ & ~new_new_n36683__;
  assign new_new_n36685__ = new_new_n36552__ & ~new_new_n36683__;
  assign ys__n29040 = new_new_n36684__ | new_new_n36685__;
  assign new_new_n36687__ = ~new_new_n23255__ & new_new_n36545__;
  assign new_new_n36688__ = ys__n30026 & ~new_new_n23415__;
  assign new_new_n36689__ = ys__n30058 & new_new_n23415__;
  assign new_new_n36690__ = ~new_new_n36688__ & ~new_new_n36689__;
  assign new_new_n36691__ = ~new_new_n23419__ & ~new_new_n36690__;
  assign new_new_n36692__ = ys__n30042 & ~new_new_n23415__;
  assign new_new_n36693__ = ys__n30074 & new_new_n23415__;
  assign new_new_n36694__ = ~new_new_n36692__ & ~new_new_n36693__;
  assign new_new_n36695__ = new_new_n23419__ & ~new_new_n36694__;
  assign new_new_n36696__ = ~new_new_n36691__ & ~new_new_n36695__;
  assign new_new_n36697__ = ~new_new_n23427__ & ~new_new_n36696__;
  assign new_new_n36698__ = ys__n30026 & new_new_n23427__;
  assign new_new_n36699__ = ~new_new_n36697__ & ~new_new_n36698__;
  assign new_new_n36700__ = ~new_new_n23431__ & ~new_new_n36699__;
  assign new_new_n36701__ = new_new_n23442__ & new_new_n36700__;
  assign new_new_n36702__ = new_new_n23247__ & ~new_new_n23442__;
  assign new_new_n36703__ = ~new_new_n36701__ & ~new_new_n36702__;
  assign new_new_n36704__ = ~new_new_n36545__ & ~new_new_n36703__;
  assign new_new_n36705__ = ~new_new_n36687__ & ~new_new_n36704__;
  assign new_new_n36706__ = new_new_n12210__ & ~new_new_n36705__;
  assign new_new_n36707__ = new_new_n36552__ & ~new_new_n36705__;
  assign ys__n29043 = new_new_n36706__ | new_new_n36707__;
  assign new_new_n36709__ = ~new_new_n22936__ & new_new_n36545__;
  assign new_new_n36710__ = ys__n14 & ~ys__n4688;
  assign new_new_n36711__ = ~ys__n14 & ys__n4688;
  assign new_new_n36712__ = ~new_new_n36710__ & ~new_new_n36711__;
  assign new_new_n36713__ = ~ys__n16 & ys__n2693;
  assign new_new_n36714__ = ys__n16 & ~ys__n2693;
  assign new_new_n36715__ = ~new_new_n36713__ & ~new_new_n36714__;
  assign new_new_n36716__ = new_new_n36712__ & ~new_new_n36715__;
  assign new_new_n36717__ = ~new_new_n36712__ & new_new_n36715__;
  assign new_new_n36718__ = ~new_new_n36716__ & ~new_new_n36717__;
  assign new_new_n36719__ = ~new_new_n23423__ & new_new_n36718__;
  assign new_new_n36720__ = ys__n14 & ~ys__n16;
  assign new_new_n36721__ = ~ys__n2693 & new_new_n36720__;
  assign new_new_n36722__ = ~ys__n2693 & ~new_new_n36721__;
  assign new_new_n36723__ = ~ys__n14 & ~ys__n16;
  assign new_new_n36724__ = ~ys__n2693 & new_new_n36723__;
  assign new_new_n36725__ = ~ys__n2693 & ~new_new_n36714__;
  assign new_new_n36726__ = ~new_new_n36721__ & new_new_n36725__;
  assign new_new_n36727__ = ~new_new_n36724__ & new_new_n36726__;
  assign new_new_n36728__ = ~new_new_n36722__ & ~new_new_n36727__;
  assign new_new_n36729__ = ~new_new_n36725__ & ~new_new_n36727__;
  assign new_new_n36730__ = new_new_n36728__ & new_new_n36729__;
  assign new_new_n36731__ = ys__n30074 & new_new_n36730__;
  assign new_new_n36732__ = ~new_new_n36728__ & new_new_n36729__;
  assign new_new_n36733__ = ys__n30058 & new_new_n36732__;
  assign new_new_n36734__ = ~new_new_n36731__ & ~new_new_n36733__;
  assign new_new_n36735__ = new_new_n36728__ & ~new_new_n36729__;
  assign new_new_n36736__ = ys__n30042 & new_new_n36735__;
  assign new_new_n36737__ = ~new_new_n36728__ & ~new_new_n36729__;
  assign new_new_n36738__ = ys__n30026 & new_new_n36737__;
  assign new_new_n36739__ = ~new_new_n36736__ & ~new_new_n36738__;
  assign new_new_n36740__ = new_new_n36734__ & new_new_n36739__;
  assign new_new_n36741__ = ~new_new_n36730__ & ~new_new_n36732__;
  assign new_new_n36742__ = ~new_new_n36735__ & ~new_new_n36737__;
  assign new_new_n36743__ = new_new_n36741__ & new_new_n36742__;
  assign new_new_n36744__ = ys__n38724 & ~new_new_n36743__;
  assign new_new_n36745__ = ~new_new_n36740__ & new_new_n36744__;
  assign new_new_n36746__ = ~new_new_n36718__ & new_new_n36745__;
  assign new_new_n36747__ = ~new_new_n36719__ & ~new_new_n36746__;
  assign new_new_n36748__ = ~new_new_n23427__ & ~new_new_n36747__;
  assign new_new_n36749__ = ys__n30028 & new_new_n23427__;
  assign new_new_n36750__ = ~new_new_n36748__ & ~new_new_n36749__;
  assign new_new_n36751__ = ~new_new_n23431__ & ~new_new_n36750__;
  assign new_new_n36752__ = new_new_n23442__ & new_new_n36751__;
  assign new_new_n36753__ = new_new_n22928__ & ~new_new_n23442__;
  assign new_new_n36754__ = ~new_new_n36752__ & ~new_new_n36753__;
  assign new_new_n36755__ = ~new_new_n36545__ & ~new_new_n36754__;
  assign new_new_n36756__ = ~new_new_n36709__ & ~new_new_n36755__;
  assign new_new_n36757__ = new_new_n12210__ & ~new_new_n36756__;
  assign new_new_n36758__ = new_new_n36552__ & ~new_new_n36756__;
  assign ys__n29046 = new_new_n36757__ | new_new_n36758__;
  assign new_new_n36760__ = ~new_new_n22954__ & new_new_n36545__;
  assign new_new_n36761__ = ~new_new_n36562__ & new_new_n36718__;
  assign new_new_n36762__ = ~new_new_n36746__ & ~new_new_n36761__;
  assign new_new_n36763__ = ~new_new_n23427__ & ~new_new_n36762__;
  assign new_new_n36764__ = ys__n30030 & new_new_n23427__;
  assign new_new_n36765__ = ~new_new_n36763__ & ~new_new_n36764__;
  assign new_new_n36766__ = ~new_new_n23431__ & ~new_new_n36765__;
  assign new_new_n36767__ = new_new_n23442__ & new_new_n36766__;
  assign new_new_n36768__ = new_new_n22946__ & ~new_new_n23442__;
  assign new_new_n36769__ = ~new_new_n36767__ & ~new_new_n36768__;
  assign new_new_n36770__ = ~new_new_n36545__ & ~new_new_n36769__;
  assign new_new_n36771__ = ~new_new_n36760__ & ~new_new_n36770__;
  assign new_new_n36772__ = new_new_n12210__ & ~new_new_n36771__;
  assign new_new_n36773__ = new_new_n36552__ & ~new_new_n36771__;
  assign ys__n29049 = new_new_n36772__ | new_new_n36773__;
  assign new_new_n36775__ = ~new_new_n22972__ & new_new_n36545__;
  assign new_new_n36776__ = ~new_new_n36584__ & new_new_n36718__;
  assign new_new_n36777__ = ~new_new_n36746__ & ~new_new_n36776__;
  assign new_new_n36778__ = ~new_new_n23427__ & ~new_new_n36777__;
  assign new_new_n36779__ = ys__n30032 & new_new_n23427__;
  assign new_new_n36780__ = ~new_new_n36778__ & ~new_new_n36779__;
  assign new_new_n36781__ = ~new_new_n23431__ & ~new_new_n36780__;
  assign new_new_n36782__ = new_new_n23442__ & new_new_n36781__;
  assign new_new_n36783__ = new_new_n22964__ & ~new_new_n23442__;
  assign new_new_n36784__ = ~new_new_n36782__ & ~new_new_n36783__;
  assign new_new_n36785__ = ~new_new_n36545__ & ~new_new_n36784__;
  assign new_new_n36786__ = ~new_new_n36775__ & ~new_new_n36785__;
  assign new_new_n36787__ = new_new_n12210__ & ~new_new_n36786__;
  assign new_new_n36788__ = new_new_n36552__ & ~new_new_n36786__;
  assign ys__n29052 = new_new_n36787__ | new_new_n36788__;
  assign new_new_n36790__ = ~new_new_n22990__ & new_new_n36545__;
  assign new_new_n36791__ = ~new_new_n36606__ & new_new_n36718__;
  assign new_new_n36792__ = ~new_new_n36746__ & ~new_new_n36791__;
  assign new_new_n36793__ = ~new_new_n23427__ & ~new_new_n36792__;
  assign new_new_n36794__ = ys__n30034 & new_new_n23427__;
  assign new_new_n36795__ = ~new_new_n36793__ & ~new_new_n36794__;
  assign new_new_n36796__ = ~new_new_n23431__ & ~new_new_n36795__;
  assign new_new_n36797__ = new_new_n23442__ & new_new_n36796__;
  assign new_new_n36798__ = new_new_n22982__ & ~new_new_n23442__;
  assign new_new_n36799__ = ~new_new_n36797__ & ~new_new_n36798__;
  assign new_new_n36800__ = ~new_new_n36545__ & ~new_new_n36799__;
  assign new_new_n36801__ = ~new_new_n36790__ & ~new_new_n36800__;
  assign new_new_n36802__ = new_new_n12210__ & ~new_new_n36801__;
  assign new_new_n36803__ = new_new_n36552__ & ~new_new_n36801__;
  assign ys__n29055 = new_new_n36802__ | new_new_n36803__;
  assign new_new_n36805__ = ~new_new_n23008__ & new_new_n36545__;
  assign new_new_n36806__ = ~new_new_n36628__ & new_new_n36718__;
  assign new_new_n36807__ = ~new_new_n36746__ & ~new_new_n36806__;
  assign new_new_n36808__ = ~new_new_n23427__ & ~new_new_n36807__;
  assign new_new_n36809__ = ys__n30036 & new_new_n23427__;
  assign new_new_n36810__ = ~new_new_n36808__ & ~new_new_n36809__;
  assign new_new_n36811__ = ~new_new_n23431__ & ~new_new_n36810__;
  assign new_new_n36812__ = new_new_n23442__ & new_new_n36811__;
  assign new_new_n36813__ = new_new_n23000__ & ~new_new_n23442__;
  assign new_new_n36814__ = ~new_new_n36812__ & ~new_new_n36813__;
  assign new_new_n36815__ = ~new_new_n36545__ & ~new_new_n36814__;
  assign new_new_n36816__ = ~new_new_n36805__ & ~new_new_n36815__;
  assign new_new_n36817__ = new_new_n12210__ & ~new_new_n36816__;
  assign new_new_n36818__ = new_new_n36552__ & ~new_new_n36816__;
  assign ys__n29058 = new_new_n36817__ | new_new_n36818__;
  assign new_new_n36820__ = ~new_new_n23026__ & new_new_n36545__;
  assign new_new_n36821__ = ~new_new_n36650__ & new_new_n36718__;
  assign new_new_n36822__ = ~new_new_n36746__ & ~new_new_n36821__;
  assign new_new_n36823__ = ~new_new_n23427__ & ~new_new_n36822__;
  assign new_new_n36824__ = ys__n30038 & new_new_n23427__;
  assign new_new_n36825__ = ~new_new_n36823__ & ~new_new_n36824__;
  assign new_new_n36826__ = ~new_new_n23431__ & ~new_new_n36825__;
  assign new_new_n36827__ = new_new_n23442__ & new_new_n36826__;
  assign new_new_n36828__ = new_new_n23018__ & ~new_new_n23442__;
  assign new_new_n36829__ = ~new_new_n36827__ & ~new_new_n36828__;
  assign new_new_n36830__ = ~new_new_n36545__ & ~new_new_n36829__;
  assign new_new_n36831__ = ~new_new_n36820__ & ~new_new_n36830__;
  assign new_new_n36832__ = new_new_n12210__ & ~new_new_n36831__;
  assign new_new_n36833__ = new_new_n36552__ & ~new_new_n36831__;
  assign ys__n29061 = new_new_n36832__ | new_new_n36833__;
  assign new_new_n36835__ = ~new_new_n23044__ & new_new_n36545__;
  assign new_new_n36836__ = ~new_new_n36672__ & new_new_n36718__;
  assign new_new_n36837__ = ~new_new_n36746__ & ~new_new_n36836__;
  assign new_new_n36838__ = ~new_new_n23427__ & ~new_new_n36837__;
  assign new_new_n36839__ = ys__n30040 & new_new_n23427__;
  assign new_new_n36840__ = ~new_new_n36838__ & ~new_new_n36839__;
  assign new_new_n36841__ = ~new_new_n23431__ & ~new_new_n36840__;
  assign new_new_n36842__ = new_new_n23442__ & new_new_n36841__;
  assign new_new_n36843__ = new_new_n23036__ & ~new_new_n23442__;
  assign new_new_n36844__ = ~new_new_n36842__ & ~new_new_n36843__;
  assign new_new_n36845__ = ~new_new_n36545__ & ~new_new_n36844__;
  assign new_new_n36846__ = ~new_new_n36835__ & ~new_new_n36845__;
  assign new_new_n36847__ = new_new_n12210__ & ~new_new_n36846__;
  assign new_new_n36848__ = new_new_n36552__ & ~new_new_n36846__;
  assign ys__n29064 = new_new_n36847__ | new_new_n36848__;
  assign new_new_n36850__ = ~new_new_n23062__ & new_new_n36545__;
  assign new_new_n36851__ = ~new_new_n36694__ & new_new_n36718__;
  assign new_new_n36852__ = ~new_new_n36746__ & ~new_new_n36851__;
  assign new_new_n36853__ = ~new_new_n23427__ & ~new_new_n36852__;
  assign new_new_n36854__ = ys__n30042 & new_new_n23427__;
  assign new_new_n36855__ = ~new_new_n36853__ & ~new_new_n36854__;
  assign new_new_n36856__ = ~new_new_n23431__ & ~new_new_n36855__;
  assign new_new_n36857__ = new_new_n23442__ & new_new_n36856__;
  assign new_new_n36858__ = new_new_n23054__ & ~new_new_n23442__;
  assign new_new_n36859__ = ~new_new_n36857__ & ~new_new_n36858__;
  assign new_new_n36860__ = ~new_new_n36545__ & ~new_new_n36859__;
  assign new_new_n36861__ = ~new_new_n36850__ & ~new_new_n36860__;
  assign new_new_n36862__ = new_new_n12210__ & ~new_new_n36861__;
  assign new_new_n36863__ = new_new_n36552__ & ~new_new_n36861__;
  assign ys__n29067 = new_new_n36862__ | new_new_n36863__;
  assign new_new_n36865__ = ~new_new_n22776__ & new_new_n36545__;
  assign new_new_n36866__ = ys__n14 & ys__n16;
  assign new_new_n36867__ = ys__n2693 & ys__n4688;
  assign new_new_n36868__ = new_new_n36866__ & new_new_n36867__;
  assign new_new_n36869__ = ys__n30044 & new_new_n36868__;
  assign new_new_n36870__ = new_new_n36745__ & ~new_new_n36868__;
  assign new_new_n36871__ = ~new_new_n36869__ & ~new_new_n36870__;
  assign new_new_n36872__ = ~new_new_n23427__ & ~new_new_n36871__;
  assign new_new_n36873__ = ys__n30044 & new_new_n23427__;
  assign new_new_n36874__ = ~new_new_n36872__ & ~new_new_n36873__;
  assign new_new_n36875__ = ~new_new_n23431__ & ~new_new_n36874__;
  assign new_new_n36876__ = new_new_n23442__ & new_new_n36875__;
  assign new_new_n36877__ = new_new_n22768__ & ~new_new_n23442__;
  assign new_new_n36878__ = ~new_new_n36876__ & ~new_new_n36877__;
  assign new_new_n36879__ = ~new_new_n36545__ & ~new_new_n36878__;
  assign new_new_n36880__ = ~new_new_n36865__ & ~new_new_n36879__;
  assign new_new_n36881__ = new_new_n12210__ & ~new_new_n36880__;
  assign new_new_n36882__ = new_new_n36552__ & ~new_new_n36880__;
  assign ys__n29070 = new_new_n36881__ | new_new_n36882__;
  assign new_new_n36884__ = ~new_new_n22791__ & new_new_n36545__;
  assign new_new_n36885__ = ys__n30046 & new_new_n36868__;
  assign new_new_n36886__ = ~new_new_n36870__ & ~new_new_n36885__;
  assign new_new_n36887__ = ~new_new_n23427__ & ~new_new_n36886__;
  assign new_new_n36888__ = ys__n30046 & new_new_n23427__;
  assign new_new_n36889__ = ~new_new_n36887__ & ~new_new_n36888__;
  assign new_new_n36890__ = ~new_new_n23431__ & ~new_new_n36889__;
  assign new_new_n36891__ = new_new_n23442__ & new_new_n36890__;
  assign new_new_n36892__ = new_new_n22783__ & ~new_new_n23442__;
  assign new_new_n36893__ = ~new_new_n36891__ & ~new_new_n36892__;
  assign new_new_n36894__ = ~new_new_n36545__ & ~new_new_n36893__;
  assign new_new_n36895__ = ~new_new_n36884__ & ~new_new_n36894__;
  assign new_new_n36896__ = new_new_n12210__ & ~new_new_n36895__;
  assign new_new_n36897__ = new_new_n36552__ & ~new_new_n36895__;
  assign ys__n29073 = new_new_n36896__ | new_new_n36897__;
  assign new_new_n36899__ = ~new_new_n22806__ & new_new_n36545__;
  assign new_new_n36900__ = ys__n30048 & new_new_n36868__;
  assign new_new_n36901__ = ~new_new_n36870__ & ~new_new_n36900__;
  assign new_new_n36902__ = ~new_new_n23427__ & ~new_new_n36901__;
  assign new_new_n36903__ = ys__n30048 & new_new_n23427__;
  assign new_new_n36904__ = ~new_new_n36902__ & ~new_new_n36903__;
  assign new_new_n36905__ = ~new_new_n23431__ & ~new_new_n36904__;
  assign new_new_n36906__ = new_new_n23442__ & new_new_n36905__;
  assign new_new_n36907__ = new_new_n22798__ & ~new_new_n23442__;
  assign new_new_n36908__ = ~new_new_n36906__ & ~new_new_n36907__;
  assign new_new_n36909__ = ~new_new_n36545__ & ~new_new_n36908__;
  assign new_new_n36910__ = ~new_new_n36899__ & ~new_new_n36909__;
  assign new_new_n36911__ = new_new_n12210__ & ~new_new_n36910__;
  assign new_new_n36912__ = new_new_n36552__ & ~new_new_n36910__;
  assign ys__n29076 = new_new_n36911__ | new_new_n36912__;
  assign new_new_n36914__ = ~new_new_n22821__ & new_new_n36545__;
  assign new_new_n36915__ = ys__n30050 & new_new_n36868__;
  assign new_new_n36916__ = ~new_new_n36870__ & ~new_new_n36915__;
  assign new_new_n36917__ = ~new_new_n23427__ & ~new_new_n36916__;
  assign new_new_n36918__ = ys__n30050 & new_new_n23427__;
  assign new_new_n36919__ = ~new_new_n36917__ & ~new_new_n36918__;
  assign new_new_n36920__ = ~new_new_n23431__ & ~new_new_n36919__;
  assign new_new_n36921__ = new_new_n23442__ & new_new_n36920__;
  assign new_new_n36922__ = new_new_n22813__ & ~new_new_n23442__;
  assign new_new_n36923__ = ~new_new_n36921__ & ~new_new_n36922__;
  assign new_new_n36924__ = ~new_new_n36545__ & ~new_new_n36923__;
  assign new_new_n36925__ = ~new_new_n36914__ & ~new_new_n36924__;
  assign new_new_n36926__ = new_new_n12210__ & ~new_new_n36925__;
  assign new_new_n36927__ = new_new_n36552__ & ~new_new_n36925__;
  assign ys__n29079 = new_new_n36926__ | new_new_n36927__;
  assign new_new_n36929__ = ~new_new_n22836__ & new_new_n36545__;
  assign new_new_n36930__ = ys__n30052 & new_new_n36868__;
  assign new_new_n36931__ = ~new_new_n36870__ & ~new_new_n36930__;
  assign new_new_n36932__ = ~new_new_n23427__ & ~new_new_n36931__;
  assign new_new_n36933__ = ys__n30052 & new_new_n23427__;
  assign new_new_n36934__ = ~new_new_n36932__ & ~new_new_n36933__;
  assign new_new_n36935__ = ~new_new_n23431__ & ~new_new_n36934__;
  assign new_new_n36936__ = new_new_n23442__ & new_new_n36935__;
  assign new_new_n36937__ = new_new_n22828__ & ~new_new_n23442__;
  assign new_new_n36938__ = ~new_new_n36936__ & ~new_new_n36937__;
  assign new_new_n36939__ = ~new_new_n36545__ & ~new_new_n36938__;
  assign new_new_n36940__ = ~new_new_n36929__ & ~new_new_n36939__;
  assign new_new_n36941__ = new_new_n12210__ & ~new_new_n36940__;
  assign new_new_n36942__ = new_new_n36552__ & ~new_new_n36940__;
  assign ys__n29082 = new_new_n36941__ | new_new_n36942__;
  assign new_new_n36944__ = ~new_new_n22851__ & new_new_n36545__;
  assign new_new_n36945__ = ys__n30054 & new_new_n36868__;
  assign new_new_n36946__ = ~new_new_n36870__ & ~new_new_n36945__;
  assign new_new_n36947__ = ~new_new_n23427__ & ~new_new_n36946__;
  assign new_new_n36948__ = ys__n30054 & new_new_n23427__;
  assign new_new_n36949__ = ~new_new_n36947__ & ~new_new_n36948__;
  assign new_new_n36950__ = ~new_new_n23431__ & ~new_new_n36949__;
  assign new_new_n36951__ = new_new_n23442__ & new_new_n36950__;
  assign new_new_n36952__ = new_new_n22843__ & ~new_new_n23442__;
  assign new_new_n36953__ = ~new_new_n36951__ & ~new_new_n36952__;
  assign new_new_n36954__ = ~new_new_n36545__ & ~new_new_n36953__;
  assign new_new_n36955__ = ~new_new_n36944__ & ~new_new_n36954__;
  assign new_new_n36956__ = new_new_n12210__ & ~new_new_n36955__;
  assign new_new_n36957__ = new_new_n36552__ & ~new_new_n36955__;
  assign ys__n29085 = new_new_n36956__ | new_new_n36957__;
  assign new_new_n36959__ = ~new_new_n22866__ & new_new_n36545__;
  assign new_new_n36960__ = ys__n30056 & new_new_n36868__;
  assign new_new_n36961__ = ~new_new_n36870__ & ~new_new_n36960__;
  assign new_new_n36962__ = ~new_new_n23427__ & ~new_new_n36961__;
  assign new_new_n36963__ = ys__n30056 & new_new_n23427__;
  assign new_new_n36964__ = ~new_new_n36962__ & ~new_new_n36963__;
  assign new_new_n36965__ = ~new_new_n23431__ & ~new_new_n36964__;
  assign new_new_n36966__ = new_new_n23442__ & new_new_n36965__;
  assign new_new_n36967__ = new_new_n22858__ & ~new_new_n23442__;
  assign new_new_n36968__ = ~new_new_n36966__ & ~new_new_n36967__;
  assign new_new_n36969__ = ~new_new_n36545__ & ~new_new_n36968__;
  assign new_new_n36970__ = ~new_new_n36959__ & ~new_new_n36969__;
  assign new_new_n36971__ = new_new_n12210__ & ~new_new_n36970__;
  assign new_new_n36972__ = new_new_n36552__ & ~new_new_n36970__;
  assign ys__n29088 = new_new_n36971__ | new_new_n36972__;
  assign new_new_n36974__ = ~new_new_n22881__ & new_new_n36545__;
  assign new_new_n36975__ = ys__n30058 & new_new_n36868__;
  assign new_new_n36976__ = ~new_new_n36870__ & ~new_new_n36975__;
  assign new_new_n36977__ = ~new_new_n23427__ & ~new_new_n36976__;
  assign new_new_n36978__ = ys__n30058 & new_new_n23427__;
  assign new_new_n36979__ = ~new_new_n36977__ & ~new_new_n36978__;
  assign new_new_n36980__ = ~new_new_n23431__ & ~new_new_n36979__;
  assign new_new_n36981__ = new_new_n23442__ & new_new_n36980__;
  assign new_new_n36982__ = new_new_n22873__ & ~new_new_n23442__;
  assign new_new_n36983__ = ~new_new_n36981__ & ~new_new_n36982__;
  assign new_new_n36984__ = ~new_new_n36545__ & ~new_new_n36983__;
  assign new_new_n36985__ = ~new_new_n36974__ & ~new_new_n36984__;
  assign new_new_n36986__ = new_new_n12210__ & ~new_new_n36985__;
  assign new_new_n36987__ = new_new_n36552__ & ~new_new_n36985__;
  assign ys__n29091 = new_new_n36986__ | new_new_n36987__;
  assign new_new_n36989__ = ~new_new_n22628__ & new_new_n36545__;
  assign new_new_n36990__ = ys__n30060 & new_new_n36868__;
  assign new_new_n36991__ = ~new_new_n36870__ & ~new_new_n36990__;
  assign new_new_n36992__ = ~new_new_n23427__ & ~new_new_n36991__;
  assign new_new_n36993__ = ys__n30060 & new_new_n23427__;
  assign new_new_n36994__ = ~new_new_n36992__ & ~new_new_n36993__;
  assign new_new_n36995__ = ~new_new_n23431__ & ~new_new_n36994__;
  assign new_new_n36996__ = new_new_n23442__ & new_new_n36995__;
  assign new_new_n36997__ = new_new_n22614__ & ~new_new_n23442__;
  assign new_new_n36998__ = ~new_new_n36996__ & ~new_new_n36997__;
  assign new_new_n36999__ = ~new_new_n36545__ & ~new_new_n36998__;
  assign new_new_n37000__ = ~new_new_n36989__ & ~new_new_n36999__;
  assign new_new_n37001__ = new_new_n12210__ & ~new_new_n37000__;
  assign new_new_n37002__ = new_new_n36552__ & ~new_new_n37000__;
  assign ys__n29094 = new_new_n37001__ | new_new_n37002__;
  assign new_new_n37004__ = ~new_new_n22643__ & new_new_n36545__;
  assign new_new_n37005__ = ys__n30062 & new_new_n36868__;
  assign new_new_n37006__ = ~new_new_n36870__ & ~new_new_n37005__;
  assign new_new_n37007__ = ~new_new_n23427__ & ~new_new_n37006__;
  assign new_new_n37008__ = ys__n30062 & new_new_n23427__;
  assign new_new_n37009__ = ~new_new_n37007__ & ~new_new_n37008__;
  assign new_new_n37010__ = ~new_new_n23431__ & ~new_new_n37009__;
  assign new_new_n37011__ = new_new_n23442__ & new_new_n37010__;
  assign new_new_n37012__ = new_new_n22635__ & ~new_new_n23442__;
  assign new_new_n37013__ = ~new_new_n37011__ & ~new_new_n37012__;
  assign new_new_n37014__ = ~new_new_n36545__ & ~new_new_n37013__;
  assign new_new_n37015__ = ~new_new_n37004__ & ~new_new_n37014__;
  assign new_new_n37016__ = new_new_n12210__ & ~new_new_n37015__;
  assign new_new_n37017__ = new_new_n36552__ & ~new_new_n37015__;
  assign ys__n29097 = new_new_n37016__ | new_new_n37017__;
  assign new_new_n37019__ = ~new_new_n22658__ & new_new_n36545__;
  assign new_new_n37020__ = ys__n30064 & new_new_n36868__;
  assign new_new_n37021__ = ~new_new_n36870__ & ~new_new_n37020__;
  assign new_new_n37022__ = ~new_new_n23427__ & ~new_new_n37021__;
  assign new_new_n37023__ = ys__n30064 & new_new_n23427__;
  assign new_new_n37024__ = ~new_new_n37022__ & ~new_new_n37023__;
  assign new_new_n37025__ = ~new_new_n23431__ & ~new_new_n37024__;
  assign new_new_n37026__ = new_new_n23442__ & new_new_n37025__;
  assign new_new_n37027__ = new_new_n22650__ & ~new_new_n23442__;
  assign new_new_n37028__ = ~new_new_n37026__ & ~new_new_n37027__;
  assign new_new_n37029__ = ~new_new_n36545__ & ~new_new_n37028__;
  assign new_new_n37030__ = ~new_new_n37019__ & ~new_new_n37029__;
  assign new_new_n37031__ = new_new_n12210__ & ~new_new_n37030__;
  assign new_new_n37032__ = new_new_n36552__ & ~new_new_n37030__;
  assign ys__n29100 = new_new_n37031__ | new_new_n37032__;
  assign new_new_n37034__ = ~new_new_n22673__ & new_new_n36545__;
  assign new_new_n37035__ = ys__n30066 & new_new_n36868__;
  assign new_new_n37036__ = ~new_new_n36870__ & ~new_new_n37035__;
  assign new_new_n37037__ = ~new_new_n23427__ & ~new_new_n37036__;
  assign new_new_n37038__ = ys__n30066 & new_new_n23427__;
  assign new_new_n37039__ = ~new_new_n37037__ & ~new_new_n37038__;
  assign new_new_n37040__ = ~new_new_n23431__ & ~new_new_n37039__;
  assign new_new_n37041__ = new_new_n23442__ & new_new_n37040__;
  assign new_new_n37042__ = new_new_n22665__ & ~new_new_n23442__;
  assign new_new_n37043__ = ~new_new_n37041__ & ~new_new_n37042__;
  assign new_new_n37044__ = ~new_new_n36545__ & ~new_new_n37043__;
  assign new_new_n37045__ = ~new_new_n37034__ & ~new_new_n37044__;
  assign new_new_n37046__ = new_new_n12210__ & ~new_new_n37045__;
  assign new_new_n37047__ = new_new_n36552__ & ~new_new_n37045__;
  assign ys__n29103 = new_new_n37046__ | new_new_n37047__;
  assign new_new_n37049__ = ~new_new_n22688__ & new_new_n36545__;
  assign new_new_n37050__ = ys__n30068 & new_new_n36868__;
  assign new_new_n37051__ = ~new_new_n36870__ & ~new_new_n37050__;
  assign new_new_n37052__ = ~new_new_n23427__ & ~new_new_n37051__;
  assign new_new_n37053__ = ys__n30068 & new_new_n23427__;
  assign new_new_n37054__ = ~new_new_n37052__ & ~new_new_n37053__;
  assign new_new_n37055__ = ~new_new_n23431__ & ~new_new_n37054__;
  assign new_new_n37056__ = new_new_n23442__ & new_new_n37055__;
  assign new_new_n37057__ = new_new_n22680__ & ~new_new_n23442__;
  assign new_new_n37058__ = ~new_new_n37056__ & ~new_new_n37057__;
  assign new_new_n37059__ = ~new_new_n36545__ & ~new_new_n37058__;
  assign new_new_n37060__ = ~new_new_n37049__ & ~new_new_n37059__;
  assign new_new_n37061__ = new_new_n12210__ & ~new_new_n37060__;
  assign new_new_n37062__ = new_new_n36552__ & ~new_new_n37060__;
  assign ys__n29106 = new_new_n37061__ | new_new_n37062__;
  assign new_new_n37064__ = ~new_new_n22703__ & new_new_n36545__;
  assign new_new_n37065__ = ys__n30070 & new_new_n36868__;
  assign new_new_n37066__ = ~new_new_n36870__ & ~new_new_n37065__;
  assign new_new_n37067__ = ~new_new_n23427__ & ~new_new_n37066__;
  assign new_new_n37068__ = ys__n30070 & new_new_n23427__;
  assign new_new_n37069__ = ~new_new_n37067__ & ~new_new_n37068__;
  assign new_new_n37070__ = ~new_new_n23431__ & ~new_new_n37069__;
  assign new_new_n37071__ = new_new_n23442__ & new_new_n37070__;
  assign new_new_n37072__ = new_new_n22695__ & ~new_new_n23442__;
  assign new_new_n37073__ = ~new_new_n37071__ & ~new_new_n37072__;
  assign new_new_n37074__ = ~new_new_n36545__ & ~new_new_n37073__;
  assign new_new_n37075__ = ~new_new_n37064__ & ~new_new_n37074__;
  assign new_new_n37076__ = new_new_n12210__ & ~new_new_n37075__;
  assign new_new_n37077__ = new_new_n36552__ & ~new_new_n37075__;
  assign ys__n29109 = new_new_n37076__ | new_new_n37077__;
  assign new_new_n37079__ = ~new_new_n22718__ & new_new_n36545__;
  assign new_new_n37080__ = ys__n30072 & new_new_n36868__;
  assign new_new_n37081__ = ~new_new_n36870__ & ~new_new_n37080__;
  assign new_new_n37082__ = ~new_new_n23427__ & ~new_new_n37081__;
  assign new_new_n37083__ = ys__n30072 & new_new_n23427__;
  assign new_new_n37084__ = ~new_new_n37082__ & ~new_new_n37083__;
  assign new_new_n37085__ = ~new_new_n23431__ & ~new_new_n37084__;
  assign new_new_n37086__ = new_new_n23442__ & new_new_n37085__;
  assign new_new_n37087__ = new_new_n22710__ & ~new_new_n23442__;
  assign new_new_n37088__ = ~new_new_n37086__ & ~new_new_n37087__;
  assign new_new_n37089__ = ~new_new_n36545__ & ~new_new_n37088__;
  assign new_new_n37090__ = ~new_new_n37079__ & ~new_new_n37089__;
  assign new_new_n37091__ = new_new_n12210__ & ~new_new_n37090__;
  assign new_new_n37092__ = new_new_n36552__ & ~new_new_n37090__;
  assign ys__n29112 = new_new_n37091__ | new_new_n37092__;
  assign new_new_n37094__ = ~new_new_n22733__ & new_new_n36545__;
  assign new_new_n37095__ = ys__n30074 & new_new_n36868__;
  assign new_new_n37096__ = ~new_new_n36870__ & ~new_new_n37095__;
  assign new_new_n37097__ = ~new_new_n23427__ & ~new_new_n37096__;
  assign new_new_n37098__ = ys__n30074 & new_new_n23427__;
  assign new_new_n37099__ = ~new_new_n37097__ & ~new_new_n37098__;
  assign new_new_n37100__ = ~new_new_n23431__ & ~new_new_n37099__;
  assign new_new_n37101__ = new_new_n23442__ & new_new_n37100__;
  assign new_new_n37102__ = new_new_n22725__ & ~new_new_n23442__;
  assign new_new_n37103__ = ~new_new_n37101__ & ~new_new_n37102__;
  assign new_new_n37104__ = ~new_new_n36545__ & ~new_new_n37103__;
  assign new_new_n37105__ = ~new_new_n37094__ & ~new_new_n37104__;
  assign new_new_n37106__ = new_new_n12210__ & ~new_new_n37105__;
  assign new_new_n37107__ = new_new_n36552__ & ~new_new_n37105__;
  assign ys__n29115 = new_new_n37106__ | new_new_n37107__;
  assign new_new_n37109__ = new_new_n21548__ & new_new_n21550__;
  assign new_new_n37110__ = new_new_n21534__ & new_new_n21538__;
  assign new_new_n37111__ = ~new_new_n37109__ & ~new_new_n37110__;
  assign new_new_n37112__ = ~new_new_n21555__ & new_new_n21561__;
  assign new_new_n37113__ = ~new_new_n37111__ & new_new_n37112__;
  assign new_new_n37114__ = ~new_new_n21561__ & new_new_n21587__;
  assign new_new_n37115__ = new_new_n21583__ & new_new_n37114__;
  assign new_new_n37116__ = ~new_new_n37113__ & ~new_new_n37115__;
  assign new_new_n37117__ = ~ys__n28243 & ~ys__n29117;
  assign ys__n29118 = ~new_new_n37116__ & new_new_n37117__;
  assign new_new_n37119__ = ~ys__n28243 & new_new_n21545__;
  assign new_new_n37120__ = new_new_n21561__ & new_new_n37119__;
  assign ys__n29217 = ~ys__n4566 & new_new_n37120__;
  assign ys__n29219 = ys__n29218 & ~ys__n4566;
  assign ys__n29221 = ys__n29220 & ~ys__n4566;
  assign new_new_n37124__ = new_new_n21542__ & new_new_n21561__;
  assign new_new_n37125__ = ~new_new_n21587__ & new_new_n21590__;
  assign new_new_n37126__ = ~new_new_n21561__ & new_new_n37125__;
  assign new_new_n37127__ = ~new_new_n37124__ & ~new_new_n37126__;
  assign new_new_n37128__ = ~ys__n28243 & ~ys__n4566;
  assign ys__n29223 = ~new_new_n37127__ & new_new_n37128__;
  assign ys__n29225 = ys__n29224 & ~ys__n4566;
  assign ys__n29226 = ys__n18114 & ~ys__n4566;
  assign ys__n29227 = ~ys__n28243 & ys__n23795;
  assign ys__n29228 = ~ys__n28243 & ys__n23798;
  assign ys__n29229 = ~ys__n28243 & ys__n23801;
  assign ys__n29230 = ~ys__n28243 & ys__n23804;
  assign ys__n29231 = ~ys__n28243 & ys__n23807;
  assign new_new_n37137__ = ~new_new_n37112__ & ~new_new_n37114__;
  assign ys__n29232 = ~ys__n28243 & ~new_new_n37137__;
  assign new_new_n37139__ = ~ys__n28243 & new_new_n21550__;
  assign new_new_n37140__ = new_new_n21561__ & new_new_n37139__;
  assign ys__n29233 = ~new_new_n21548__ & new_new_n37140__;
  assign new_new_n37142__ = new_new_n21538__ & new_new_n21561__;
  assign new_new_n37143__ = ~new_new_n21534__ & new_new_n37142__;
  assign new_new_n37144__ = ~new_new_n21583__ & new_new_n37114__;
  assign new_new_n37145__ = ~new_new_n37143__ & ~new_new_n37144__;
  assign ys__n29234 = ~ys__n28243 & ~new_new_n37145__;
  assign new_new_n37147__ = ~new_new_n21587__ & ~new_new_n37125__;
  assign new_new_n37148__ = ~ys__n28243 & ~new_new_n21561__;
  assign ys__n29235 = ~new_new_n37147__ & new_new_n37148__;
  assign new_new_n37150__ = ~ys__n4625 & ~ys__n38502;
  assign new_new_n37151__ = new_new_n12225__ & new_new_n37150__;
  assign new_new_n37152__ = ~new_new_n23120__ & new_new_n37151__;
  assign new_new_n37153__ = ~new_new_n22619__ & ~new_new_n36548__;
  assign new_new_n37154__ = ~new_new_n23116__ & ~new_new_n37153__;
  assign new_new_n37155__ = ~new_new_n37151__ & ~new_new_n37154__;
  assign new_new_n37156__ = ~new_new_n37152__ & ~new_new_n37155__;
  assign new_new_n37157__ = new_new_n12188__ & ~new_new_n37156__;
  assign new_new_n37158__ = ~ys__n740 & ~new_new_n12188__;
  assign new_new_n37159__ = ~new_new_n37156__ & new_new_n37158__;
  assign ys__n29336 = new_new_n37157__ | new_new_n37159__;
  assign new_new_n37161__ = ~new_new_n23139__ & new_new_n37151__;
  assign new_new_n37162__ = ~new_new_n22619__ & ~new_new_n36571__;
  assign new_new_n37163__ = ~new_new_n23135__ & ~new_new_n37162__;
  assign new_new_n37164__ = ~new_new_n37151__ & ~new_new_n37163__;
  assign new_new_n37165__ = ~new_new_n37161__ & ~new_new_n37164__;
  assign new_new_n37166__ = new_new_n12188__ & ~new_new_n37165__;
  assign new_new_n37167__ = new_new_n37158__ & ~new_new_n37165__;
  assign ys__n29339 = new_new_n37166__ | new_new_n37167__;
  assign new_new_n37169__ = ~new_new_n23158__ & new_new_n37151__;
  assign new_new_n37170__ = ~new_new_n22619__ & ~new_new_n36593__;
  assign new_new_n37171__ = ~new_new_n23154__ & ~new_new_n37170__;
  assign new_new_n37172__ = ~new_new_n37151__ & ~new_new_n37171__;
  assign new_new_n37173__ = ~new_new_n37169__ & ~new_new_n37172__;
  assign new_new_n37174__ = new_new_n12188__ & ~new_new_n37173__;
  assign new_new_n37175__ = new_new_n37158__ & ~new_new_n37173__;
  assign ys__n29342 = new_new_n37174__ | new_new_n37175__;
  assign new_new_n37177__ = ~new_new_n23177__ & new_new_n37151__;
  assign new_new_n37178__ = ~new_new_n22619__ & ~new_new_n36615__;
  assign new_new_n37179__ = ~new_new_n23173__ & ~new_new_n37178__;
  assign new_new_n37180__ = ~new_new_n37151__ & ~new_new_n37179__;
  assign new_new_n37181__ = ~new_new_n37177__ & ~new_new_n37180__;
  assign new_new_n37182__ = new_new_n12188__ & ~new_new_n37181__;
  assign new_new_n37183__ = new_new_n37158__ & ~new_new_n37181__;
  assign ys__n29345 = new_new_n37182__ | new_new_n37183__;
  assign new_new_n37185__ = ~new_new_n23196__ & new_new_n37151__;
  assign new_new_n37186__ = ~new_new_n22619__ & ~new_new_n36637__;
  assign new_new_n37187__ = ~new_new_n23192__ & ~new_new_n37186__;
  assign new_new_n37188__ = ~new_new_n37151__ & ~new_new_n37187__;
  assign new_new_n37189__ = ~new_new_n37185__ & ~new_new_n37188__;
  assign new_new_n37190__ = new_new_n12188__ & ~new_new_n37189__;
  assign new_new_n37191__ = new_new_n37158__ & ~new_new_n37189__;
  assign ys__n29348 = new_new_n37190__ | new_new_n37191__;
  assign new_new_n37193__ = ~new_new_n23215__ & new_new_n37151__;
  assign new_new_n37194__ = ~new_new_n22619__ & ~new_new_n36659__;
  assign new_new_n37195__ = ~new_new_n23211__ & ~new_new_n37194__;
  assign new_new_n37196__ = ~new_new_n37151__ & ~new_new_n37195__;
  assign new_new_n37197__ = ~new_new_n37193__ & ~new_new_n37196__;
  assign new_new_n37198__ = new_new_n12188__ & ~new_new_n37197__;
  assign new_new_n37199__ = new_new_n37158__ & ~new_new_n37197__;
  assign ys__n29351 = new_new_n37198__ | new_new_n37199__;
  assign new_new_n37201__ = ~new_new_n23234__ & new_new_n37151__;
  assign new_new_n37202__ = ~new_new_n22619__ & ~new_new_n36681__;
  assign new_new_n37203__ = ~new_new_n23230__ & ~new_new_n37202__;
  assign new_new_n37204__ = ~new_new_n37151__ & ~new_new_n37203__;
  assign new_new_n37205__ = ~new_new_n37201__ & ~new_new_n37204__;
  assign new_new_n37206__ = new_new_n12188__ & ~new_new_n37205__;
  assign new_new_n37207__ = new_new_n37158__ & ~new_new_n37205__;
  assign ys__n29354 = new_new_n37206__ | new_new_n37207__;
  assign new_new_n37209__ = ~new_new_n23253__ & new_new_n37151__;
  assign new_new_n37210__ = ~new_new_n22619__ & ~new_new_n36703__;
  assign new_new_n37211__ = ~new_new_n23249__ & ~new_new_n37210__;
  assign new_new_n37212__ = ~new_new_n37151__ & ~new_new_n37211__;
  assign new_new_n37213__ = ~new_new_n37209__ & ~new_new_n37212__;
  assign new_new_n37214__ = new_new_n12188__ & ~new_new_n37213__;
  assign new_new_n37215__ = new_new_n37158__ & ~new_new_n37213__;
  assign ys__n29357 = new_new_n37214__ | new_new_n37215__;
  assign new_new_n37217__ = ~new_new_n22934__ & new_new_n37151__;
  assign new_new_n37218__ = ~new_new_n22619__ & ~new_new_n36754__;
  assign new_new_n37219__ = ~new_new_n22930__ & ~new_new_n37218__;
  assign new_new_n37220__ = ~new_new_n37151__ & ~new_new_n37219__;
  assign new_new_n37221__ = ~new_new_n37217__ & ~new_new_n37220__;
  assign new_new_n37222__ = new_new_n12188__ & ~new_new_n37221__;
  assign new_new_n37223__ = new_new_n37158__ & ~new_new_n37221__;
  assign ys__n29360 = new_new_n37222__ | new_new_n37223__;
  assign new_new_n37225__ = ~new_new_n22952__ & new_new_n37151__;
  assign new_new_n37226__ = ~new_new_n22619__ & ~new_new_n36769__;
  assign new_new_n37227__ = ~new_new_n22948__ & ~new_new_n37226__;
  assign new_new_n37228__ = ~new_new_n37151__ & ~new_new_n37227__;
  assign new_new_n37229__ = ~new_new_n37225__ & ~new_new_n37228__;
  assign new_new_n37230__ = new_new_n12188__ & ~new_new_n37229__;
  assign new_new_n37231__ = new_new_n37158__ & ~new_new_n37229__;
  assign ys__n29363 = new_new_n37230__ | new_new_n37231__;
  assign new_new_n37233__ = ~new_new_n22970__ & new_new_n37151__;
  assign new_new_n37234__ = ~new_new_n22619__ & ~new_new_n36784__;
  assign new_new_n37235__ = ~new_new_n22966__ & ~new_new_n37234__;
  assign new_new_n37236__ = ~new_new_n37151__ & ~new_new_n37235__;
  assign new_new_n37237__ = ~new_new_n37233__ & ~new_new_n37236__;
  assign new_new_n37238__ = new_new_n12188__ & ~new_new_n37237__;
  assign new_new_n37239__ = new_new_n37158__ & ~new_new_n37237__;
  assign ys__n29366 = new_new_n37238__ | new_new_n37239__;
  assign new_new_n37241__ = ~new_new_n22988__ & new_new_n37151__;
  assign new_new_n37242__ = ~new_new_n22619__ & ~new_new_n36799__;
  assign new_new_n37243__ = ~new_new_n22984__ & ~new_new_n37242__;
  assign new_new_n37244__ = ~new_new_n37151__ & ~new_new_n37243__;
  assign new_new_n37245__ = ~new_new_n37241__ & ~new_new_n37244__;
  assign new_new_n37246__ = new_new_n12188__ & ~new_new_n37245__;
  assign new_new_n37247__ = new_new_n37158__ & ~new_new_n37245__;
  assign ys__n29369 = new_new_n37246__ | new_new_n37247__;
  assign new_new_n37249__ = ~new_new_n23006__ & new_new_n37151__;
  assign new_new_n37250__ = ~new_new_n22619__ & ~new_new_n36814__;
  assign new_new_n37251__ = ~new_new_n23002__ & ~new_new_n37250__;
  assign new_new_n37252__ = ~new_new_n37151__ & ~new_new_n37251__;
  assign new_new_n37253__ = ~new_new_n37249__ & ~new_new_n37252__;
  assign new_new_n37254__ = new_new_n12188__ & ~new_new_n37253__;
  assign new_new_n37255__ = new_new_n37158__ & ~new_new_n37253__;
  assign ys__n29372 = new_new_n37254__ | new_new_n37255__;
  assign new_new_n37257__ = ~new_new_n23024__ & new_new_n37151__;
  assign new_new_n37258__ = ~new_new_n22619__ & ~new_new_n36829__;
  assign new_new_n37259__ = ~new_new_n23020__ & ~new_new_n37258__;
  assign new_new_n37260__ = ~new_new_n37151__ & ~new_new_n37259__;
  assign new_new_n37261__ = ~new_new_n37257__ & ~new_new_n37260__;
  assign new_new_n37262__ = new_new_n12188__ & ~new_new_n37261__;
  assign new_new_n37263__ = new_new_n37158__ & ~new_new_n37261__;
  assign ys__n29375 = new_new_n37262__ | new_new_n37263__;
  assign new_new_n37265__ = ~new_new_n23042__ & new_new_n37151__;
  assign new_new_n37266__ = ~new_new_n22619__ & ~new_new_n36844__;
  assign new_new_n37267__ = ~new_new_n23038__ & ~new_new_n37266__;
  assign new_new_n37268__ = ~new_new_n37151__ & ~new_new_n37267__;
  assign new_new_n37269__ = ~new_new_n37265__ & ~new_new_n37268__;
  assign new_new_n37270__ = new_new_n12188__ & ~new_new_n37269__;
  assign new_new_n37271__ = new_new_n37158__ & ~new_new_n37269__;
  assign ys__n29378 = new_new_n37270__ | new_new_n37271__;
  assign new_new_n37273__ = ~new_new_n23060__ & new_new_n37151__;
  assign new_new_n37274__ = ~new_new_n22619__ & ~new_new_n36859__;
  assign new_new_n37275__ = ~new_new_n23056__ & ~new_new_n37274__;
  assign new_new_n37276__ = ~new_new_n37151__ & ~new_new_n37275__;
  assign new_new_n37277__ = ~new_new_n37273__ & ~new_new_n37276__;
  assign new_new_n37278__ = new_new_n12188__ & ~new_new_n37277__;
  assign new_new_n37279__ = new_new_n37158__ & ~new_new_n37277__;
  assign ys__n29381 = new_new_n37278__ | new_new_n37279__;
  assign new_new_n37281__ = ~new_new_n22774__ & new_new_n37151__;
  assign new_new_n37282__ = ~new_new_n22619__ & ~new_new_n36878__;
  assign new_new_n37283__ = ~new_new_n22770__ & ~new_new_n37282__;
  assign new_new_n37284__ = ~new_new_n37151__ & ~new_new_n37283__;
  assign new_new_n37285__ = ~new_new_n37281__ & ~new_new_n37284__;
  assign new_new_n37286__ = new_new_n12188__ & ~new_new_n37285__;
  assign new_new_n37287__ = new_new_n37158__ & ~new_new_n37285__;
  assign ys__n29384 = new_new_n37286__ | new_new_n37287__;
  assign new_new_n37289__ = ~new_new_n22789__ & new_new_n37151__;
  assign new_new_n37290__ = ~new_new_n22619__ & ~new_new_n36893__;
  assign new_new_n37291__ = ~new_new_n22785__ & ~new_new_n37290__;
  assign new_new_n37292__ = ~new_new_n37151__ & ~new_new_n37291__;
  assign new_new_n37293__ = ~new_new_n37289__ & ~new_new_n37292__;
  assign new_new_n37294__ = new_new_n12188__ & ~new_new_n37293__;
  assign new_new_n37295__ = new_new_n37158__ & ~new_new_n37293__;
  assign ys__n29387 = new_new_n37294__ | new_new_n37295__;
  assign new_new_n37297__ = ~new_new_n22804__ & new_new_n37151__;
  assign new_new_n37298__ = ~new_new_n22619__ & ~new_new_n36908__;
  assign new_new_n37299__ = ~new_new_n22800__ & ~new_new_n37298__;
  assign new_new_n37300__ = ~new_new_n37151__ & ~new_new_n37299__;
  assign new_new_n37301__ = ~new_new_n37297__ & ~new_new_n37300__;
  assign new_new_n37302__ = new_new_n12188__ & ~new_new_n37301__;
  assign new_new_n37303__ = new_new_n37158__ & ~new_new_n37301__;
  assign ys__n29390 = new_new_n37302__ | new_new_n37303__;
  assign new_new_n37305__ = ~new_new_n22819__ & new_new_n37151__;
  assign new_new_n37306__ = ~new_new_n22619__ & ~new_new_n36923__;
  assign new_new_n37307__ = ~new_new_n22815__ & ~new_new_n37306__;
  assign new_new_n37308__ = ~new_new_n37151__ & ~new_new_n37307__;
  assign new_new_n37309__ = ~new_new_n37305__ & ~new_new_n37308__;
  assign new_new_n37310__ = new_new_n12188__ & ~new_new_n37309__;
  assign new_new_n37311__ = new_new_n37158__ & ~new_new_n37309__;
  assign ys__n29393 = new_new_n37310__ | new_new_n37311__;
  assign new_new_n37313__ = ~new_new_n22834__ & new_new_n37151__;
  assign new_new_n37314__ = ~new_new_n22619__ & ~new_new_n36938__;
  assign new_new_n37315__ = ~new_new_n22830__ & ~new_new_n37314__;
  assign new_new_n37316__ = ~new_new_n37151__ & ~new_new_n37315__;
  assign new_new_n37317__ = ~new_new_n37313__ & ~new_new_n37316__;
  assign new_new_n37318__ = new_new_n12188__ & ~new_new_n37317__;
  assign new_new_n37319__ = new_new_n37158__ & ~new_new_n37317__;
  assign ys__n29396 = new_new_n37318__ | new_new_n37319__;
  assign new_new_n37321__ = ~new_new_n22849__ & new_new_n37151__;
  assign new_new_n37322__ = ~new_new_n22619__ & ~new_new_n36953__;
  assign new_new_n37323__ = ~new_new_n22845__ & ~new_new_n37322__;
  assign new_new_n37324__ = ~new_new_n37151__ & ~new_new_n37323__;
  assign new_new_n37325__ = ~new_new_n37321__ & ~new_new_n37324__;
  assign new_new_n37326__ = new_new_n12188__ & ~new_new_n37325__;
  assign new_new_n37327__ = new_new_n37158__ & ~new_new_n37325__;
  assign ys__n29399 = new_new_n37326__ | new_new_n37327__;
  assign new_new_n37329__ = ~new_new_n22864__ & new_new_n37151__;
  assign new_new_n37330__ = ~new_new_n22619__ & ~new_new_n36968__;
  assign new_new_n37331__ = ~new_new_n22860__ & ~new_new_n37330__;
  assign new_new_n37332__ = ~new_new_n37151__ & ~new_new_n37331__;
  assign new_new_n37333__ = ~new_new_n37329__ & ~new_new_n37332__;
  assign new_new_n37334__ = new_new_n12188__ & ~new_new_n37333__;
  assign new_new_n37335__ = new_new_n37158__ & ~new_new_n37333__;
  assign ys__n29402 = new_new_n37334__ | new_new_n37335__;
  assign new_new_n37337__ = ~new_new_n22879__ & new_new_n37151__;
  assign new_new_n37338__ = ~new_new_n22619__ & ~new_new_n36983__;
  assign new_new_n37339__ = ~new_new_n22875__ & ~new_new_n37338__;
  assign new_new_n37340__ = ~new_new_n37151__ & ~new_new_n37339__;
  assign new_new_n37341__ = ~new_new_n37337__ & ~new_new_n37340__;
  assign new_new_n37342__ = new_new_n12188__ & ~new_new_n37341__;
  assign new_new_n37343__ = new_new_n37158__ & ~new_new_n37341__;
  assign ys__n29405 = new_new_n37342__ | new_new_n37343__;
  assign new_new_n37345__ = ~new_new_n22626__ & new_new_n37151__;
  assign new_new_n37346__ = ~new_new_n22619__ & ~new_new_n36998__;
  assign new_new_n37347__ = ~new_new_n22620__ & ~new_new_n37346__;
  assign new_new_n37348__ = ~new_new_n37151__ & ~new_new_n37347__;
  assign new_new_n37349__ = ~new_new_n37345__ & ~new_new_n37348__;
  assign new_new_n37350__ = new_new_n12188__ & ~new_new_n37349__;
  assign new_new_n37351__ = new_new_n37158__ & ~new_new_n37349__;
  assign ys__n29408 = new_new_n37350__ | new_new_n37351__;
  assign new_new_n37353__ = ~new_new_n22641__ & new_new_n37151__;
  assign new_new_n37354__ = ~new_new_n22619__ & ~new_new_n37013__;
  assign new_new_n37355__ = ~new_new_n22637__ & ~new_new_n37354__;
  assign new_new_n37356__ = ~new_new_n37151__ & ~new_new_n37355__;
  assign new_new_n37357__ = ~new_new_n37353__ & ~new_new_n37356__;
  assign new_new_n37358__ = new_new_n12188__ & ~new_new_n37357__;
  assign new_new_n37359__ = new_new_n37158__ & ~new_new_n37357__;
  assign ys__n29411 = new_new_n37358__ | new_new_n37359__;
  assign new_new_n37361__ = ~new_new_n22656__ & new_new_n37151__;
  assign new_new_n37362__ = ~new_new_n22619__ & ~new_new_n37028__;
  assign new_new_n37363__ = ~new_new_n22652__ & ~new_new_n37362__;
  assign new_new_n37364__ = ~new_new_n37151__ & ~new_new_n37363__;
  assign new_new_n37365__ = ~new_new_n37361__ & ~new_new_n37364__;
  assign new_new_n37366__ = new_new_n12188__ & ~new_new_n37365__;
  assign new_new_n37367__ = new_new_n37158__ & ~new_new_n37365__;
  assign ys__n29414 = new_new_n37366__ | new_new_n37367__;
  assign new_new_n37369__ = ~new_new_n22671__ & new_new_n37151__;
  assign new_new_n37370__ = ~new_new_n22619__ & ~new_new_n37043__;
  assign new_new_n37371__ = ~new_new_n22667__ & ~new_new_n37370__;
  assign new_new_n37372__ = ~new_new_n37151__ & ~new_new_n37371__;
  assign new_new_n37373__ = ~new_new_n37369__ & ~new_new_n37372__;
  assign new_new_n37374__ = new_new_n12188__ & ~new_new_n37373__;
  assign new_new_n37375__ = new_new_n37158__ & ~new_new_n37373__;
  assign ys__n29417 = new_new_n37374__ | new_new_n37375__;
  assign new_new_n37377__ = ~new_new_n22686__ & new_new_n37151__;
  assign new_new_n37378__ = ~new_new_n22619__ & ~new_new_n37058__;
  assign new_new_n37379__ = ~new_new_n22682__ & ~new_new_n37378__;
  assign new_new_n37380__ = ~new_new_n37151__ & ~new_new_n37379__;
  assign new_new_n37381__ = ~new_new_n37377__ & ~new_new_n37380__;
  assign new_new_n37382__ = new_new_n12188__ & ~new_new_n37381__;
  assign new_new_n37383__ = new_new_n37158__ & ~new_new_n37381__;
  assign ys__n29420 = new_new_n37382__ | new_new_n37383__;
  assign new_new_n37385__ = ~new_new_n22701__ & new_new_n37151__;
  assign new_new_n37386__ = ~new_new_n22619__ & ~new_new_n37073__;
  assign new_new_n37387__ = ~new_new_n22697__ & ~new_new_n37386__;
  assign new_new_n37388__ = ~new_new_n37151__ & ~new_new_n37387__;
  assign new_new_n37389__ = ~new_new_n37385__ & ~new_new_n37388__;
  assign new_new_n37390__ = new_new_n12188__ & ~new_new_n37389__;
  assign new_new_n37391__ = new_new_n37158__ & ~new_new_n37389__;
  assign ys__n29423 = new_new_n37390__ | new_new_n37391__;
  assign new_new_n37393__ = ~new_new_n22716__ & new_new_n37151__;
  assign new_new_n37394__ = ~new_new_n22619__ & ~new_new_n37088__;
  assign new_new_n37395__ = ~new_new_n22712__ & ~new_new_n37394__;
  assign new_new_n37396__ = ~new_new_n37151__ & ~new_new_n37395__;
  assign new_new_n37397__ = ~new_new_n37393__ & ~new_new_n37396__;
  assign new_new_n37398__ = new_new_n12188__ & ~new_new_n37397__;
  assign new_new_n37399__ = new_new_n37158__ & ~new_new_n37397__;
  assign ys__n29426 = new_new_n37398__ | new_new_n37399__;
  assign new_new_n37401__ = ~new_new_n22731__ & new_new_n37151__;
  assign new_new_n37402__ = ~new_new_n22619__ & ~new_new_n37103__;
  assign new_new_n37403__ = ~new_new_n22727__ & ~new_new_n37402__;
  assign new_new_n37404__ = ~new_new_n37151__ & ~new_new_n37403__;
  assign new_new_n37405__ = ~new_new_n37401__ & ~new_new_n37404__;
  assign new_new_n37406__ = new_new_n12188__ & ~new_new_n37405__;
  assign new_new_n37407__ = new_new_n37158__ & ~new_new_n37405__;
  assign ys__n29429 = new_new_n37406__ | new_new_n37407__;
  assign new_new_n37409__ = new_new_n21695__ & new_new_n21697__;
  assign new_new_n37410__ = new_new_n21681__ & new_new_n21685__;
  assign new_new_n37411__ = ~new_new_n37409__ & ~new_new_n37410__;
  assign new_new_n37412__ = ~new_new_n21702__ & new_new_n21708__;
  assign new_new_n37413__ = ~new_new_n37411__ & new_new_n37412__;
  assign new_new_n37414__ = ~new_new_n21708__ & new_new_n21734__;
  assign new_new_n37415__ = new_new_n21730__ & new_new_n37414__;
  assign new_new_n37416__ = ~new_new_n37413__ & ~new_new_n37415__;
  assign ys__n29431 = new_new_n37117__ & ~new_new_n37416__;
  assign new_new_n37418__ = ~ys__n28243 & new_new_n21692__;
  assign new_new_n37419__ = new_new_n21708__ & new_new_n37418__;
  assign ys__n29530 = ~ys__n4566 & new_new_n37419__;
  assign ys__n29532 = ys__n29531 & ~ys__n4566;
  assign ys__n29534 = ys__n29533 & ~ys__n4566;
  assign new_new_n37423__ = new_new_n21689__ & new_new_n21708__;
  assign new_new_n37424__ = ~new_new_n21734__ & new_new_n21737__;
  assign new_new_n37425__ = ~new_new_n21708__ & new_new_n37424__;
  assign new_new_n37426__ = ~new_new_n37423__ & ~new_new_n37425__;
  assign ys__n29536 = new_new_n37128__ & ~new_new_n37426__;
  assign ys__n29538 = ys__n29537 & ~ys__n4566;
  assign ys__n29539 = ys__n18116 & ~ys__n4566;
  assign ys__n29540 = ~ys__n28243 & ys__n23865;
  assign ys__n29541 = ~ys__n28243 & ys__n23868;
  assign ys__n29542 = ~ys__n28243 & ys__n23871;
  assign ys__n29543 = ~ys__n28243 & ys__n23874;
  assign ys__n29544 = ~ys__n28243 & ys__n23877;
  assign new_new_n37435__ = ~new_new_n37412__ & ~new_new_n37414__;
  assign ys__n29545 = ~ys__n28243 & ~new_new_n37435__;
  assign new_new_n37437__ = ~ys__n28243 & new_new_n21697__;
  assign new_new_n37438__ = new_new_n21708__ & new_new_n37437__;
  assign ys__n29546 = ~new_new_n21695__ & new_new_n37438__;
  assign new_new_n37440__ = new_new_n21685__ & new_new_n21708__;
  assign new_new_n37441__ = ~new_new_n21681__ & new_new_n37440__;
  assign new_new_n37442__ = ~new_new_n21730__ & new_new_n37414__;
  assign new_new_n37443__ = ~new_new_n37441__ & ~new_new_n37442__;
  assign ys__n29547 = ~ys__n28243 & ~new_new_n37443__;
  assign new_new_n37445__ = ~new_new_n21734__ & ~new_new_n37424__;
  assign new_new_n37446__ = ~ys__n28243 & ~new_new_n21708__;
  assign ys__n29548 = ~new_new_n37445__ & new_new_n37446__;
  assign new_new_n37448__ = ~ys__n4625 & ~ys__n38513;
  assign new_new_n37449__ = new_new_n12225__ & new_new_n37448__;
  assign new_new_n37450__ = ys__n28462 & new_new_n37449__;
  assign new_new_n37451__ = ~new_new_n22621__ & ~new_new_n37154__;
  assign new_new_n37452__ = ~new_new_n23117__ & ~new_new_n37451__;
  assign new_new_n37453__ = ~new_new_n37449__ & ~new_new_n37452__;
  assign new_new_n37454__ = ~new_new_n37450__ & ~new_new_n37453__;
  assign new_new_n37455__ = new_new_n12177__ & ~new_new_n37454__;
  assign new_new_n37456__ = ~ys__n740 & ~new_new_n12177__;
  assign new_new_n37457__ = ~new_new_n37454__ & new_new_n37456__;
  assign ys__n29611 = new_new_n37455__ | new_new_n37457__;
  assign new_new_n37459__ = ys__n28464 & new_new_n37449__;
  assign new_new_n37460__ = ~new_new_n22621__ & ~new_new_n37163__;
  assign new_new_n37461__ = ~new_new_n23136__ & ~new_new_n37460__;
  assign new_new_n37462__ = ~new_new_n37449__ & ~new_new_n37461__;
  assign new_new_n37463__ = ~new_new_n37459__ & ~new_new_n37462__;
  assign new_new_n37464__ = new_new_n12177__ & ~new_new_n37463__;
  assign new_new_n37465__ = new_new_n37456__ & ~new_new_n37463__;
  assign ys__n29614 = new_new_n37464__ | new_new_n37465__;
  assign new_new_n37467__ = ys__n28466 & new_new_n37449__;
  assign new_new_n37468__ = ~new_new_n22621__ & ~new_new_n37171__;
  assign new_new_n37469__ = ~new_new_n23155__ & ~new_new_n37468__;
  assign new_new_n37470__ = ~new_new_n37449__ & ~new_new_n37469__;
  assign new_new_n37471__ = ~new_new_n37467__ & ~new_new_n37470__;
  assign new_new_n37472__ = new_new_n12177__ & ~new_new_n37471__;
  assign new_new_n37473__ = new_new_n37456__ & ~new_new_n37471__;
  assign ys__n29617 = new_new_n37472__ | new_new_n37473__;
  assign new_new_n37475__ = ys__n28468 & new_new_n37449__;
  assign new_new_n37476__ = ~new_new_n22621__ & ~new_new_n37179__;
  assign new_new_n37477__ = ~new_new_n23174__ & ~new_new_n37476__;
  assign new_new_n37478__ = ~new_new_n37449__ & ~new_new_n37477__;
  assign new_new_n37479__ = ~new_new_n37475__ & ~new_new_n37478__;
  assign new_new_n37480__ = new_new_n12177__ & ~new_new_n37479__;
  assign new_new_n37481__ = new_new_n37456__ & ~new_new_n37479__;
  assign ys__n29620 = new_new_n37480__ | new_new_n37481__;
  assign new_new_n37483__ = ys__n28470 & new_new_n37449__;
  assign new_new_n37484__ = ~new_new_n22621__ & ~new_new_n37187__;
  assign new_new_n37485__ = ~new_new_n23193__ & ~new_new_n37484__;
  assign new_new_n37486__ = ~new_new_n37449__ & ~new_new_n37485__;
  assign new_new_n37487__ = ~new_new_n37483__ & ~new_new_n37486__;
  assign new_new_n37488__ = new_new_n12177__ & ~new_new_n37487__;
  assign new_new_n37489__ = new_new_n37456__ & ~new_new_n37487__;
  assign ys__n29623 = new_new_n37488__ | new_new_n37489__;
  assign new_new_n37491__ = ys__n28472 & new_new_n37449__;
  assign new_new_n37492__ = ~new_new_n22621__ & ~new_new_n37195__;
  assign new_new_n37493__ = ~new_new_n23212__ & ~new_new_n37492__;
  assign new_new_n37494__ = ~new_new_n37449__ & ~new_new_n37493__;
  assign new_new_n37495__ = ~new_new_n37491__ & ~new_new_n37494__;
  assign new_new_n37496__ = new_new_n12177__ & ~new_new_n37495__;
  assign new_new_n37497__ = new_new_n37456__ & ~new_new_n37495__;
  assign ys__n29626 = new_new_n37496__ | new_new_n37497__;
  assign new_new_n37499__ = ys__n29558 & new_new_n37449__;
  assign new_new_n37500__ = ~new_new_n22621__ & ~new_new_n37203__;
  assign new_new_n37501__ = ~new_new_n23231__ & ~new_new_n37500__;
  assign new_new_n37502__ = ~new_new_n37449__ & ~new_new_n37501__;
  assign new_new_n37503__ = ~new_new_n37499__ & ~new_new_n37502__;
  assign new_new_n37504__ = new_new_n12177__ & ~new_new_n37503__;
  assign new_new_n37505__ = new_new_n37456__ & ~new_new_n37503__;
  assign ys__n29629 = new_new_n37504__ | new_new_n37505__;
  assign new_new_n37507__ = ys__n29560 & new_new_n37449__;
  assign new_new_n37508__ = ~new_new_n22621__ & ~new_new_n37211__;
  assign new_new_n37509__ = ~new_new_n23250__ & ~new_new_n37508__;
  assign new_new_n37510__ = ~new_new_n37449__ & ~new_new_n37509__;
  assign new_new_n37511__ = ~new_new_n37507__ & ~new_new_n37510__;
  assign new_new_n37512__ = new_new_n12177__ & ~new_new_n37511__;
  assign new_new_n37513__ = new_new_n37456__ & ~new_new_n37511__;
  assign ys__n29632 = new_new_n37512__ | new_new_n37513__;
  assign new_new_n37515__ = ys__n29562 & new_new_n37449__;
  assign new_new_n37516__ = ~new_new_n22621__ & ~new_new_n37219__;
  assign new_new_n37517__ = ~new_new_n22931__ & ~new_new_n37516__;
  assign new_new_n37518__ = ~new_new_n37449__ & ~new_new_n37517__;
  assign new_new_n37519__ = ~new_new_n37515__ & ~new_new_n37518__;
  assign new_new_n37520__ = new_new_n12177__ & ~new_new_n37519__;
  assign new_new_n37521__ = new_new_n37456__ & ~new_new_n37519__;
  assign ys__n29635 = new_new_n37520__ | new_new_n37521__;
  assign new_new_n37523__ = ys__n29564 & new_new_n37449__;
  assign new_new_n37524__ = ~new_new_n22621__ & ~new_new_n37227__;
  assign new_new_n37525__ = ~new_new_n22949__ & ~new_new_n37524__;
  assign new_new_n37526__ = ~new_new_n37449__ & ~new_new_n37525__;
  assign new_new_n37527__ = ~new_new_n37523__ & ~new_new_n37526__;
  assign new_new_n37528__ = new_new_n12177__ & ~new_new_n37527__;
  assign new_new_n37529__ = new_new_n37456__ & ~new_new_n37527__;
  assign ys__n29638 = new_new_n37528__ | new_new_n37529__;
  assign new_new_n37531__ = ys__n29566 & new_new_n37449__;
  assign new_new_n37532__ = ~new_new_n22621__ & ~new_new_n37235__;
  assign new_new_n37533__ = ~new_new_n22967__ & ~new_new_n37532__;
  assign new_new_n37534__ = ~new_new_n37449__ & ~new_new_n37533__;
  assign new_new_n37535__ = ~new_new_n37531__ & ~new_new_n37534__;
  assign new_new_n37536__ = new_new_n12177__ & ~new_new_n37535__;
  assign new_new_n37537__ = new_new_n37456__ & ~new_new_n37535__;
  assign ys__n29641 = new_new_n37536__ | new_new_n37537__;
  assign new_new_n37539__ = ys__n29568 & new_new_n37449__;
  assign new_new_n37540__ = ~new_new_n22621__ & ~new_new_n37243__;
  assign new_new_n37541__ = ~new_new_n22985__ & ~new_new_n37540__;
  assign new_new_n37542__ = ~new_new_n37449__ & ~new_new_n37541__;
  assign new_new_n37543__ = ~new_new_n37539__ & ~new_new_n37542__;
  assign new_new_n37544__ = new_new_n12177__ & ~new_new_n37543__;
  assign new_new_n37545__ = new_new_n37456__ & ~new_new_n37543__;
  assign ys__n29644 = new_new_n37544__ | new_new_n37545__;
  assign new_new_n37547__ = ys__n29570 & new_new_n37449__;
  assign new_new_n37548__ = ~new_new_n22621__ & ~new_new_n37251__;
  assign new_new_n37549__ = ~new_new_n23003__ & ~new_new_n37548__;
  assign new_new_n37550__ = ~new_new_n37449__ & ~new_new_n37549__;
  assign new_new_n37551__ = ~new_new_n37547__ & ~new_new_n37550__;
  assign new_new_n37552__ = new_new_n12177__ & ~new_new_n37551__;
  assign new_new_n37553__ = new_new_n37456__ & ~new_new_n37551__;
  assign ys__n29647 = new_new_n37552__ | new_new_n37553__;
  assign new_new_n37555__ = ys__n29572 & new_new_n37449__;
  assign new_new_n37556__ = ~new_new_n22621__ & ~new_new_n37259__;
  assign new_new_n37557__ = ~new_new_n23021__ & ~new_new_n37556__;
  assign new_new_n37558__ = ~new_new_n37449__ & ~new_new_n37557__;
  assign new_new_n37559__ = ~new_new_n37555__ & ~new_new_n37558__;
  assign new_new_n37560__ = new_new_n12177__ & ~new_new_n37559__;
  assign new_new_n37561__ = new_new_n37456__ & ~new_new_n37559__;
  assign ys__n29650 = new_new_n37560__ | new_new_n37561__;
  assign new_new_n37563__ = ys__n29574 & new_new_n37449__;
  assign new_new_n37564__ = ~new_new_n22621__ & ~new_new_n37267__;
  assign new_new_n37565__ = ~new_new_n23039__ & ~new_new_n37564__;
  assign new_new_n37566__ = ~new_new_n37449__ & ~new_new_n37565__;
  assign new_new_n37567__ = ~new_new_n37563__ & ~new_new_n37566__;
  assign new_new_n37568__ = new_new_n12177__ & ~new_new_n37567__;
  assign new_new_n37569__ = new_new_n37456__ & ~new_new_n37567__;
  assign ys__n29653 = new_new_n37568__ | new_new_n37569__;
  assign new_new_n37571__ = ys__n29576 & new_new_n37449__;
  assign new_new_n37572__ = ~new_new_n22621__ & ~new_new_n37275__;
  assign new_new_n37573__ = ~new_new_n23057__ & ~new_new_n37572__;
  assign new_new_n37574__ = ~new_new_n37449__ & ~new_new_n37573__;
  assign new_new_n37575__ = ~new_new_n37571__ & ~new_new_n37574__;
  assign new_new_n37576__ = new_new_n12177__ & ~new_new_n37575__;
  assign new_new_n37577__ = new_new_n37456__ & ~new_new_n37575__;
  assign ys__n29656 = new_new_n37576__ | new_new_n37577__;
  assign new_new_n37579__ = ys__n29578 & new_new_n37449__;
  assign new_new_n37580__ = ~new_new_n22621__ & ~new_new_n37283__;
  assign new_new_n37581__ = ~new_new_n22771__ & ~new_new_n37580__;
  assign new_new_n37582__ = ~new_new_n37449__ & ~new_new_n37581__;
  assign new_new_n37583__ = ~new_new_n37579__ & ~new_new_n37582__;
  assign new_new_n37584__ = new_new_n12177__ & ~new_new_n37583__;
  assign new_new_n37585__ = new_new_n37456__ & ~new_new_n37583__;
  assign ys__n29659 = new_new_n37584__ | new_new_n37585__;
  assign new_new_n37587__ = ys__n29580 & new_new_n37449__;
  assign new_new_n37588__ = ~new_new_n22621__ & ~new_new_n37291__;
  assign new_new_n37589__ = ~new_new_n22786__ & ~new_new_n37588__;
  assign new_new_n37590__ = ~new_new_n37449__ & ~new_new_n37589__;
  assign new_new_n37591__ = ~new_new_n37587__ & ~new_new_n37590__;
  assign new_new_n37592__ = new_new_n12177__ & ~new_new_n37591__;
  assign new_new_n37593__ = new_new_n37456__ & ~new_new_n37591__;
  assign ys__n29662 = new_new_n37592__ | new_new_n37593__;
  assign new_new_n37595__ = ys__n29582 & new_new_n37449__;
  assign new_new_n37596__ = ~new_new_n22621__ & ~new_new_n37299__;
  assign new_new_n37597__ = ~new_new_n22801__ & ~new_new_n37596__;
  assign new_new_n37598__ = ~new_new_n37449__ & ~new_new_n37597__;
  assign new_new_n37599__ = ~new_new_n37595__ & ~new_new_n37598__;
  assign new_new_n37600__ = new_new_n12177__ & ~new_new_n37599__;
  assign new_new_n37601__ = new_new_n37456__ & ~new_new_n37599__;
  assign ys__n29665 = new_new_n37600__ | new_new_n37601__;
  assign new_new_n37603__ = ys__n29584 & new_new_n37449__;
  assign new_new_n37604__ = ~new_new_n22621__ & ~new_new_n37307__;
  assign new_new_n37605__ = ~new_new_n22816__ & ~new_new_n37604__;
  assign new_new_n37606__ = ~new_new_n37449__ & ~new_new_n37605__;
  assign new_new_n37607__ = ~new_new_n37603__ & ~new_new_n37606__;
  assign new_new_n37608__ = new_new_n12177__ & ~new_new_n37607__;
  assign new_new_n37609__ = new_new_n37456__ & ~new_new_n37607__;
  assign ys__n29668 = new_new_n37608__ | new_new_n37609__;
  assign new_new_n37611__ = ys__n29586 & new_new_n37449__;
  assign new_new_n37612__ = ~new_new_n22621__ & ~new_new_n37315__;
  assign new_new_n37613__ = ~new_new_n22831__ & ~new_new_n37612__;
  assign new_new_n37614__ = ~new_new_n37449__ & ~new_new_n37613__;
  assign new_new_n37615__ = ~new_new_n37611__ & ~new_new_n37614__;
  assign new_new_n37616__ = new_new_n12177__ & ~new_new_n37615__;
  assign new_new_n37617__ = new_new_n37456__ & ~new_new_n37615__;
  assign ys__n29671 = new_new_n37616__ | new_new_n37617__;
  assign new_new_n37619__ = ys__n29588 & new_new_n37449__;
  assign new_new_n37620__ = ~new_new_n22621__ & ~new_new_n37323__;
  assign new_new_n37621__ = ~new_new_n22846__ & ~new_new_n37620__;
  assign new_new_n37622__ = ~new_new_n37449__ & ~new_new_n37621__;
  assign new_new_n37623__ = ~new_new_n37619__ & ~new_new_n37622__;
  assign new_new_n37624__ = new_new_n12177__ & ~new_new_n37623__;
  assign new_new_n37625__ = new_new_n37456__ & ~new_new_n37623__;
  assign ys__n29674 = new_new_n37624__ | new_new_n37625__;
  assign new_new_n37627__ = ys__n29590 & new_new_n37449__;
  assign new_new_n37628__ = ~new_new_n22621__ & ~new_new_n37331__;
  assign new_new_n37629__ = ~new_new_n22861__ & ~new_new_n37628__;
  assign new_new_n37630__ = ~new_new_n37449__ & ~new_new_n37629__;
  assign new_new_n37631__ = ~new_new_n37627__ & ~new_new_n37630__;
  assign new_new_n37632__ = new_new_n12177__ & ~new_new_n37631__;
  assign new_new_n37633__ = new_new_n37456__ & ~new_new_n37631__;
  assign ys__n29677 = new_new_n37632__ | new_new_n37633__;
  assign new_new_n37635__ = ys__n29592 & new_new_n37449__;
  assign new_new_n37636__ = ~new_new_n22621__ & ~new_new_n37339__;
  assign new_new_n37637__ = ~new_new_n22876__ & ~new_new_n37636__;
  assign new_new_n37638__ = ~new_new_n37449__ & ~new_new_n37637__;
  assign new_new_n37639__ = ~new_new_n37635__ & ~new_new_n37638__;
  assign new_new_n37640__ = new_new_n12177__ & ~new_new_n37639__;
  assign new_new_n37641__ = new_new_n37456__ & ~new_new_n37639__;
  assign ys__n29680 = new_new_n37640__ | new_new_n37641__;
  assign new_new_n37643__ = ys__n29594 & new_new_n37449__;
  assign new_new_n37644__ = ~new_new_n22621__ & ~new_new_n37347__;
  assign new_new_n37645__ = ~new_new_n22622__ & ~new_new_n37644__;
  assign new_new_n37646__ = ~new_new_n37449__ & ~new_new_n37645__;
  assign new_new_n37647__ = ~new_new_n37643__ & ~new_new_n37646__;
  assign new_new_n37648__ = new_new_n12177__ & ~new_new_n37647__;
  assign new_new_n37649__ = new_new_n37456__ & ~new_new_n37647__;
  assign ys__n29683 = new_new_n37648__ | new_new_n37649__;
  assign new_new_n37651__ = ys__n29596 & new_new_n37449__;
  assign new_new_n37652__ = ~new_new_n22621__ & ~new_new_n37355__;
  assign new_new_n37653__ = ~new_new_n22638__ & ~new_new_n37652__;
  assign new_new_n37654__ = ~new_new_n37449__ & ~new_new_n37653__;
  assign new_new_n37655__ = ~new_new_n37651__ & ~new_new_n37654__;
  assign new_new_n37656__ = new_new_n12177__ & ~new_new_n37655__;
  assign new_new_n37657__ = new_new_n37456__ & ~new_new_n37655__;
  assign ys__n29686 = new_new_n37656__ | new_new_n37657__;
  assign new_new_n37659__ = ys__n29598 & new_new_n37449__;
  assign new_new_n37660__ = ~new_new_n22621__ & ~new_new_n37363__;
  assign new_new_n37661__ = ~new_new_n22653__ & ~new_new_n37660__;
  assign new_new_n37662__ = ~new_new_n37449__ & ~new_new_n37661__;
  assign new_new_n37663__ = ~new_new_n37659__ & ~new_new_n37662__;
  assign new_new_n37664__ = new_new_n12177__ & ~new_new_n37663__;
  assign new_new_n37665__ = new_new_n37456__ & ~new_new_n37663__;
  assign ys__n29689 = new_new_n37664__ | new_new_n37665__;
  assign new_new_n37667__ = ys__n29600 & new_new_n37449__;
  assign new_new_n37668__ = ~new_new_n22621__ & ~new_new_n37371__;
  assign new_new_n37669__ = ~new_new_n22668__ & ~new_new_n37668__;
  assign new_new_n37670__ = ~new_new_n37449__ & ~new_new_n37669__;
  assign new_new_n37671__ = ~new_new_n37667__ & ~new_new_n37670__;
  assign new_new_n37672__ = new_new_n12177__ & ~new_new_n37671__;
  assign new_new_n37673__ = new_new_n37456__ & ~new_new_n37671__;
  assign ys__n29692 = new_new_n37672__ | new_new_n37673__;
  assign new_new_n37675__ = ys__n29602 & new_new_n37449__;
  assign new_new_n37676__ = ~new_new_n22621__ & ~new_new_n37379__;
  assign new_new_n37677__ = ~new_new_n22683__ & ~new_new_n37676__;
  assign new_new_n37678__ = ~new_new_n37449__ & ~new_new_n37677__;
  assign new_new_n37679__ = ~new_new_n37675__ & ~new_new_n37678__;
  assign new_new_n37680__ = new_new_n12177__ & ~new_new_n37679__;
  assign new_new_n37681__ = new_new_n37456__ & ~new_new_n37679__;
  assign ys__n29695 = new_new_n37680__ | new_new_n37681__;
  assign new_new_n37683__ = ys__n29604 & new_new_n37449__;
  assign new_new_n37684__ = ~new_new_n22621__ & ~new_new_n37387__;
  assign new_new_n37685__ = ~new_new_n22698__ & ~new_new_n37684__;
  assign new_new_n37686__ = ~new_new_n37449__ & ~new_new_n37685__;
  assign new_new_n37687__ = ~new_new_n37683__ & ~new_new_n37686__;
  assign new_new_n37688__ = new_new_n12177__ & ~new_new_n37687__;
  assign new_new_n37689__ = new_new_n37456__ & ~new_new_n37687__;
  assign ys__n29698 = new_new_n37688__ | new_new_n37689__;
  assign new_new_n37691__ = ys__n29606 & new_new_n37449__;
  assign new_new_n37692__ = ~new_new_n22621__ & ~new_new_n37395__;
  assign new_new_n37693__ = ~new_new_n22713__ & ~new_new_n37692__;
  assign new_new_n37694__ = ~new_new_n37449__ & ~new_new_n37693__;
  assign new_new_n37695__ = ~new_new_n37691__ & ~new_new_n37694__;
  assign new_new_n37696__ = new_new_n12177__ & ~new_new_n37695__;
  assign new_new_n37697__ = new_new_n37456__ & ~new_new_n37695__;
  assign ys__n29701 = new_new_n37696__ | new_new_n37697__;
  assign new_new_n37699__ = ys__n29608 & new_new_n37449__;
  assign new_new_n37700__ = ~new_new_n22621__ & ~new_new_n37403__;
  assign new_new_n37701__ = ~new_new_n22728__ & ~new_new_n37700__;
  assign new_new_n37702__ = ~new_new_n37449__ & ~new_new_n37701__;
  assign new_new_n37703__ = ~new_new_n37699__ & ~new_new_n37702__;
  assign new_new_n37704__ = new_new_n12177__ & ~new_new_n37703__;
  assign new_new_n37705__ = new_new_n37456__ & ~new_new_n37703__;
  assign ys__n29704 = new_new_n37704__ | new_new_n37705__;
  assign new_new_n37707__ = new_new_n21842__ & new_new_n21844__;
  assign new_new_n37708__ = new_new_n21828__ & new_new_n21832__;
  assign new_new_n37709__ = ~new_new_n37707__ & ~new_new_n37708__;
  assign new_new_n37710__ = ~new_new_n21849__ & new_new_n21855__;
  assign new_new_n37711__ = ~new_new_n37709__ & new_new_n37710__;
  assign new_new_n37712__ = ~new_new_n21855__ & new_new_n21881__;
  assign new_new_n37713__ = new_new_n21877__ & new_new_n37712__;
  assign new_new_n37714__ = ~new_new_n37711__ & ~new_new_n37713__;
  assign ys__n29706 = new_new_n37117__ & ~new_new_n37714__;
  assign new_new_n37716__ = ~ys__n28243 & new_new_n21839__;
  assign new_new_n37717__ = new_new_n21855__ & new_new_n37716__;
  assign ys__n29805 = ~ys__n4566 & new_new_n37717__;
  assign ys__n29807 = ys__n29806 & ~ys__n4566;
  assign ys__n29809 = ys__n29808 & ~ys__n4566;
  assign new_new_n37721__ = new_new_n21836__ & new_new_n21855__;
  assign new_new_n37722__ = ~new_new_n21881__ & new_new_n21884__;
  assign new_new_n37723__ = ~new_new_n21855__ & new_new_n37722__;
  assign new_new_n37724__ = ~new_new_n37721__ & ~new_new_n37723__;
  assign ys__n29811 = new_new_n37128__ & ~new_new_n37724__;
  assign ys__n29813 = ys__n29812 & ~ys__n4566;
  assign ys__n29814 = ys__n18118 & ~ys__n4566;
  assign ys__n29815 = ~ys__n28243 & ys__n23933;
  assign ys__n29816 = ~ys__n28243 & ys__n23936;
  assign ys__n29817 = ~ys__n28243 & ys__n23939;
  assign ys__n29818 = ~ys__n28243 & ys__n23942;
  assign ys__n29819 = ~ys__n28243 & ys__n23945;
  assign new_new_n37733__ = ~new_new_n37710__ & ~new_new_n37712__;
  assign ys__n29820 = ~ys__n28243 & ~new_new_n37733__;
  assign new_new_n37735__ = ~ys__n28243 & new_new_n21844__;
  assign new_new_n37736__ = new_new_n21855__ & new_new_n37735__;
  assign ys__n29821 = ~new_new_n21842__ & new_new_n37736__;
  assign new_new_n37738__ = new_new_n21832__ & new_new_n21855__;
  assign new_new_n37739__ = ~new_new_n21828__ & new_new_n37738__;
  assign new_new_n37740__ = ~new_new_n21877__ & new_new_n37712__;
  assign new_new_n37741__ = ~new_new_n37739__ & ~new_new_n37740__;
  assign ys__n29822 = ~ys__n28243 & ~new_new_n37741__;
  assign new_new_n37743__ = ~new_new_n21881__ & ~new_new_n37722__;
  assign new_new_n37744__ = ~ys__n28243 & ~new_new_n21855__;
  assign ys__n29823 = ~new_new_n37743__ & new_new_n37744__;
  assign new_new_n37746__ = ys__n29880 & ~new_new_n10603__;
  assign new_new_n37747__ = ys__n29881 & new_new_n10603__;
  assign ys__n29847 = new_new_n37746__ | new_new_n37747__;
  assign new_new_n37749__ = ys__n24389 & ~new_new_n12473__;
  assign new_new_n37750__ = new_new_n12473__ & ys__n24408;
  assign ys__n30010 = new_new_n37749__ | new_new_n37750__;
  assign new_new_n37752__ = ~new_new_n22613__ & ~new_new_n23445__;
  assign ys__n30080 = new_new_n23102__ | new_new_n37752__;
  assign new_new_n37754__ = ~new_new_n23143__ & ~new_new_n23442__;
  assign new_new_n37755__ = ~new_new_n36569__ & ~new_new_n37754__;
  assign ys__n30081 = ~new_new_n22613__ & ~new_new_n37755__;
  assign new_new_n37757__ = ~new_new_n23162__ & ~new_new_n23442__;
  assign new_new_n37758__ = ~new_new_n36591__ & ~new_new_n37757__;
  assign ys__n30082 = ~new_new_n22613__ & ~new_new_n37758__;
  assign new_new_n37760__ = ~new_new_n23181__ & ~new_new_n23442__;
  assign new_new_n37761__ = ~new_new_n36613__ & ~new_new_n37760__;
  assign ys__n30083 = ~new_new_n22613__ & ~new_new_n37761__;
  assign new_new_n37763__ = ~new_new_n23200__ & ~new_new_n23442__;
  assign new_new_n37764__ = ~new_new_n36635__ & ~new_new_n37763__;
  assign ys__n30084 = ~new_new_n22613__ & ~new_new_n37764__;
  assign new_new_n37766__ = ~new_new_n23219__ & ~new_new_n23442__;
  assign new_new_n37767__ = ~new_new_n36657__ & ~new_new_n37766__;
  assign ys__n30085 = ~new_new_n22613__ & ~new_new_n37767__;
  assign new_new_n37769__ = ~new_new_n23238__ & ~new_new_n23442__;
  assign new_new_n37770__ = ~new_new_n36679__ & ~new_new_n37769__;
  assign ys__n30086 = ~new_new_n22613__ & ~new_new_n37770__;
  assign new_new_n37772__ = ~new_new_n23257__ & ~new_new_n23442__;
  assign new_new_n37773__ = ~new_new_n36701__ & ~new_new_n37772__;
  assign ys__n30087 = ~new_new_n22613__ & ~new_new_n37773__;
  assign new_new_n37775__ = ~new_new_n22938__ & ~new_new_n23442__;
  assign new_new_n37776__ = ~new_new_n36752__ & ~new_new_n37775__;
  assign ys__n30089 = ~new_new_n22613__ & ~new_new_n37776__;
  assign new_new_n37778__ = ~new_new_n22956__ & ~new_new_n23442__;
  assign new_new_n37779__ = ~new_new_n36767__ & ~new_new_n37778__;
  assign ys__n30090 = ~new_new_n22613__ & ~new_new_n37779__;
  assign new_new_n37781__ = ~new_new_n22974__ & ~new_new_n23442__;
  assign new_new_n37782__ = ~new_new_n36782__ & ~new_new_n37781__;
  assign ys__n30091 = ~new_new_n22613__ & ~new_new_n37782__;
  assign new_new_n37784__ = ~new_new_n22992__ & ~new_new_n23442__;
  assign new_new_n37785__ = ~new_new_n36797__ & ~new_new_n37784__;
  assign ys__n30092 = ~new_new_n22613__ & ~new_new_n37785__;
  assign new_new_n37787__ = ~new_new_n23010__ & ~new_new_n23442__;
  assign new_new_n37788__ = ~new_new_n36812__ & ~new_new_n37787__;
  assign ys__n30093 = ~new_new_n22613__ & ~new_new_n37788__;
  assign new_new_n37790__ = ~new_new_n23028__ & ~new_new_n23442__;
  assign new_new_n37791__ = ~new_new_n36827__ & ~new_new_n37790__;
  assign ys__n30094 = ~new_new_n22613__ & ~new_new_n37791__;
  assign new_new_n37793__ = ~new_new_n23046__ & ~new_new_n23442__;
  assign new_new_n37794__ = ~new_new_n36842__ & ~new_new_n37793__;
  assign ys__n30095 = ~new_new_n22613__ & ~new_new_n37794__;
  assign new_new_n37796__ = ~new_new_n23064__ & ~new_new_n23442__;
  assign new_new_n37797__ = ~new_new_n36857__ & ~new_new_n37796__;
  assign ys__n30096 = ~new_new_n22613__ & ~new_new_n37797__;
  assign new_new_n37799__ = ~new_new_n22778__ & ~new_new_n23442__;
  assign new_new_n37800__ = ~new_new_n36876__ & ~new_new_n37799__;
  assign ys__n30098 = ~new_new_n22613__ & ~new_new_n37800__;
  assign new_new_n37802__ = ~new_new_n22793__ & ~new_new_n23442__;
  assign new_new_n37803__ = ~new_new_n36891__ & ~new_new_n37802__;
  assign ys__n30099 = ~new_new_n22613__ & ~new_new_n37803__;
  assign new_new_n37805__ = ~new_new_n22808__ & ~new_new_n23442__;
  assign new_new_n37806__ = ~new_new_n36906__ & ~new_new_n37805__;
  assign ys__n30100 = ~new_new_n22613__ & ~new_new_n37806__;
  assign new_new_n37808__ = ~new_new_n22823__ & ~new_new_n23442__;
  assign new_new_n37809__ = ~new_new_n36921__ & ~new_new_n37808__;
  assign ys__n30101 = ~new_new_n22613__ & ~new_new_n37809__;
  assign new_new_n37811__ = ~new_new_n22838__ & ~new_new_n23442__;
  assign new_new_n37812__ = ~new_new_n36936__ & ~new_new_n37811__;
  assign ys__n30102 = ~new_new_n22613__ & ~new_new_n37812__;
  assign new_new_n37814__ = ~new_new_n22853__ & ~new_new_n23442__;
  assign new_new_n37815__ = ~new_new_n36951__ & ~new_new_n37814__;
  assign ys__n30103 = ~new_new_n22613__ & ~new_new_n37815__;
  assign new_new_n37817__ = ~new_new_n22868__ & ~new_new_n23442__;
  assign new_new_n37818__ = ~new_new_n36966__ & ~new_new_n37817__;
  assign ys__n30104 = ~new_new_n22613__ & ~new_new_n37818__;
  assign new_new_n37820__ = ~new_new_n22883__ & ~new_new_n23442__;
  assign new_new_n37821__ = ~new_new_n36981__ & ~new_new_n37820__;
  assign ys__n30105 = ~new_new_n22613__ & ~new_new_n37821__;
  assign new_new_n37823__ = ~new_new_n22630__ & ~new_new_n23442__;
  assign new_new_n37824__ = ~new_new_n36996__ & ~new_new_n37823__;
  assign ys__n30106 = ~new_new_n22613__ & ~new_new_n37824__;
  assign new_new_n37826__ = ~new_new_n22645__ & ~new_new_n23442__;
  assign new_new_n37827__ = ~new_new_n37011__ & ~new_new_n37826__;
  assign ys__n30107 = ~new_new_n22613__ & ~new_new_n37827__;
  assign new_new_n37829__ = ~new_new_n22660__ & ~new_new_n23442__;
  assign new_new_n37830__ = ~new_new_n37026__ & ~new_new_n37829__;
  assign ys__n30108 = ~new_new_n22613__ & ~new_new_n37830__;
  assign new_new_n37832__ = ~new_new_n22675__ & ~new_new_n23442__;
  assign new_new_n37833__ = ~new_new_n37041__ & ~new_new_n37832__;
  assign ys__n30109 = ~new_new_n22613__ & ~new_new_n37833__;
  assign new_new_n37835__ = ~new_new_n22690__ & ~new_new_n23442__;
  assign new_new_n37836__ = ~new_new_n37056__ & ~new_new_n37835__;
  assign ys__n30110 = ~new_new_n22613__ & ~new_new_n37836__;
  assign new_new_n37838__ = ~new_new_n22705__ & ~new_new_n23442__;
  assign new_new_n37839__ = ~new_new_n37071__ & ~new_new_n37838__;
  assign ys__n30111 = ~new_new_n22613__ & ~new_new_n37839__;
  assign new_new_n37841__ = ~new_new_n22720__ & ~new_new_n23442__;
  assign new_new_n37842__ = ~new_new_n37086__ & ~new_new_n37841__;
  assign ys__n30112 = ~new_new_n22613__ & ~new_new_n37842__;
  assign new_new_n37844__ = ~new_new_n22735__ & ~new_new_n23442__;
  assign new_new_n37845__ = ~new_new_n37101__ & ~new_new_n37844__;
  assign ys__n30113 = ~new_new_n22613__ & ~new_new_n37845__;
  assign new_new_n37847__ = ~ys__n3039 & ys__n30080;
  assign new_new_n37848__ = ys__n3039 & ~new_new_n23112__;
  assign new_new_n37849__ = ~new_new_n37847__ & ~new_new_n37848__;
  assign new_new_n37850__ = ~ys__n740 & ~ys__n3039;
  assign new_new_n37851__ = ~new_new_n37849__ & new_new_n37850__;
  assign new_new_n37852__ = ys__n3039 & ~new_new_n37849__;
  assign ys__n30119 = new_new_n37851__ | new_new_n37852__;
  assign new_new_n37854__ = ~ys__n3039 & ys__n30081;
  assign new_new_n37855__ = ys__n3039 & ~new_new_n23132__;
  assign new_new_n37856__ = ~new_new_n37854__ & ~new_new_n37855__;
  assign new_new_n37857__ = new_new_n37850__ & ~new_new_n37856__;
  assign new_new_n37858__ = ys__n3039 & ~new_new_n37856__;
  assign ys__n30122 = new_new_n37857__ | new_new_n37858__;
  assign new_new_n37860__ = ~ys__n3039 & ys__n30082;
  assign new_new_n37861__ = ys__n3039 & ~new_new_n23151__;
  assign new_new_n37862__ = ~new_new_n37860__ & ~new_new_n37861__;
  assign new_new_n37863__ = new_new_n37850__ & ~new_new_n37862__;
  assign new_new_n37864__ = ys__n3039 & ~new_new_n37862__;
  assign ys__n30125 = new_new_n37863__ | new_new_n37864__;
  assign new_new_n37866__ = ~ys__n3039 & ys__n30083;
  assign new_new_n37867__ = ys__n3039 & ~new_new_n23170__;
  assign new_new_n37868__ = ~new_new_n37866__ & ~new_new_n37867__;
  assign new_new_n37869__ = new_new_n37850__ & ~new_new_n37868__;
  assign new_new_n37870__ = ys__n3039 & ~new_new_n37868__;
  assign ys__n30128 = new_new_n37869__ | new_new_n37870__;
  assign new_new_n37872__ = ~ys__n3039 & ys__n30084;
  assign new_new_n37873__ = ys__n3039 & ~new_new_n23189__;
  assign new_new_n37874__ = ~new_new_n37872__ & ~new_new_n37873__;
  assign new_new_n37875__ = new_new_n37850__ & ~new_new_n37874__;
  assign new_new_n37876__ = ys__n3039 & ~new_new_n37874__;
  assign ys__n30131 = new_new_n37875__ | new_new_n37876__;
  assign new_new_n37878__ = ~ys__n3039 & ys__n30085;
  assign new_new_n37879__ = ys__n3039 & ~new_new_n23208__;
  assign new_new_n37880__ = ~new_new_n37878__ & ~new_new_n37879__;
  assign new_new_n37881__ = new_new_n37850__ & ~new_new_n37880__;
  assign new_new_n37882__ = ys__n3039 & ~new_new_n37880__;
  assign ys__n30134 = new_new_n37881__ | new_new_n37882__;
  assign new_new_n37884__ = ~ys__n3039 & ys__n30086;
  assign new_new_n37885__ = ys__n3039 & ~new_new_n23227__;
  assign new_new_n37886__ = ~new_new_n37884__ & ~new_new_n37885__;
  assign new_new_n37887__ = new_new_n37850__ & ~new_new_n37886__;
  assign new_new_n37888__ = ys__n3039 & ~new_new_n37886__;
  assign ys__n30137 = new_new_n37887__ | new_new_n37888__;
  assign new_new_n37890__ = ~ys__n3039 & ys__n30087;
  assign new_new_n37891__ = ys__n3039 & ~new_new_n23246__;
  assign new_new_n37892__ = ~new_new_n37890__ & ~new_new_n37891__;
  assign new_new_n37893__ = new_new_n37850__ & ~new_new_n37892__;
  assign new_new_n37894__ = ys__n3039 & ~new_new_n37892__;
  assign ys__n30140 = new_new_n37893__ | new_new_n37894__;
  assign new_new_n37896__ = ~ys__n3039 & ys__n30089;
  assign new_new_n37897__ = ys__n3039 & ~new_new_n22927__;
  assign new_new_n37898__ = ~new_new_n37896__ & ~new_new_n37897__;
  assign new_new_n37899__ = new_new_n37850__ & ~new_new_n37898__;
  assign new_new_n37900__ = ys__n3039 & ~new_new_n37898__;
  assign ys__n30143 = new_new_n37899__ | new_new_n37900__;
  assign new_new_n37902__ = ~ys__n3039 & ys__n30090;
  assign new_new_n37903__ = ys__n3039 & ~new_new_n22945__;
  assign new_new_n37904__ = ~new_new_n37902__ & ~new_new_n37903__;
  assign new_new_n37905__ = new_new_n37850__ & ~new_new_n37904__;
  assign new_new_n37906__ = ys__n3039 & ~new_new_n37904__;
  assign ys__n30146 = new_new_n37905__ | new_new_n37906__;
  assign new_new_n37908__ = ~ys__n3039 & ys__n30091;
  assign new_new_n37909__ = ys__n3039 & ~new_new_n22963__;
  assign new_new_n37910__ = ~new_new_n37908__ & ~new_new_n37909__;
  assign new_new_n37911__ = new_new_n37850__ & ~new_new_n37910__;
  assign new_new_n37912__ = ys__n3039 & ~new_new_n37910__;
  assign ys__n30149 = new_new_n37911__ | new_new_n37912__;
  assign new_new_n37914__ = ~ys__n3039 & ys__n30092;
  assign new_new_n37915__ = ys__n3039 & ~new_new_n22981__;
  assign new_new_n37916__ = ~new_new_n37914__ & ~new_new_n37915__;
  assign new_new_n37917__ = new_new_n37850__ & ~new_new_n37916__;
  assign new_new_n37918__ = ys__n3039 & ~new_new_n37916__;
  assign ys__n30152 = new_new_n37917__ | new_new_n37918__;
  assign new_new_n37920__ = ~ys__n3039 & ys__n30093;
  assign new_new_n37921__ = ys__n3039 & ~new_new_n22999__;
  assign new_new_n37922__ = ~new_new_n37920__ & ~new_new_n37921__;
  assign new_new_n37923__ = new_new_n37850__ & ~new_new_n37922__;
  assign new_new_n37924__ = ys__n3039 & ~new_new_n37922__;
  assign ys__n30155 = new_new_n37923__ | new_new_n37924__;
  assign new_new_n37926__ = ~ys__n3039 & ys__n30094;
  assign new_new_n37927__ = ys__n3039 & ~new_new_n23017__;
  assign new_new_n37928__ = ~new_new_n37926__ & ~new_new_n37927__;
  assign new_new_n37929__ = new_new_n37850__ & ~new_new_n37928__;
  assign new_new_n37930__ = ys__n3039 & ~new_new_n37928__;
  assign ys__n30158 = new_new_n37929__ | new_new_n37930__;
  assign new_new_n37932__ = ~ys__n3039 & ys__n30095;
  assign new_new_n37933__ = ys__n3039 & ~new_new_n23035__;
  assign new_new_n37934__ = ~new_new_n37932__ & ~new_new_n37933__;
  assign new_new_n37935__ = new_new_n37850__ & ~new_new_n37934__;
  assign new_new_n37936__ = ys__n3039 & ~new_new_n37934__;
  assign ys__n30161 = new_new_n37935__ | new_new_n37936__;
  assign new_new_n37938__ = ~ys__n3039 & ys__n30096;
  assign new_new_n37939__ = ys__n3039 & ~new_new_n23053__;
  assign new_new_n37940__ = ~new_new_n37938__ & ~new_new_n37939__;
  assign new_new_n37941__ = new_new_n37850__ & ~new_new_n37940__;
  assign new_new_n37942__ = ys__n3039 & ~new_new_n37940__;
  assign ys__n30164 = new_new_n37941__ | new_new_n37942__;
  assign new_new_n37944__ = ~ys__n3039 & ys__n30098;
  assign new_new_n37945__ = ys__n3039 & ~new_new_n22767__;
  assign new_new_n37946__ = ~new_new_n37944__ & ~new_new_n37945__;
  assign new_new_n37947__ = new_new_n37850__ & ~new_new_n37946__;
  assign new_new_n37948__ = ys__n3039 & ~new_new_n37946__;
  assign ys__n30167 = new_new_n37947__ | new_new_n37948__;
  assign new_new_n37950__ = ~ys__n3039 & ys__n30099;
  assign new_new_n37951__ = ys__n3039 & ~new_new_n22782__;
  assign new_new_n37952__ = ~new_new_n37950__ & ~new_new_n37951__;
  assign new_new_n37953__ = new_new_n37850__ & ~new_new_n37952__;
  assign new_new_n37954__ = ys__n3039 & ~new_new_n37952__;
  assign ys__n30170 = new_new_n37953__ | new_new_n37954__;
  assign new_new_n37956__ = ~ys__n3039 & ys__n30100;
  assign new_new_n37957__ = ys__n3039 & ~new_new_n22797__;
  assign new_new_n37958__ = ~new_new_n37956__ & ~new_new_n37957__;
  assign new_new_n37959__ = new_new_n37850__ & ~new_new_n37958__;
  assign new_new_n37960__ = ys__n3039 & ~new_new_n37958__;
  assign ys__n30173 = new_new_n37959__ | new_new_n37960__;
  assign new_new_n37962__ = ~ys__n3039 & ys__n30101;
  assign new_new_n37963__ = ys__n3039 & ~new_new_n22812__;
  assign new_new_n37964__ = ~new_new_n37962__ & ~new_new_n37963__;
  assign new_new_n37965__ = new_new_n37850__ & ~new_new_n37964__;
  assign new_new_n37966__ = ys__n3039 & ~new_new_n37964__;
  assign ys__n30176 = new_new_n37965__ | new_new_n37966__;
  assign new_new_n37968__ = ~ys__n3039 & ys__n30102;
  assign new_new_n37969__ = ys__n3039 & ~new_new_n22827__;
  assign new_new_n37970__ = ~new_new_n37968__ & ~new_new_n37969__;
  assign new_new_n37971__ = new_new_n37850__ & ~new_new_n37970__;
  assign new_new_n37972__ = ys__n3039 & ~new_new_n37970__;
  assign ys__n30179 = new_new_n37971__ | new_new_n37972__;
  assign new_new_n37974__ = ~ys__n3039 & ys__n30103;
  assign new_new_n37975__ = ys__n3039 & ~new_new_n22842__;
  assign new_new_n37976__ = ~new_new_n37974__ & ~new_new_n37975__;
  assign new_new_n37977__ = new_new_n37850__ & ~new_new_n37976__;
  assign new_new_n37978__ = ys__n3039 & ~new_new_n37976__;
  assign ys__n30182 = new_new_n37977__ | new_new_n37978__;
  assign new_new_n37980__ = ~ys__n3039 & ys__n30104;
  assign new_new_n37981__ = ys__n3039 & ~new_new_n22857__;
  assign new_new_n37982__ = ~new_new_n37980__ & ~new_new_n37981__;
  assign new_new_n37983__ = new_new_n37850__ & ~new_new_n37982__;
  assign new_new_n37984__ = ys__n3039 & ~new_new_n37982__;
  assign ys__n30185 = new_new_n37983__ | new_new_n37984__;
  assign new_new_n37986__ = ~ys__n3039 & ys__n30105;
  assign new_new_n37987__ = ys__n3039 & ~new_new_n22872__;
  assign new_new_n37988__ = ~new_new_n37986__ & ~new_new_n37987__;
  assign new_new_n37989__ = new_new_n37850__ & ~new_new_n37988__;
  assign new_new_n37990__ = ys__n3039 & ~new_new_n37988__;
  assign ys__n30188 = new_new_n37989__ | new_new_n37990__;
  assign new_new_n37992__ = ~ys__n3039 & ys__n30106;
  assign new_new_n37993__ = ys__n3039 & ~new_new_n22608__;
  assign new_new_n37994__ = ~new_new_n37992__ & ~new_new_n37993__;
  assign new_new_n37995__ = new_new_n37850__ & ~new_new_n37994__;
  assign new_new_n37996__ = ys__n3039 & ~new_new_n37994__;
  assign ys__n30191 = new_new_n37995__ | new_new_n37996__;
  assign new_new_n37998__ = ~ys__n3039 & ys__n30107;
  assign new_new_n37999__ = ys__n3039 & ~new_new_n22634__;
  assign new_new_n38000__ = ~new_new_n37998__ & ~new_new_n37999__;
  assign new_new_n38001__ = new_new_n37850__ & ~new_new_n38000__;
  assign new_new_n38002__ = ys__n3039 & ~new_new_n38000__;
  assign ys__n30194 = new_new_n38001__ | new_new_n38002__;
  assign new_new_n38004__ = ~ys__n3039 & ys__n30108;
  assign new_new_n38005__ = ys__n3039 & ~new_new_n22649__;
  assign new_new_n38006__ = ~new_new_n38004__ & ~new_new_n38005__;
  assign new_new_n38007__ = new_new_n37850__ & ~new_new_n38006__;
  assign new_new_n38008__ = ys__n3039 & ~new_new_n38006__;
  assign ys__n30197 = new_new_n38007__ | new_new_n38008__;
  assign new_new_n38010__ = ~ys__n3039 & ys__n30109;
  assign new_new_n38011__ = ys__n3039 & ~new_new_n22664__;
  assign new_new_n38012__ = ~new_new_n38010__ & ~new_new_n38011__;
  assign new_new_n38013__ = new_new_n37850__ & ~new_new_n38012__;
  assign new_new_n38014__ = ys__n3039 & ~new_new_n38012__;
  assign ys__n30200 = new_new_n38013__ | new_new_n38014__;
  assign new_new_n38016__ = ~ys__n3039 & ys__n30110;
  assign new_new_n38017__ = ys__n3039 & ~new_new_n22679__;
  assign new_new_n38018__ = ~new_new_n38016__ & ~new_new_n38017__;
  assign new_new_n38019__ = new_new_n37850__ & ~new_new_n38018__;
  assign new_new_n38020__ = ys__n3039 & ~new_new_n38018__;
  assign ys__n30203 = new_new_n38019__ | new_new_n38020__;
  assign new_new_n38022__ = ~ys__n3039 & ys__n30111;
  assign new_new_n38023__ = ys__n3039 & ~new_new_n22694__;
  assign new_new_n38024__ = ~new_new_n38022__ & ~new_new_n38023__;
  assign new_new_n38025__ = new_new_n37850__ & ~new_new_n38024__;
  assign new_new_n38026__ = ys__n3039 & ~new_new_n38024__;
  assign ys__n30206 = new_new_n38025__ | new_new_n38026__;
  assign new_new_n38028__ = ~ys__n3039 & ys__n30112;
  assign new_new_n38029__ = ys__n3039 & ~new_new_n22709__;
  assign new_new_n38030__ = ~new_new_n38028__ & ~new_new_n38029__;
  assign new_new_n38031__ = new_new_n37850__ & ~new_new_n38030__;
  assign new_new_n38032__ = ys__n3039 & ~new_new_n38030__;
  assign ys__n30209 = new_new_n38031__ | new_new_n38032__;
  assign new_new_n38034__ = ~ys__n3039 & ys__n30113;
  assign new_new_n38035__ = ys__n3039 & ~new_new_n22724__;
  assign new_new_n38036__ = ~new_new_n38034__ & ~new_new_n38035__;
  assign new_new_n38037__ = new_new_n37850__ & ~new_new_n38036__;
  assign new_new_n38038__ = ys__n3039 & ~new_new_n38036__;
  assign ys__n30212 = new_new_n38037__ | new_new_n38038__;
  assign new_new_n38040__ = ys__n30220 & ~ys__n740;
  assign new_new_n38041__ = ~ys__n4566 & new_new_n38040__;
  assign new_new_n38042__ = ys__n30214 & ys__n740;
  assign ys__n30215 = new_new_n38041__ | new_new_n38042__;
  assign ys__n33414 = ~ys__n18120 & ~ys__n740;
  assign new_new_n38045__ = ys__n30225 & ys__n740;
  assign ys__n30226 = ys__n33414 | new_new_n38045__;
  assign new_new_n38047__ = ys__n352 & ys__n23335;
  assign new_new_n38048__ = new_new_n14002__ & new_new_n38047__;
  assign new_new_n38049__ = ~ys__n17867 & ~ys__n30334;
  assign new_new_n38050__ = ys__n17867 & ys__n30334;
  assign new_new_n38051__ = ~new_new_n38049__ & ~new_new_n38050__;
  assign new_new_n38052__ = ~ys__n17869 & ~ys__n30334;
  assign new_new_n38053__ = ys__n17869 & ys__n30334;
  assign new_new_n38054__ = ~new_new_n38052__ & ~new_new_n38053__;
  assign new_new_n38055__ = ~ys__n17803 & ~new_new_n38054__;
  assign new_new_n38056__ = ys__n17803 & new_new_n38054__;
  assign new_new_n38057__ = ~new_new_n38055__ & ~new_new_n38056__;
  assign new_new_n38058__ = ~new_new_n38051__ & new_new_n38057__;
  assign new_new_n38059__ = new_new_n38051__ & ~new_new_n38057__;
  assign new_new_n38060__ = ~new_new_n38058__ & ~new_new_n38059__;
  assign new_new_n38061__ = ~ys__n33581 & ~new_new_n38051__;
  assign new_new_n38062__ = ~ys__n17866 & ~ys__n30334;
  assign new_new_n38063__ = ys__n17866 & ys__n30334;
  assign new_new_n38064__ = ~new_new_n38062__ & ~new_new_n38063__;
  assign new_new_n38065__ = new_new_n38061__ & ~new_new_n38064__;
  assign new_new_n38066__ = new_new_n38051__ & new_new_n38064__;
  assign new_new_n38067__ = ys__n33581 & ~new_new_n38066__;
  assign new_new_n38068__ = ~new_new_n38065__ & ~new_new_n38067__;
  assign new_new_n38069__ = ~new_new_n38060__ & ~new_new_n38068__;
  assign new_new_n38070__ = new_new_n38060__ & ~new_new_n38068__;
  assign new_new_n38071__ = ~new_new_n38060__ & new_new_n38068__;
  assign new_new_n38072__ = ~new_new_n38070__ & ~new_new_n38071__;
  assign new_new_n38073__ = ys__n33581 & new_new_n38051__;
  assign new_new_n38074__ = ~new_new_n38061__ & ~new_new_n38073__;
  assign new_new_n38075__ = ~new_new_n38064__ & new_new_n38074__;
  assign new_new_n38076__ = new_new_n38064__ & ~new_new_n38074__;
  assign new_new_n38077__ = ~new_new_n38075__ & ~new_new_n38076__;
  assign new_new_n38078__ = ~ys__n33579 & ~new_new_n38064__;
  assign new_new_n38079__ = ~ys__n30334 & new_new_n38078__;
  assign new_new_n38080__ = ys__n30334 & new_new_n38064__;
  assign new_new_n38081__ = ys__n33579 & ~new_new_n38080__;
  assign new_new_n38082__ = ~new_new_n38079__ & ~new_new_n38081__;
  assign new_new_n38083__ = ~new_new_n38077__ & ~new_new_n38082__;
  assign new_new_n38084__ = ~new_new_n38072__ & new_new_n38083__;
  assign new_new_n38085__ = ~new_new_n38069__ & ~new_new_n38084__;
  assign new_new_n38086__ = ~ys__n17870 & ~ys__n30334;
  assign new_new_n38087__ = ys__n17870 & ys__n30334;
  assign new_new_n38088__ = ~new_new_n38086__ & ~new_new_n38087__;
  assign new_new_n38089__ = ~ys__n17872 & ~ys__n30334;
  assign new_new_n38090__ = ys__n17872 & ys__n30334;
  assign new_new_n38091__ = ~new_new_n38089__ & ~new_new_n38090__;
  assign new_new_n38092__ = ~ys__n17806 & ~new_new_n38091__;
  assign new_new_n38093__ = ys__n17806 & new_new_n38091__;
  assign new_new_n38094__ = ~new_new_n38092__ & ~new_new_n38093__;
  assign new_new_n38095__ = ~new_new_n38088__ & new_new_n38094__;
  assign new_new_n38096__ = new_new_n38088__ & ~new_new_n38094__;
  assign new_new_n38097__ = ~new_new_n38095__ & ~new_new_n38096__;
  assign new_new_n38098__ = ~ys__n17804 & ~new_new_n38088__;
  assign new_new_n38099__ = ~new_new_n38054__ & new_new_n38098__;
  assign new_new_n38100__ = new_new_n38054__ & new_new_n38088__;
  assign new_new_n38101__ = ys__n17804 & ~new_new_n38100__;
  assign new_new_n38102__ = ~new_new_n38099__ & ~new_new_n38101__;
  assign new_new_n38103__ = new_new_n38097__ & ~new_new_n38102__;
  assign new_new_n38104__ = ~new_new_n38097__ & new_new_n38102__;
  assign new_new_n38105__ = ~new_new_n38103__ & ~new_new_n38104__;
  assign new_new_n38106__ = ys__n17804 & new_new_n38088__;
  assign new_new_n38107__ = ~new_new_n38098__ & ~new_new_n38106__;
  assign new_new_n38108__ = ~new_new_n38054__ & new_new_n38107__;
  assign new_new_n38109__ = new_new_n38054__ & ~new_new_n38107__;
  assign new_new_n38110__ = ~new_new_n38108__ & ~new_new_n38109__;
  assign new_new_n38111__ = ~new_new_n38051__ & new_new_n38055__;
  assign new_new_n38112__ = new_new_n38051__ & new_new_n38054__;
  assign new_new_n38113__ = ys__n17803 & ~new_new_n38112__;
  assign new_new_n38114__ = ~new_new_n38111__ & ~new_new_n38113__;
  assign new_new_n38115__ = new_new_n38110__ & ~new_new_n38114__;
  assign new_new_n38116__ = ~new_new_n38110__ & new_new_n38114__;
  assign new_new_n38117__ = ~new_new_n38115__ & ~new_new_n38116__;
  assign new_new_n38118__ = ~new_new_n38105__ & ~new_new_n38117__;
  assign new_new_n38119__ = ~new_new_n38085__ & new_new_n38118__;
  assign new_new_n38120__ = ~new_new_n38097__ & ~new_new_n38102__;
  assign new_new_n38121__ = ~new_new_n38110__ & ~new_new_n38114__;
  assign new_new_n38122__ = ~new_new_n38105__ & new_new_n38121__;
  assign new_new_n38123__ = ~new_new_n38120__ & ~new_new_n38122__;
  assign new_new_n38124__ = ~new_new_n38119__ & new_new_n38123__;
  assign new_new_n38125__ = ~ys__n17876 & ~ys__n30334;
  assign new_new_n38126__ = ys__n17876 & ys__n30334;
  assign new_new_n38127__ = ~new_new_n38125__ & ~new_new_n38126__;
  assign new_new_n38128__ = ~ys__n17878 & ~ys__n30334;
  assign new_new_n38129__ = ys__n17878 & ys__n30334;
  assign new_new_n38130__ = ~new_new_n38128__ & ~new_new_n38129__;
  assign new_new_n38131__ = ~ys__n17812 & ~new_new_n38130__;
  assign new_new_n38132__ = ys__n17812 & new_new_n38130__;
  assign new_new_n38133__ = ~new_new_n38131__ & ~new_new_n38132__;
  assign new_new_n38134__ = ~new_new_n38127__ & new_new_n38133__;
  assign new_new_n38135__ = new_new_n38127__ & ~new_new_n38133__;
  assign new_new_n38136__ = ~new_new_n38134__ & ~new_new_n38135__;
  assign new_new_n38137__ = ~ys__n17810 & ~new_new_n38127__;
  assign new_new_n38138__ = ~ys__n17875 & ~ys__n30334;
  assign new_new_n38139__ = ys__n17875 & ys__n30334;
  assign new_new_n38140__ = ~new_new_n38138__ & ~new_new_n38139__;
  assign new_new_n38141__ = new_new_n38137__ & ~new_new_n38140__;
  assign new_new_n38142__ = new_new_n38127__ & new_new_n38140__;
  assign new_new_n38143__ = ys__n17810 & ~new_new_n38142__;
  assign new_new_n38144__ = ~new_new_n38141__ & ~new_new_n38143__;
  assign new_new_n38145__ = new_new_n38136__ & ~new_new_n38144__;
  assign new_new_n38146__ = ~new_new_n38136__ & new_new_n38144__;
  assign new_new_n38147__ = ~new_new_n38145__ & ~new_new_n38146__;
  assign new_new_n38148__ = ys__n17810 & new_new_n38127__;
  assign new_new_n38149__ = ~new_new_n38137__ & ~new_new_n38148__;
  assign new_new_n38150__ = ~new_new_n38140__ & new_new_n38149__;
  assign new_new_n38151__ = new_new_n38140__ & ~new_new_n38149__;
  assign new_new_n38152__ = ~new_new_n38150__ & ~new_new_n38151__;
  assign new_new_n38153__ = ~ys__n17809 & ~new_new_n38140__;
  assign new_new_n38154__ = ~ys__n17873 & ~ys__n30334;
  assign new_new_n38155__ = ys__n17873 & ys__n30334;
  assign new_new_n38156__ = ~new_new_n38154__ & ~new_new_n38155__;
  assign new_new_n38157__ = new_new_n38153__ & ~new_new_n38156__;
  assign new_new_n38158__ = new_new_n38140__ & new_new_n38156__;
  assign new_new_n38159__ = ys__n17809 & ~new_new_n38158__;
  assign new_new_n38160__ = ~new_new_n38157__ & ~new_new_n38159__;
  assign new_new_n38161__ = new_new_n38152__ & ~new_new_n38160__;
  assign new_new_n38162__ = ~new_new_n38152__ & new_new_n38160__;
  assign new_new_n38163__ = ~new_new_n38161__ & ~new_new_n38162__;
  assign new_new_n38164__ = ~new_new_n38147__ & ~new_new_n38163__;
  assign new_new_n38165__ = ys__n17809 & new_new_n38140__;
  assign new_new_n38166__ = ~new_new_n38153__ & ~new_new_n38165__;
  assign new_new_n38167__ = ~new_new_n38156__ & new_new_n38166__;
  assign new_new_n38168__ = new_new_n38156__ & ~new_new_n38166__;
  assign new_new_n38169__ = ~new_new_n38167__ & ~new_new_n38168__;
  assign new_new_n38170__ = ~ys__n17807 & ~new_new_n38156__;
  assign new_new_n38171__ = ~new_new_n38091__ & new_new_n38170__;
  assign new_new_n38172__ = new_new_n38091__ & new_new_n38156__;
  assign new_new_n38173__ = ys__n17807 & ~new_new_n38172__;
  assign new_new_n38174__ = ~new_new_n38171__ & ~new_new_n38173__;
  assign new_new_n38175__ = new_new_n38169__ & ~new_new_n38174__;
  assign new_new_n38176__ = ~new_new_n38169__ & new_new_n38174__;
  assign new_new_n38177__ = ~new_new_n38175__ & ~new_new_n38176__;
  assign new_new_n38178__ = ys__n17807 & new_new_n38156__;
  assign new_new_n38179__ = ~new_new_n38170__ & ~new_new_n38178__;
  assign new_new_n38180__ = ~new_new_n38091__ & new_new_n38179__;
  assign new_new_n38181__ = new_new_n38091__ & ~new_new_n38179__;
  assign new_new_n38182__ = ~new_new_n38180__ & ~new_new_n38181__;
  assign new_new_n38183__ = ~new_new_n38088__ & new_new_n38092__;
  assign new_new_n38184__ = new_new_n38088__ & new_new_n38091__;
  assign new_new_n38185__ = ys__n17806 & ~new_new_n38184__;
  assign new_new_n38186__ = ~new_new_n38183__ & ~new_new_n38185__;
  assign new_new_n38187__ = new_new_n38182__ & ~new_new_n38186__;
  assign new_new_n38188__ = ~new_new_n38182__ & new_new_n38186__;
  assign new_new_n38189__ = ~new_new_n38187__ & ~new_new_n38188__;
  assign new_new_n38190__ = ~new_new_n38177__ & ~new_new_n38189__;
  assign new_new_n38191__ = new_new_n38164__ & new_new_n38190__;
  assign new_new_n38192__ = ~new_new_n38124__ & new_new_n38191__;
  assign new_new_n38193__ = ~new_new_n38169__ & ~new_new_n38174__;
  assign new_new_n38194__ = ~new_new_n38182__ & ~new_new_n38186__;
  assign new_new_n38195__ = ~new_new_n38177__ & new_new_n38194__;
  assign new_new_n38196__ = ~new_new_n38193__ & ~new_new_n38195__;
  assign new_new_n38197__ = new_new_n38164__ & ~new_new_n38196__;
  assign new_new_n38198__ = ~new_new_n38136__ & ~new_new_n38144__;
  assign new_new_n38199__ = ~new_new_n38152__ & ~new_new_n38160__;
  assign new_new_n38200__ = ~new_new_n38147__ & new_new_n38199__;
  assign new_new_n38201__ = ~new_new_n38198__ & ~new_new_n38200__;
  assign new_new_n38202__ = ~new_new_n38197__ & new_new_n38201__;
  assign new_new_n38203__ = ~new_new_n38192__ & new_new_n38202__;
  assign new_new_n38204__ = ~ys__n17888 & ~ys__n30334;
  assign new_new_n38205__ = ys__n17888 & ys__n30334;
  assign new_new_n38206__ = ~new_new_n38204__ & ~new_new_n38205__;
  assign new_new_n38207__ = ~ys__n17890 & ~ys__n30334;
  assign new_new_n38208__ = ys__n17890 & ys__n30334;
  assign new_new_n38209__ = ~new_new_n38207__ & ~new_new_n38208__;
  assign new_new_n38210__ = ~ys__n17824 & ~new_new_n38209__;
  assign new_new_n38211__ = ys__n17824 & new_new_n38209__;
  assign new_new_n38212__ = ~new_new_n38210__ & ~new_new_n38211__;
  assign new_new_n38213__ = ~new_new_n38206__ & new_new_n38212__;
  assign new_new_n38214__ = new_new_n38206__ & ~new_new_n38212__;
  assign new_new_n38215__ = ~new_new_n38213__ & ~new_new_n38214__;
  assign new_new_n38216__ = ~ys__n17822 & ~new_new_n38206__;
  assign new_new_n38217__ = ~ys__n17887 & ~ys__n30334;
  assign new_new_n38218__ = ys__n17887 & ys__n30334;
  assign new_new_n38219__ = ~new_new_n38217__ & ~new_new_n38218__;
  assign new_new_n38220__ = new_new_n38216__ & ~new_new_n38219__;
  assign new_new_n38221__ = new_new_n38206__ & new_new_n38219__;
  assign new_new_n38222__ = ys__n17822 & ~new_new_n38221__;
  assign new_new_n38223__ = ~new_new_n38220__ & ~new_new_n38222__;
  assign new_new_n38224__ = new_new_n38215__ & ~new_new_n38223__;
  assign new_new_n38225__ = ~new_new_n38215__ & new_new_n38223__;
  assign new_new_n38226__ = ~new_new_n38224__ & ~new_new_n38225__;
  assign new_new_n38227__ = ys__n17822 & new_new_n38206__;
  assign new_new_n38228__ = ~new_new_n38216__ & ~new_new_n38227__;
  assign new_new_n38229__ = ~new_new_n38219__ & new_new_n38228__;
  assign new_new_n38230__ = new_new_n38219__ & ~new_new_n38228__;
  assign new_new_n38231__ = ~new_new_n38229__ & ~new_new_n38230__;
  assign new_new_n38232__ = ~ys__n17821 & ~new_new_n38219__;
  assign new_new_n38233__ = ~ys__n17885 & ~ys__n30334;
  assign new_new_n38234__ = ys__n17885 & ys__n30334;
  assign new_new_n38235__ = ~new_new_n38233__ & ~new_new_n38234__;
  assign new_new_n38236__ = new_new_n38232__ & ~new_new_n38235__;
  assign new_new_n38237__ = new_new_n38219__ & new_new_n38235__;
  assign new_new_n38238__ = ys__n17821 & ~new_new_n38237__;
  assign new_new_n38239__ = ~new_new_n38236__ & ~new_new_n38238__;
  assign new_new_n38240__ = new_new_n38231__ & ~new_new_n38239__;
  assign new_new_n38241__ = ~new_new_n38231__ & new_new_n38239__;
  assign new_new_n38242__ = ~new_new_n38240__ & ~new_new_n38241__;
  assign new_new_n38243__ = ~new_new_n38226__ & ~new_new_n38242__;
  assign new_new_n38244__ = ys__n17821 & new_new_n38219__;
  assign new_new_n38245__ = ~new_new_n38232__ & ~new_new_n38244__;
  assign new_new_n38246__ = ~new_new_n38235__ & new_new_n38245__;
  assign new_new_n38247__ = new_new_n38235__ & ~new_new_n38245__;
  assign new_new_n38248__ = ~new_new_n38246__ & ~new_new_n38247__;
  assign new_new_n38249__ = ~ys__n17819 & ~new_new_n38235__;
  assign new_new_n38250__ = ~ys__n17884 & ~ys__n30334;
  assign new_new_n38251__ = ys__n17884 & ys__n30334;
  assign new_new_n38252__ = ~new_new_n38250__ & ~new_new_n38251__;
  assign new_new_n38253__ = new_new_n38249__ & ~new_new_n38252__;
  assign new_new_n38254__ = new_new_n38235__ & new_new_n38252__;
  assign new_new_n38255__ = ys__n17819 & ~new_new_n38254__;
  assign new_new_n38256__ = ~new_new_n38253__ & ~new_new_n38255__;
  assign new_new_n38257__ = new_new_n38248__ & ~new_new_n38256__;
  assign new_new_n38258__ = ~new_new_n38248__ & new_new_n38256__;
  assign new_new_n38259__ = ~new_new_n38257__ & ~new_new_n38258__;
  assign new_new_n38260__ = ys__n17819 & new_new_n38235__;
  assign new_new_n38261__ = ~new_new_n38249__ & ~new_new_n38260__;
  assign new_new_n38262__ = ~new_new_n38252__ & new_new_n38261__;
  assign new_new_n38263__ = new_new_n38252__ & ~new_new_n38261__;
  assign new_new_n38264__ = ~new_new_n38262__ & ~new_new_n38263__;
  assign new_new_n38265__ = ~ys__n17818 & ~new_new_n38252__;
  assign new_new_n38266__ = ~ys__n17882 & ~ys__n30334;
  assign new_new_n38267__ = ys__n17882 & ys__n30334;
  assign new_new_n38268__ = ~new_new_n38266__ & ~new_new_n38267__;
  assign new_new_n38269__ = new_new_n38265__ & ~new_new_n38268__;
  assign new_new_n38270__ = new_new_n38252__ & new_new_n38268__;
  assign new_new_n38271__ = ys__n17818 & ~new_new_n38270__;
  assign new_new_n38272__ = ~new_new_n38269__ & ~new_new_n38271__;
  assign new_new_n38273__ = new_new_n38264__ & ~new_new_n38272__;
  assign new_new_n38274__ = ~new_new_n38264__ & new_new_n38272__;
  assign new_new_n38275__ = ~new_new_n38273__ & ~new_new_n38274__;
  assign new_new_n38276__ = ~new_new_n38259__ & ~new_new_n38275__;
  assign new_new_n38277__ = new_new_n38243__ & new_new_n38276__;
  assign new_new_n38278__ = ys__n17818 & new_new_n38252__;
  assign new_new_n38279__ = ~new_new_n38265__ & ~new_new_n38278__;
  assign new_new_n38280__ = ~new_new_n38268__ & new_new_n38279__;
  assign new_new_n38281__ = new_new_n38268__ & ~new_new_n38279__;
  assign new_new_n38282__ = ~new_new_n38280__ & ~new_new_n38281__;
  assign new_new_n38283__ = ~ys__n17816 & ~new_new_n38268__;
  assign new_new_n38284__ = ~ys__n17881 & ~ys__n30334;
  assign new_new_n38285__ = ys__n17881 & ys__n30334;
  assign new_new_n38286__ = ~new_new_n38284__ & ~new_new_n38285__;
  assign new_new_n38287__ = new_new_n38283__ & ~new_new_n38286__;
  assign new_new_n38288__ = new_new_n38268__ & new_new_n38286__;
  assign new_new_n38289__ = ys__n17816 & ~new_new_n38288__;
  assign new_new_n38290__ = ~new_new_n38287__ & ~new_new_n38289__;
  assign new_new_n38291__ = new_new_n38282__ & ~new_new_n38290__;
  assign new_new_n38292__ = ~new_new_n38282__ & new_new_n38290__;
  assign new_new_n38293__ = ~new_new_n38291__ & ~new_new_n38292__;
  assign new_new_n38294__ = ys__n17816 & new_new_n38268__;
  assign new_new_n38295__ = ~new_new_n38283__ & ~new_new_n38294__;
  assign new_new_n38296__ = ~new_new_n38286__ & new_new_n38295__;
  assign new_new_n38297__ = new_new_n38286__ & ~new_new_n38295__;
  assign new_new_n38298__ = ~new_new_n38296__ & ~new_new_n38297__;
  assign new_new_n38299__ = ~ys__n17815 & ~new_new_n38286__;
  assign new_new_n38300__ = ~ys__n17879 & ~ys__n30334;
  assign new_new_n38301__ = ys__n17879 & ys__n30334;
  assign new_new_n38302__ = ~new_new_n38300__ & ~new_new_n38301__;
  assign new_new_n38303__ = new_new_n38299__ & ~new_new_n38302__;
  assign new_new_n38304__ = new_new_n38286__ & new_new_n38302__;
  assign new_new_n38305__ = ys__n17815 & ~new_new_n38304__;
  assign new_new_n38306__ = ~new_new_n38303__ & ~new_new_n38305__;
  assign new_new_n38307__ = new_new_n38298__ & ~new_new_n38306__;
  assign new_new_n38308__ = ~new_new_n38298__ & new_new_n38306__;
  assign new_new_n38309__ = ~new_new_n38307__ & ~new_new_n38308__;
  assign new_new_n38310__ = ~new_new_n38293__ & ~new_new_n38309__;
  assign new_new_n38311__ = ys__n17815 & new_new_n38286__;
  assign new_new_n38312__ = ~new_new_n38299__ & ~new_new_n38311__;
  assign new_new_n38313__ = ~new_new_n38302__ & new_new_n38312__;
  assign new_new_n38314__ = new_new_n38302__ & ~new_new_n38312__;
  assign new_new_n38315__ = ~new_new_n38313__ & ~new_new_n38314__;
  assign new_new_n38316__ = ~ys__n17813 & ~new_new_n38302__;
  assign new_new_n38317__ = ~new_new_n38130__ & new_new_n38316__;
  assign new_new_n38318__ = new_new_n38130__ & new_new_n38302__;
  assign new_new_n38319__ = ys__n17813 & ~new_new_n38318__;
  assign new_new_n38320__ = ~new_new_n38317__ & ~new_new_n38319__;
  assign new_new_n38321__ = new_new_n38315__ & ~new_new_n38320__;
  assign new_new_n38322__ = ~new_new_n38315__ & new_new_n38320__;
  assign new_new_n38323__ = ~new_new_n38321__ & ~new_new_n38322__;
  assign new_new_n38324__ = ys__n17813 & new_new_n38302__;
  assign new_new_n38325__ = ~new_new_n38316__ & ~new_new_n38324__;
  assign new_new_n38326__ = ~new_new_n38130__ & new_new_n38325__;
  assign new_new_n38327__ = new_new_n38130__ & ~new_new_n38325__;
  assign new_new_n38328__ = ~new_new_n38326__ & ~new_new_n38327__;
  assign new_new_n38329__ = ~new_new_n38127__ & new_new_n38131__;
  assign new_new_n38330__ = new_new_n38127__ & new_new_n38130__;
  assign new_new_n38331__ = ys__n17812 & ~new_new_n38330__;
  assign new_new_n38332__ = ~new_new_n38329__ & ~new_new_n38331__;
  assign new_new_n38333__ = new_new_n38328__ & ~new_new_n38332__;
  assign new_new_n38334__ = ~new_new_n38328__ & new_new_n38332__;
  assign new_new_n38335__ = ~new_new_n38333__ & ~new_new_n38334__;
  assign new_new_n38336__ = ~new_new_n38323__ & ~new_new_n38335__;
  assign new_new_n38337__ = new_new_n38310__ & new_new_n38336__;
  assign new_new_n38338__ = new_new_n38277__ & new_new_n38337__;
  assign new_new_n38339__ = ~new_new_n38203__ & new_new_n38338__;
  assign new_new_n38340__ = ~new_new_n38315__ & ~new_new_n38320__;
  assign new_new_n38341__ = ~new_new_n38328__ & ~new_new_n38332__;
  assign new_new_n38342__ = ~new_new_n38323__ & new_new_n38341__;
  assign new_new_n38343__ = ~new_new_n38340__ & ~new_new_n38342__;
  assign new_new_n38344__ = new_new_n38310__ & ~new_new_n38343__;
  assign new_new_n38345__ = ~new_new_n38282__ & ~new_new_n38290__;
  assign new_new_n38346__ = ~new_new_n38298__ & ~new_new_n38306__;
  assign new_new_n38347__ = ~new_new_n38293__ & new_new_n38346__;
  assign new_new_n38348__ = ~new_new_n38345__ & ~new_new_n38347__;
  assign new_new_n38349__ = ~new_new_n38344__ & new_new_n38348__;
  assign new_new_n38350__ = new_new_n38277__ & ~new_new_n38349__;
  assign new_new_n38351__ = ~new_new_n38248__ & ~new_new_n38256__;
  assign new_new_n38352__ = ~new_new_n38264__ & ~new_new_n38272__;
  assign new_new_n38353__ = ~new_new_n38259__ & new_new_n38352__;
  assign new_new_n38354__ = ~new_new_n38351__ & ~new_new_n38353__;
  assign new_new_n38355__ = new_new_n38243__ & ~new_new_n38354__;
  assign new_new_n38356__ = ~new_new_n38215__ & ~new_new_n38223__;
  assign new_new_n38357__ = ~new_new_n38231__ & ~new_new_n38239__;
  assign new_new_n38358__ = ~new_new_n38226__ & new_new_n38357__;
  assign new_new_n38359__ = ~new_new_n38356__ & ~new_new_n38358__;
  assign new_new_n38360__ = ~new_new_n38355__ & new_new_n38359__;
  assign new_new_n38361__ = ~new_new_n38350__ & new_new_n38360__;
  assign new_new_n38362__ = ~new_new_n38339__ & new_new_n38361__;
  assign new_new_n38363__ = ~new_new_n38203__ & new_new_n38337__;
  assign new_new_n38364__ = new_new_n38349__ & ~new_new_n38363__;
  assign new_new_n38365__ = new_new_n38276__ & ~new_new_n38364__;
  assign new_new_n38366__ = new_new_n38354__ & ~new_new_n38365__;
  assign new_new_n38367__ = ~new_new_n38242__ & ~new_new_n38366__;
  assign new_new_n38368__ = ~new_new_n38357__ & ~new_new_n38367__;
  assign new_new_n38369__ = new_new_n38226__ & ~new_new_n38368__;
  assign new_new_n38370__ = ~new_new_n38226__ & new_new_n38368__;
  assign new_new_n38371__ = ~new_new_n38369__ & ~new_new_n38370__;
  assign new_new_n38372__ = ~new_new_n38203__ & new_new_n38336__;
  assign new_new_n38373__ = new_new_n38343__ & ~new_new_n38372__;
  assign new_new_n38374__ = ~new_new_n38309__ & ~new_new_n38373__;
  assign new_new_n38375__ = ~new_new_n38346__ & ~new_new_n38374__;
  assign new_new_n38376__ = new_new_n38293__ & ~new_new_n38375__;
  assign new_new_n38377__ = ~new_new_n38293__ & new_new_n38375__;
  assign new_new_n38378__ = ~new_new_n38376__ & ~new_new_n38377__;
  assign new_new_n38379__ = new_new_n38309__ & ~new_new_n38373__;
  assign new_new_n38380__ = ~new_new_n38309__ & new_new_n38373__;
  assign new_new_n38381__ = ~new_new_n38379__ & ~new_new_n38380__;
  assign new_new_n38382__ = ~new_new_n38203__ & ~new_new_n38335__;
  assign new_new_n38383__ = ~new_new_n38341__ & ~new_new_n38382__;
  assign new_new_n38384__ = new_new_n38323__ & ~new_new_n38383__;
  assign new_new_n38385__ = ~new_new_n38323__ & new_new_n38383__;
  assign new_new_n38386__ = ~new_new_n38384__ & ~new_new_n38385__;
  assign new_new_n38387__ = ~new_new_n38203__ & new_new_n38335__;
  assign new_new_n38388__ = new_new_n38203__ & ~new_new_n38335__;
  assign new_new_n38389__ = ~new_new_n38387__ & ~new_new_n38388__;
  assign new_new_n38390__ = ~new_new_n38386__ & ~new_new_n38389__;
  assign new_new_n38391__ = ~new_new_n38381__ & new_new_n38390__;
  assign new_new_n38392__ = ~new_new_n38378__ & new_new_n38391__;
  assign new_new_n38393__ = ~new_new_n38275__ & ~new_new_n38364__;
  assign new_new_n38394__ = ~new_new_n38352__ & ~new_new_n38393__;
  assign new_new_n38395__ = new_new_n38259__ & ~new_new_n38394__;
  assign new_new_n38396__ = ~new_new_n38259__ & new_new_n38394__;
  assign new_new_n38397__ = ~new_new_n38395__ & ~new_new_n38396__;
  assign new_new_n38398__ = new_new_n38275__ & ~new_new_n38364__;
  assign new_new_n38399__ = ~new_new_n38275__ & new_new_n38364__;
  assign new_new_n38400__ = ~new_new_n38398__ & ~new_new_n38399__;
  assign new_new_n38401__ = ~new_new_n38397__ & ~new_new_n38400__;
  assign new_new_n38402__ = new_new_n38242__ & ~new_new_n38366__;
  assign new_new_n38403__ = ~new_new_n38242__ & new_new_n38366__;
  assign new_new_n38404__ = ~new_new_n38402__ & ~new_new_n38403__;
  assign new_new_n38405__ = ~new_new_n38124__ & new_new_n38190__;
  assign new_new_n38406__ = new_new_n38196__ & ~new_new_n38405__;
  assign new_new_n38407__ = ~new_new_n38163__ & ~new_new_n38406__;
  assign new_new_n38408__ = ~new_new_n38199__ & ~new_new_n38407__;
  assign new_new_n38409__ = new_new_n38147__ & ~new_new_n38408__;
  assign new_new_n38410__ = ~new_new_n38147__ & new_new_n38408__;
  assign new_new_n38411__ = ~new_new_n38409__ & ~new_new_n38410__;
  assign new_new_n38412__ = ~new_new_n38124__ & ~new_new_n38189__;
  assign new_new_n38413__ = ~new_new_n38194__ & ~new_new_n38412__;
  assign new_new_n38414__ = new_new_n38177__ & ~new_new_n38413__;
  assign new_new_n38415__ = ~new_new_n38177__ & new_new_n38413__;
  assign new_new_n38416__ = ~new_new_n38414__ & ~new_new_n38415__;
  assign new_new_n38417__ = ~new_new_n38124__ & new_new_n38189__;
  assign new_new_n38418__ = new_new_n38124__ & ~new_new_n38189__;
  assign new_new_n38419__ = ~new_new_n38417__ & ~new_new_n38418__;
  assign new_new_n38420__ = ~new_new_n38416__ & ~new_new_n38419__;
  assign new_new_n38421__ = new_new_n38163__ & ~new_new_n38406__;
  assign new_new_n38422__ = ~new_new_n38163__ & new_new_n38406__;
  assign new_new_n38423__ = ~new_new_n38421__ & ~new_new_n38422__;
  assign new_new_n38424__ = ~new_new_n38085__ & ~new_new_n38117__;
  assign new_new_n38425__ = ~new_new_n38121__ & ~new_new_n38424__;
  assign new_new_n38426__ = new_new_n38105__ & ~new_new_n38425__;
  assign new_new_n38427__ = ~new_new_n38105__ & new_new_n38425__;
  assign new_new_n38428__ = ~new_new_n38426__ & ~new_new_n38427__;
  assign new_new_n38429__ = ~new_new_n38085__ & new_new_n38117__;
  assign new_new_n38430__ = new_new_n38085__ & ~new_new_n38117__;
  assign new_new_n38431__ = ~new_new_n38429__ & ~new_new_n38430__;
  assign new_new_n38432__ = new_new_n38072__ & new_new_n38083__;
  assign new_new_n38433__ = ~new_new_n38072__ & ~new_new_n38083__;
  assign new_new_n38434__ = ~new_new_n38432__ & ~new_new_n38433__;
  assign new_new_n38435__ = new_new_n38077__ & ~new_new_n38082__;
  assign new_new_n38436__ = ~new_new_n38077__ & new_new_n38082__;
  assign new_new_n38437__ = ~new_new_n38435__ & ~new_new_n38436__;
  assign new_new_n38438__ = ~ys__n30334 & ~new_new_n38437__;
  assign new_new_n38439__ = ~new_new_n38434__ & new_new_n38438__;
  assign new_new_n38440__ = ~new_new_n38431__ & new_new_n38439__;
  assign new_new_n38441__ = ~new_new_n38428__ & new_new_n38440__;
  assign new_new_n38442__ = ~new_new_n38423__ & new_new_n38441__;
  assign new_new_n38443__ = new_new_n38420__ & new_new_n38442__;
  assign new_new_n38444__ = ~new_new_n38411__ & new_new_n38443__;
  assign new_new_n38445__ = ~new_new_n38404__ & new_new_n38444__;
  assign new_new_n38446__ = new_new_n38401__ & new_new_n38445__;
  assign new_new_n38447__ = new_new_n38392__ & new_new_n38446__;
  assign new_new_n38448__ = ~new_new_n38371__ & new_new_n38447__;
  assign new_new_n38449__ = new_new_n38362__ & new_new_n38448__;
  assign new_new_n38450__ = ~new_new_n38362__ & ~new_new_n38448__;
  assign new_new_n38451__ = ~new_new_n38449__ & ~new_new_n38450__;
  assign new_new_n38452__ = ~ys__n17912 & ~ys__n30334;
  assign new_new_n38453__ = ys__n17912 & ys__n30334;
  assign new_new_n38454__ = ~new_new_n38452__ & ~new_new_n38453__;
  assign new_new_n38455__ = ~ys__n30333 & ~ys__n30334;
  assign new_new_n38456__ = ys__n30333 & ys__n30334;
  assign new_new_n38457__ = ~new_new_n38455__ & ~new_new_n38456__;
  assign new_new_n38458__ = ~ys__n17848 & ~new_new_n38457__;
  assign new_new_n38459__ = ys__n17848 & new_new_n38457__;
  assign new_new_n38460__ = ~new_new_n38458__ & ~new_new_n38459__;
  assign new_new_n38461__ = ~new_new_n38454__ & new_new_n38460__;
  assign new_new_n38462__ = new_new_n38454__ & ~new_new_n38460__;
  assign new_new_n38463__ = ~new_new_n38461__ & ~new_new_n38462__;
  assign new_new_n38464__ = ~ys__n17846 & ~new_new_n38454__;
  assign new_new_n38465__ = ~ys__n17911 & ~ys__n30334;
  assign new_new_n38466__ = ys__n17911 & ys__n30334;
  assign new_new_n38467__ = ~new_new_n38465__ & ~new_new_n38466__;
  assign new_new_n38468__ = new_new_n38464__ & ~new_new_n38467__;
  assign new_new_n38469__ = new_new_n38454__ & new_new_n38467__;
  assign new_new_n38470__ = ys__n17846 & ~new_new_n38469__;
  assign new_new_n38471__ = ~new_new_n38468__ & ~new_new_n38470__;
  assign new_new_n38472__ = new_new_n38463__ & ~new_new_n38471__;
  assign new_new_n38473__ = ~new_new_n38463__ & new_new_n38471__;
  assign new_new_n38474__ = ~new_new_n38472__ & ~new_new_n38473__;
  assign new_new_n38475__ = ys__n17846 & new_new_n38454__;
  assign new_new_n38476__ = ~new_new_n38464__ & ~new_new_n38475__;
  assign new_new_n38477__ = ~new_new_n38467__ & new_new_n38476__;
  assign new_new_n38478__ = new_new_n38467__ & ~new_new_n38476__;
  assign new_new_n38479__ = ~new_new_n38477__ & ~new_new_n38478__;
  assign new_new_n38480__ = ~ys__n17845 & ~new_new_n38467__;
  assign new_new_n38481__ = ~ys__n17909 & ~ys__n30334;
  assign new_new_n38482__ = ys__n17909 & ys__n30334;
  assign new_new_n38483__ = ~new_new_n38481__ & ~new_new_n38482__;
  assign new_new_n38484__ = new_new_n38480__ & ~new_new_n38483__;
  assign new_new_n38485__ = new_new_n38467__ & new_new_n38483__;
  assign new_new_n38486__ = ys__n17845 & ~new_new_n38485__;
  assign new_new_n38487__ = ~new_new_n38484__ & ~new_new_n38486__;
  assign new_new_n38488__ = ~new_new_n38479__ & ~new_new_n38487__;
  assign new_new_n38489__ = new_new_n38479__ & ~new_new_n38487__;
  assign new_new_n38490__ = ~new_new_n38479__ & new_new_n38487__;
  assign new_new_n38491__ = ~new_new_n38489__ & ~new_new_n38490__;
  assign new_new_n38492__ = ys__n17845 & new_new_n38467__;
  assign new_new_n38493__ = ~new_new_n38480__ & ~new_new_n38492__;
  assign new_new_n38494__ = ~new_new_n38483__ & new_new_n38493__;
  assign new_new_n38495__ = new_new_n38483__ & ~new_new_n38493__;
  assign new_new_n38496__ = ~new_new_n38494__ & ~new_new_n38495__;
  assign new_new_n38497__ = ~ys__n17843 & ~new_new_n38483__;
  assign new_new_n38498__ = ~ys__n17908 & ~ys__n30334;
  assign new_new_n38499__ = ys__n17908 & ys__n30334;
  assign new_new_n38500__ = ~new_new_n38498__ & ~new_new_n38499__;
  assign new_new_n38501__ = new_new_n38497__ & ~new_new_n38500__;
  assign new_new_n38502__ = new_new_n38483__ & new_new_n38500__;
  assign new_new_n38503__ = ys__n17843 & ~new_new_n38502__;
  assign new_new_n38504__ = ~new_new_n38501__ & ~new_new_n38503__;
  assign new_new_n38505__ = ~new_new_n38496__ & ~new_new_n38504__;
  assign new_new_n38506__ = new_new_n38496__ & ~new_new_n38504__;
  assign new_new_n38507__ = ~new_new_n38496__ & new_new_n38504__;
  assign new_new_n38508__ = ~new_new_n38506__ & ~new_new_n38507__;
  assign new_new_n38509__ = ys__n17843 & new_new_n38483__;
  assign new_new_n38510__ = ~new_new_n38497__ & ~new_new_n38509__;
  assign new_new_n38511__ = ~new_new_n38500__ & new_new_n38510__;
  assign new_new_n38512__ = new_new_n38500__ & ~new_new_n38510__;
  assign new_new_n38513__ = ~new_new_n38511__ & ~new_new_n38512__;
  assign new_new_n38514__ = ~ys__n17842 & ~new_new_n38500__;
  assign new_new_n38515__ = ~ys__n17906 & ~ys__n30334;
  assign new_new_n38516__ = ys__n17906 & ys__n30334;
  assign new_new_n38517__ = ~new_new_n38515__ & ~new_new_n38516__;
  assign new_new_n38518__ = new_new_n38514__ & ~new_new_n38517__;
  assign new_new_n38519__ = new_new_n38500__ & new_new_n38517__;
  assign new_new_n38520__ = ys__n17842 & ~new_new_n38519__;
  assign new_new_n38521__ = ~new_new_n38518__ & ~new_new_n38520__;
  assign new_new_n38522__ = ~new_new_n38513__ & ~new_new_n38521__;
  assign new_new_n38523__ = ~new_new_n38508__ & new_new_n38522__;
  assign new_new_n38524__ = ~new_new_n38505__ & ~new_new_n38523__;
  assign new_new_n38525__ = new_new_n38513__ & ~new_new_n38521__;
  assign new_new_n38526__ = ~new_new_n38513__ & new_new_n38521__;
  assign new_new_n38527__ = ~new_new_n38525__ & ~new_new_n38526__;
  assign new_new_n38528__ = ~new_new_n38508__ & ~new_new_n38527__;
  assign new_new_n38529__ = ys__n17842 & new_new_n38500__;
  assign new_new_n38530__ = ~new_new_n38514__ & ~new_new_n38529__;
  assign new_new_n38531__ = ~new_new_n38517__ & new_new_n38530__;
  assign new_new_n38532__ = new_new_n38517__ & ~new_new_n38530__;
  assign new_new_n38533__ = ~new_new_n38531__ & ~new_new_n38532__;
  assign new_new_n38534__ = ~ys__n17840 & ~new_new_n38517__;
  assign new_new_n38535__ = ~ys__n17905 & ~ys__n30334;
  assign new_new_n38536__ = ys__n17905 & ys__n30334;
  assign new_new_n38537__ = ~new_new_n38535__ & ~new_new_n38536__;
  assign new_new_n38538__ = new_new_n38534__ & ~new_new_n38537__;
  assign new_new_n38539__ = new_new_n38517__ & new_new_n38537__;
  assign new_new_n38540__ = ys__n17840 & ~new_new_n38539__;
  assign new_new_n38541__ = ~new_new_n38538__ & ~new_new_n38540__;
  assign new_new_n38542__ = new_new_n38533__ & ~new_new_n38541__;
  assign new_new_n38543__ = ~new_new_n38533__ & new_new_n38541__;
  assign new_new_n38544__ = ~new_new_n38542__ & ~new_new_n38543__;
  assign new_new_n38545__ = ys__n17840 & new_new_n38517__;
  assign new_new_n38546__ = ~new_new_n38534__ & ~new_new_n38545__;
  assign new_new_n38547__ = ~new_new_n38537__ & new_new_n38546__;
  assign new_new_n38548__ = new_new_n38537__ & ~new_new_n38546__;
  assign new_new_n38549__ = ~new_new_n38547__ & ~new_new_n38548__;
  assign new_new_n38550__ = ~ys__n17839 & ~new_new_n38537__;
  assign new_new_n38551__ = ~ys__n17903 & ~ys__n30334;
  assign new_new_n38552__ = ys__n17903 & ys__n30334;
  assign new_new_n38553__ = ~new_new_n38551__ & ~new_new_n38552__;
  assign new_new_n38554__ = new_new_n38550__ & ~new_new_n38553__;
  assign new_new_n38555__ = new_new_n38537__ & new_new_n38553__;
  assign new_new_n38556__ = ys__n17839 & ~new_new_n38555__;
  assign new_new_n38557__ = ~new_new_n38554__ & ~new_new_n38556__;
  assign new_new_n38558__ = new_new_n38549__ & ~new_new_n38557__;
  assign new_new_n38559__ = ~new_new_n38549__ & new_new_n38557__;
  assign new_new_n38560__ = ~new_new_n38558__ & ~new_new_n38559__;
  assign new_new_n38561__ = ~new_new_n38544__ & ~new_new_n38560__;
  assign new_new_n38562__ = ys__n17839 & new_new_n38537__;
  assign new_new_n38563__ = ~new_new_n38550__ & ~new_new_n38562__;
  assign new_new_n38564__ = ~new_new_n38553__ & new_new_n38563__;
  assign new_new_n38565__ = new_new_n38553__ & ~new_new_n38563__;
  assign new_new_n38566__ = ~new_new_n38564__ & ~new_new_n38565__;
  assign new_new_n38567__ = ~ys__n17837 & ~new_new_n38553__;
  assign new_new_n38568__ = ~ys__n17902 & ~ys__n30334;
  assign new_new_n38569__ = ys__n17902 & ys__n30334;
  assign new_new_n38570__ = ~new_new_n38568__ & ~new_new_n38569__;
  assign new_new_n38571__ = new_new_n38567__ & ~new_new_n38570__;
  assign new_new_n38572__ = new_new_n38553__ & new_new_n38570__;
  assign new_new_n38573__ = ys__n17837 & ~new_new_n38572__;
  assign new_new_n38574__ = ~new_new_n38571__ & ~new_new_n38573__;
  assign new_new_n38575__ = ~new_new_n38566__ & ~new_new_n38574__;
  assign new_new_n38576__ = new_new_n38566__ & ~new_new_n38574__;
  assign new_new_n38577__ = ~new_new_n38566__ & new_new_n38574__;
  assign new_new_n38578__ = ~new_new_n38576__ & ~new_new_n38577__;
  assign new_new_n38579__ = ys__n17837 & new_new_n38553__;
  assign new_new_n38580__ = ~new_new_n38567__ & ~new_new_n38579__;
  assign new_new_n38581__ = ~new_new_n38570__ & new_new_n38580__;
  assign new_new_n38582__ = new_new_n38570__ & ~new_new_n38580__;
  assign new_new_n38583__ = ~new_new_n38581__ & ~new_new_n38582__;
  assign new_new_n38584__ = ~ys__n17836 & ~new_new_n38570__;
  assign new_new_n38585__ = ~ys__n17900 & ~ys__n30334;
  assign new_new_n38586__ = ys__n17900 & ys__n30334;
  assign new_new_n38587__ = ~new_new_n38585__ & ~new_new_n38586__;
  assign new_new_n38588__ = new_new_n38584__ & ~new_new_n38587__;
  assign new_new_n38589__ = new_new_n38570__ & new_new_n38587__;
  assign new_new_n38590__ = ys__n17836 & ~new_new_n38589__;
  assign new_new_n38591__ = ~new_new_n38588__ & ~new_new_n38590__;
  assign new_new_n38592__ = ~new_new_n38583__ & ~new_new_n38591__;
  assign new_new_n38593__ = ~new_new_n38578__ & new_new_n38592__;
  assign new_new_n38594__ = ~new_new_n38575__ & ~new_new_n38593__;
  assign new_new_n38595__ = new_new_n38561__ & ~new_new_n38594__;
  assign new_new_n38596__ = ~new_new_n38533__ & ~new_new_n38541__;
  assign new_new_n38597__ = ~new_new_n38549__ & ~new_new_n38557__;
  assign new_new_n38598__ = ~new_new_n38544__ & new_new_n38597__;
  assign new_new_n38599__ = ~new_new_n38596__ & ~new_new_n38598__;
  assign new_new_n38600__ = ~new_new_n38595__ & new_new_n38599__;
  assign new_new_n38601__ = new_new_n38583__ & ~new_new_n38591__;
  assign new_new_n38602__ = ~new_new_n38583__ & new_new_n38591__;
  assign new_new_n38603__ = ~new_new_n38601__ & ~new_new_n38602__;
  assign new_new_n38604__ = ~new_new_n38578__ & ~new_new_n38603__;
  assign new_new_n38605__ = new_new_n38561__ & new_new_n38604__;
  assign new_new_n38606__ = ~ys__n17891 & ~ys__n30334;
  assign new_new_n38607__ = ys__n17891 & ys__n30334;
  assign new_new_n38608__ = ~new_new_n38606__ & ~new_new_n38607__;
  assign new_new_n38609__ = ~ys__n17893 & ~ys__n30334;
  assign new_new_n38610__ = ys__n17893 & ys__n30334;
  assign new_new_n38611__ = ~new_new_n38609__ & ~new_new_n38610__;
  assign new_new_n38612__ = ~ys__n17827 & ~new_new_n38611__;
  assign new_new_n38613__ = ys__n17827 & new_new_n38611__;
  assign new_new_n38614__ = ~new_new_n38612__ & ~new_new_n38613__;
  assign new_new_n38615__ = ~new_new_n38608__ & new_new_n38614__;
  assign new_new_n38616__ = new_new_n38608__ & ~new_new_n38614__;
  assign new_new_n38617__ = ~new_new_n38615__ & ~new_new_n38616__;
  assign new_new_n38618__ = ~ys__n17825 & ~new_new_n38608__;
  assign new_new_n38619__ = ~new_new_n38209__ & new_new_n38618__;
  assign new_new_n38620__ = new_new_n38209__ & new_new_n38608__;
  assign new_new_n38621__ = ys__n17825 & ~new_new_n38620__;
  assign new_new_n38622__ = ~new_new_n38619__ & ~new_new_n38621__;
  assign new_new_n38623__ = ~new_new_n38617__ & ~new_new_n38622__;
  assign new_new_n38624__ = new_new_n38617__ & ~new_new_n38622__;
  assign new_new_n38625__ = ~new_new_n38617__ & new_new_n38622__;
  assign new_new_n38626__ = ~new_new_n38624__ & ~new_new_n38625__;
  assign new_new_n38627__ = ys__n17825 & new_new_n38608__;
  assign new_new_n38628__ = ~new_new_n38618__ & ~new_new_n38627__;
  assign new_new_n38629__ = ~new_new_n38209__ & new_new_n38628__;
  assign new_new_n38630__ = new_new_n38209__ & ~new_new_n38628__;
  assign new_new_n38631__ = ~new_new_n38629__ & ~new_new_n38630__;
  assign new_new_n38632__ = ~new_new_n38206__ & new_new_n38210__;
  assign new_new_n38633__ = new_new_n38206__ & new_new_n38209__;
  assign new_new_n38634__ = ys__n17824 & ~new_new_n38633__;
  assign new_new_n38635__ = ~new_new_n38632__ & ~new_new_n38634__;
  assign new_new_n38636__ = ~new_new_n38631__ & ~new_new_n38635__;
  assign new_new_n38637__ = ~new_new_n38626__ & new_new_n38636__;
  assign new_new_n38638__ = ~new_new_n38623__ & ~new_new_n38637__;
  assign new_new_n38639__ = ~ys__n17894 & ~ys__n30334;
  assign new_new_n38640__ = ys__n17894 & ys__n30334;
  assign new_new_n38641__ = ~new_new_n38639__ & ~new_new_n38640__;
  assign new_new_n38642__ = ~ys__n17896 & ~ys__n30334;
  assign new_new_n38643__ = ys__n17896 & ys__n30334;
  assign new_new_n38644__ = ~new_new_n38642__ & ~new_new_n38643__;
  assign new_new_n38645__ = ~ys__n17830 & ~new_new_n38644__;
  assign new_new_n38646__ = ys__n17830 & new_new_n38644__;
  assign new_new_n38647__ = ~new_new_n38645__ & ~new_new_n38646__;
  assign new_new_n38648__ = ~new_new_n38641__ & new_new_n38647__;
  assign new_new_n38649__ = new_new_n38641__ & ~new_new_n38647__;
  assign new_new_n38650__ = ~new_new_n38648__ & ~new_new_n38649__;
  assign new_new_n38651__ = ~ys__n17828 & ~new_new_n38641__;
  assign new_new_n38652__ = ~new_new_n38611__ & new_new_n38651__;
  assign new_new_n38653__ = new_new_n38611__ & new_new_n38641__;
  assign new_new_n38654__ = ys__n17828 & ~new_new_n38653__;
  assign new_new_n38655__ = ~new_new_n38652__ & ~new_new_n38654__;
  assign new_new_n38656__ = new_new_n38650__ & ~new_new_n38655__;
  assign new_new_n38657__ = ~new_new_n38650__ & new_new_n38655__;
  assign new_new_n38658__ = ~new_new_n38656__ & ~new_new_n38657__;
  assign new_new_n38659__ = ys__n17828 & new_new_n38641__;
  assign new_new_n38660__ = ~new_new_n38651__ & ~new_new_n38659__;
  assign new_new_n38661__ = ~new_new_n38611__ & new_new_n38660__;
  assign new_new_n38662__ = new_new_n38611__ & ~new_new_n38660__;
  assign new_new_n38663__ = ~new_new_n38661__ & ~new_new_n38662__;
  assign new_new_n38664__ = ~new_new_n38608__ & new_new_n38612__;
  assign new_new_n38665__ = new_new_n38608__ & new_new_n38611__;
  assign new_new_n38666__ = ys__n17827 & ~new_new_n38665__;
  assign new_new_n38667__ = ~new_new_n38664__ & ~new_new_n38666__;
  assign new_new_n38668__ = new_new_n38663__ & ~new_new_n38667__;
  assign new_new_n38669__ = ~new_new_n38663__ & new_new_n38667__;
  assign new_new_n38670__ = ~new_new_n38668__ & ~new_new_n38669__;
  assign new_new_n38671__ = ~new_new_n38658__ & ~new_new_n38670__;
  assign new_new_n38672__ = ~new_new_n38638__ & new_new_n38671__;
  assign new_new_n38673__ = ~new_new_n38650__ & ~new_new_n38655__;
  assign new_new_n38674__ = ~new_new_n38663__ & ~new_new_n38667__;
  assign new_new_n38675__ = ~new_new_n38658__ & new_new_n38674__;
  assign new_new_n38676__ = ~new_new_n38673__ & ~new_new_n38675__;
  assign new_new_n38677__ = ~new_new_n38672__ & new_new_n38676__;
  assign new_new_n38678__ = ys__n17836 & new_new_n38570__;
  assign new_new_n38679__ = ~new_new_n38584__ & ~new_new_n38678__;
  assign new_new_n38680__ = ~new_new_n38587__ & new_new_n38679__;
  assign new_new_n38681__ = new_new_n38587__ & ~new_new_n38679__;
  assign new_new_n38682__ = ~new_new_n38680__ & ~new_new_n38681__;
  assign new_new_n38683__ = ~ys__n17834 & ~new_new_n38587__;
  assign new_new_n38684__ = ~ys__n17899 & ~ys__n30334;
  assign new_new_n38685__ = ys__n17899 & ys__n30334;
  assign new_new_n38686__ = ~new_new_n38684__ & ~new_new_n38685__;
  assign new_new_n38687__ = new_new_n38683__ & ~new_new_n38686__;
  assign new_new_n38688__ = new_new_n38587__ & new_new_n38686__;
  assign new_new_n38689__ = ys__n17834 & ~new_new_n38688__;
  assign new_new_n38690__ = ~new_new_n38687__ & ~new_new_n38689__;
  assign new_new_n38691__ = new_new_n38682__ & ~new_new_n38690__;
  assign new_new_n38692__ = ~new_new_n38682__ & new_new_n38690__;
  assign new_new_n38693__ = ~new_new_n38691__ & ~new_new_n38692__;
  assign new_new_n38694__ = ys__n17834 & new_new_n38587__;
  assign new_new_n38695__ = ~new_new_n38683__ & ~new_new_n38694__;
  assign new_new_n38696__ = ~new_new_n38686__ & new_new_n38695__;
  assign new_new_n38697__ = new_new_n38686__ & ~new_new_n38695__;
  assign new_new_n38698__ = ~new_new_n38696__ & ~new_new_n38697__;
  assign new_new_n38699__ = ~ys__n17833 & ~new_new_n38686__;
  assign new_new_n38700__ = ~ys__n17897 & ~ys__n30334;
  assign new_new_n38701__ = ys__n17897 & ys__n30334;
  assign new_new_n38702__ = ~new_new_n38700__ & ~new_new_n38701__;
  assign new_new_n38703__ = new_new_n38699__ & ~new_new_n38702__;
  assign new_new_n38704__ = new_new_n38686__ & new_new_n38702__;
  assign new_new_n38705__ = ys__n17833 & ~new_new_n38704__;
  assign new_new_n38706__ = ~new_new_n38703__ & ~new_new_n38705__;
  assign new_new_n38707__ = new_new_n38698__ & ~new_new_n38706__;
  assign new_new_n38708__ = ~new_new_n38698__ & new_new_n38706__;
  assign new_new_n38709__ = ~new_new_n38707__ & ~new_new_n38708__;
  assign new_new_n38710__ = ~new_new_n38693__ & ~new_new_n38709__;
  assign new_new_n38711__ = ys__n17833 & new_new_n38686__;
  assign new_new_n38712__ = ~new_new_n38699__ & ~new_new_n38711__;
  assign new_new_n38713__ = ~new_new_n38702__ & new_new_n38712__;
  assign new_new_n38714__ = new_new_n38702__ & ~new_new_n38712__;
  assign new_new_n38715__ = ~new_new_n38713__ & ~new_new_n38714__;
  assign new_new_n38716__ = ~ys__n17831 & ~new_new_n38702__;
  assign new_new_n38717__ = ~new_new_n38644__ & new_new_n38716__;
  assign new_new_n38718__ = new_new_n38644__ & new_new_n38702__;
  assign new_new_n38719__ = ys__n17831 & ~new_new_n38718__;
  assign new_new_n38720__ = ~new_new_n38717__ & ~new_new_n38719__;
  assign new_new_n38721__ = new_new_n38715__ & ~new_new_n38720__;
  assign new_new_n38722__ = ~new_new_n38715__ & new_new_n38720__;
  assign new_new_n38723__ = ~new_new_n38721__ & ~new_new_n38722__;
  assign new_new_n38724__ = ys__n17831 & new_new_n38702__;
  assign new_new_n38725__ = ~new_new_n38716__ & ~new_new_n38724__;
  assign new_new_n38726__ = ~new_new_n38644__ & new_new_n38725__;
  assign new_new_n38727__ = new_new_n38644__ & ~new_new_n38725__;
  assign new_new_n38728__ = ~new_new_n38726__ & ~new_new_n38727__;
  assign new_new_n38729__ = ~new_new_n38641__ & new_new_n38645__;
  assign new_new_n38730__ = new_new_n38641__ & new_new_n38644__;
  assign new_new_n38731__ = ys__n17830 & ~new_new_n38730__;
  assign new_new_n38732__ = ~new_new_n38729__ & ~new_new_n38731__;
  assign new_new_n38733__ = new_new_n38728__ & ~new_new_n38732__;
  assign new_new_n38734__ = ~new_new_n38728__ & new_new_n38732__;
  assign new_new_n38735__ = ~new_new_n38733__ & ~new_new_n38734__;
  assign new_new_n38736__ = ~new_new_n38723__ & ~new_new_n38735__;
  assign new_new_n38737__ = new_new_n38710__ & new_new_n38736__;
  assign new_new_n38738__ = ~new_new_n38677__ & new_new_n38737__;
  assign new_new_n38739__ = ~new_new_n38715__ & ~new_new_n38720__;
  assign new_new_n38740__ = ~new_new_n38728__ & ~new_new_n38732__;
  assign new_new_n38741__ = ~new_new_n38723__ & new_new_n38740__;
  assign new_new_n38742__ = ~new_new_n38739__ & ~new_new_n38741__;
  assign new_new_n38743__ = new_new_n38710__ & ~new_new_n38742__;
  assign new_new_n38744__ = ~new_new_n38682__ & ~new_new_n38690__;
  assign new_new_n38745__ = ~new_new_n38698__ & ~new_new_n38706__;
  assign new_new_n38746__ = ~new_new_n38693__ & new_new_n38745__;
  assign new_new_n38747__ = ~new_new_n38744__ & ~new_new_n38746__;
  assign new_new_n38748__ = ~new_new_n38743__ & new_new_n38747__;
  assign new_new_n38749__ = ~new_new_n38738__ & new_new_n38748__;
  assign new_new_n38750__ = new_new_n38605__ & ~new_new_n38749__;
  assign new_new_n38751__ = new_new_n38600__ & ~new_new_n38750__;
  assign new_new_n38752__ = new_new_n38528__ & ~new_new_n38751__;
  assign new_new_n38753__ = new_new_n38524__ & ~new_new_n38752__;
  assign new_new_n38754__ = ~new_new_n38491__ & ~new_new_n38753__;
  assign new_new_n38755__ = ~new_new_n38488__ & ~new_new_n38754__;
  assign new_new_n38756__ = new_new_n38474__ & ~new_new_n38755__;
  assign new_new_n38757__ = ~new_new_n38474__ & new_new_n38755__;
  assign new_new_n38758__ = ~new_new_n38756__ & ~new_new_n38757__;
  assign new_new_n38759__ = new_new_n38451__ & ~new_new_n38758__;
  assign new_new_n38760__ = new_new_n38491__ & ~new_new_n38753__;
  assign new_new_n38761__ = ~new_new_n38491__ & new_new_n38753__;
  assign new_new_n38762__ = ~new_new_n38760__ & ~new_new_n38761__;
  assign new_new_n38763__ = ~new_new_n38527__ & ~new_new_n38751__;
  assign new_new_n38764__ = ~new_new_n38522__ & ~new_new_n38763__;
  assign new_new_n38765__ = new_new_n38508__ & ~new_new_n38764__;
  assign new_new_n38766__ = ~new_new_n38508__ & new_new_n38764__;
  assign new_new_n38767__ = ~new_new_n38765__ & ~new_new_n38766__;
  assign new_new_n38768__ = new_new_n38527__ & ~new_new_n38751__;
  assign new_new_n38769__ = ~new_new_n38527__ & new_new_n38751__;
  assign new_new_n38770__ = ~new_new_n38768__ & ~new_new_n38769__;
  assign new_new_n38771__ = ~new_new_n38767__ & ~new_new_n38770__;
  assign new_new_n38772__ = new_new_n38604__ & ~new_new_n38749__;
  assign new_new_n38773__ = new_new_n38594__ & ~new_new_n38772__;
  assign new_new_n38774__ = ~new_new_n38560__ & ~new_new_n38773__;
  assign new_new_n38775__ = ~new_new_n38597__ & ~new_new_n38774__;
  assign new_new_n38776__ = new_new_n38544__ & ~new_new_n38775__;
  assign new_new_n38777__ = ~new_new_n38544__ & new_new_n38775__;
  assign new_new_n38778__ = ~new_new_n38776__ & ~new_new_n38777__;
  assign new_new_n38779__ = new_new_n38560__ & ~new_new_n38773__;
  assign new_new_n38780__ = ~new_new_n38560__ & new_new_n38773__;
  assign new_new_n38781__ = ~new_new_n38779__ & ~new_new_n38780__;
  assign new_new_n38782__ = ~new_new_n38603__ & ~new_new_n38749__;
  assign new_new_n38783__ = ~new_new_n38592__ & ~new_new_n38782__;
  assign new_new_n38784__ = new_new_n38578__ & ~new_new_n38783__;
  assign new_new_n38785__ = ~new_new_n38578__ & new_new_n38783__;
  assign new_new_n38786__ = ~new_new_n38784__ & ~new_new_n38785__;
  assign new_new_n38787__ = new_new_n38603__ & ~new_new_n38749__;
  assign new_new_n38788__ = ~new_new_n38603__ & new_new_n38749__;
  assign new_new_n38789__ = ~new_new_n38787__ & ~new_new_n38788__;
  assign new_new_n38790__ = ~new_new_n38786__ & ~new_new_n38789__;
  assign new_new_n38791__ = ~new_new_n38781__ & new_new_n38790__;
  assign new_new_n38792__ = ~new_new_n38778__ & new_new_n38791__;
  assign new_new_n38793__ = ~new_new_n38677__ & new_new_n38736__;
  assign new_new_n38794__ = new_new_n38742__ & ~new_new_n38793__;
  assign new_new_n38795__ = ~new_new_n38709__ & ~new_new_n38794__;
  assign new_new_n38796__ = ~new_new_n38745__ & ~new_new_n38795__;
  assign new_new_n38797__ = new_new_n38693__ & ~new_new_n38796__;
  assign new_new_n38798__ = ~new_new_n38693__ & new_new_n38796__;
  assign new_new_n38799__ = ~new_new_n38797__ & ~new_new_n38798__;
  assign new_new_n38800__ = ~new_new_n38677__ & ~new_new_n38735__;
  assign new_new_n38801__ = ~new_new_n38740__ & ~new_new_n38800__;
  assign new_new_n38802__ = new_new_n38723__ & ~new_new_n38801__;
  assign new_new_n38803__ = ~new_new_n38723__ & new_new_n38801__;
  assign new_new_n38804__ = ~new_new_n38802__ & ~new_new_n38803__;
  assign new_new_n38805__ = ~new_new_n38677__ & new_new_n38735__;
  assign new_new_n38806__ = new_new_n38677__ & ~new_new_n38735__;
  assign new_new_n38807__ = ~new_new_n38805__ & ~new_new_n38806__;
  assign new_new_n38808__ = ~new_new_n38804__ & ~new_new_n38807__;
  assign new_new_n38809__ = new_new_n38709__ & ~new_new_n38794__;
  assign new_new_n38810__ = ~new_new_n38709__ & new_new_n38794__;
  assign new_new_n38811__ = ~new_new_n38809__ & ~new_new_n38810__;
  assign new_new_n38812__ = ~new_new_n38638__ & ~new_new_n38670__;
  assign new_new_n38813__ = ~new_new_n38674__ & ~new_new_n38812__;
  assign new_new_n38814__ = new_new_n38658__ & ~new_new_n38813__;
  assign new_new_n38815__ = ~new_new_n38658__ & new_new_n38813__;
  assign new_new_n38816__ = ~new_new_n38814__ & ~new_new_n38815__;
  assign new_new_n38817__ = ~new_new_n38638__ & new_new_n38670__;
  assign new_new_n38818__ = new_new_n38638__ & ~new_new_n38670__;
  assign new_new_n38819__ = ~new_new_n38817__ & ~new_new_n38818__;
  assign new_new_n38820__ = new_new_n38626__ & new_new_n38636__;
  assign new_new_n38821__ = ~new_new_n38626__ & ~new_new_n38636__;
  assign new_new_n38822__ = ~new_new_n38820__ & ~new_new_n38821__;
  assign new_new_n38823__ = new_new_n38631__ & ~new_new_n38635__;
  assign new_new_n38824__ = ~new_new_n38631__ & new_new_n38635__;
  assign new_new_n38825__ = ~new_new_n38823__ & ~new_new_n38824__;
  assign new_new_n38826__ = ~new_new_n38822__ & ~new_new_n38825__;
  assign new_new_n38827__ = ~new_new_n38819__ & new_new_n38826__;
  assign new_new_n38828__ = ~new_new_n38816__ & new_new_n38827__;
  assign new_new_n38829__ = ~new_new_n38811__ & new_new_n38828__;
  assign new_new_n38830__ = new_new_n38808__ & new_new_n38829__;
  assign new_new_n38831__ = ~new_new_n38799__ & new_new_n38830__;
  assign new_new_n38832__ = new_new_n38792__ & new_new_n38831__;
  assign new_new_n38833__ = new_new_n38771__ & new_new_n38832__;
  assign new_new_n38834__ = ~new_new_n38762__ & new_new_n38833__;
  assign new_new_n38835__ = new_new_n38758__ & new_new_n38834__;
  assign new_new_n38836__ = ~new_new_n38758__ & ~new_new_n38834__;
  assign new_new_n38837__ = ~new_new_n38835__ & ~new_new_n38836__;
  assign new_new_n38838__ = ~new_new_n38451__ & ~new_new_n38837__;
  assign new_new_n38839__ = ~new_new_n38759__ & ~new_new_n38838__;
  assign new_new_n38840__ = ys__n18156 & ~new_new_n38839__;
  assign new_new_n38841__ = ~ys__n17849 & ~new_new_n38457__;
  assign new_new_n38842__ = ys__n17849 & new_new_n38457__;
  assign new_new_n38843__ = ~new_new_n38841__ & ~new_new_n38842__;
  assign new_new_n38844__ = ~new_new_n38457__ & new_new_n38843__;
  assign new_new_n38845__ = new_new_n38457__ & ~new_new_n38843__;
  assign new_new_n38846__ = ~new_new_n38844__ & ~new_new_n38845__;
  assign new_new_n38847__ = ~new_new_n38454__ & new_new_n38458__;
  assign new_new_n38848__ = new_new_n38454__ & new_new_n38457__;
  assign new_new_n38849__ = ys__n17848 & ~new_new_n38848__;
  assign new_new_n38850__ = ~new_new_n38847__ & ~new_new_n38849__;
  assign new_new_n38851__ = new_new_n38846__ & ~new_new_n38850__;
  assign new_new_n38852__ = ~new_new_n38846__ & new_new_n38850__;
  assign new_new_n38853__ = ~new_new_n38851__ & ~new_new_n38852__;
  assign new_new_n38854__ = ~new_new_n38474__ & ~new_new_n38491__;
  assign new_new_n38855__ = new_new_n38528__ & new_new_n38854__;
  assign new_new_n38856__ = new_new_n38605__ & new_new_n38855__;
  assign new_new_n38857__ = ~new_new_n38749__ & new_new_n38856__;
  assign new_new_n38858__ = ~new_new_n38600__ & new_new_n38855__;
  assign new_new_n38859__ = ~new_new_n38524__ & new_new_n38854__;
  assign new_new_n38860__ = ~new_new_n38463__ & ~new_new_n38471__;
  assign new_new_n38861__ = ~new_new_n38474__ & new_new_n38488__;
  assign new_new_n38862__ = ~new_new_n38860__ & ~new_new_n38861__;
  assign new_new_n38863__ = ~new_new_n38859__ & new_new_n38862__;
  assign new_new_n38864__ = ~new_new_n38858__ & new_new_n38863__;
  assign new_new_n38865__ = ~new_new_n38857__ & new_new_n38864__;
  assign new_new_n38866__ = new_new_n38853__ & ~new_new_n38865__;
  assign new_new_n38867__ = ~new_new_n38853__ & new_new_n38865__;
  assign new_new_n38868__ = ~new_new_n38866__ & ~new_new_n38867__;
  assign new_new_n38869__ = new_new_n38451__ & ~new_new_n38868__;
  assign new_new_n38870__ = ~new_new_n38762__ & new_new_n38831__;
  assign new_new_n38871__ = new_new_n38771__ & new_new_n38870__;
  assign new_new_n38872__ = new_new_n38792__ & new_new_n38871__;
  assign new_new_n38873__ = ~new_new_n38758__ & new_new_n38872__;
  assign new_new_n38874__ = new_new_n38868__ & new_new_n38873__;
  assign new_new_n38875__ = ~new_new_n38868__ & ~new_new_n38873__;
  assign new_new_n38876__ = ~new_new_n38874__ & ~new_new_n38875__;
  assign new_new_n38877__ = ~new_new_n38451__ & ~new_new_n38876__;
  assign new_new_n38878__ = ~new_new_n38869__ & ~new_new_n38877__;
  assign new_new_n38879__ = ~new_new_n38840__ & new_new_n38878__;
  assign new_new_n38880__ = ys__n33581 & ~new_new_n38064__;
  assign new_new_n38881__ = ~ys__n33581 & ~new_new_n38064__;
  assign new_new_n38882__ = ys__n33581 & new_new_n38064__;
  assign new_new_n38883__ = ~new_new_n38881__ & ~new_new_n38882__;
  assign new_new_n38884__ = ~ys__n30334 & ys__n33579;
  assign new_new_n38885__ = ~new_new_n38883__ & new_new_n38884__;
  assign new_new_n38886__ = ~new_new_n38880__ & ~new_new_n38885__;
  assign new_new_n38887__ = ~ys__n17804 & ~new_new_n38054__;
  assign new_new_n38888__ = ys__n17804 & new_new_n38054__;
  assign new_new_n38889__ = ~new_new_n38887__ & ~new_new_n38888__;
  assign new_new_n38890__ = ~ys__n17803 & ~new_new_n38051__;
  assign new_new_n38891__ = ys__n17803 & new_new_n38051__;
  assign new_new_n38892__ = ~new_new_n38890__ & ~new_new_n38891__;
  assign new_new_n38893__ = ~new_new_n38889__ & ~new_new_n38892__;
  assign new_new_n38894__ = ~new_new_n38886__ & new_new_n38893__;
  assign new_new_n38895__ = ys__n17804 & ~new_new_n38054__;
  assign new_new_n38896__ = ys__n17803 & ~new_new_n38051__;
  assign new_new_n38897__ = ~new_new_n38889__ & new_new_n38896__;
  assign new_new_n38898__ = ~new_new_n38895__ & ~new_new_n38897__;
  assign new_new_n38899__ = ~new_new_n38894__ & new_new_n38898__;
  assign new_new_n38900__ = ~ys__n17810 & ~new_new_n38140__;
  assign new_new_n38901__ = ys__n17810 & new_new_n38140__;
  assign new_new_n38902__ = ~new_new_n38900__ & ~new_new_n38901__;
  assign new_new_n38903__ = ~ys__n17809 & ~new_new_n38156__;
  assign new_new_n38904__ = ys__n17809 & new_new_n38156__;
  assign new_new_n38905__ = ~new_new_n38903__ & ~new_new_n38904__;
  assign new_new_n38906__ = ~new_new_n38902__ & ~new_new_n38905__;
  assign new_new_n38907__ = ~ys__n17807 & ~new_new_n38091__;
  assign new_new_n38908__ = ys__n17807 & new_new_n38091__;
  assign new_new_n38909__ = ~new_new_n38907__ & ~new_new_n38908__;
  assign new_new_n38910__ = ~ys__n17806 & ~new_new_n38088__;
  assign new_new_n38911__ = ys__n17806 & new_new_n38088__;
  assign new_new_n38912__ = ~new_new_n38910__ & ~new_new_n38911__;
  assign new_new_n38913__ = ~new_new_n38909__ & ~new_new_n38912__;
  assign new_new_n38914__ = new_new_n38906__ & new_new_n38913__;
  assign new_new_n38915__ = ~new_new_n38899__ & new_new_n38914__;
  assign new_new_n38916__ = ys__n17807 & ~new_new_n38091__;
  assign new_new_n38917__ = ys__n17806 & ~new_new_n38088__;
  assign new_new_n38918__ = ~new_new_n38909__ & new_new_n38917__;
  assign new_new_n38919__ = ~new_new_n38916__ & ~new_new_n38918__;
  assign new_new_n38920__ = new_new_n38906__ & ~new_new_n38919__;
  assign new_new_n38921__ = ys__n17810 & ~new_new_n38140__;
  assign new_new_n38922__ = ys__n17809 & ~new_new_n38156__;
  assign new_new_n38923__ = ~new_new_n38902__ & new_new_n38922__;
  assign new_new_n38924__ = ~new_new_n38921__ & ~new_new_n38923__;
  assign new_new_n38925__ = ~new_new_n38920__ & new_new_n38924__;
  assign new_new_n38926__ = ~new_new_n38915__ & new_new_n38925__;
  assign new_new_n38927__ = ~ys__n17822 & ~new_new_n38219__;
  assign new_new_n38928__ = ys__n17822 & new_new_n38219__;
  assign new_new_n38929__ = ~new_new_n38927__ & ~new_new_n38928__;
  assign new_new_n38930__ = ~ys__n17821 & ~new_new_n38235__;
  assign new_new_n38931__ = ys__n17821 & new_new_n38235__;
  assign new_new_n38932__ = ~new_new_n38930__ & ~new_new_n38931__;
  assign new_new_n38933__ = ~new_new_n38929__ & ~new_new_n38932__;
  assign new_new_n38934__ = ~ys__n17819 & ~new_new_n38252__;
  assign new_new_n38935__ = ys__n17819 & new_new_n38252__;
  assign new_new_n38936__ = ~new_new_n38934__ & ~new_new_n38935__;
  assign new_new_n38937__ = ~ys__n17818 & ~new_new_n38268__;
  assign new_new_n38938__ = ys__n17818 & new_new_n38268__;
  assign new_new_n38939__ = ~new_new_n38937__ & ~new_new_n38938__;
  assign new_new_n38940__ = ~new_new_n38936__ & ~new_new_n38939__;
  assign new_new_n38941__ = new_new_n38933__ & new_new_n38940__;
  assign new_new_n38942__ = ~ys__n17816 & ~new_new_n38286__;
  assign new_new_n38943__ = ys__n17816 & new_new_n38286__;
  assign new_new_n38944__ = ~new_new_n38942__ & ~new_new_n38943__;
  assign new_new_n38945__ = ~ys__n17815 & ~new_new_n38302__;
  assign new_new_n38946__ = ys__n17815 & new_new_n38302__;
  assign new_new_n38947__ = ~new_new_n38945__ & ~new_new_n38946__;
  assign new_new_n38948__ = ~new_new_n38944__ & ~new_new_n38947__;
  assign new_new_n38949__ = ~ys__n17813 & ~new_new_n38130__;
  assign new_new_n38950__ = ys__n17813 & new_new_n38130__;
  assign new_new_n38951__ = ~new_new_n38949__ & ~new_new_n38950__;
  assign new_new_n38952__ = ~ys__n17812 & ~new_new_n38127__;
  assign new_new_n38953__ = ys__n17812 & new_new_n38127__;
  assign new_new_n38954__ = ~new_new_n38952__ & ~new_new_n38953__;
  assign new_new_n38955__ = ~new_new_n38951__ & ~new_new_n38954__;
  assign new_new_n38956__ = new_new_n38948__ & new_new_n38955__;
  assign new_new_n38957__ = new_new_n38941__ & new_new_n38956__;
  assign new_new_n38958__ = ~new_new_n38926__ & new_new_n38957__;
  assign new_new_n38959__ = ys__n17813 & ~new_new_n38130__;
  assign new_new_n38960__ = ys__n17812 & ~new_new_n38127__;
  assign new_new_n38961__ = ~new_new_n38951__ & new_new_n38960__;
  assign new_new_n38962__ = ~new_new_n38959__ & ~new_new_n38961__;
  assign new_new_n38963__ = new_new_n38948__ & ~new_new_n38962__;
  assign new_new_n38964__ = ys__n17816 & ~new_new_n38286__;
  assign new_new_n38965__ = ys__n17815 & ~new_new_n38302__;
  assign new_new_n38966__ = ~new_new_n38944__ & new_new_n38965__;
  assign new_new_n38967__ = ~new_new_n38964__ & ~new_new_n38966__;
  assign new_new_n38968__ = ~new_new_n38963__ & new_new_n38967__;
  assign new_new_n38969__ = new_new_n38941__ & ~new_new_n38968__;
  assign new_new_n38970__ = ys__n17819 & ~new_new_n38252__;
  assign new_new_n38971__ = ys__n17818 & ~new_new_n38268__;
  assign new_new_n38972__ = ~new_new_n38936__ & new_new_n38971__;
  assign new_new_n38973__ = ~new_new_n38970__ & ~new_new_n38972__;
  assign new_new_n38974__ = new_new_n38933__ & ~new_new_n38973__;
  assign new_new_n38975__ = ys__n17822 & ~new_new_n38219__;
  assign new_new_n38976__ = ys__n17821 & ~new_new_n38235__;
  assign new_new_n38977__ = ~new_new_n38929__ & new_new_n38976__;
  assign new_new_n38978__ = ~new_new_n38975__ & ~new_new_n38977__;
  assign new_new_n38979__ = ~new_new_n38974__ & new_new_n38978__;
  assign new_new_n38980__ = ~new_new_n38969__ & new_new_n38979__;
  assign new_new_n38981__ = ~new_new_n38958__ & new_new_n38980__;
  assign new_new_n38982__ = ~new_new_n38926__ & new_new_n38956__;
  assign new_new_n38983__ = new_new_n38968__ & ~new_new_n38982__;
  assign new_new_n38984__ = new_new_n38940__ & ~new_new_n38983__;
  assign new_new_n38985__ = new_new_n38973__ & ~new_new_n38984__;
  assign new_new_n38986__ = ~new_new_n38932__ & ~new_new_n38985__;
  assign new_new_n38987__ = ~new_new_n38976__ & ~new_new_n38986__;
  assign new_new_n38988__ = new_new_n38929__ & ~new_new_n38987__;
  assign new_new_n38989__ = ~new_new_n38929__ & new_new_n38987__;
  assign new_new_n38990__ = ~new_new_n38988__ & ~new_new_n38989__;
  assign new_new_n38991__ = ~new_new_n38926__ & new_new_n38955__;
  assign new_new_n38992__ = new_new_n38962__ & ~new_new_n38991__;
  assign new_new_n38993__ = ~new_new_n38947__ & ~new_new_n38992__;
  assign new_new_n38994__ = ~new_new_n38965__ & ~new_new_n38993__;
  assign new_new_n38995__ = new_new_n38944__ & ~new_new_n38994__;
  assign new_new_n38996__ = ~new_new_n38944__ & new_new_n38994__;
  assign new_new_n38997__ = ~new_new_n38995__ & ~new_new_n38996__;
  assign new_new_n38998__ = new_new_n38947__ & ~new_new_n38992__;
  assign new_new_n38999__ = ~new_new_n38947__ & new_new_n38992__;
  assign new_new_n39000__ = ~new_new_n38998__ & ~new_new_n38999__;
  assign new_new_n39001__ = ~new_new_n38926__ & ~new_new_n38954__;
  assign new_new_n39002__ = ~new_new_n38960__ & ~new_new_n39001__;
  assign new_new_n39003__ = new_new_n38951__ & ~new_new_n39002__;
  assign new_new_n39004__ = ~new_new_n38951__ & new_new_n39002__;
  assign new_new_n39005__ = ~new_new_n39003__ & ~new_new_n39004__;
  assign new_new_n39006__ = ~new_new_n38926__ & new_new_n38954__;
  assign new_new_n39007__ = new_new_n38926__ & ~new_new_n38954__;
  assign new_new_n39008__ = ~new_new_n39006__ & ~new_new_n39007__;
  assign new_new_n39009__ = ~new_new_n39005__ & ~new_new_n39008__;
  assign new_new_n39010__ = ~new_new_n39000__ & new_new_n39009__;
  assign new_new_n39011__ = ~new_new_n38997__ & new_new_n39010__;
  assign new_new_n39012__ = ~new_new_n38939__ & ~new_new_n38983__;
  assign new_new_n39013__ = ~new_new_n38971__ & ~new_new_n39012__;
  assign new_new_n39014__ = new_new_n38936__ & ~new_new_n39013__;
  assign new_new_n39015__ = ~new_new_n38936__ & new_new_n39013__;
  assign new_new_n39016__ = ~new_new_n39014__ & ~new_new_n39015__;
  assign new_new_n39017__ = new_new_n38939__ & ~new_new_n38983__;
  assign new_new_n39018__ = ~new_new_n38939__ & new_new_n38983__;
  assign new_new_n39019__ = ~new_new_n39017__ & ~new_new_n39018__;
  assign new_new_n39020__ = ~new_new_n39016__ & ~new_new_n39019__;
  assign new_new_n39021__ = new_new_n38932__ & ~new_new_n38985__;
  assign new_new_n39022__ = ~new_new_n38932__ & new_new_n38985__;
  assign new_new_n39023__ = ~new_new_n39021__ & ~new_new_n39022__;
  assign new_new_n39024__ = ~new_new_n38899__ & new_new_n38913__;
  assign new_new_n39025__ = new_new_n38919__ & ~new_new_n39024__;
  assign new_new_n39026__ = ~new_new_n38905__ & ~new_new_n39025__;
  assign new_new_n39027__ = ~new_new_n38922__ & ~new_new_n39026__;
  assign new_new_n39028__ = new_new_n38902__ & ~new_new_n39027__;
  assign new_new_n39029__ = ~new_new_n38902__ & new_new_n39027__;
  assign new_new_n39030__ = ~new_new_n39028__ & ~new_new_n39029__;
  assign new_new_n39031__ = ~new_new_n38899__ & ~new_new_n38912__;
  assign new_new_n39032__ = ~new_new_n38917__ & ~new_new_n39031__;
  assign new_new_n39033__ = new_new_n38909__ & ~new_new_n39032__;
  assign new_new_n39034__ = ~new_new_n38909__ & new_new_n39032__;
  assign new_new_n39035__ = ~new_new_n39033__ & ~new_new_n39034__;
  assign new_new_n39036__ = ~new_new_n38899__ & new_new_n38912__;
  assign new_new_n39037__ = new_new_n38899__ & ~new_new_n38912__;
  assign new_new_n39038__ = ~new_new_n39036__ & ~new_new_n39037__;
  assign new_new_n39039__ = ~new_new_n39035__ & ~new_new_n39038__;
  assign new_new_n39040__ = new_new_n38905__ & ~new_new_n39025__;
  assign new_new_n39041__ = ~new_new_n38905__ & new_new_n39025__;
  assign new_new_n39042__ = ~new_new_n39040__ & ~new_new_n39041__;
  assign new_new_n39043__ = ~new_new_n38886__ & ~new_new_n38892__;
  assign new_new_n39044__ = ~new_new_n38896__ & ~new_new_n39043__;
  assign new_new_n39045__ = new_new_n38889__ & ~new_new_n39044__;
  assign new_new_n39046__ = ~new_new_n38889__ & new_new_n39044__;
  assign new_new_n39047__ = ~new_new_n39045__ & ~new_new_n39046__;
  assign new_new_n39048__ = ~new_new_n38886__ & new_new_n38892__;
  assign new_new_n39049__ = new_new_n38886__ & ~new_new_n38892__;
  assign new_new_n39050__ = ~new_new_n39048__ & ~new_new_n39049__;
  assign new_new_n39051__ = new_new_n38883__ & new_new_n38884__;
  assign new_new_n39052__ = ~new_new_n38883__ & ~new_new_n38884__;
  assign new_new_n39053__ = ~new_new_n39051__ & ~new_new_n39052__;
  assign new_new_n39054__ = ~ys__n30334 & ~ys__n33579;
  assign new_new_n39055__ = ys__n30334 & ys__n33579;
  assign new_new_n39056__ = ~new_new_n39054__ & ~new_new_n39055__;
  assign new_new_n39057__ = ~ys__n30334 & ~new_new_n39056__;
  assign new_new_n39058__ = ~new_new_n39053__ & new_new_n39057__;
  assign new_new_n39059__ = ~new_new_n39050__ & new_new_n39058__;
  assign new_new_n39060__ = ~new_new_n39047__ & new_new_n39059__;
  assign new_new_n39061__ = ~new_new_n39042__ & new_new_n39060__;
  assign new_new_n39062__ = new_new_n39039__ & new_new_n39061__;
  assign new_new_n39063__ = ~new_new_n39030__ & new_new_n39062__;
  assign new_new_n39064__ = ~new_new_n39023__ & new_new_n39063__;
  assign new_new_n39065__ = new_new_n39020__ & new_new_n39064__;
  assign new_new_n39066__ = new_new_n39011__ & new_new_n39065__;
  assign new_new_n39067__ = ~new_new_n38990__ & new_new_n39066__;
  assign new_new_n39068__ = new_new_n38981__ & new_new_n39067__;
  assign new_new_n39069__ = ~new_new_n38981__ & ~new_new_n39067__;
  assign new_new_n39070__ = ~new_new_n39068__ & ~new_new_n39069__;
  assign new_new_n39071__ = ~ys__n17848 & ~new_new_n38454__;
  assign new_new_n39072__ = ys__n17848 & new_new_n38454__;
  assign new_new_n39073__ = ~new_new_n39071__ & ~new_new_n39072__;
  assign new_new_n39074__ = ys__n17825 & ~new_new_n38209__;
  assign new_new_n39075__ = ~ys__n17825 & ~new_new_n38209__;
  assign new_new_n39076__ = ys__n17825 & new_new_n38209__;
  assign new_new_n39077__ = ~new_new_n39075__ & ~new_new_n39076__;
  assign new_new_n39078__ = ys__n17824 & ~new_new_n38206__;
  assign new_new_n39079__ = ~new_new_n39077__ & new_new_n39078__;
  assign new_new_n39080__ = ~new_new_n39074__ & ~new_new_n39079__;
  assign new_new_n39081__ = ~ys__n17828 & ~new_new_n38611__;
  assign new_new_n39082__ = ys__n17828 & new_new_n38611__;
  assign new_new_n39083__ = ~new_new_n39081__ & ~new_new_n39082__;
  assign new_new_n39084__ = ~ys__n17827 & ~new_new_n38608__;
  assign new_new_n39085__ = ys__n17827 & new_new_n38608__;
  assign new_new_n39086__ = ~new_new_n39084__ & ~new_new_n39085__;
  assign new_new_n39087__ = ~new_new_n39083__ & ~new_new_n39086__;
  assign new_new_n39088__ = ~new_new_n39080__ & new_new_n39087__;
  assign new_new_n39089__ = ys__n17828 & ~new_new_n38611__;
  assign new_new_n39090__ = ys__n17827 & ~new_new_n38608__;
  assign new_new_n39091__ = ~new_new_n39083__ & new_new_n39090__;
  assign new_new_n39092__ = ~new_new_n39089__ & ~new_new_n39091__;
  assign new_new_n39093__ = ~new_new_n39088__ & new_new_n39092__;
  assign new_new_n39094__ = ~ys__n17834 & ~new_new_n38686__;
  assign new_new_n39095__ = ys__n17834 & new_new_n38686__;
  assign new_new_n39096__ = ~new_new_n39094__ & ~new_new_n39095__;
  assign new_new_n39097__ = ~ys__n17833 & ~new_new_n38702__;
  assign new_new_n39098__ = ys__n17833 & new_new_n38702__;
  assign new_new_n39099__ = ~new_new_n39097__ & ~new_new_n39098__;
  assign new_new_n39100__ = ~new_new_n39096__ & ~new_new_n39099__;
  assign new_new_n39101__ = ~ys__n17831 & ~new_new_n38644__;
  assign new_new_n39102__ = ys__n17831 & new_new_n38644__;
  assign new_new_n39103__ = ~new_new_n39101__ & ~new_new_n39102__;
  assign new_new_n39104__ = ~ys__n17830 & ~new_new_n38641__;
  assign new_new_n39105__ = ys__n17830 & new_new_n38641__;
  assign new_new_n39106__ = ~new_new_n39104__ & ~new_new_n39105__;
  assign new_new_n39107__ = ~new_new_n39103__ & ~new_new_n39106__;
  assign new_new_n39108__ = new_new_n39100__ & new_new_n39107__;
  assign new_new_n39109__ = ~new_new_n39093__ & new_new_n39108__;
  assign new_new_n39110__ = ys__n17831 & ~new_new_n38644__;
  assign new_new_n39111__ = ys__n17830 & ~new_new_n38641__;
  assign new_new_n39112__ = ~new_new_n39103__ & new_new_n39111__;
  assign new_new_n39113__ = ~new_new_n39110__ & ~new_new_n39112__;
  assign new_new_n39114__ = new_new_n39100__ & ~new_new_n39113__;
  assign new_new_n39115__ = ys__n17834 & ~new_new_n38686__;
  assign new_new_n39116__ = ys__n17833 & ~new_new_n38702__;
  assign new_new_n39117__ = ~new_new_n39096__ & new_new_n39116__;
  assign new_new_n39118__ = ~new_new_n39115__ & ~new_new_n39117__;
  assign new_new_n39119__ = ~new_new_n39114__ & new_new_n39118__;
  assign new_new_n39120__ = ~new_new_n39109__ & new_new_n39119__;
  assign new_new_n39121__ = ~ys__n17846 & ~new_new_n38467__;
  assign new_new_n39122__ = ys__n17846 & new_new_n38467__;
  assign new_new_n39123__ = ~new_new_n39121__ & ~new_new_n39122__;
  assign new_new_n39124__ = ~ys__n17845 & ~new_new_n38483__;
  assign new_new_n39125__ = ys__n17845 & new_new_n38483__;
  assign new_new_n39126__ = ~new_new_n39124__ & ~new_new_n39125__;
  assign new_new_n39127__ = ~new_new_n39123__ & ~new_new_n39126__;
  assign new_new_n39128__ = ~ys__n17843 & ~new_new_n38500__;
  assign new_new_n39129__ = ys__n17843 & new_new_n38500__;
  assign new_new_n39130__ = ~new_new_n39128__ & ~new_new_n39129__;
  assign new_new_n39131__ = ~ys__n17842 & ~new_new_n38517__;
  assign new_new_n39132__ = ys__n17842 & new_new_n38517__;
  assign new_new_n39133__ = ~new_new_n39131__ & ~new_new_n39132__;
  assign new_new_n39134__ = ~new_new_n39130__ & ~new_new_n39133__;
  assign new_new_n39135__ = new_new_n39127__ & new_new_n39134__;
  assign new_new_n39136__ = ~ys__n17840 & ~new_new_n38537__;
  assign new_new_n39137__ = ys__n17840 & new_new_n38537__;
  assign new_new_n39138__ = ~new_new_n39136__ & ~new_new_n39137__;
  assign new_new_n39139__ = ~ys__n17839 & ~new_new_n38553__;
  assign new_new_n39140__ = ys__n17839 & new_new_n38553__;
  assign new_new_n39141__ = ~new_new_n39139__ & ~new_new_n39140__;
  assign new_new_n39142__ = ~new_new_n39138__ & ~new_new_n39141__;
  assign new_new_n39143__ = ~ys__n17837 & ~new_new_n38570__;
  assign new_new_n39144__ = ys__n17837 & new_new_n38570__;
  assign new_new_n39145__ = ~new_new_n39143__ & ~new_new_n39144__;
  assign new_new_n39146__ = ~ys__n17836 & ~new_new_n38587__;
  assign new_new_n39147__ = ys__n17836 & new_new_n38587__;
  assign new_new_n39148__ = ~new_new_n39146__ & ~new_new_n39147__;
  assign new_new_n39149__ = ~new_new_n39145__ & ~new_new_n39148__;
  assign new_new_n39150__ = new_new_n39142__ & new_new_n39149__;
  assign new_new_n39151__ = new_new_n39135__ & new_new_n39150__;
  assign new_new_n39152__ = ~new_new_n39120__ & new_new_n39151__;
  assign new_new_n39153__ = ys__n17837 & ~new_new_n38570__;
  assign new_new_n39154__ = ys__n17836 & ~new_new_n38587__;
  assign new_new_n39155__ = ~new_new_n39145__ & new_new_n39154__;
  assign new_new_n39156__ = ~new_new_n39153__ & ~new_new_n39155__;
  assign new_new_n39157__ = new_new_n39142__ & ~new_new_n39156__;
  assign new_new_n39158__ = ys__n17840 & ~new_new_n38537__;
  assign new_new_n39159__ = ys__n17839 & ~new_new_n38553__;
  assign new_new_n39160__ = ~new_new_n39138__ & new_new_n39159__;
  assign new_new_n39161__ = ~new_new_n39158__ & ~new_new_n39160__;
  assign new_new_n39162__ = ~new_new_n39157__ & new_new_n39161__;
  assign new_new_n39163__ = new_new_n39135__ & ~new_new_n39162__;
  assign new_new_n39164__ = ys__n17843 & ~new_new_n38500__;
  assign new_new_n39165__ = ys__n17842 & ~new_new_n38517__;
  assign new_new_n39166__ = ~new_new_n39130__ & new_new_n39165__;
  assign new_new_n39167__ = ~new_new_n39164__ & ~new_new_n39166__;
  assign new_new_n39168__ = new_new_n39127__ & ~new_new_n39167__;
  assign new_new_n39169__ = ys__n17846 & ~new_new_n38467__;
  assign new_new_n39170__ = ys__n17845 & ~new_new_n38483__;
  assign new_new_n39171__ = ~new_new_n39123__ & new_new_n39170__;
  assign new_new_n39172__ = ~new_new_n39169__ & ~new_new_n39171__;
  assign new_new_n39173__ = ~new_new_n39168__ & new_new_n39172__;
  assign new_new_n39174__ = ~new_new_n39163__ & new_new_n39173__;
  assign new_new_n39175__ = ~new_new_n39152__ & new_new_n39174__;
  assign new_new_n39176__ = new_new_n39073__ & ~new_new_n39175__;
  assign new_new_n39177__ = ~new_new_n39073__ & new_new_n39175__;
  assign new_new_n39178__ = ~new_new_n39176__ & ~new_new_n39177__;
  assign new_new_n39179__ = new_new_n39070__ & ~new_new_n39178__;
  assign new_new_n39180__ = ~new_new_n39120__ & new_new_n39150__;
  assign new_new_n39181__ = new_new_n39162__ & ~new_new_n39180__;
  assign new_new_n39182__ = new_new_n39134__ & ~new_new_n39181__;
  assign new_new_n39183__ = new_new_n39167__ & ~new_new_n39182__;
  assign new_new_n39184__ = ~new_new_n39126__ & ~new_new_n39183__;
  assign new_new_n39185__ = ~new_new_n39170__ & ~new_new_n39184__;
  assign new_new_n39186__ = new_new_n39123__ & ~new_new_n39185__;
  assign new_new_n39187__ = ~new_new_n39123__ & new_new_n39185__;
  assign new_new_n39188__ = ~new_new_n39186__ & ~new_new_n39187__;
  assign new_new_n39189__ = ~new_new_n39120__ & new_new_n39149__;
  assign new_new_n39190__ = new_new_n39156__ & ~new_new_n39189__;
  assign new_new_n39191__ = ~new_new_n39141__ & ~new_new_n39190__;
  assign new_new_n39192__ = ~new_new_n39159__ & ~new_new_n39191__;
  assign new_new_n39193__ = new_new_n39138__ & ~new_new_n39192__;
  assign new_new_n39194__ = ~new_new_n39138__ & new_new_n39192__;
  assign new_new_n39195__ = ~new_new_n39193__ & ~new_new_n39194__;
  assign new_new_n39196__ = new_new_n39141__ & ~new_new_n39190__;
  assign new_new_n39197__ = ~new_new_n39141__ & new_new_n39190__;
  assign new_new_n39198__ = ~new_new_n39196__ & ~new_new_n39197__;
  assign new_new_n39199__ = ~new_new_n39120__ & ~new_new_n39148__;
  assign new_new_n39200__ = ~new_new_n39154__ & ~new_new_n39199__;
  assign new_new_n39201__ = new_new_n39145__ & ~new_new_n39200__;
  assign new_new_n39202__ = ~new_new_n39145__ & new_new_n39200__;
  assign new_new_n39203__ = ~new_new_n39201__ & ~new_new_n39202__;
  assign new_new_n39204__ = ~new_new_n39120__ & new_new_n39148__;
  assign new_new_n39205__ = new_new_n39120__ & ~new_new_n39148__;
  assign new_new_n39206__ = ~new_new_n39204__ & ~new_new_n39205__;
  assign new_new_n39207__ = ~new_new_n39203__ & ~new_new_n39206__;
  assign new_new_n39208__ = ~new_new_n39198__ & new_new_n39207__;
  assign new_new_n39209__ = ~new_new_n39195__ & new_new_n39208__;
  assign new_new_n39210__ = ~new_new_n39133__ & ~new_new_n39181__;
  assign new_new_n39211__ = ~new_new_n39165__ & ~new_new_n39210__;
  assign new_new_n39212__ = new_new_n39130__ & ~new_new_n39211__;
  assign new_new_n39213__ = ~new_new_n39130__ & new_new_n39211__;
  assign new_new_n39214__ = ~new_new_n39212__ & ~new_new_n39213__;
  assign new_new_n39215__ = new_new_n39133__ & ~new_new_n39181__;
  assign new_new_n39216__ = ~new_new_n39133__ & new_new_n39181__;
  assign new_new_n39217__ = ~new_new_n39215__ & ~new_new_n39216__;
  assign new_new_n39218__ = ~new_new_n39214__ & ~new_new_n39217__;
  assign new_new_n39219__ = new_new_n39126__ & ~new_new_n39183__;
  assign new_new_n39220__ = ~new_new_n39126__ & new_new_n39183__;
  assign new_new_n39221__ = ~new_new_n39219__ & ~new_new_n39220__;
  assign new_new_n39222__ = ~new_new_n39093__ & new_new_n39107__;
  assign new_new_n39223__ = new_new_n39113__ & ~new_new_n39222__;
  assign new_new_n39224__ = ~new_new_n39099__ & ~new_new_n39223__;
  assign new_new_n39225__ = ~new_new_n39116__ & ~new_new_n39224__;
  assign new_new_n39226__ = new_new_n39096__ & ~new_new_n39225__;
  assign new_new_n39227__ = ~new_new_n39096__ & new_new_n39225__;
  assign new_new_n39228__ = ~new_new_n39226__ & ~new_new_n39227__;
  assign new_new_n39229__ = ~new_new_n39093__ & ~new_new_n39106__;
  assign new_new_n39230__ = ~new_new_n39111__ & ~new_new_n39229__;
  assign new_new_n39231__ = new_new_n39103__ & ~new_new_n39230__;
  assign new_new_n39232__ = ~new_new_n39103__ & new_new_n39230__;
  assign new_new_n39233__ = ~new_new_n39231__ & ~new_new_n39232__;
  assign new_new_n39234__ = ~new_new_n39093__ & new_new_n39106__;
  assign new_new_n39235__ = new_new_n39093__ & ~new_new_n39106__;
  assign new_new_n39236__ = ~new_new_n39234__ & ~new_new_n39235__;
  assign new_new_n39237__ = ~new_new_n39233__ & ~new_new_n39236__;
  assign new_new_n39238__ = new_new_n39099__ & ~new_new_n39223__;
  assign new_new_n39239__ = ~new_new_n39099__ & new_new_n39223__;
  assign new_new_n39240__ = ~new_new_n39238__ & ~new_new_n39239__;
  assign new_new_n39241__ = ~new_new_n39080__ & ~new_new_n39086__;
  assign new_new_n39242__ = ~new_new_n39090__ & ~new_new_n39241__;
  assign new_new_n39243__ = new_new_n39083__ & ~new_new_n39242__;
  assign new_new_n39244__ = ~new_new_n39083__ & new_new_n39242__;
  assign new_new_n39245__ = ~new_new_n39243__ & ~new_new_n39244__;
  assign new_new_n39246__ = ~new_new_n39080__ & new_new_n39086__;
  assign new_new_n39247__ = new_new_n39080__ & ~new_new_n39086__;
  assign new_new_n39248__ = ~new_new_n39246__ & ~new_new_n39247__;
  assign new_new_n39249__ = new_new_n39077__ & new_new_n39078__;
  assign new_new_n39250__ = ~new_new_n39077__ & ~new_new_n39078__;
  assign new_new_n39251__ = ~new_new_n39249__ & ~new_new_n39250__;
  assign new_new_n39252__ = ~ys__n17824 & ~new_new_n38206__;
  assign new_new_n39253__ = ys__n17824 & new_new_n38206__;
  assign new_new_n39254__ = ~new_new_n39252__ & ~new_new_n39253__;
  assign new_new_n39255__ = ~new_new_n39251__ & ~new_new_n39254__;
  assign new_new_n39256__ = ~new_new_n39248__ & new_new_n39255__;
  assign new_new_n39257__ = ~new_new_n39245__ & new_new_n39256__;
  assign new_new_n39258__ = ~new_new_n39240__ & new_new_n39257__;
  assign new_new_n39259__ = new_new_n39237__ & new_new_n39258__;
  assign new_new_n39260__ = ~new_new_n39228__ & new_new_n39259__;
  assign new_new_n39261__ = ~new_new_n39221__ & new_new_n39260__;
  assign new_new_n39262__ = new_new_n39218__ & new_new_n39261__;
  assign new_new_n39263__ = new_new_n39209__ & new_new_n39262__;
  assign new_new_n39264__ = ~new_new_n39188__ & new_new_n39263__;
  assign new_new_n39265__ = new_new_n39178__ & new_new_n39264__;
  assign new_new_n39266__ = ~new_new_n39178__ & ~new_new_n39264__;
  assign new_new_n39267__ = ~new_new_n39265__ & ~new_new_n39266__;
  assign new_new_n39268__ = ~new_new_n39070__ & ~new_new_n39267__;
  assign new_new_n39269__ = ~new_new_n39179__ & ~new_new_n39268__;
  assign new_new_n39270__ = ys__n18156 & ~new_new_n39269__;
  assign new_new_n39271__ = ys__n17848 & ~new_new_n38454__;
  assign new_new_n39272__ = ~new_new_n39073__ & ~new_new_n39175__;
  assign new_new_n39273__ = ~new_new_n39271__ & ~new_new_n39272__;
  assign new_new_n39274__ = new_new_n38843__ & ~new_new_n39273__;
  assign new_new_n39275__ = ~new_new_n38843__ & new_new_n39273__;
  assign new_new_n39276__ = ~new_new_n39274__ & ~new_new_n39275__;
  assign new_new_n39277__ = new_new_n39070__ & ~new_new_n39276__;
  assign new_new_n39278__ = ~new_new_n39178__ & new_new_n39264__;
  assign new_new_n39279__ = new_new_n39276__ & new_new_n39278__;
  assign new_new_n39280__ = ~new_new_n39276__ & ~new_new_n39278__;
  assign new_new_n39281__ = ~new_new_n39279__ & ~new_new_n39280__;
  assign new_new_n39282__ = ~new_new_n39070__ & ~new_new_n39281__;
  assign new_new_n39283__ = ~new_new_n39277__ & ~new_new_n39282__;
  assign new_new_n39284__ = ~new_new_n39270__ & new_new_n39283__;
  assign new_new_n39285__ = ~new_new_n38879__ & ~new_new_n39284__;
  assign new_new_n39286__ = ys__n33581 & ~new_new_n38051__;
  assign new_new_n39287__ = ys__n33579 & ~new_new_n38064__;
  assign new_new_n39288__ = ~new_new_n38074__ & new_new_n39287__;
  assign new_new_n39289__ = ~new_new_n39286__ & ~new_new_n39288__;
  assign new_new_n39290__ = ~new_new_n38057__ & ~new_new_n38107__;
  assign new_new_n39291__ = ~new_new_n39289__ & new_new_n39290__;
  assign new_new_n39292__ = ys__n17804 & ~new_new_n38088__;
  assign new_new_n39293__ = ys__n17803 & ~new_new_n38054__;
  assign new_new_n39294__ = ~new_new_n38107__ & new_new_n39293__;
  assign new_new_n39295__ = ~new_new_n39292__ & ~new_new_n39294__;
  assign new_new_n39296__ = ~new_new_n39291__ & new_new_n39295__;
  assign new_new_n39297__ = ~new_new_n38149__ & ~new_new_n38166__;
  assign new_new_n39298__ = ~new_new_n38094__ & ~new_new_n38179__;
  assign new_new_n39299__ = new_new_n39297__ & new_new_n39298__;
  assign new_new_n39300__ = ~new_new_n39296__ & new_new_n39299__;
  assign new_new_n39301__ = ys__n17807 & ~new_new_n38156__;
  assign new_new_n39302__ = ys__n17806 & ~new_new_n38091__;
  assign new_new_n39303__ = ~new_new_n38179__ & new_new_n39302__;
  assign new_new_n39304__ = ~new_new_n39301__ & ~new_new_n39303__;
  assign new_new_n39305__ = new_new_n39297__ & ~new_new_n39304__;
  assign new_new_n39306__ = ys__n17810 & ~new_new_n38127__;
  assign new_new_n39307__ = ys__n17809 & ~new_new_n38140__;
  assign new_new_n39308__ = ~new_new_n38149__ & new_new_n39307__;
  assign new_new_n39309__ = ~new_new_n39306__ & ~new_new_n39308__;
  assign new_new_n39310__ = ~new_new_n39305__ & new_new_n39309__;
  assign new_new_n39311__ = ~new_new_n39300__ & new_new_n39310__;
  assign new_new_n39312__ = ~new_new_n38228__ & ~new_new_n38245__;
  assign new_new_n39313__ = ~new_new_n38261__ & ~new_new_n38279__;
  assign new_new_n39314__ = new_new_n39312__ & new_new_n39313__;
  assign new_new_n39315__ = ~new_new_n38295__ & ~new_new_n38312__;
  assign new_new_n39316__ = ~new_new_n38133__ & ~new_new_n38325__;
  assign new_new_n39317__ = new_new_n39315__ & new_new_n39316__;
  assign new_new_n39318__ = new_new_n39314__ & new_new_n39317__;
  assign new_new_n39319__ = ~new_new_n39311__ & new_new_n39318__;
  assign new_new_n39320__ = ys__n17813 & ~new_new_n38302__;
  assign new_new_n39321__ = ys__n17812 & ~new_new_n38130__;
  assign new_new_n39322__ = ~new_new_n38325__ & new_new_n39321__;
  assign new_new_n39323__ = ~new_new_n39320__ & ~new_new_n39322__;
  assign new_new_n39324__ = new_new_n39315__ & ~new_new_n39323__;
  assign new_new_n39325__ = ys__n17816 & ~new_new_n38268__;
  assign new_new_n39326__ = ys__n17815 & ~new_new_n38286__;
  assign new_new_n39327__ = ~new_new_n38295__ & new_new_n39326__;
  assign new_new_n39328__ = ~new_new_n39325__ & ~new_new_n39327__;
  assign new_new_n39329__ = ~new_new_n39324__ & new_new_n39328__;
  assign new_new_n39330__ = new_new_n39314__ & ~new_new_n39329__;
  assign new_new_n39331__ = ys__n17819 & ~new_new_n38235__;
  assign new_new_n39332__ = ys__n17818 & ~new_new_n38252__;
  assign new_new_n39333__ = ~new_new_n38261__ & new_new_n39332__;
  assign new_new_n39334__ = ~new_new_n39331__ & ~new_new_n39333__;
  assign new_new_n39335__ = new_new_n39312__ & ~new_new_n39334__;
  assign new_new_n39336__ = ys__n17822 & ~new_new_n38206__;
  assign new_new_n39337__ = ys__n17821 & ~new_new_n38219__;
  assign new_new_n39338__ = ~new_new_n38228__ & new_new_n39337__;
  assign new_new_n39339__ = ~new_new_n39336__ & ~new_new_n39338__;
  assign new_new_n39340__ = ~new_new_n39335__ & new_new_n39339__;
  assign new_new_n39341__ = ~new_new_n39330__ & new_new_n39340__;
  assign new_new_n39342__ = ~new_new_n39319__ & new_new_n39341__;
  assign new_new_n39343__ = ~new_new_n39311__ & new_new_n39317__;
  assign new_new_n39344__ = new_new_n39329__ & ~new_new_n39343__;
  assign new_new_n39345__ = new_new_n39313__ & ~new_new_n39344__;
  assign new_new_n39346__ = new_new_n39334__ & ~new_new_n39345__;
  assign new_new_n39347__ = ~new_new_n38245__ & ~new_new_n39346__;
  assign new_new_n39348__ = ~new_new_n39337__ & ~new_new_n39347__;
  assign new_new_n39349__ = new_new_n38228__ & ~new_new_n39348__;
  assign new_new_n39350__ = ~new_new_n38228__ & new_new_n39348__;
  assign new_new_n39351__ = ~new_new_n39349__ & ~new_new_n39350__;
  assign new_new_n39352__ = ~new_new_n39311__ & new_new_n39316__;
  assign new_new_n39353__ = new_new_n39323__ & ~new_new_n39352__;
  assign new_new_n39354__ = ~new_new_n38312__ & ~new_new_n39353__;
  assign new_new_n39355__ = ~new_new_n39326__ & ~new_new_n39354__;
  assign new_new_n39356__ = new_new_n38295__ & ~new_new_n39355__;
  assign new_new_n39357__ = ~new_new_n38295__ & new_new_n39355__;
  assign new_new_n39358__ = ~new_new_n39356__ & ~new_new_n39357__;
  assign new_new_n39359__ = new_new_n38312__ & ~new_new_n39353__;
  assign new_new_n39360__ = ~new_new_n38312__ & new_new_n39353__;
  assign new_new_n39361__ = ~new_new_n39359__ & ~new_new_n39360__;
  assign new_new_n39362__ = ~new_new_n38133__ & ~new_new_n39311__;
  assign new_new_n39363__ = ~new_new_n39321__ & ~new_new_n39362__;
  assign new_new_n39364__ = new_new_n38325__ & ~new_new_n39363__;
  assign new_new_n39365__ = ~new_new_n38325__ & new_new_n39363__;
  assign new_new_n39366__ = ~new_new_n39364__ & ~new_new_n39365__;
  assign new_new_n39367__ = new_new_n38133__ & ~new_new_n39311__;
  assign new_new_n39368__ = ~new_new_n38133__ & new_new_n39311__;
  assign new_new_n39369__ = ~new_new_n39367__ & ~new_new_n39368__;
  assign new_new_n39370__ = ~new_new_n39366__ & ~new_new_n39369__;
  assign new_new_n39371__ = ~new_new_n39361__ & new_new_n39370__;
  assign new_new_n39372__ = ~new_new_n39358__ & new_new_n39371__;
  assign new_new_n39373__ = ~new_new_n38279__ & ~new_new_n39344__;
  assign new_new_n39374__ = ~new_new_n39332__ & ~new_new_n39373__;
  assign new_new_n39375__ = new_new_n38261__ & ~new_new_n39374__;
  assign new_new_n39376__ = ~new_new_n38261__ & new_new_n39374__;
  assign new_new_n39377__ = ~new_new_n39375__ & ~new_new_n39376__;
  assign new_new_n39378__ = new_new_n38279__ & ~new_new_n39344__;
  assign new_new_n39379__ = ~new_new_n38279__ & new_new_n39344__;
  assign new_new_n39380__ = ~new_new_n39378__ & ~new_new_n39379__;
  assign new_new_n39381__ = ~new_new_n39377__ & ~new_new_n39380__;
  assign new_new_n39382__ = new_new_n38245__ & ~new_new_n39346__;
  assign new_new_n39383__ = ~new_new_n38245__ & new_new_n39346__;
  assign new_new_n39384__ = ~new_new_n39382__ & ~new_new_n39383__;
  assign new_new_n39385__ = ~new_new_n39296__ & new_new_n39298__;
  assign new_new_n39386__ = new_new_n39304__ & ~new_new_n39385__;
  assign new_new_n39387__ = ~new_new_n38166__ & ~new_new_n39386__;
  assign new_new_n39388__ = ~new_new_n39307__ & ~new_new_n39387__;
  assign new_new_n39389__ = new_new_n38149__ & ~new_new_n39388__;
  assign new_new_n39390__ = ~new_new_n38149__ & new_new_n39388__;
  assign new_new_n39391__ = ~new_new_n39389__ & ~new_new_n39390__;
  assign new_new_n39392__ = ~new_new_n38094__ & ~new_new_n39296__;
  assign new_new_n39393__ = ~new_new_n39302__ & ~new_new_n39392__;
  assign new_new_n39394__ = new_new_n38179__ & ~new_new_n39393__;
  assign new_new_n39395__ = ~new_new_n38179__ & new_new_n39393__;
  assign new_new_n39396__ = ~new_new_n39394__ & ~new_new_n39395__;
  assign new_new_n39397__ = new_new_n38094__ & ~new_new_n39296__;
  assign new_new_n39398__ = ~new_new_n38094__ & new_new_n39296__;
  assign new_new_n39399__ = ~new_new_n39397__ & ~new_new_n39398__;
  assign new_new_n39400__ = ~new_new_n39396__ & ~new_new_n39399__;
  assign new_new_n39401__ = new_new_n38166__ & ~new_new_n39386__;
  assign new_new_n39402__ = ~new_new_n38166__ & new_new_n39386__;
  assign new_new_n39403__ = ~new_new_n39401__ & ~new_new_n39402__;
  assign new_new_n39404__ = ~new_new_n38057__ & ~new_new_n39289__;
  assign new_new_n39405__ = ~new_new_n39293__ & ~new_new_n39404__;
  assign new_new_n39406__ = new_new_n38107__ & ~new_new_n39405__;
  assign new_new_n39407__ = ~new_new_n38107__ & new_new_n39405__;
  assign new_new_n39408__ = ~new_new_n39406__ & ~new_new_n39407__;
  assign new_new_n39409__ = new_new_n38057__ & ~new_new_n39289__;
  assign new_new_n39410__ = ~new_new_n38057__ & new_new_n39289__;
  assign new_new_n39411__ = ~new_new_n39409__ & ~new_new_n39410__;
  assign new_new_n39412__ = new_new_n38074__ & new_new_n39287__;
  assign new_new_n39413__ = ~new_new_n38074__ & ~new_new_n39287__;
  assign new_new_n39414__ = ~new_new_n39412__ & ~new_new_n39413__;
  assign new_new_n39415__ = ys__n33579 & new_new_n38064__;
  assign new_new_n39416__ = ~new_new_n38078__ & ~new_new_n39415__;
  assign new_new_n39417__ = ~ys__n402 & ~ys__n30334;
  assign new_new_n39418__ = ~ys__n402 & ~new_new_n39417__;
  assign new_new_n39419__ = ~new_new_n39416__ & ~new_new_n39418__;
  assign new_new_n39420__ = ~new_new_n39414__ & new_new_n39419__;
  assign new_new_n39421__ = ~new_new_n39411__ & new_new_n39420__;
  assign new_new_n39422__ = ~new_new_n39408__ & new_new_n39421__;
  assign new_new_n39423__ = ~new_new_n39403__ & new_new_n39422__;
  assign new_new_n39424__ = new_new_n39400__ & new_new_n39423__;
  assign new_new_n39425__ = ~new_new_n39391__ & new_new_n39424__;
  assign new_new_n39426__ = ~new_new_n39384__ & new_new_n39425__;
  assign new_new_n39427__ = new_new_n39381__ & new_new_n39426__;
  assign new_new_n39428__ = new_new_n39372__ & new_new_n39427__;
  assign new_new_n39429__ = ~new_new_n39351__ & new_new_n39428__;
  assign new_new_n39430__ = new_new_n39342__ & new_new_n39429__;
  assign new_new_n39431__ = ~new_new_n39342__ & ~new_new_n39429__;
  assign new_new_n39432__ = ~new_new_n39430__ & ~new_new_n39431__;
  assign new_new_n39433__ = ys__n17825 & ~new_new_n38608__;
  assign new_new_n39434__ = ys__n17824 & ~new_new_n38209__;
  assign new_new_n39435__ = ~new_new_n38628__ & new_new_n39434__;
  assign new_new_n39436__ = ~new_new_n39433__ & ~new_new_n39435__;
  assign new_new_n39437__ = ~new_new_n38614__ & ~new_new_n38660__;
  assign new_new_n39438__ = ~new_new_n39436__ & new_new_n39437__;
  assign new_new_n39439__ = ys__n17828 & ~new_new_n38641__;
  assign new_new_n39440__ = ys__n17827 & ~new_new_n38611__;
  assign new_new_n39441__ = ~new_new_n38660__ & new_new_n39440__;
  assign new_new_n39442__ = ~new_new_n39439__ & ~new_new_n39441__;
  assign new_new_n39443__ = ~new_new_n39438__ & new_new_n39442__;
  assign new_new_n39444__ = ~new_new_n38695__ & ~new_new_n38712__;
  assign new_new_n39445__ = ~new_new_n38647__ & ~new_new_n38725__;
  assign new_new_n39446__ = new_new_n39444__ & new_new_n39445__;
  assign new_new_n39447__ = ~new_new_n39443__ & new_new_n39446__;
  assign new_new_n39448__ = ys__n17831 & ~new_new_n38702__;
  assign new_new_n39449__ = ys__n17830 & ~new_new_n38644__;
  assign new_new_n39450__ = ~new_new_n38725__ & new_new_n39449__;
  assign new_new_n39451__ = ~new_new_n39448__ & ~new_new_n39450__;
  assign new_new_n39452__ = new_new_n39444__ & ~new_new_n39451__;
  assign new_new_n39453__ = ys__n17834 & ~new_new_n38587__;
  assign new_new_n39454__ = ys__n17833 & ~new_new_n38686__;
  assign new_new_n39455__ = ~new_new_n38695__ & new_new_n39454__;
  assign new_new_n39456__ = ~new_new_n39453__ & ~new_new_n39455__;
  assign new_new_n39457__ = ~new_new_n39452__ & new_new_n39456__;
  assign new_new_n39458__ = ~new_new_n39447__ & new_new_n39457__;
  assign new_new_n39459__ = ~new_new_n38476__ & ~new_new_n38493__;
  assign new_new_n39460__ = ~new_new_n38510__ & ~new_new_n38530__;
  assign new_new_n39461__ = new_new_n39459__ & new_new_n39460__;
  assign new_new_n39462__ = ~new_new_n38546__ & ~new_new_n38563__;
  assign new_new_n39463__ = ~new_new_n38580__ & ~new_new_n38679__;
  assign new_new_n39464__ = new_new_n39462__ & new_new_n39463__;
  assign new_new_n39465__ = new_new_n39461__ & new_new_n39464__;
  assign new_new_n39466__ = ~new_new_n39458__ & new_new_n39465__;
  assign new_new_n39467__ = ys__n17837 & ~new_new_n38553__;
  assign new_new_n39468__ = ys__n17836 & ~new_new_n38570__;
  assign new_new_n39469__ = ~new_new_n38580__ & new_new_n39468__;
  assign new_new_n39470__ = ~new_new_n39467__ & ~new_new_n39469__;
  assign new_new_n39471__ = new_new_n39462__ & ~new_new_n39470__;
  assign new_new_n39472__ = ys__n17840 & ~new_new_n38517__;
  assign new_new_n39473__ = ys__n17839 & ~new_new_n38537__;
  assign new_new_n39474__ = ~new_new_n38546__ & new_new_n39473__;
  assign new_new_n39475__ = ~new_new_n39472__ & ~new_new_n39474__;
  assign new_new_n39476__ = ~new_new_n39471__ & new_new_n39475__;
  assign new_new_n39477__ = new_new_n39461__ & ~new_new_n39476__;
  assign new_new_n39478__ = ys__n17843 & ~new_new_n38483__;
  assign new_new_n39479__ = ys__n17842 & ~new_new_n38500__;
  assign new_new_n39480__ = ~new_new_n38510__ & new_new_n39479__;
  assign new_new_n39481__ = ~new_new_n39478__ & ~new_new_n39480__;
  assign new_new_n39482__ = new_new_n39459__ & ~new_new_n39481__;
  assign new_new_n39483__ = ys__n17846 & ~new_new_n38454__;
  assign new_new_n39484__ = ys__n17845 & ~new_new_n38467__;
  assign new_new_n39485__ = ~new_new_n38476__ & new_new_n39484__;
  assign new_new_n39486__ = ~new_new_n39483__ & ~new_new_n39485__;
  assign new_new_n39487__ = ~new_new_n39482__ & new_new_n39486__;
  assign new_new_n39488__ = ~new_new_n39477__ & new_new_n39487__;
  assign new_new_n39489__ = ~new_new_n39466__ & new_new_n39488__;
  assign new_new_n39490__ = new_new_n38460__ & ~new_new_n39489__;
  assign new_new_n39491__ = ~new_new_n38460__ & new_new_n39489__;
  assign new_new_n39492__ = ~new_new_n39490__ & ~new_new_n39491__;
  assign new_new_n39493__ = new_new_n39432__ & ~new_new_n39492__;
  assign new_new_n39494__ = ~new_new_n39458__ & new_new_n39464__;
  assign new_new_n39495__ = new_new_n39476__ & ~new_new_n39494__;
  assign new_new_n39496__ = new_new_n39460__ & ~new_new_n39495__;
  assign new_new_n39497__ = new_new_n39481__ & ~new_new_n39496__;
  assign new_new_n39498__ = ~new_new_n38493__ & ~new_new_n39497__;
  assign new_new_n39499__ = ~new_new_n39484__ & ~new_new_n39498__;
  assign new_new_n39500__ = new_new_n38476__ & ~new_new_n39499__;
  assign new_new_n39501__ = ~new_new_n38476__ & new_new_n39499__;
  assign new_new_n39502__ = ~new_new_n39500__ & ~new_new_n39501__;
  assign new_new_n39503__ = ~new_new_n39458__ & new_new_n39463__;
  assign new_new_n39504__ = new_new_n39470__ & ~new_new_n39503__;
  assign new_new_n39505__ = ~new_new_n38563__ & ~new_new_n39504__;
  assign new_new_n39506__ = ~new_new_n39473__ & ~new_new_n39505__;
  assign new_new_n39507__ = new_new_n38546__ & ~new_new_n39506__;
  assign new_new_n39508__ = ~new_new_n38546__ & new_new_n39506__;
  assign new_new_n39509__ = ~new_new_n39507__ & ~new_new_n39508__;
  assign new_new_n39510__ = new_new_n38563__ & ~new_new_n39504__;
  assign new_new_n39511__ = ~new_new_n38563__ & new_new_n39504__;
  assign new_new_n39512__ = ~new_new_n39510__ & ~new_new_n39511__;
  assign new_new_n39513__ = ~new_new_n38679__ & ~new_new_n39458__;
  assign new_new_n39514__ = ~new_new_n39468__ & ~new_new_n39513__;
  assign new_new_n39515__ = new_new_n38580__ & ~new_new_n39514__;
  assign new_new_n39516__ = ~new_new_n38580__ & new_new_n39514__;
  assign new_new_n39517__ = ~new_new_n39515__ & ~new_new_n39516__;
  assign new_new_n39518__ = new_new_n38679__ & ~new_new_n39458__;
  assign new_new_n39519__ = ~new_new_n38679__ & new_new_n39458__;
  assign new_new_n39520__ = ~new_new_n39518__ & ~new_new_n39519__;
  assign new_new_n39521__ = ~new_new_n39517__ & ~new_new_n39520__;
  assign new_new_n39522__ = ~new_new_n39512__ & new_new_n39521__;
  assign new_new_n39523__ = ~new_new_n39509__ & new_new_n39522__;
  assign new_new_n39524__ = ~new_new_n38530__ & ~new_new_n39495__;
  assign new_new_n39525__ = ~new_new_n39479__ & ~new_new_n39524__;
  assign new_new_n39526__ = new_new_n38510__ & ~new_new_n39525__;
  assign new_new_n39527__ = ~new_new_n38510__ & new_new_n39525__;
  assign new_new_n39528__ = ~new_new_n39526__ & ~new_new_n39527__;
  assign new_new_n39529__ = new_new_n38530__ & ~new_new_n39495__;
  assign new_new_n39530__ = ~new_new_n38530__ & new_new_n39495__;
  assign new_new_n39531__ = ~new_new_n39529__ & ~new_new_n39530__;
  assign new_new_n39532__ = ~new_new_n39528__ & ~new_new_n39531__;
  assign new_new_n39533__ = new_new_n38493__ & ~new_new_n39497__;
  assign new_new_n39534__ = ~new_new_n38493__ & new_new_n39497__;
  assign new_new_n39535__ = ~new_new_n39533__ & ~new_new_n39534__;
  assign new_new_n39536__ = ~new_new_n39443__ & new_new_n39445__;
  assign new_new_n39537__ = new_new_n39451__ & ~new_new_n39536__;
  assign new_new_n39538__ = ~new_new_n38712__ & ~new_new_n39537__;
  assign new_new_n39539__ = ~new_new_n39454__ & ~new_new_n39538__;
  assign new_new_n39540__ = new_new_n38695__ & ~new_new_n39539__;
  assign new_new_n39541__ = ~new_new_n38695__ & new_new_n39539__;
  assign new_new_n39542__ = ~new_new_n39540__ & ~new_new_n39541__;
  assign new_new_n39543__ = ~new_new_n38647__ & ~new_new_n39443__;
  assign new_new_n39544__ = ~new_new_n39449__ & ~new_new_n39543__;
  assign new_new_n39545__ = new_new_n38725__ & ~new_new_n39544__;
  assign new_new_n39546__ = ~new_new_n38725__ & new_new_n39544__;
  assign new_new_n39547__ = ~new_new_n39545__ & ~new_new_n39546__;
  assign new_new_n39548__ = new_new_n38647__ & ~new_new_n39443__;
  assign new_new_n39549__ = ~new_new_n38647__ & new_new_n39443__;
  assign new_new_n39550__ = ~new_new_n39548__ & ~new_new_n39549__;
  assign new_new_n39551__ = ~new_new_n39547__ & ~new_new_n39550__;
  assign new_new_n39552__ = new_new_n38712__ & ~new_new_n39537__;
  assign new_new_n39553__ = ~new_new_n38712__ & new_new_n39537__;
  assign new_new_n39554__ = ~new_new_n39552__ & ~new_new_n39553__;
  assign new_new_n39555__ = ~new_new_n38614__ & ~new_new_n39436__;
  assign new_new_n39556__ = ~new_new_n39440__ & ~new_new_n39555__;
  assign new_new_n39557__ = new_new_n38660__ & ~new_new_n39556__;
  assign new_new_n39558__ = ~new_new_n38660__ & new_new_n39556__;
  assign new_new_n39559__ = ~new_new_n39557__ & ~new_new_n39558__;
  assign new_new_n39560__ = new_new_n38614__ & ~new_new_n39436__;
  assign new_new_n39561__ = ~new_new_n38614__ & new_new_n39436__;
  assign new_new_n39562__ = ~new_new_n39560__ & ~new_new_n39561__;
  assign new_new_n39563__ = new_new_n38628__ & new_new_n39434__;
  assign new_new_n39564__ = ~new_new_n38628__ & ~new_new_n39434__;
  assign new_new_n39565__ = ~new_new_n39563__ & ~new_new_n39564__;
  assign new_new_n39566__ = ~new_new_n38212__ & ~new_new_n39565__;
  assign new_new_n39567__ = ~new_new_n39562__ & new_new_n39566__;
  assign new_new_n39568__ = ~new_new_n39559__ & new_new_n39567__;
  assign new_new_n39569__ = ~new_new_n39554__ & new_new_n39568__;
  assign new_new_n39570__ = new_new_n39551__ & new_new_n39569__;
  assign new_new_n39571__ = ~new_new_n39542__ & new_new_n39570__;
  assign new_new_n39572__ = ~new_new_n39535__ & new_new_n39571__;
  assign new_new_n39573__ = new_new_n39532__ & new_new_n39572__;
  assign new_new_n39574__ = new_new_n39523__ & new_new_n39573__;
  assign new_new_n39575__ = ~new_new_n39502__ & new_new_n39574__;
  assign new_new_n39576__ = new_new_n39492__ & new_new_n39575__;
  assign new_new_n39577__ = ~new_new_n39492__ & ~new_new_n39575__;
  assign new_new_n39578__ = ~new_new_n39576__ & ~new_new_n39577__;
  assign new_new_n39579__ = ~new_new_n39432__ & ~new_new_n39578__;
  assign new_new_n39580__ = ~new_new_n39493__ & ~new_new_n39579__;
  assign new_new_n39581__ = ys__n18156 & ~new_new_n39580__;
  assign new_new_n39582__ = ys__n17848 & ~new_new_n38457__;
  assign new_new_n39583__ = ~new_new_n38460__ & ~new_new_n39489__;
  assign new_new_n39584__ = ~new_new_n39582__ & ~new_new_n39583__;
  assign new_new_n39585__ = new_new_n38843__ & ~new_new_n39584__;
  assign new_new_n39586__ = ~new_new_n38843__ & new_new_n39584__;
  assign new_new_n39587__ = ~new_new_n39585__ & ~new_new_n39586__;
  assign new_new_n39588__ = new_new_n39432__ & ~new_new_n39587__;
  assign new_new_n39589__ = ~new_new_n39492__ & new_new_n39575__;
  assign new_new_n39590__ = new_new_n39587__ & new_new_n39589__;
  assign new_new_n39591__ = ~new_new_n39587__ & ~new_new_n39589__;
  assign new_new_n39592__ = ~new_new_n39590__ & ~new_new_n39591__;
  assign new_new_n39593__ = ~new_new_n39432__ & ~new_new_n39592__;
  assign new_new_n39594__ = ~new_new_n39588__ & ~new_new_n39593__;
  assign new_new_n39595__ = ~new_new_n39581__ & new_new_n39594__;
  assign new_new_n39596__ = ys__n408 & ~new_new_n39595__;
  assign new_new_n39597__ = new_new_n39285__ & new_new_n39596__;
  assign new_new_n39598__ = ys__n33579 & new_new_n39597__;
  assign new_new_n39599__ = ~ys__n30334 & new_new_n39416__;
  assign new_new_n39600__ = ys__n30334 & ~new_new_n39416__;
  assign new_new_n39601__ = ~new_new_n39599__ & ~new_new_n39600__;
  assign new_new_n39602__ = ys__n408 & new_new_n38879__;
  assign new_new_n39603__ = ~new_new_n39601__ & new_new_n39602__;
  assign new_new_n39604__ = ys__n402 & ys__n404;
  assign new_new_n39605__ = ys__n402 & ~new_new_n39604__;
  assign new_new_n39606__ = ~ys__n408 & ys__n17803;
  assign new_new_n39607__ = new_new_n39604__ & new_new_n39606__;
  assign new_new_n39608__ = ~new_new_n39605__ & new_new_n39607__;
  assign new_new_n39609__ = ~new_new_n39603__ & ~new_new_n39608__;
  assign new_new_n39610__ = ~new_new_n39598__ & new_new_n39609__;
  assign new_new_n39611__ = new_new_n39416__ & ~new_new_n39418__;
  assign new_new_n39612__ = ~new_new_n39416__ & new_new_n39418__;
  assign new_new_n39613__ = ~new_new_n39611__ & ~new_new_n39612__;
  assign new_new_n39614__ = ys__n408 & new_new_n39595__;
  assign new_new_n39615__ = new_new_n39285__ & new_new_n39614__;
  assign new_new_n39616__ = ~new_new_n39613__ & new_new_n39615__;
  assign new_new_n39617__ = ~ys__n30334 & new_new_n39056__;
  assign new_new_n39618__ = ys__n30334 & ~new_new_n39056__;
  assign new_new_n39619__ = ~new_new_n39617__ & ~new_new_n39618__;
  assign new_new_n39620__ = ~new_new_n38879__ & new_new_n39284__;
  assign new_new_n39621__ = ys__n408 & new_new_n39620__;
  assign new_new_n39622__ = ~new_new_n39619__ & new_new_n39621__;
  assign new_new_n39623__ = ~new_new_n39616__ & ~new_new_n39622__;
  assign new_new_n39624__ = new_new_n39610__ & new_new_n39623__;
  assign new_new_n39625__ = ys__n408 & ~new_new_n39602__;
  assign new_new_n39626__ = ~new_new_n39597__ & new_new_n39625__;
  assign new_new_n39627__ = ~new_new_n39615__ & ~new_new_n39621__;
  assign new_new_n39628__ = new_new_n39626__ & new_new_n39627__;
  assign new_new_n39629__ = ~new_new_n14002__ & ~new_new_n39628__;
  assign new_new_n39630__ = ~new_new_n39624__ & new_new_n39629__;
  assign ys__n30235 = new_new_n38048__ | new_new_n39630__;
  assign new_new_n39632__ = ys__n352 & ys__n23272;
  assign new_new_n39633__ = new_new_n14002__ & new_new_n39632__;
  assign new_new_n39634__ = ys__n33581 & new_new_n39597__;
  assign new_new_n39635__ = ~ys__n30334 & new_new_n38437__;
  assign new_new_n39636__ = ys__n30334 & ~new_new_n38437__;
  assign new_new_n39637__ = ~new_new_n39635__ & ~new_new_n39636__;
  assign new_new_n39638__ = new_new_n39602__ & ~new_new_n39637__;
  assign new_new_n39639__ = ~ys__n17803 & ys__n17804;
  assign new_new_n39640__ = ys__n17803 & ~ys__n17804;
  assign new_new_n39641__ = ~new_new_n39639__ & ~new_new_n39640__;
  assign new_new_n39642__ = ~ys__n408 & new_new_n39604__;
  assign new_new_n39643__ = ~new_new_n39641__ & new_new_n39642__;
  assign new_new_n39644__ = ~new_new_n39605__ & new_new_n39643__;
  assign new_new_n39645__ = ~new_new_n39638__ & ~new_new_n39644__;
  assign new_new_n39646__ = ~new_new_n39634__ & new_new_n39645__;
  assign new_new_n39647__ = new_new_n39414__ & new_new_n39419__;
  assign new_new_n39648__ = ~new_new_n39414__ & ~new_new_n39419__;
  assign new_new_n39649__ = ~new_new_n39647__ & ~new_new_n39648__;
  assign new_new_n39650__ = new_new_n39615__ & ~new_new_n39649__;
  assign new_new_n39651__ = new_new_n39053__ & new_new_n39057__;
  assign new_new_n39652__ = ~new_new_n39053__ & ~new_new_n39057__;
  assign new_new_n39653__ = ~new_new_n39651__ & ~new_new_n39652__;
  assign new_new_n39654__ = new_new_n39621__ & ~new_new_n39653__;
  assign new_new_n39655__ = ~new_new_n39650__ & ~new_new_n39654__;
  assign new_new_n39656__ = new_new_n39646__ & new_new_n39655__;
  assign new_new_n39657__ = new_new_n39629__ & ~new_new_n39656__;
  assign ys__n30238 = new_new_n39633__ | new_new_n39657__;
  assign new_new_n39659__ = ys__n352 & ys__n23274;
  assign new_new_n39660__ = new_new_n14002__ & new_new_n39659__;
  assign new_new_n39661__ = ys__n17803 & new_new_n39597__;
  assign new_new_n39662__ = new_new_n38434__ & new_new_n38438__;
  assign new_new_n39663__ = ~new_new_n38434__ & ~new_new_n38438__;
  assign new_new_n39664__ = ~new_new_n39662__ & ~new_new_n39663__;
  assign new_new_n39665__ = new_new_n39602__ & ~new_new_n39664__;
  assign new_new_n39666__ = ys__n17806 & new_new_n16672__;
  assign new_new_n39667__ = ~ys__n17806 & ~new_new_n16672__;
  assign new_new_n39668__ = ~new_new_n39666__ & ~new_new_n39667__;
  assign new_new_n39669__ = ~new_new_n39605__ & new_new_n39642__;
  assign new_new_n39670__ = ~new_new_n39668__ & new_new_n39669__;
  assign new_new_n39671__ = ~new_new_n39665__ & ~new_new_n39670__;
  assign new_new_n39672__ = ~new_new_n39661__ & new_new_n39671__;
  assign new_new_n39673__ = new_new_n39411__ & new_new_n39420__;
  assign new_new_n39674__ = ~new_new_n39411__ & ~new_new_n39420__;
  assign new_new_n39675__ = ~new_new_n39673__ & ~new_new_n39674__;
  assign new_new_n39676__ = new_new_n39615__ & ~new_new_n39675__;
  assign new_new_n39677__ = new_new_n39050__ & new_new_n39058__;
  assign new_new_n39678__ = ~new_new_n39050__ & ~new_new_n39058__;
  assign new_new_n39679__ = ~new_new_n39677__ & ~new_new_n39678__;
  assign new_new_n39680__ = new_new_n39621__ & ~new_new_n39679__;
  assign new_new_n39681__ = ~new_new_n39676__ & ~new_new_n39680__;
  assign new_new_n39682__ = new_new_n39672__ & new_new_n39681__;
  assign new_new_n39683__ = new_new_n39629__ & ~new_new_n39682__;
  assign ys__n30241 = new_new_n39660__ | new_new_n39683__;
  assign new_new_n39685__ = ys__n352 & ys__n23276;
  assign new_new_n39686__ = new_new_n14002__ & new_new_n39685__;
  assign new_new_n39687__ = ys__n17804 & new_new_n39597__;
  assign new_new_n39688__ = new_new_n38431__ & new_new_n38439__;
  assign new_new_n39689__ = ~new_new_n38431__ & ~new_new_n38439__;
  assign new_new_n39690__ = ~new_new_n39688__ & ~new_new_n39689__;
  assign new_new_n39691__ = new_new_n39602__ & ~new_new_n39690__;
  assign new_new_n39692__ = ~ys__n17806 & new_new_n16672__;
  assign new_new_n39693__ = ys__n17807 & new_new_n39692__;
  assign new_new_n39694__ = ~ys__n17807 & ~new_new_n39692__;
  assign new_new_n39695__ = ~new_new_n39693__ & ~new_new_n39694__;
  assign new_new_n39696__ = new_new_n39669__ & ~new_new_n39695__;
  assign new_new_n39697__ = ~new_new_n39691__ & ~new_new_n39696__;
  assign new_new_n39698__ = ~new_new_n39687__ & new_new_n39697__;
  assign new_new_n39699__ = new_new_n39408__ & new_new_n39421__;
  assign new_new_n39700__ = ~new_new_n39408__ & ~new_new_n39421__;
  assign new_new_n39701__ = ~new_new_n39699__ & ~new_new_n39700__;
  assign new_new_n39702__ = new_new_n39615__ & ~new_new_n39701__;
  assign new_new_n39703__ = new_new_n39047__ & new_new_n39059__;
  assign new_new_n39704__ = ~new_new_n39047__ & ~new_new_n39059__;
  assign new_new_n39705__ = ~new_new_n39703__ & ~new_new_n39704__;
  assign new_new_n39706__ = new_new_n39621__ & ~new_new_n39705__;
  assign new_new_n39707__ = ~new_new_n39702__ & ~new_new_n39706__;
  assign new_new_n39708__ = new_new_n39698__ & new_new_n39707__;
  assign new_new_n39709__ = new_new_n39629__ & ~new_new_n39708__;
  assign ys__n30244 = new_new_n39686__ | new_new_n39709__;
  assign new_new_n39711__ = ys__n352 & ys__n23278;
  assign new_new_n39712__ = new_new_n14002__ & new_new_n39711__;
  assign new_new_n39713__ = ys__n17806 & new_new_n39597__;
  assign new_new_n39714__ = new_new_n38428__ & new_new_n38440__;
  assign new_new_n39715__ = ~new_new_n38428__ & ~new_new_n38440__;
  assign new_new_n39716__ = ~new_new_n39714__ & ~new_new_n39715__;
  assign new_new_n39717__ = new_new_n39602__ & ~new_new_n39716__;
  assign new_new_n39718__ = ys__n17809 & new_new_n16674__;
  assign new_new_n39719__ = ~ys__n17809 & ~new_new_n16674__;
  assign new_new_n39720__ = ~new_new_n39718__ & ~new_new_n39719__;
  assign new_new_n39721__ = new_new_n39669__ & ~new_new_n39720__;
  assign new_new_n39722__ = ~new_new_n39717__ & ~new_new_n39721__;
  assign new_new_n39723__ = ~new_new_n39713__ & new_new_n39722__;
  assign new_new_n39724__ = new_new_n39399__ & new_new_n39422__;
  assign new_new_n39725__ = ~new_new_n39399__ & ~new_new_n39422__;
  assign new_new_n39726__ = ~new_new_n39724__ & ~new_new_n39725__;
  assign new_new_n39727__ = new_new_n39615__ & ~new_new_n39726__;
  assign new_new_n39728__ = new_new_n39038__ & new_new_n39060__;
  assign new_new_n39729__ = ~new_new_n39038__ & ~new_new_n39060__;
  assign new_new_n39730__ = ~new_new_n39728__ & ~new_new_n39729__;
  assign new_new_n39731__ = new_new_n39621__ & ~new_new_n39730__;
  assign new_new_n39732__ = ~new_new_n39727__ & ~new_new_n39731__;
  assign new_new_n39733__ = new_new_n39723__ & new_new_n39732__;
  assign new_new_n39734__ = new_new_n39629__ & ~new_new_n39733__;
  assign ys__n30247 = new_new_n39712__ | new_new_n39734__;
  assign new_new_n39736__ = ys__n352 & ys__n23280;
  assign new_new_n39737__ = new_new_n14002__ & new_new_n39736__;
  assign new_new_n39738__ = ys__n17807 & new_new_n39597__;
  assign new_new_n39739__ = new_new_n38419__ & new_new_n38441__;
  assign new_new_n39740__ = ~new_new_n38419__ & ~new_new_n38441__;
  assign new_new_n39741__ = ~new_new_n39739__ & ~new_new_n39740__;
  assign new_new_n39742__ = new_new_n39602__ & ~new_new_n39741__;
  assign new_new_n39743__ = ~ys__n17809 & new_new_n16674__;
  assign new_new_n39744__ = ys__n17810 & new_new_n39743__;
  assign new_new_n39745__ = ~ys__n17810 & ~new_new_n39743__;
  assign new_new_n39746__ = ~new_new_n39744__ & ~new_new_n39745__;
  assign new_new_n39747__ = new_new_n39669__ & ~new_new_n39746__;
  assign new_new_n39748__ = ~new_new_n39742__ & ~new_new_n39747__;
  assign new_new_n39749__ = ~new_new_n39738__ & new_new_n39748__;
  assign new_new_n39750__ = ~new_new_n39399__ & new_new_n39422__;
  assign new_new_n39751__ = new_new_n39396__ & new_new_n39750__;
  assign new_new_n39752__ = ~new_new_n39396__ & ~new_new_n39750__;
  assign new_new_n39753__ = ~new_new_n39751__ & ~new_new_n39752__;
  assign new_new_n39754__ = new_new_n39615__ & ~new_new_n39753__;
  assign new_new_n39755__ = ~new_new_n39038__ & new_new_n39060__;
  assign new_new_n39756__ = new_new_n39035__ & new_new_n39755__;
  assign new_new_n39757__ = ~new_new_n39035__ & ~new_new_n39755__;
  assign new_new_n39758__ = ~new_new_n39756__ & ~new_new_n39757__;
  assign new_new_n39759__ = new_new_n39621__ & ~new_new_n39758__;
  assign new_new_n39760__ = ~new_new_n39754__ & ~new_new_n39759__;
  assign new_new_n39761__ = new_new_n39749__ & new_new_n39760__;
  assign new_new_n39762__ = new_new_n39629__ & ~new_new_n39761__;
  assign ys__n30250 = new_new_n39737__ | new_new_n39762__;
  assign new_new_n39764__ = ys__n352 & ys__n23282;
  assign new_new_n39765__ = new_new_n14002__ & new_new_n39764__;
  assign new_new_n39766__ = ys__n17809 & new_new_n39597__;
  assign new_new_n39767__ = ~new_new_n38419__ & new_new_n38441__;
  assign new_new_n39768__ = new_new_n38416__ & new_new_n39767__;
  assign new_new_n39769__ = ~new_new_n38416__ & ~new_new_n39767__;
  assign new_new_n39770__ = ~new_new_n39768__ & ~new_new_n39769__;
  assign new_new_n39771__ = new_new_n39602__ & ~new_new_n39770__;
  assign new_new_n39772__ = new_new_n16674__ & new_new_n16675__;
  assign new_new_n39773__ = ys__n17812 & new_new_n39772__;
  assign new_new_n39774__ = ~ys__n17812 & ~new_new_n39772__;
  assign new_new_n39775__ = ~new_new_n39773__ & ~new_new_n39774__;
  assign new_new_n39776__ = new_new_n39669__ & ~new_new_n39775__;
  assign new_new_n39777__ = ~new_new_n39771__ & ~new_new_n39776__;
  assign new_new_n39778__ = ~new_new_n39766__ & new_new_n39777__;
  assign new_new_n39779__ = new_new_n39400__ & new_new_n39422__;
  assign new_new_n39780__ = new_new_n39403__ & new_new_n39779__;
  assign new_new_n39781__ = ~new_new_n39403__ & ~new_new_n39779__;
  assign new_new_n39782__ = ~new_new_n39780__ & ~new_new_n39781__;
  assign new_new_n39783__ = new_new_n39615__ & ~new_new_n39782__;
  assign new_new_n39784__ = new_new_n39039__ & new_new_n39060__;
  assign new_new_n39785__ = new_new_n39042__ & new_new_n39784__;
  assign new_new_n39786__ = ~new_new_n39042__ & ~new_new_n39784__;
  assign new_new_n39787__ = ~new_new_n39785__ & ~new_new_n39786__;
  assign new_new_n39788__ = new_new_n39621__ & ~new_new_n39787__;
  assign new_new_n39789__ = ~new_new_n39783__ & ~new_new_n39788__;
  assign new_new_n39790__ = new_new_n39778__ & new_new_n39789__;
  assign new_new_n39791__ = new_new_n39629__ & ~new_new_n39790__;
  assign ys__n30253 = new_new_n39765__ | new_new_n39791__;
  assign new_new_n39793__ = ys__n352 & ys__n23284;
  assign new_new_n39794__ = new_new_n14002__ & new_new_n39793__;
  assign new_new_n39795__ = ys__n17810 & new_new_n39597__;
  assign new_new_n39796__ = new_new_n38420__ & new_new_n38441__;
  assign new_new_n39797__ = new_new_n38423__ & new_new_n39796__;
  assign new_new_n39798__ = ~new_new_n38423__ & ~new_new_n39796__;
  assign new_new_n39799__ = ~new_new_n39797__ & ~new_new_n39798__;
  assign new_new_n39800__ = new_new_n39602__ & ~new_new_n39799__;
  assign new_new_n39801__ = ~ys__n17812 & new_new_n39772__;
  assign new_new_n39802__ = ys__n17813 & new_new_n39801__;
  assign new_new_n39803__ = ~ys__n17813 & ~new_new_n39801__;
  assign new_new_n39804__ = ~new_new_n39802__ & ~new_new_n39803__;
  assign new_new_n39805__ = new_new_n39669__ & ~new_new_n39804__;
  assign new_new_n39806__ = ~new_new_n39800__ & ~new_new_n39805__;
  assign new_new_n39807__ = ~new_new_n39795__ & new_new_n39806__;
  assign new_new_n39808__ = ~new_new_n39403__ & new_new_n39779__;
  assign new_new_n39809__ = new_new_n39391__ & new_new_n39808__;
  assign new_new_n39810__ = ~new_new_n39391__ & ~new_new_n39808__;
  assign new_new_n39811__ = ~new_new_n39809__ & ~new_new_n39810__;
  assign new_new_n39812__ = new_new_n39615__ & ~new_new_n39811__;
  assign new_new_n39813__ = ~new_new_n39042__ & new_new_n39784__;
  assign new_new_n39814__ = new_new_n39030__ & new_new_n39813__;
  assign new_new_n39815__ = ~new_new_n39030__ & ~new_new_n39813__;
  assign new_new_n39816__ = ~new_new_n39814__ & ~new_new_n39815__;
  assign new_new_n39817__ = new_new_n39621__ & ~new_new_n39816__;
  assign new_new_n39818__ = ~new_new_n39812__ & ~new_new_n39817__;
  assign new_new_n39819__ = new_new_n39807__ & new_new_n39818__;
  assign new_new_n39820__ = new_new_n39629__ & ~new_new_n39819__;
  assign ys__n30256 = new_new_n39794__ | new_new_n39820__;
  assign new_new_n39822__ = ys__n352 & ys__n23286;
  assign new_new_n39823__ = new_new_n14002__ & new_new_n39822__;
  assign new_new_n39824__ = ys__n17812 & new_new_n39597__;
  assign new_new_n39825__ = ~new_new_n38423__ & new_new_n39796__;
  assign new_new_n39826__ = new_new_n38411__ & new_new_n39825__;
  assign new_new_n39827__ = ~new_new_n38411__ & ~new_new_n39825__;
  assign new_new_n39828__ = ~new_new_n39826__ & ~new_new_n39827__;
  assign new_new_n39829__ = new_new_n39602__ & ~new_new_n39828__;
  assign new_new_n39830__ = ys__n17815 & new_new_n16678__;
  assign new_new_n39831__ = ~ys__n17815 & ~new_new_n16678__;
  assign new_new_n39832__ = ~new_new_n39830__ & ~new_new_n39831__;
  assign new_new_n39833__ = new_new_n39669__ & ~new_new_n39832__;
  assign new_new_n39834__ = ~new_new_n39829__ & ~new_new_n39833__;
  assign new_new_n39835__ = ~new_new_n39824__ & new_new_n39834__;
  assign new_new_n39836__ = new_new_n39369__ & new_new_n39425__;
  assign new_new_n39837__ = ~new_new_n39369__ & ~new_new_n39425__;
  assign new_new_n39838__ = ~new_new_n39836__ & ~new_new_n39837__;
  assign new_new_n39839__ = new_new_n39615__ & ~new_new_n39838__;
  assign new_new_n39840__ = new_new_n39008__ & new_new_n39063__;
  assign new_new_n39841__ = ~new_new_n39008__ & ~new_new_n39063__;
  assign new_new_n39842__ = ~new_new_n39840__ & ~new_new_n39841__;
  assign new_new_n39843__ = new_new_n39621__ & ~new_new_n39842__;
  assign new_new_n39844__ = ~new_new_n39839__ & ~new_new_n39843__;
  assign new_new_n39845__ = new_new_n39835__ & new_new_n39844__;
  assign new_new_n39846__ = new_new_n39629__ & ~new_new_n39845__;
  assign ys__n30259 = new_new_n39823__ | new_new_n39846__;
  assign new_new_n39848__ = ys__n352 & ys__n23288;
  assign new_new_n39849__ = new_new_n14002__ & new_new_n39848__;
  assign new_new_n39850__ = ys__n17813 & new_new_n39597__;
  assign new_new_n39851__ = new_new_n38389__ & new_new_n38444__;
  assign new_new_n39852__ = ~new_new_n38389__ & ~new_new_n38444__;
  assign new_new_n39853__ = ~new_new_n39851__ & ~new_new_n39852__;
  assign new_new_n39854__ = new_new_n39602__ & ~new_new_n39853__;
  assign new_new_n39855__ = ~ys__n17815 & new_new_n16678__;
  assign new_new_n39856__ = ys__n17816 & new_new_n39855__;
  assign new_new_n39857__ = ~ys__n17816 & ~new_new_n39855__;
  assign new_new_n39858__ = ~new_new_n39856__ & ~new_new_n39857__;
  assign new_new_n39859__ = new_new_n39669__ & ~new_new_n39858__;
  assign new_new_n39860__ = ~new_new_n39854__ & ~new_new_n39859__;
  assign new_new_n39861__ = ~new_new_n39850__ & new_new_n39860__;
  assign new_new_n39862__ = ~new_new_n39369__ & new_new_n39425__;
  assign new_new_n39863__ = new_new_n39366__ & new_new_n39862__;
  assign new_new_n39864__ = ~new_new_n39366__ & ~new_new_n39862__;
  assign new_new_n39865__ = ~new_new_n39863__ & ~new_new_n39864__;
  assign new_new_n39866__ = new_new_n39615__ & ~new_new_n39865__;
  assign new_new_n39867__ = ~new_new_n39008__ & new_new_n39063__;
  assign new_new_n39868__ = new_new_n39005__ & new_new_n39867__;
  assign new_new_n39869__ = ~new_new_n39005__ & ~new_new_n39867__;
  assign new_new_n39870__ = ~new_new_n39868__ & ~new_new_n39869__;
  assign new_new_n39871__ = new_new_n39621__ & ~new_new_n39870__;
  assign new_new_n39872__ = ~new_new_n39866__ & ~new_new_n39871__;
  assign new_new_n39873__ = new_new_n39861__ & new_new_n39872__;
  assign new_new_n39874__ = new_new_n39629__ & ~new_new_n39873__;
  assign ys__n30262 = new_new_n39849__ | new_new_n39874__;
  assign new_new_n39876__ = ys__n352 & ys__n23290;
  assign new_new_n39877__ = new_new_n14002__ & new_new_n39876__;
  assign new_new_n39878__ = ys__n17815 & new_new_n39597__;
  assign new_new_n39879__ = ~new_new_n38389__ & new_new_n38444__;
  assign new_new_n39880__ = new_new_n38386__ & new_new_n39879__;
  assign new_new_n39881__ = ~new_new_n38386__ & ~new_new_n39879__;
  assign new_new_n39882__ = ~new_new_n39880__ & ~new_new_n39881__;
  assign new_new_n39883__ = new_new_n39602__ & ~new_new_n39882__;
  assign new_new_n39884__ = new_new_n16678__ & new_new_n16679__;
  assign new_new_n39885__ = ys__n17818 & new_new_n39884__;
  assign new_new_n39886__ = ~ys__n17818 & ~new_new_n39884__;
  assign new_new_n39887__ = ~new_new_n39885__ & ~new_new_n39886__;
  assign new_new_n39888__ = new_new_n39669__ & ~new_new_n39887__;
  assign new_new_n39889__ = ~new_new_n39883__ & ~new_new_n39888__;
  assign new_new_n39890__ = ~new_new_n39878__ & new_new_n39889__;
  assign new_new_n39891__ = new_new_n39370__ & new_new_n39425__;
  assign new_new_n39892__ = new_new_n39361__ & new_new_n39891__;
  assign new_new_n39893__ = ~new_new_n39361__ & ~new_new_n39891__;
  assign new_new_n39894__ = ~new_new_n39892__ & ~new_new_n39893__;
  assign new_new_n39895__ = new_new_n39615__ & ~new_new_n39894__;
  assign new_new_n39896__ = new_new_n39009__ & new_new_n39063__;
  assign new_new_n39897__ = new_new_n39000__ & new_new_n39896__;
  assign new_new_n39898__ = ~new_new_n39000__ & ~new_new_n39896__;
  assign new_new_n39899__ = ~new_new_n39897__ & ~new_new_n39898__;
  assign new_new_n39900__ = new_new_n39621__ & ~new_new_n39899__;
  assign new_new_n39901__ = ~new_new_n39895__ & ~new_new_n39900__;
  assign new_new_n39902__ = new_new_n39890__ & new_new_n39901__;
  assign new_new_n39903__ = new_new_n39629__ & ~new_new_n39902__;
  assign ys__n30265 = new_new_n39877__ | new_new_n39903__;
  assign new_new_n39905__ = ys__n352 & ys__n23292;
  assign new_new_n39906__ = new_new_n14002__ & new_new_n39905__;
  assign new_new_n39907__ = ys__n17816 & new_new_n39597__;
  assign new_new_n39908__ = new_new_n38390__ & new_new_n38444__;
  assign new_new_n39909__ = new_new_n38381__ & new_new_n39908__;
  assign new_new_n39910__ = ~new_new_n38381__ & ~new_new_n39908__;
  assign new_new_n39911__ = ~new_new_n39909__ & ~new_new_n39910__;
  assign new_new_n39912__ = new_new_n39602__ & ~new_new_n39911__;
  assign new_new_n39913__ = ~ys__n17818 & new_new_n39884__;
  assign new_new_n39914__ = ys__n17819 & new_new_n39913__;
  assign new_new_n39915__ = ~ys__n17819 & ~new_new_n39913__;
  assign new_new_n39916__ = ~new_new_n39914__ & ~new_new_n39915__;
  assign new_new_n39917__ = new_new_n39669__ & ~new_new_n39916__;
  assign new_new_n39918__ = ~new_new_n39912__ & ~new_new_n39917__;
  assign new_new_n39919__ = ~new_new_n39907__ & new_new_n39918__;
  assign new_new_n39920__ = ~new_new_n39361__ & new_new_n39891__;
  assign new_new_n39921__ = new_new_n39358__ & new_new_n39920__;
  assign new_new_n39922__ = ~new_new_n39358__ & ~new_new_n39920__;
  assign new_new_n39923__ = ~new_new_n39921__ & ~new_new_n39922__;
  assign new_new_n39924__ = new_new_n39615__ & ~new_new_n39923__;
  assign new_new_n39925__ = ~new_new_n39000__ & new_new_n39896__;
  assign new_new_n39926__ = new_new_n38997__ & new_new_n39925__;
  assign new_new_n39927__ = ~new_new_n38997__ & ~new_new_n39925__;
  assign new_new_n39928__ = ~new_new_n39926__ & ~new_new_n39927__;
  assign new_new_n39929__ = new_new_n39621__ & ~new_new_n39928__;
  assign new_new_n39930__ = ~new_new_n39924__ & ~new_new_n39929__;
  assign new_new_n39931__ = new_new_n39919__ & new_new_n39930__;
  assign new_new_n39932__ = new_new_n39629__ & ~new_new_n39931__;
  assign ys__n30268 = new_new_n39906__ | new_new_n39932__;
  assign new_new_n39934__ = ys__n352 & ys__n23294;
  assign new_new_n39935__ = new_new_n14002__ & new_new_n39934__;
  assign new_new_n39936__ = ys__n17818 & new_new_n39597__;
  assign new_new_n39937__ = ~new_new_n38381__ & new_new_n39908__;
  assign new_new_n39938__ = new_new_n38378__ & new_new_n39937__;
  assign new_new_n39939__ = ~new_new_n38378__ & ~new_new_n39937__;
  assign new_new_n39940__ = ~new_new_n39938__ & ~new_new_n39939__;
  assign new_new_n39941__ = new_new_n39602__ & ~new_new_n39940__;
  assign new_new_n39942__ = new_new_n16678__ & new_new_n16681__;
  assign new_new_n39943__ = ys__n17821 & new_new_n39942__;
  assign new_new_n39944__ = ~ys__n17821 & ~new_new_n39942__;
  assign new_new_n39945__ = ~new_new_n39943__ & ~new_new_n39944__;
  assign new_new_n39946__ = new_new_n39669__ & ~new_new_n39945__;
  assign new_new_n39947__ = ~new_new_n39941__ & ~new_new_n39946__;
  assign new_new_n39948__ = ~new_new_n39936__ & new_new_n39947__;
  assign new_new_n39949__ = new_new_n39372__ & new_new_n39425__;
  assign new_new_n39950__ = new_new_n39380__ & new_new_n39949__;
  assign new_new_n39951__ = ~new_new_n39380__ & ~new_new_n39949__;
  assign new_new_n39952__ = ~new_new_n39950__ & ~new_new_n39951__;
  assign new_new_n39953__ = new_new_n39615__ & ~new_new_n39952__;
  assign new_new_n39954__ = new_new_n39011__ & new_new_n39063__;
  assign new_new_n39955__ = new_new_n39019__ & new_new_n39954__;
  assign new_new_n39956__ = ~new_new_n39019__ & ~new_new_n39954__;
  assign new_new_n39957__ = ~new_new_n39955__ & ~new_new_n39956__;
  assign new_new_n39958__ = new_new_n39621__ & ~new_new_n39957__;
  assign new_new_n39959__ = ~new_new_n39953__ & ~new_new_n39958__;
  assign new_new_n39960__ = new_new_n39948__ & new_new_n39959__;
  assign new_new_n39961__ = new_new_n39629__ & ~new_new_n39960__;
  assign ys__n30271 = new_new_n39935__ | new_new_n39961__;
  assign new_new_n39963__ = ys__n352 & ys__n23296;
  assign new_new_n39964__ = new_new_n14002__ & new_new_n39963__;
  assign new_new_n39965__ = ys__n17819 & new_new_n39597__;
  assign new_new_n39966__ = new_new_n38392__ & new_new_n38444__;
  assign new_new_n39967__ = new_new_n38400__ & new_new_n39966__;
  assign new_new_n39968__ = ~new_new_n38400__ & ~new_new_n39966__;
  assign new_new_n39969__ = ~new_new_n39967__ & ~new_new_n39968__;
  assign new_new_n39970__ = new_new_n39602__ & ~new_new_n39969__;
  assign new_new_n39971__ = ~ys__n17821 & new_new_n39942__;
  assign new_new_n39972__ = ys__n17822 & new_new_n39971__;
  assign new_new_n39973__ = ~ys__n17822 & ~new_new_n39971__;
  assign new_new_n39974__ = ~new_new_n39972__ & ~new_new_n39973__;
  assign new_new_n39975__ = new_new_n39669__ & ~new_new_n39974__;
  assign new_new_n39976__ = ~new_new_n39970__ & ~new_new_n39975__;
  assign new_new_n39977__ = ~new_new_n39965__ & new_new_n39976__;
  assign new_new_n39978__ = ~new_new_n39380__ & new_new_n39949__;
  assign new_new_n39979__ = new_new_n39377__ & new_new_n39978__;
  assign new_new_n39980__ = ~new_new_n39377__ & ~new_new_n39978__;
  assign new_new_n39981__ = ~new_new_n39979__ & ~new_new_n39980__;
  assign new_new_n39982__ = new_new_n39615__ & ~new_new_n39981__;
  assign new_new_n39983__ = ~new_new_n39019__ & new_new_n39954__;
  assign new_new_n39984__ = new_new_n39016__ & new_new_n39983__;
  assign new_new_n39985__ = ~new_new_n39016__ & ~new_new_n39983__;
  assign new_new_n39986__ = ~new_new_n39984__ & ~new_new_n39985__;
  assign new_new_n39987__ = new_new_n39621__ & ~new_new_n39986__;
  assign new_new_n39988__ = ~new_new_n39982__ & ~new_new_n39987__;
  assign new_new_n39989__ = new_new_n39977__ & new_new_n39988__;
  assign new_new_n39990__ = new_new_n39629__ & ~new_new_n39989__;
  assign ys__n30274 = new_new_n39964__ | new_new_n39990__;
  assign new_new_n39992__ = ys__n352 & ys__n23298;
  assign new_new_n39993__ = new_new_n14002__ & new_new_n39992__;
  assign new_new_n39994__ = ys__n17821 & new_new_n39597__;
  assign new_new_n39995__ = ~new_new_n38400__ & new_new_n39966__;
  assign new_new_n39996__ = new_new_n38397__ & new_new_n39995__;
  assign new_new_n39997__ = ~new_new_n38397__ & ~new_new_n39995__;
  assign new_new_n39998__ = ~new_new_n39996__ & ~new_new_n39997__;
  assign new_new_n39999__ = new_new_n39602__ & ~new_new_n39998__;
  assign new_new_n40000__ = new_new_n16682__ & new_new_n39942__;
  assign new_new_n40001__ = ys__n17824 & new_new_n40000__;
  assign new_new_n40002__ = ~ys__n17824 & ~new_new_n40000__;
  assign new_new_n40003__ = ~new_new_n40001__ & ~new_new_n40002__;
  assign new_new_n40004__ = new_new_n39669__ & ~new_new_n40003__;
  assign new_new_n40005__ = ~new_new_n39999__ & ~new_new_n40004__;
  assign new_new_n40006__ = ~new_new_n39994__ & new_new_n40005__;
  assign new_new_n40007__ = new_new_n39381__ & new_new_n39949__;
  assign new_new_n40008__ = new_new_n39384__ & new_new_n40007__;
  assign new_new_n40009__ = ~new_new_n39384__ & ~new_new_n40007__;
  assign new_new_n40010__ = ~new_new_n40008__ & ~new_new_n40009__;
  assign new_new_n40011__ = new_new_n39615__ & ~new_new_n40010__;
  assign new_new_n40012__ = new_new_n39020__ & new_new_n39954__;
  assign new_new_n40013__ = new_new_n39023__ & new_new_n40012__;
  assign new_new_n40014__ = ~new_new_n39023__ & ~new_new_n40012__;
  assign new_new_n40015__ = ~new_new_n40013__ & ~new_new_n40014__;
  assign new_new_n40016__ = new_new_n39621__ & ~new_new_n40015__;
  assign new_new_n40017__ = ~new_new_n40011__ & ~new_new_n40016__;
  assign new_new_n40018__ = new_new_n40006__ & new_new_n40017__;
  assign new_new_n40019__ = new_new_n39629__ & ~new_new_n40018__;
  assign ys__n30277 = new_new_n39993__ | new_new_n40019__;
  assign new_new_n40021__ = ys__n352 & ys__n23300;
  assign new_new_n40022__ = new_new_n14002__ & new_new_n40021__;
  assign new_new_n40023__ = ys__n17822 & new_new_n39597__;
  assign new_new_n40024__ = new_new_n38401__ & new_new_n39966__;
  assign new_new_n40025__ = new_new_n38404__ & new_new_n40024__;
  assign new_new_n40026__ = ~new_new_n38404__ & ~new_new_n40024__;
  assign new_new_n40027__ = ~new_new_n40025__ & ~new_new_n40026__;
  assign new_new_n40028__ = new_new_n39602__ & ~new_new_n40027__;
  assign new_new_n40029__ = ~ys__n17824 & new_new_n40000__;
  assign new_new_n40030__ = ys__n17825 & new_new_n40029__;
  assign new_new_n40031__ = ~ys__n17825 & ~new_new_n40029__;
  assign new_new_n40032__ = ~new_new_n40030__ & ~new_new_n40031__;
  assign new_new_n40033__ = new_new_n39669__ & ~new_new_n40032__;
  assign new_new_n40034__ = ~new_new_n40028__ & ~new_new_n40033__;
  assign new_new_n40035__ = ~new_new_n40023__ & new_new_n40034__;
  assign new_new_n40036__ = ~new_new_n39384__ & new_new_n40007__;
  assign new_new_n40037__ = new_new_n39351__ & new_new_n40036__;
  assign new_new_n40038__ = ~new_new_n39351__ & ~new_new_n40036__;
  assign new_new_n40039__ = ~new_new_n40037__ & ~new_new_n40038__;
  assign new_new_n40040__ = new_new_n39615__ & ~new_new_n40039__;
  assign new_new_n40041__ = ~new_new_n39023__ & new_new_n40012__;
  assign new_new_n40042__ = new_new_n38990__ & new_new_n40041__;
  assign new_new_n40043__ = ~new_new_n38990__ & ~new_new_n40041__;
  assign new_new_n40044__ = ~new_new_n40042__ & ~new_new_n40043__;
  assign new_new_n40045__ = new_new_n39621__ & ~new_new_n40044__;
  assign new_new_n40046__ = ~new_new_n40040__ & ~new_new_n40045__;
  assign new_new_n40047__ = new_new_n40035__ & new_new_n40046__;
  assign new_new_n40048__ = new_new_n39629__ & ~new_new_n40047__;
  assign ys__n30280 = new_new_n40022__ | new_new_n40048__;
  assign new_new_n40050__ = ys__n352 & ys__n23302;
  assign new_new_n40051__ = new_new_n14002__ & new_new_n40050__;
  assign new_new_n40052__ = ys__n17824 & new_new_n39597__;
  assign new_new_n40053__ = ~new_new_n38404__ & new_new_n40024__;
  assign new_new_n40054__ = new_new_n38371__ & new_new_n40053__;
  assign new_new_n40055__ = ~new_new_n38371__ & ~new_new_n40053__;
  assign new_new_n40056__ = ~new_new_n40054__ & ~new_new_n40055__;
  assign new_new_n40057__ = new_new_n39602__ & ~new_new_n40056__;
  assign new_new_n40058__ = ys__n17827 & new_new_n16686__;
  assign new_new_n40059__ = ~ys__n17827 & ~new_new_n16686__;
  assign new_new_n40060__ = ~new_new_n40058__ & ~new_new_n40059__;
  assign new_new_n40061__ = new_new_n39669__ & ~new_new_n40060__;
  assign new_new_n40062__ = ~new_new_n40057__ & ~new_new_n40061__;
  assign new_new_n40063__ = ~new_new_n40052__ & new_new_n40062__;
  assign new_new_n40064__ = ~new_new_n38212__ & new_new_n39432__;
  assign new_new_n40065__ = new_new_n38212__ & ~new_new_n39432__;
  assign new_new_n40066__ = ~new_new_n40064__ & ~new_new_n40065__;
  assign new_new_n40067__ = new_new_n39615__ & ~new_new_n40066__;
  assign new_new_n40068__ = new_new_n39070__ & ~new_new_n39254__;
  assign new_new_n40069__ = ~new_new_n39070__ & new_new_n39254__;
  assign new_new_n40070__ = ~new_new_n40068__ & ~new_new_n40069__;
  assign new_new_n40071__ = new_new_n39621__ & ~new_new_n40070__;
  assign new_new_n40072__ = ~new_new_n40067__ & ~new_new_n40071__;
  assign new_new_n40073__ = new_new_n40063__ & new_new_n40072__;
  assign new_new_n40074__ = new_new_n39629__ & ~new_new_n40073__;
  assign ys__n30283 = new_new_n40051__ | new_new_n40074__;
  assign new_new_n40076__ = ys__n352 & ys__n23304;
  assign new_new_n40077__ = new_new_n14002__ & new_new_n40076__;
  assign new_new_n40078__ = ys__n17825 & new_new_n39597__;
  assign new_new_n40079__ = new_new_n38451__ & ~new_new_n38825__;
  assign new_new_n40080__ = ~new_new_n38451__ & new_new_n38825__;
  assign new_new_n40081__ = ~new_new_n40079__ & ~new_new_n40080__;
  assign new_new_n40082__ = new_new_n39602__ & ~new_new_n40081__;
  assign new_new_n40083__ = ~ys__n17827 & new_new_n16686__;
  assign new_new_n40084__ = ys__n17828 & new_new_n40083__;
  assign new_new_n40085__ = ~ys__n17828 & ~new_new_n40083__;
  assign new_new_n40086__ = ~new_new_n40084__ & ~new_new_n40085__;
  assign new_new_n40087__ = new_new_n39669__ & ~new_new_n40086__;
  assign new_new_n40088__ = ~new_new_n40082__ & ~new_new_n40087__;
  assign new_new_n40089__ = ~new_new_n40078__ & new_new_n40088__;
  assign new_new_n40090__ = new_new_n39432__ & ~new_new_n39565__;
  assign new_new_n40091__ = ~new_new_n38212__ & new_new_n39565__;
  assign new_new_n40092__ = new_new_n38212__ & ~new_new_n39565__;
  assign new_new_n40093__ = ~new_new_n40091__ & ~new_new_n40092__;
  assign new_new_n40094__ = ~new_new_n39432__ & ~new_new_n40093__;
  assign new_new_n40095__ = ~new_new_n40090__ & ~new_new_n40094__;
  assign new_new_n40096__ = new_new_n39615__ & ~new_new_n40095__;
  assign new_new_n40097__ = new_new_n39070__ & ~new_new_n39251__;
  assign new_new_n40098__ = new_new_n39251__ & ~new_new_n39254__;
  assign new_new_n40099__ = ~new_new_n39251__ & new_new_n39254__;
  assign new_new_n40100__ = ~new_new_n40098__ & ~new_new_n40099__;
  assign new_new_n40101__ = ~new_new_n39070__ & ~new_new_n40100__;
  assign new_new_n40102__ = ~new_new_n40097__ & ~new_new_n40101__;
  assign new_new_n40103__ = new_new_n39621__ & ~new_new_n40102__;
  assign new_new_n40104__ = ~new_new_n40096__ & ~new_new_n40103__;
  assign new_new_n40105__ = new_new_n40089__ & new_new_n40104__;
  assign new_new_n40106__ = new_new_n39629__ & ~new_new_n40105__;
  assign ys__n30286 = new_new_n40077__ | new_new_n40106__;
  assign new_new_n40108__ = ys__n352 & ys__n23306;
  assign new_new_n40109__ = new_new_n14002__ & new_new_n40108__;
  assign new_new_n40110__ = ys__n17827 & new_new_n39597__;
  assign new_new_n40111__ = new_new_n38451__ & ~new_new_n38822__;
  assign new_new_n40112__ = new_new_n38822__ & ~new_new_n38825__;
  assign new_new_n40113__ = ~new_new_n38822__ & new_new_n38825__;
  assign new_new_n40114__ = ~new_new_n40112__ & ~new_new_n40113__;
  assign new_new_n40115__ = ~new_new_n38451__ & ~new_new_n40114__;
  assign new_new_n40116__ = ~new_new_n40111__ & ~new_new_n40115__;
  assign new_new_n40117__ = new_new_n39602__ & ~new_new_n40116__;
  assign new_new_n40118__ = new_new_n16656__ & new_new_n16686__;
  assign new_new_n40119__ = ys__n17830 & new_new_n40118__;
  assign new_new_n40120__ = ~ys__n17830 & ~new_new_n40118__;
  assign new_new_n40121__ = ~new_new_n40119__ & ~new_new_n40120__;
  assign new_new_n40122__ = new_new_n39669__ & ~new_new_n40121__;
  assign new_new_n40123__ = ~new_new_n40117__ & ~new_new_n40122__;
  assign new_new_n40124__ = ~new_new_n40110__ & new_new_n40123__;
  assign new_new_n40125__ = new_new_n39432__ & ~new_new_n39562__;
  assign new_new_n40126__ = new_new_n39562__ & new_new_n39566__;
  assign new_new_n40127__ = ~new_new_n39562__ & ~new_new_n39566__;
  assign new_new_n40128__ = ~new_new_n40126__ & ~new_new_n40127__;
  assign new_new_n40129__ = ~new_new_n39432__ & ~new_new_n40128__;
  assign new_new_n40130__ = ~new_new_n40125__ & ~new_new_n40129__;
  assign new_new_n40131__ = new_new_n39615__ & ~new_new_n40130__;
  assign new_new_n40132__ = new_new_n39070__ & ~new_new_n39248__;
  assign new_new_n40133__ = new_new_n39248__ & new_new_n39255__;
  assign new_new_n40134__ = ~new_new_n39248__ & ~new_new_n39255__;
  assign new_new_n40135__ = ~new_new_n40133__ & ~new_new_n40134__;
  assign new_new_n40136__ = ~new_new_n39070__ & ~new_new_n40135__;
  assign new_new_n40137__ = ~new_new_n40132__ & ~new_new_n40136__;
  assign new_new_n40138__ = new_new_n39621__ & ~new_new_n40137__;
  assign new_new_n40139__ = ~new_new_n40131__ & ~new_new_n40138__;
  assign new_new_n40140__ = new_new_n40124__ & new_new_n40139__;
  assign new_new_n40141__ = new_new_n39629__ & ~new_new_n40140__;
  assign ys__n30289 = new_new_n40109__ | new_new_n40141__;
  assign new_new_n40143__ = ys__n352 & ys__n23308;
  assign new_new_n40144__ = new_new_n14002__ & new_new_n40143__;
  assign new_new_n40145__ = ys__n17828 & new_new_n39597__;
  assign new_new_n40146__ = new_new_n38451__ & ~new_new_n38819__;
  assign new_new_n40147__ = new_new_n38819__ & new_new_n38826__;
  assign new_new_n40148__ = ~new_new_n38819__ & ~new_new_n38826__;
  assign new_new_n40149__ = ~new_new_n40147__ & ~new_new_n40148__;
  assign new_new_n40150__ = ~new_new_n38451__ & ~new_new_n40149__;
  assign new_new_n40151__ = ~new_new_n40146__ & ~new_new_n40150__;
  assign new_new_n40152__ = new_new_n39602__ & ~new_new_n40151__;
  assign new_new_n40153__ = ~ys__n17830 & new_new_n40118__;
  assign new_new_n40154__ = ys__n17831 & new_new_n40153__;
  assign new_new_n40155__ = ~ys__n17831 & ~new_new_n40153__;
  assign new_new_n40156__ = ~new_new_n40154__ & ~new_new_n40155__;
  assign new_new_n40157__ = new_new_n39669__ & ~new_new_n40156__;
  assign new_new_n40158__ = ~new_new_n40152__ & ~new_new_n40157__;
  assign new_new_n40159__ = ~new_new_n40145__ & new_new_n40158__;
  assign new_new_n40160__ = new_new_n39432__ & ~new_new_n39559__;
  assign new_new_n40161__ = new_new_n39559__ & new_new_n39567__;
  assign new_new_n40162__ = ~new_new_n39559__ & ~new_new_n39567__;
  assign new_new_n40163__ = ~new_new_n40161__ & ~new_new_n40162__;
  assign new_new_n40164__ = ~new_new_n39432__ & ~new_new_n40163__;
  assign new_new_n40165__ = ~new_new_n40160__ & ~new_new_n40164__;
  assign new_new_n40166__ = new_new_n39615__ & ~new_new_n40165__;
  assign new_new_n40167__ = new_new_n39070__ & ~new_new_n39245__;
  assign new_new_n40168__ = new_new_n39245__ & new_new_n39256__;
  assign new_new_n40169__ = ~new_new_n39245__ & ~new_new_n39256__;
  assign new_new_n40170__ = ~new_new_n40168__ & ~new_new_n40169__;
  assign new_new_n40171__ = ~new_new_n39070__ & ~new_new_n40170__;
  assign new_new_n40172__ = ~new_new_n40167__ & ~new_new_n40171__;
  assign new_new_n40173__ = new_new_n39621__ & ~new_new_n40172__;
  assign new_new_n40174__ = ~new_new_n40166__ & ~new_new_n40173__;
  assign new_new_n40175__ = new_new_n40159__ & new_new_n40174__;
  assign new_new_n40176__ = new_new_n39629__ & ~new_new_n40175__;
  assign ys__n30292 = new_new_n40144__ | new_new_n40176__;
  assign new_new_n40178__ = ys__n352 & ys__n23310;
  assign new_new_n40179__ = new_new_n14002__ & new_new_n40178__;
  assign new_new_n40180__ = ys__n17830 & new_new_n39597__;
  assign new_new_n40181__ = new_new_n38451__ & ~new_new_n38816__;
  assign new_new_n40182__ = new_new_n38816__ & new_new_n38827__;
  assign new_new_n40183__ = ~new_new_n38816__ & ~new_new_n38827__;
  assign new_new_n40184__ = ~new_new_n40182__ & ~new_new_n40183__;
  assign new_new_n40185__ = ~new_new_n38451__ & ~new_new_n40184__;
  assign new_new_n40186__ = ~new_new_n40181__ & ~new_new_n40185__;
  assign new_new_n40187__ = new_new_n39602__ & ~new_new_n40186__;
  assign new_new_n40188__ = new_new_n16658__ & new_new_n16686__;
  assign new_new_n40189__ = ys__n17833 & new_new_n40188__;
  assign new_new_n40190__ = ~ys__n17833 & ~new_new_n40188__;
  assign new_new_n40191__ = ~new_new_n40189__ & ~new_new_n40190__;
  assign new_new_n40192__ = new_new_n39669__ & ~new_new_n40191__;
  assign new_new_n40193__ = ~new_new_n40187__ & ~new_new_n40192__;
  assign new_new_n40194__ = ~new_new_n40180__ & new_new_n40193__;
  assign new_new_n40195__ = new_new_n39432__ & ~new_new_n39550__;
  assign new_new_n40196__ = new_new_n39550__ & new_new_n39568__;
  assign new_new_n40197__ = ~new_new_n39550__ & ~new_new_n39568__;
  assign new_new_n40198__ = ~new_new_n40196__ & ~new_new_n40197__;
  assign new_new_n40199__ = ~new_new_n39432__ & ~new_new_n40198__;
  assign new_new_n40200__ = ~new_new_n40195__ & ~new_new_n40199__;
  assign new_new_n40201__ = new_new_n39615__ & ~new_new_n40200__;
  assign new_new_n40202__ = new_new_n39070__ & ~new_new_n39236__;
  assign new_new_n40203__ = new_new_n39236__ & new_new_n39257__;
  assign new_new_n40204__ = ~new_new_n39236__ & ~new_new_n39257__;
  assign new_new_n40205__ = ~new_new_n40203__ & ~new_new_n40204__;
  assign new_new_n40206__ = ~new_new_n39070__ & ~new_new_n40205__;
  assign new_new_n40207__ = ~new_new_n40202__ & ~new_new_n40206__;
  assign new_new_n40208__ = new_new_n39621__ & ~new_new_n40207__;
  assign new_new_n40209__ = ~new_new_n40201__ & ~new_new_n40208__;
  assign new_new_n40210__ = new_new_n40194__ & new_new_n40209__;
  assign new_new_n40211__ = new_new_n39629__ & ~new_new_n40210__;
  assign ys__n30295 = new_new_n40179__ | new_new_n40211__;
  assign new_new_n40213__ = ys__n352 & ys__n23312;
  assign new_new_n40214__ = new_new_n14002__ & new_new_n40213__;
  assign new_new_n40215__ = ys__n17831 & new_new_n39597__;
  assign new_new_n40216__ = new_new_n38451__ & ~new_new_n38807__;
  assign new_new_n40217__ = new_new_n38807__ & new_new_n38828__;
  assign new_new_n40218__ = ~new_new_n38807__ & ~new_new_n38828__;
  assign new_new_n40219__ = ~new_new_n40217__ & ~new_new_n40218__;
  assign new_new_n40220__ = ~new_new_n38451__ & ~new_new_n40219__;
  assign new_new_n40221__ = ~new_new_n40216__ & ~new_new_n40220__;
  assign new_new_n40222__ = new_new_n39602__ & ~new_new_n40221__;
  assign new_new_n40223__ = ~ys__n17833 & new_new_n40188__;
  assign new_new_n40224__ = ys__n17834 & new_new_n40223__;
  assign new_new_n40225__ = ~ys__n17834 & ~new_new_n40223__;
  assign new_new_n40226__ = ~new_new_n40224__ & ~new_new_n40225__;
  assign new_new_n40227__ = new_new_n39669__ & ~new_new_n40226__;
  assign new_new_n40228__ = ~new_new_n40222__ & ~new_new_n40227__;
  assign new_new_n40229__ = ~new_new_n40215__ & new_new_n40228__;
  assign new_new_n40230__ = new_new_n39432__ & ~new_new_n39547__;
  assign new_new_n40231__ = ~new_new_n39550__ & new_new_n39568__;
  assign new_new_n40232__ = new_new_n39547__ & new_new_n40231__;
  assign new_new_n40233__ = ~new_new_n39547__ & ~new_new_n40231__;
  assign new_new_n40234__ = ~new_new_n40232__ & ~new_new_n40233__;
  assign new_new_n40235__ = ~new_new_n39432__ & ~new_new_n40234__;
  assign new_new_n40236__ = ~new_new_n40230__ & ~new_new_n40235__;
  assign new_new_n40237__ = new_new_n39615__ & ~new_new_n40236__;
  assign new_new_n40238__ = new_new_n39070__ & ~new_new_n39233__;
  assign new_new_n40239__ = ~new_new_n39236__ & new_new_n39257__;
  assign new_new_n40240__ = new_new_n39233__ & new_new_n40239__;
  assign new_new_n40241__ = ~new_new_n39233__ & ~new_new_n40239__;
  assign new_new_n40242__ = ~new_new_n40240__ & ~new_new_n40241__;
  assign new_new_n40243__ = ~new_new_n39070__ & ~new_new_n40242__;
  assign new_new_n40244__ = ~new_new_n40238__ & ~new_new_n40243__;
  assign new_new_n40245__ = new_new_n39621__ & ~new_new_n40244__;
  assign new_new_n40246__ = ~new_new_n40237__ & ~new_new_n40245__;
  assign new_new_n40247__ = new_new_n40229__ & new_new_n40246__;
  assign new_new_n40248__ = new_new_n39629__ & ~new_new_n40247__;
  assign ys__n30298 = new_new_n40214__ | new_new_n40248__;
  assign new_new_n40250__ = ys__n352 & ys__n23314;
  assign new_new_n40251__ = new_new_n14002__ & new_new_n40250__;
  assign new_new_n40252__ = ys__n17833 & new_new_n39597__;
  assign new_new_n40253__ = new_new_n38451__ & ~new_new_n38804__;
  assign new_new_n40254__ = ~new_new_n38807__ & new_new_n38828__;
  assign new_new_n40255__ = new_new_n38804__ & new_new_n40254__;
  assign new_new_n40256__ = ~new_new_n38804__ & ~new_new_n40254__;
  assign new_new_n40257__ = ~new_new_n40255__ & ~new_new_n40256__;
  assign new_new_n40258__ = ~new_new_n38451__ & ~new_new_n40257__;
  assign new_new_n40259__ = ~new_new_n40253__ & ~new_new_n40258__;
  assign new_new_n40260__ = new_new_n39602__ & ~new_new_n40259__;
  assign new_new_n40261__ = new_new_n16659__ & new_new_n40188__;
  assign new_new_n40262__ = ys__n17836 & new_new_n40261__;
  assign new_new_n40263__ = ~ys__n17836 & ~new_new_n40261__;
  assign new_new_n40264__ = ~new_new_n40262__ & ~new_new_n40263__;
  assign new_new_n40265__ = new_new_n39669__ & ~new_new_n40264__;
  assign new_new_n40266__ = ~new_new_n40260__ & ~new_new_n40265__;
  assign new_new_n40267__ = ~new_new_n40252__ & new_new_n40266__;
  assign new_new_n40268__ = new_new_n39432__ & ~new_new_n39554__;
  assign new_new_n40269__ = new_new_n39551__ & new_new_n39568__;
  assign new_new_n40270__ = new_new_n39554__ & new_new_n40269__;
  assign new_new_n40271__ = ~new_new_n39554__ & ~new_new_n40269__;
  assign new_new_n40272__ = ~new_new_n40270__ & ~new_new_n40271__;
  assign new_new_n40273__ = ~new_new_n39432__ & ~new_new_n40272__;
  assign new_new_n40274__ = ~new_new_n40268__ & ~new_new_n40273__;
  assign new_new_n40275__ = new_new_n39615__ & ~new_new_n40274__;
  assign new_new_n40276__ = new_new_n39070__ & ~new_new_n39240__;
  assign new_new_n40277__ = new_new_n39237__ & new_new_n39257__;
  assign new_new_n40278__ = new_new_n39240__ & new_new_n40277__;
  assign new_new_n40279__ = ~new_new_n39240__ & ~new_new_n40277__;
  assign new_new_n40280__ = ~new_new_n40278__ & ~new_new_n40279__;
  assign new_new_n40281__ = ~new_new_n39070__ & ~new_new_n40280__;
  assign new_new_n40282__ = ~new_new_n40276__ & ~new_new_n40281__;
  assign new_new_n40283__ = new_new_n39621__ & ~new_new_n40282__;
  assign new_new_n40284__ = ~new_new_n40275__ & ~new_new_n40283__;
  assign new_new_n40285__ = new_new_n40267__ & new_new_n40284__;
  assign new_new_n40286__ = new_new_n39629__ & ~new_new_n40285__;
  assign ys__n30301 = new_new_n40251__ | new_new_n40286__;
  assign new_new_n40288__ = ys__n352 & ys__n23316;
  assign new_new_n40289__ = new_new_n14002__ & new_new_n40288__;
  assign new_new_n40290__ = ys__n17834 & new_new_n39597__;
  assign new_new_n40291__ = new_new_n38451__ & ~new_new_n38811__;
  assign new_new_n40292__ = new_new_n38808__ & new_new_n38828__;
  assign new_new_n40293__ = new_new_n38811__ & new_new_n40292__;
  assign new_new_n40294__ = ~new_new_n38811__ & ~new_new_n40292__;
  assign new_new_n40295__ = ~new_new_n40293__ & ~new_new_n40294__;
  assign new_new_n40296__ = ~new_new_n38451__ & ~new_new_n40295__;
  assign new_new_n40297__ = ~new_new_n40291__ & ~new_new_n40296__;
  assign new_new_n40298__ = new_new_n39602__ & ~new_new_n40297__;
  assign new_new_n40299__ = ~ys__n17836 & new_new_n40261__;
  assign new_new_n40300__ = ys__n17837 & new_new_n40299__;
  assign new_new_n40301__ = ~ys__n17837 & ~new_new_n40299__;
  assign new_new_n40302__ = ~new_new_n40300__ & ~new_new_n40301__;
  assign new_new_n40303__ = new_new_n39669__ & ~new_new_n40302__;
  assign new_new_n40304__ = ~new_new_n40298__ & ~new_new_n40303__;
  assign new_new_n40305__ = ~new_new_n40290__ & new_new_n40304__;
  assign new_new_n40306__ = new_new_n39432__ & ~new_new_n39542__;
  assign new_new_n40307__ = ~new_new_n39554__ & new_new_n40269__;
  assign new_new_n40308__ = new_new_n39542__ & new_new_n40307__;
  assign new_new_n40309__ = ~new_new_n39542__ & ~new_new_n40307__;
  assign new_new_n40310__ = ~new_new_n40308__ & ~new_new_n40309__;
  assign new_new_n40311__ = ~new_new_n39432__ & ~new_new_n40310__;
  assign new_new_n40312__ = ~new_new_n40306__ & ~new_new_n40311__;
  assign new_new_n40313__ = new_new_n39615__ & ~new_new_n40312__;
  assign new_new_n40314__ = new_new_n39070__ & ~new_new_n39228__;
  assign new_new_n40315__ = ~new_new_n39240__ & new_new_n40277__;
  assign new_new_n40316__ = new_new_n39228__ & new_new_n40315__;
  assign new_new_n40317__ = ~new_new_n39228__ & ~new_new_n40315__;
  assign new_new_n40318__ = ~new_new_n40316__ & ~new_new_n40317__;
  assign new_new_n40319__ = ~new_new_n39070__ & ~new_new_n40318__;
  assign new_new_n40320__ = ~new_new_n40314__ & ~new_new_n40319__;
  assign new_new_n40321__ = new_new_n39621__ & ~new_new_n40320__;
  assign new_new_n40322__ = ~new_new_n40313__ & ~new_new_n40321__;
  assign new_new_n40323__ = new_new_n40305__ & new_new_n40322__;
  assign new_new_n40324__ = new_new_n39629__ & ~new_new_n40323__;
  assign ys__n30304 = new_new_n40289__ | new_new_n40324__;
  assign new_new_n40326__ = ys__n352 & ys__n23318;
  assign new_new_n40327__ = new_new_n14002__ & new_new_n40326__;
  assign new_new_n40328__ = ys__n17836 & new_new_n39597__;
  assign new_new_n40329__ = new_new_n38451__ & ~new_new_n38799__;
  assign new_new_n40330__ = ~new_new_n38811__ & new_new_n40292__;
  assign new_new_n40331__ = new_new_n38799__ & new_new_n40330__;
  assign new_new_n40332__ = ~new_new_n38799__ & ~new_new_n40330__;
  assign new_new_n40333__ = ~new_new_n40331__ & ~new_new_n40332__;
  assign new_new_n40334__ = ~new_new_n38451__ & ~new_new_n40333__;
  assign new_new_n40335__ = ~new_new_n40329__ & ~new_new_n40334__;
  assign new_new_n40336__ = new_new_n39602__ & ~new_new_n40335__;
  assign new_new_n40337__ = new_new_n16662__ & new_new_n16686__;
  assign new_new_n40338__ = ys__n17839 & new_new_n40337__;
  assign new_new_n40339__ = ~ys__n17839 & ~new_new_n40337__;
  assign new_new_n40340__ = ~new_new_n40338__ & ~new_new_n40339__;
  assign new_new_n40341__ = new_new_n39669__ & ~new_new_n40340__;
  assign new_new_n40342__ = ~new_new_n40336__ & ~new_new_n40341__;
  assign new_new_n40343__ = ~new_new_n40328__ & new_new_n40342__;
  assign new_new_n40344__ = new_new_n39432__ & ~new_new_n39520__;
  assign new_new_n40345__ = new_new_n39520__ & new_new_n39571__;
  assign new_new_n40346__ = ~new_new_n39520__ & ~new_new_n39571__;
  assign new_new_n40347__ = ~new_new_n40345__ & ~new_new_n40346__;
  assign new_new_n40348__ = ~new_new_n39432__ & ~new_new_n40347__;
  assign new_new_n40349__ = ~new_new_n40344__ & ~new_new_n40348__;
  assign new_new_n40350__ = new_new_n39615__ & ~new_new_n40349__;
  assign new_new_n40351__ = new_new_n39070__ & ~new_new_n39206__;
  assign new_new_n40352__ = new_new_n39206__ & new_new_n39260__;
  assign new_new_n40353__ = ~new_new_n39206__ & ~new_new_n39260__;
  assign new_new_n40354__ = ~new_new_n40352__ & ~new_new_n40353__;
  assign new_new_n40355__ = ~new_new_n39070__ & ~new_new_n40354__;
  assign new_new_n40356__ = ~new_new_n40351__ & ~new_new_n40355__;
  assign new_new_n40357__ = new_new_n39621__ & ~new_new_n40356__;
  assign new_new_n40358__ = ~new_new_n40350__ & ~new_new_n40357__;
  assign new_new_n40359__ = new_new_n40343__ & new_new_n40358__;
  assign new_new_n40360__ = new_new_n39629__ & ~new_new_n40359__;
  assign ys__n30307 = new_new_n40327__ | new_new_n40360__;
  assign new_new_n40362__ = ys__n352 & ys__n23320;
  assign new_new_n40363__ = new_new_n14002__ & new_new_n40362__;
  assign new_new_n40364__ = ys__n17837 & new_new_n39597__;
  assign new_new_n40365__ = new_new_n38451__ & ~new_new_n38789__;
  assign new_new_n40366__ = new_new_n38789__ & new_new_n38831__;
  assign new_new_n40367__ = ~new_new_n38789__ & ~new_new_n38831__;
  assign new_new_n40368__ = ~new_new_n40366__ & ~new_new_n40367__;
  assign new_new_n40369__ = ~new_new_n38451__ & ~new_new_n40368__;
  assign new_new_n40370__ = ~new_new_n40365__ & ~new_new_n40369__;
  assign new_new_n40371__ = new_new_n39602__ & ~new_new_n40370__;
  assign new_new_n40372__ = ~ys__n17839 & new_new_n40337__;
  assign new_new_n40373__ = ys__n17840 & new_new_n40372__;
  assign new_new_n40374__ = ~ys__n17840 & ~new_new_n40372__;
  assign new_new_n40375__ = ~new_new_n40373__ & ~new_new_n40374__;
  assign new_new_n40376__ = new_new_n39669__ & ~new_new_n40375__;
  assign new_new_n40377__ = ~new_new_n40371__ & ~new_new_n40376__;
  assign new_new_n40378__ = ~new_new_n40364__ & new_new_n40377__;
  assign new_new_n40379__ = new_new_n39432__ & ~new_new_n39517__;
  assign new_new_n40380__ = ~new_new_n39520__ & new_new_n39571__;
  assign new_new_n40381__ = new_new_n39517__ & new_new_n40380__;
  assign new_new_n40382__ = ~new_new_n39517__ & ~new_new_n40380__;
  assign new_new_n40383__ = ~new_new_n40381__ & ~new_new_n40382__;
  assign new_new_n40384__ = ~new_new_n39432__ & ~new_new_n40383__;
  assign new_new_n40385__ = ~new_new_n40379__ & ~new_new_n40384__;
  assign new_new_n40386__ = new_new_n39615__ & ~new_new_n40385__;
  assign new_new_n40387__ = new_new_n39070__ & ~new_new_n39203__;
  assign new_new_n40388__ = ~new_new_n39206__ & new_new_n39260__;
  assign new_new_n40389__ = new_new_n39203__ & new_new_n40388__;
  assign new_new_n40390__ = ~new_new_n39203__ & ~new_new_n40388__;
  assign new_new_n40391__ = ~new_new_n40389__ & ~new_new_n40390__;
  assign new_new_n40392__ = ~new_new_n39070__ & ~new_new_n40391__;
  assign new_new_n40393__ = ~new_new_n40387__ & ~new_new_n40392__;
  assign new_new_n40394__ = new_new_n39621__ & ~new_new_n40393__;
  assign new_new_n40395__ = ~new_new_n40386__ & ~new_new_n40394__;
  assign new_new_n40396__ = new_new_n40378__ & new_new_n40395__;
  assign new_new_n40397__ = new_new_n39629__ & ~new_new_n40396__;
  assign ys__n30310 = new_new_n40363__ | new_new_n40397__;
  assign new_new_n40399__ = ys__n352 & ys__n23322;
  assign new_new_n40400__ = new_new_n14002__ & new_new_n40399__;
  assign new_new_n40401__ = ys__n17839 & new_new_n39597__;
  assign new_new_n40402__ = new_new_n38451__ & ~new_new_n38786__;
  assign new_new_n40403__ = ~new_new_n38789__ & new_new_n38831__;
  assign new_new_n40404__ = new_new_n38786__ & new_new_n40403__;
  assign new_new_n40405__ = ~new_new_n38786__ & ~new_new_n40403__;
  assign new_new_n40406__ = ~new_new_n40404__ & ~new_new_n40405__;
  assign new_new_n40407__ = ~new_new_n38451__ & ~new_new_n40406__;
  assign new_new_n40408__ = ~new_new_n40402__ & ~new_new_n40407__;
  assign new_new_n40409__ = new_new_n39602__ & ~new_new_n40408__;
  assign new_new_n40410__ = new_new_n16694__ & new_new_n40337__;
  assign new_new_n40411__ = ys__n17842 & new_new_n40410__;
  assign new_new_n40412__ = ~ys__n17842 & ~new_new_n40410__;
  assign new_new_n40413__ = ~new_new_n40411__ & ~new_new_n40412__;
  assign new_new_n40414__ = new_new_n39669__ & ~new_new_n40413__;
  assign new_new_n40415__ = ~new_new_n40409__ & ~new_new_n40414__;
  assign new_new_n40416__ = ~new_new_n40401__ & new_new_n40415__;
  assign new_new_n40417__ = new_new_n39432__ & ~new_new_n39512__;
  assign new_new_n40418__ = new_new_n39521__ & new_new_n39571__;
  assign new_new_n40419__ = new_new_n39512__ & new_new_n40418__;
  assign new_new_n40420__ = ~new_new_n39512__ & ~new_new_n40418__;
  assign new_new_n40421__ = ~new_new_n40419__ & ~new_new_n40420__;
  assign new_new_n40422__ = ~new_new_n39432__ & ~new_new_n40421__;
  assign new_new_n40423__ = ~new_new_n40417__ & ~new_new_n40422__;
  assign new_new_n40424__ = new_new_n39615__ & ~new_new_n40423__;
  assign new_new_n40425__ = new_new_n39070__ & ~new_new_n39198__;
  assign new_new_n40426__ = new_new_n39207__ & new_new_n39260__;
  assign new_new_n40427__ = new_new_n39198__ & new_new_n40426__;
  assign new_new_n40428__ = ~new_new_n39198__ & ~new_new_n40426__;
  assign new_new_n40429__ = ~new_new_n40427__ & ~new_new_n40428__;
  assign new_new_n40430__ = ~new_new_n39070__ & ~new_new_n40429__;
  assign new_new_n40431__ = ~new_new_n40425__ & ~new_new_n40430__;
  assign new_new_n40432__ = new_new_n39621__ & ~new_new_n40431__;
  assign new_new_n40433__ = ~new_new_n40424__ & ~new_new_n40432__;
  assign new_new_n40434__ = new_new_n40416__ & new_new_n40433__;
  assign new_new_n40435__ = new_new_n39629__ & ~new_new_n40434__;
  assign ys__n30313 = new_new_n40400__ | new_new_n40435__;
  assign new_new_n40437__ = ys__n352 & ys__n23324;
  assign new_new_n40438__ = new_new_n14002__ & new_new_n40437__;
  assign new_new_n40439__ = ys__n17840 & new_new_n39597__;
  assign new_new_n40440__ = new_new_n38451__ & ~new_new_n38781__;
  assign new_new_n40441__ = new_new_n38790__ & new_new_n38831__;
  assign new_new_n40442__ = new_new_n38781__ & new_new_n40441__;
  assign new_new_n40443__ = ~new_new_n38781__ & ~new_new_n40441__;
  assign new_new_n40444__ = ~new_new_n40442__ & ~new_new_n40443__;
  assign new_new_n40445__ = ~new_new_n38451__ & ~new_new_n40444__;
  assign new_new_n40446__ = ~new_new_n40440__ & ~new_new_n40445__;
  assign new_new_n40447__ = new_new_n39602__ & ~new_new_n40446__;
  assign new_new_n40448__ = ~ys__n17842 & new_new_n40410__;
  assign new_new_n40449__ = ys__n17843 & new_new_n40448__;
  assign new_new_n40450__ = ~ys__n17843 & ~new_new_n40448__;
  assign new_new_n40451__ = ~new_new_n40449__ & ~new_new_n40450__;
  assign new_new_n40452__ = new_new_n39669__ & ~new_new_n40451__;
  assign new_new_n40453__ = ~new_new_n40447__ & ~new_new_n40452__;
  assign new_new_n40454__ = ~new_new_n40439__ & new_new_n40453__;
  assign new_new_n40455__ = new_new_n39432__ & ~new_new_n39509__;
  assign new_new_n40456__ = ~new_new_n39512__ & new_new_n40418__;
  assign new_new_n40457__ = new_new_n39509__ & new_new_n40456__;
  assign new_new_n40458__ = ~new_new_n39509__ & ~new_new_n40456__;
  assign new_new_n40459__ = ~new_new_n40457__ & ~new_new_n40458__;
  assign new_new_n40460__ = ~new_new_n39432__ & ~new_new_n40459__;
  assign new_new_n40461__ = ~new_new_n40455__ & ~new_new_n40460__;
  assign new_new_n40462__ = new_new_n39615__ & ~new_new_n40461__;
  assign new_new_n40463__ = new_new_n39070__ & ~new_new_n39195__;
  assign new_new_n40464__ = ~new_new_n39198__ & new_new_n40426__;
  assign new_new_n40465__ = new_new_n39195__ & new_new_n40464__;
  assign new_new_n40466__ = ~new_new_n39195__ & ~new_new_n40464__;
  assign new_new_n40467__ = ~new_new_n40465__ & ~new_new_n40466__;
  assign new_new_n40468__ = ~new_new_n39070__ & ~new_new_n40467__;
  assign new_new_n40469__ = ~new_new_n40463__ & ~new_new_n40468__;
  assign new_new_n40470__ = new_new_n39621__ & ~new_new_n40469__;
  assign new_new_n40471__ = ~new_new_n40462__ & ~new_new_n40470__;
  assign new_new_n40472__ = new_new_n40454__ & new_new_n40471__;
  assign new_new_n40473__ = new_new_n39629__ & ~new_new_n40472__;
  assign ys__n30316 = new_new_n40438__ | new_new_n40473__;
  assign new_new_n40475__ = ys__n352 & ys__n23326;
  assign new_new_n40476__ = new_new_n14002__ & new_new_n40475__;
  assign new_new_n40477__ = ys__n17842 & new_new_n39597__;
  assign new_new_n40478__ = new_new_n38451__ & ~new_new_n38778__;
  assign new_new_n40479__ = ~new_new_n38781__ & new_new_n40441__;
  assign new_new_n40480__ = new_new_n38778__ & new_new_n40479__;
  assign new_new_n40481__ = ~new_new_n38778__ & ~new_new_n40479__;
  assign new_new_n40482__ = ~new_new_n40480__ & ~new_new_n40481__;
  assign new_new_n40483__ = ~new_new_n38451__ & ~new_new_n40482__;
  assign new_new_n40484__ = ~new_new_n40478__ & ~new_new_n40483__;
  assign new_new_n40485__ = new_new_n39602__ & ~new_new_n40484__;
  assign new_new_n40486__ = new_new_n16696__ & new_new_n40337__;
  assign new_new_n40487__ = ys__n17845 & new_new_n40486__;
  assign new_new_n40488__ = ~ys__n17845 & ~new_new_n40486__;
  assign new_new_n40489__ = ~new_new_n40487__ & ~new_new_n40488__;
  assign new_new_n40490__ = new_new_n39669__ & ~new_new_n40489__;
  assign new_new_n40491__ = ~new_new_n40485__ & ~new_new_n40490__;
  assign new_new_n40492__ = ~new_new_n40477__ & new_new_n40491__;
  assign new_new_n40493__ = new_new_n39432__ & ~new_new_n39531__;
  assign new_new_n40494__ = new_new_n39523__ & new_new_n39571__;
  assign new_new_n40495__ = new_new_n39531__ & new_new_n40494__;
  assign new_new_n40496__ = ~new_new_n39531__ & ~new_new_n40494__;
  assign new_new_n40497__ = ~new_new_n40495__ & ~new_new_n40496__;
  assign new_new_n40498__ = ~new_new_n39432__ & ~new_new_n40497__;
  assign new_new_n40499__ = ~new_new_n40493__ & ~new_new_n40498__;
  assign new_new_n40500__ = new_new_n39615__ & ~new_new_n40499__;
  assign new_new_n40501__ = new_new_n39070__ & ~new_new_n39217__;
  assign new_new_n40502__ = new_new_n39209__ & new_new_n39260__;
  assign new_new_n40503__ = new_new_n39217__ & new_new_n40502__;
  assign new_new_n40504__ = ~new_new_n39217__ & ~new_new_n40502__;
  assign new_new_n40505__ = ~new_new_n40503__ & ~new_new_n40504__;
  assign new_new_n40506__ = ~new_new_n39070__ & ~new_new_n40505__;
  assign new_new_n40507__ = ~new_new_n40501__ & ~new_new_n40506__;
  assign new_new_n40508__ = new_new_n39621__ & ~new_new_n40507__;
  assign new_new_n40509__ = ~new_new_n40500__ & ~new_new_n40508__;
  assign new_new_n40510__ = new_new_n40492__ & new_new_n40509__;
  assign new_new_n40511__ = new_new_n39629__ & ~new_new_n40510__;
  assign ys__n30319 = new_new_n40476__ | new_new_n40511__;
  assign new_new_n40513__ = ys__n352 & ys__n23328;
  assign new_new_n40514__ = new_new_n14002__ & new_new_n40513__;
  assign new_new_n40515__ = ys__n17843 & new_new_n39597__;
  assign new_new_n40516__ = new_new_n38451__ & ~new_new_n38770__;
  assign new_new_n40517__ = new_new_n38770__ & new_new_n38832__;
  assign new_new_n40518__ = ~new_new_n38770__ & ~new_new_n38832__;
  assign new_new_n40519__ = ~new_new_n40517__ & ~new_new_n40518__;
  assign new_new_n40520__ = ~new_new_n38451__ & ~new_new_n40519__;
  assign new_new_n40521__ = ~new_new_n40516__ & ~new_new_n40520__;
  assign new_new_n40522__ = new_new_n39602__ & ~new_new_n40521__;
  assign new_new_n40523__ = ~ys__n17845 & new_new_n40486__;
  assign new_new_n40524__ = ys__n17846 & new_new_n40523__;
  assign new_new_n40525__ = ~ys__n17846 & ~new_new_n40523__;
  assign new_new_n40526__ = ~new_new_n40524__ & ~new_new_n40525__;
  assign new_new_n40527__ = new_new_n39669__ & ~new_new_n40526__;
  assign new_new_n40528__ = ~new_new_n40522__ & ~new_new_n40527__;
  assign new_new_n40529__ = ~new_new_n40515__ & new_new_n40528__;
  assign new_new_n40530__ = new_new_n39432__ & ~new_new_n39528__;
  assign new_new_n40531__ = ~new_new_n39531__ & new_new_n40494__;
  assign new_new_n40532__ = new_new_n39528__ & new_new_n40531__;
  assign new_new_n40533__ = ~new_new_n39528__ & ~new_new_n40531__;
  assign new_new_n40534__ = ~new_new_n40532__ & ~new_new_n40533__;
  assign new_new_n40535__ = ~new_new_n39432__ & ~new_new_n40534__;
  assign new_new_n40536__ = ~new_new_n40530__ & ~new_new_n40535__;
  assign new_new_n40537__ = new_new_n39615__ & ~new_new_n40536__;
  assign new_new_n40538__ = new_new_n39070__ & ~new_new_n39214__;
  assign new_new_n40539__ = ~new_new_n39217__ & new_new_n40502__;
  assign new_new_n40540__ = new_new_n39214__ & new_new_n40539__;
  assign new_new_n40541__ = ~new_new_n39214__ & ~new_new_n40539__;
  assign new_new_n40542__ = ~new_new_n40540__ & ~new_new_n40541__;
  assign new_new_n40543__ = ~new_new_n39070__ & ~new_new_n40542__;
  assign new_new_n40544__ = ~new_new_n40538__ & ~new_new_n40543__;
  assign new_new_n40545__ = new_new_n39621__ & ~new_new_n40544__;
  assign new_new_n40546__ = ~new_new_n40537__ & ~new_new_n40545__;
  assign new_new_n40547__ = new_new_n40529__ & new_new_n40546__;
  assign new_new_n40548__ = new_new_n39629__ & ~new_new_n40547__;
  assign ys__n30322 = new_new_n40514__ | new_new_n40548__;
  assign new_new_n40550__ = ys__n352 & ys__n23330;
  assign new_new_n40551__ = new_new_n14002__ & new_new_n40550__;
  assign new_new_n40552__ = ys__n17845 & new_new_n39597__;
  assign new_new_n40553__ = new_new_n38451__ & ~new_new_n38767__;
  assign new_new_n40554__ = ~new_new_n38770__ & new_new_n38832__;
  assign new_new_n40555__ = new_new_n38767__ & new_new_n40554__;
  assign new_new_n40556__ = ~new_new_n38767__ & ~new_new_n40554__;
  assign new_new_n40557__ = ~new_new_n40555__ & ~new_new_n40556__;
  assign new_new_n40558__ = ~new_new_n38451__ & ~new_new_n40557__;
  assign new_new_n40559__ = ~new_new_n40553__ & ~new_new_n40558__;
  assign new_new_n40560__ = new_new_n39602__ & ~new_new_n40559__;
  assign new_new_n40561__ = new_new_n16666__ & new_new_n40486__;
  assign new_new_n40562__ = ys__n17848 & new_new_n40561__;
  assign new_new_n40563__ = ~ys__n17848 & ~new_new_n40561__;
  assign new_new_n40564__ = ~new_new_n40562__ & ~new_new_n40563__;
  assign new_new_n40565__ = new_new_n39669__ & ~new_new_n40564__;
  assign new_new_n40566__ = ~new_new_n40560__ & ~new_new_n40565__;
  assign new_new_n40567__ = ~new_new_n40552__ & new_new_n40566__;
  assign new_new_n40568__ = new_new_n39432__ & ~new_new_n39535__;
  assign new_new_n40569__ = new_new_n39532__ & new_new_n40494__;
  assign new_new_n40570__ = new_new_n39535__ & new_new_n40569__;
  assign new_new_n40571__ = ~new_new_n39535__ & ~new_new_n40569__;
  assign new_new_n40572__ = ~new_new_n40570__ & ~new_new_n40571__;
  assign new_new_n40573__ = ~new_new_n39432__ & ~new_new_n40572__;
  assign new_new_n40574__ = ~new_new_n40568__ & ~new_new_n40573__;
  assign new_new_n40575__ = new_new_n39615__ & ~new_new_n40574__;
  assign new_new_n40576__ = new_new_n39070__ & ~new_new_n39221__;
  assign new_new_n40577__ = new_new_n39218__ & new_new_n40502__;
  assign new_new_n40578__ = new_new_n39221__ & new_new_n40577__;
  assign new_new_n40579__ = ~new_new_n39221__ & ~new_new_n40577__;
  assign new_new_n40580__ = ~new_new_n40578__ & ~new_new_n40579__;
  assign new_new_n40581__ = ~new_new_n39070__ & ~new_new_n40580__;
  assign new_new_n40582__ = ~new_new_n40576__ & ~new_new_n40581__;
  assign new_new_n40583__ = new_new_n39621__ & ~new_new_n40582__;
  assign new_new_n40584__ = ~new_new_n40575__ & ~new_new_n40583__;
  assign new_new_n40585__ = new_new_n40567__ & new_new_n40584__;
  assign new_new_n40586__ = new_new_n39629__ & ~new_new_n40585__;
  assign ys__n30325 = new_new_n40551__ | new_new_n40586__;
  assign new_new_n40588__ = ys__n352 & ys__n23332;
  assign new_new_n40589__ = new_new_n14002__ & new_new_n40588__;
  assign new_new_n40590__ = ys__n17846 & new_new_n39597__;
  assign new_new_n40591__ = new_new_n38451__ & ~new_new_n38762__;
  assign new_new_n40592__ = new_new_n38762__ & new_new_n38833__;
  assign new_new_n40593__ = ~new_new_n38762__ & ~new_new_n38833__;
  assign new_new_n40594__ = ~new_new_n40592__ & ~new_new_n40593__;
  assign new_new_n40595__ = ~new_new_n38451__ & ~new_new_n40594__;
  assign new_new_n40596__ = ~new_new_n40591__ & ~new_new_n40595__;
  assign new_new_n40597__ = new_new_n39602__ & ~new_new_n40596__;
  assign new_new_n40598__ = ~ys__n17848 & new_new_n40561__;
  assign new_new_n40599__ = ys__n17849 & new_new_n40598__;
  assign new_new_n40600__ = ~ys__n17849 & ~new_new_n40598__;
  assign new_new_n40601__ = ~new_new_n40599__ & ~new_new_n40600__;
  assign new_new_n40602__ = new_new_n39669__ & ~new_new_n40601__;
  assign new_new_n40603__ = ~new_new_n40597__ & ~new_new_n40602__;
  assign new_new_n40604__ = ~new_new_n40590__ & new_new_n40603__;
  assign new_new_n40605__ = new_new_n39432__ & ~new_new_n39502__;
  assign new_new_n40606__ = ~new_new_n39535__ & new_new_n40569__;
  assign new_new_n40607__ = new_new_n39502__ & new_new_n40606__;
  assign new_new_n40608__ = ~new_new_n39502__ & ~new_new_n40606__;
  assign new_new_n40609__ = ~new_new_n40607__ & ~new_new_n40608__;
  assign new_new_n40610__ = ~new_new_n39432__ & ~new_new_n40609__;
  assign new_new_n40611__ = ~new_new_n40605__ & ~new_new_n40610__;
  assign new_new_n40612__ = new_new_n39615__ & ~new_new_n40611__;
  assign new_new_n40613__ = new_new_n39070__ & ~new_new_n39188__;
  assign new_new_n40614__ = ~new_new_n39221__ & new_new_n40577__;
  assign new_new_n40615__ = new_new_n39188__ & new_new_n40614__;
  assign new_new_n40616__ = ~new_new_n39188__ & ~new_new_n40614__;
  assign new_new_n40617__ = ~new_new_n40615__ & ~new_new_n40616__;
  assign new_new_n40618__ = ~new_new_n39070__ & ~new_new_n40617__;
  assign new_new_n40619__ = ~new_new_n40613__ & ~new_new_n40618__;
  assign new_new_n40620__ = new_new_n39621__ & ~new_new_n40619__;
  assign new_new_n40621__ = ~new_new_n40612__ & ~new_new_n40620__;
  assign new_new_n40622__ = new_new_n40604__ & new_new_n40621__;
  assign new_new_n40623__ = new_new_n39629__ & ~new_new_n40622__;
  assign ys__n30328 = new_new_n40589__ | new_new_n40623__;
  assign ys__n30331 = ys__n2652 & ys__n30330;
  assign new_new_n40626__ = ys__n174 & ~ys__n196;
  assign new_new_n40627__ = ys__n2830 & new_new_n40626__;
  assign new_new_n40628__ = new_new_n40021__ & new_new_n40627__;
  assign new_new_n40629__ = ys__n174 & ys__n196;
  assign new_new_n40630__ = ys__n24786 & new_new_n40629__;
  assign new_new_n40631__ = ~ys__n2830 & new_new_n40626__;
  assign new_new_n40632__ = new_new_n40021__ & new_new_n40631__;
  assign new_new_n40633__ = ~new_new_n40630__ & ~new_new_n40632__;
  assign new_new_n40634__ = ~new_new_n40628__ & new_new_n40633__;
  assign new_new_n40635__ = ~ys__n174 & ys__n196;
  assign new_new_n40636__ = ~new_new_n40629__ & ~new_new_n40635__;
  assign new_new_n40637__ = ~new_new_n40631__ & new_new_n40636__;
  assign new_new_n40638__ = ~ys__n196 & ys__n2830;
  assign new_new_n40639__ = ~ys__n174 & new_new_n40638__;
  assign new_new_n40640__ = ~ys__n174 & ~ys__n196;
  assign new_new_n40641__ = ~ys__n2830 & new_new_n40640__;
  assign new_new_n40642__ = ~new_new_n40627__ & ~new_new_n40641__;
  assign new_new_n40643__ = ~new_new_n40639__ & new_new_n40642__;
  assign new_new_n40644__ = new_new_n40637__ & new_new_n40643__;
  assign ys__n33095 = ~new_new_n40634__ & ~new_new_n40644__;
  assign new_new_n40646__ = ys__n24789 & new_new_n40629__;
  assign new_new_n40647__ = new_new_n40050__ & new_new_n40631__;
  assign new_new_n40648__ = ~new_new_n40646__ & ~new_new_n40647__;
  assign new_new_n40649__ = new_new_n38047__ & new_new_n40639__;
  assign new_new_n40650__ = new_new_n38047__ & new_new_n40641__;
  assign new_new_n40651__ = new_new_n40050__ & new_new_n40627__;
  assign new_new_n40652__ = ~new_new_n40650__ & ~new_new_n40651__;
  assign new_new_n40653__ = ~new_new_n40649__ & new_new_n40652__;
  assign new_new_n40654__ = new_new_n40648__ & new_new_n40653__;
  assign ys__n33096 = ~new_new_n40644__ & ~new_new_n40654__;
  assign new_new_n40656__ = ~ys__n33095 & ys__n33096;
  assign new_new_n40657__ = ys__n33095 & ~ys__n33096;
  assign new_new_n40658__ = ~new_new_n40656__ & ~new_new_n40657__;
  assign new_new_n40659__ = new_new_n39659__ & new_new_n40627__;
  assign new_new_n40660__ = ys__n24747 & new_new_n40629__;
  assign new_new_n40661__ = new_new_n39659__ & new_new_n40631__;
  assign new_new_n40662__ = ~new_new_n40660__ & ~new_new_n40661__;
  assign new_new_n40663__ = ~new_new_n40659__ & new_new_n40662__;
  assign ys__n33082 = ~new_new_n40644__ & ~new_new_n40663__;
  assign new_new_n40665__ = new_new_n39632__ & new_new_n40627__;
  assign new_new_n40666__ = ys__n24744 & new_new_n40629__;
  assign new_new_n40667__ = new_new_n39632__ & new_new_n40631__;
  assign new_new_n40668__ = ~new_new_n40666__ & ~new_new_n40667__;
  assign new_new_n40669__ = ~new_new_n40665__ & new_new_n40668__;
  assign ys__n33081 = ~new_new_n40644__ & ~new_new_n40669__;
  assign new_new_n40671__ = ~ys__n33082 & ys__n33081;
  assign new_new_n40672__ = ys__n33082 & ~ys__n33081;
  assign new_new_n40673__ = ~new_new_n40671__ & ~new_new_n40672__;
  assign new_new_n40674__ = new_new_n39685__ & new_new_n40627__;
  assign new_new_n40675__ = ys__n24750 & new_new_n40629__;
  assign new_new_n40676__ = new_new_n39685__ & new_new_n40631__;
  assign new_new_n40677__ = ~new_new_n40675__ & ~new_new_n40676__;
  assign new_new_n40678__ = ~new_new_n40674__ & new_new_n40677__;
  assign ys__n33083 = ~new_new_n40644__ & ~new_new_n40678__;
  assign new_new_n40680__ = ys__n33082 & ~ys__n33083;
  assign new_new_n40681__ = ~ys__n33082 & ys__n33083;
  assign new_new_n40682__ = ~new_new_n40680__ & ~new_new_n40681__;
  assign new_new_n40683__ = new_new_n38047__ & new_new_n40627__;
  assign new_new_n40684__ = ys__n24741 & new_new_n40629__;
  assign new_new_n40685__ = new_new_n38047__ & new_new_n40631__;
  assign new_new_n40686__ = ~new_new_n40684__ & ~new_new_n40685__;
  assign new_new_n40687__ = ~new_new_n40683__ & new_new_n40686__;
  assign ys__n33080 = ~new_new_n40644__ & ~new_new_n40687__;
  assign new_new_n40689__ = ys__n33081 & ys__n33080;
  assign new_new_n40690__ = ~new_new_n40682__ & new_new_n40689__;
  assign new_new_n40691__ = ~new_new_n40673__ & new_new_n40690__;
  assign new_new_n40692__ = ys__n33082 & ys__n33083;
  assign new_new_n40693__ = ys__n33082 & ys__n33081;
  assign new_new_n40694__ = ~new_new_n40682__ & new_new_n40693__;
  assign new_new_n40695__ = ~new_new_n40692__ & ~new_new_n40694__;
  assign new_new_n40696__ = ~new_new_n40691__ & new_new_n40695__;
  assign new_new_n40697__ = new_new_n39793__ & new_new_n40627__;
  assign new_new_n40698__ = ys__n24762 & new_new_n40629__;
  assign new_new_n40699__ = new_new_n39793__ & new_new_n40631__;
  assign new_new_n40700__ = ~new_new_n40698__ & ~new_new_n40699__;
  assign new_new_n40701__ = ~new_new_n40697__ & new_new_n40700__;
  assign ys__n33087 = ~new_new_n40644__ & ~new_new_n40701__;
  assign new_new_n40703__ = new_new_n39764__ & new_new_n40627__;
  assign new_new_n40704__ = ys__n24759 & new_new_n40629__;
  assign new_new_n40705__ = new_new_n39764__ & new_new_n40631__;
  assign new_new_n40706__ = ~new_new_n40704__ & ~new_new_n40705__;
  assign new_new_n40707__ = ~new_new_n40703__ & new_new_n40706__;
  assign ys__n33086 = ~new_new_n40644__ & ~new_new_n40707__;
  assign new_new_n40709__ = ~ys__n33087 & ys__n33086;
  assign new_new_n40710__ = ys__n33087 & ~ys__n33086;
  assign new_new_n40711__ = ~new_new_n40709__ & ~new_new_n40710__;
  assign new_new_n40712__ = new_new_n39736__ & new_new_n40627__;
  assign new_new_n40713__ = ys__n24756 & new_new_n40629__;
  assign new_new_n40714__ = new_new_n39736__ & new_new_n40631__;
  assign new_new_n40715__ = ~new_new_n40713__ & ~new_new_n40714__;
  assign new_new_n40716__ = ~new_new_n40712__ & new_new_n40715__;
  assign ys__n33085 = ~new_new_n40644__ & ~new_new_n40716__;
  assign new_new_n40718__ = ~ys__n33086 & ys__n33085;
  assign new_new_n40719__ = ys__n33086 & ~ys__n33085;
  assign new_new_n40720__ = ~new_new_n40718__ & ~new_new_n40719__;
  assign new_new_n40721__ = ~new_new_n40711__ & ~new_new_n40720__;
  assign new_new_n40722__ = new_new_n39711__ & new_new_n40627__;
  assign new_new_n40723__ = ys__n24753 & new_new_n40629__;
  assign new_new_n40724__ = new_new_n39711__ & new_new_n40631__;
  assign new_new_n40725__ = ~new_new_n40723__ & ~new_new_n40724__;
  assign new_new_n40726__ = ~new_new_n40722__ & new_new_n40725__;
  assign ys__n33084 = ~new_new_n40644__ & ~new_new_n40726__;
  assign new_new_n40728__ = ~ys__n33085 & ys__n33084;
  assign new_new_n40729__ = ys__n33085 & ~ys__n33084;
  assign new_new_n40730__ = ~new_new_n40728__ & ~new_new_n40729__;
  assign new_new_n40731__ = ys__n33083 & ~ys__n33084;
  assign new_new_n40732__ = ~ys__n33083 & ys__n33084;
  assign new_new_n40733__ = ~new_new_n40731__ & ~new_new_n40732__;
  assign new_new_n40734__ = ~new_new_n40730__ & ~new_new_n40733__;
  assign new_new_n40735__ = new_new_n40721__ & new_new_n40734__;
  assign new_new_n40736__ = ~new_new_n40696__ & new_new_n40735__;
  assign new_new_n40737__ = ys__n33085 & ys__n33084;
  assign new_new_n40738__ = ys__n33083 & ys__n33084;
  assign new_new_n40739__ = ~new_new_n40730__ & new_new_n40738__;
  assign new_new_n40740__ = ~new_new_n40737__ & ~new_new_n40739__;
  assign new_new_n40741__ = new_new_n40721__ & ~new_new_n40740__;
  assign new_new_n40742__ = ys__n33087 & ys__n33086;
  assign new_new_n40743__ = ys__n33086 & ys__n33085;
  assign new_new_n40744__ = ~new_new_n40711__ & new_new_n40743__;
  assign new_new_n40745__ = ~new_new_n40742__ & ~new_new_n40744__;
  assign new_new_n40746__ = ~new_new_n40741__ & new_new_n40745__;
  assign new_new_n40747__ = ~new_new_n40736__ & new_new_n40746__;
  assign new_new_n40748__ = new_new_n39992__ & new_new_n40627__;
  assign new_new_n40749__ = ys__n24783 & new_new_n40629__;
  assign new_new_n40750__ = new_new_n39992__ & new_new_n40631__;
  assign new_new_n40751__ = ~new_new_n40749__ & ~new_new_n40750__;
  assign new_new_n40752__ = ~new_new_n40748__ & new_new_n40751__;
  assign ys__n33094 = ~new_new_n40644__ & ~new_new_n40752__;
  assign new_new_n40754__ = ~ys__n33095 & ys__n33094;
  assign new_new_n40755__ = ys__n33095 & ~ys__n33094;
  assign new_new_n40756__ = ~new_new_n40754__ & ~new_new_n40755__;
  assign new_new_n40757__ = new_new_n39963__ & new_new_n40627__;
  assign new_new_n40758__ = ys__n24780 & new_new_n40629__;
  assign new_new_n40759__ = new_new_n39963__ & new_new_n40631__;
  assign new_new_n40760__ = ~new_new_n40758__ & ~new_new_n40759__;
  assign new_new_n40761__ = ~new_new_n40757__ & new_new_n40760__;
  assign ys__n33093 = ~new_new_n40644__ & ~new_new_n40761__;
  assign new_new_n40763__ = ~ys__n33094 & ys__n33093;
  assign new_new_n40764__ = ys__n33094 & ~ys__n33093;
  assign new_new_n40765__ = ~new_new_n40763__ & ~new_new_n40764__;
  assign new_new_n40766__ = ~new_new_n40756__ & ~new_new_n40765__;
  assign new_new_n40767__ = new_new_n39934__ & new_new_n40627__;
  assign new_new_n40768__ = ys__n24777 & new_new_n40629__;
  assign new_new_n40769__ = new_new_n39934__ & new_new_n40631__;
  assign new_new_n40770__ = ~new_new_n40768__ & ~new_new_n40769__;
  assign new_new_n40771__ = ~new_new_n40767__ & new_new_n40770__;
  assign ys__n33092 = ~new_new_n40644__ & ~new_new_n40771__;
  assign new_new_n40773__ = ~ys__n33093 & ys__n33092;
  assign new_new_n40774__ = ys__n33093 & ~ys__n33092;
  assign new_new_n40775__ = ~new_new_n40773__ & ~new_new_n40774__;
  assign new_new_n40776__ = new_new_n39905__ & new_new_n40627__;
  assign new_new_n40777__ = ys__n24774 & new_new_n40629__;
  assign new_new_n40778__ = new_new_n39905__ & new_new_n40631__;
  assign new_new_n40779__ = ~new_new_n40777__ & ~new_new_n40778__;
  assign new_new_n40780__ = ~new_new_n40776__ & new_new_n40779__;
  assign ys__n33091 = ~new_new_n40644__ & ~new_new_n40780__;
  assign new_new_n40782__ = ~ys__n33092 & ys__n33091;
  assign new_new_n40783__ = ys__n33092 & ~ys__n33091;
  assign new_new_n40784__ = ~new_new_n40782__ & ~new_new_n40783__;
  assign new_new_n40785__ = ~new_new_n40775__ & ~new_new_n40784__;
  assign new_new_n40786__ = new_new_n40766__ & new_new_n40785__;
  assign new_new_n40787__ = new_new_n39876__ & new_new_n40627__;
  assign new_new_n40788__ = ys__n24771 & new_new_n40629__;
  assign new_new_n40789__ = new_new_n39876__ & new_new_n40631__;
  assign new_new_n40790__ = ~new_new_n40788__ & ~new_new_n40789__;
  assign new_new_n40791__ = ~new_new_n40787__ & new_new_n40790__;
  assign ys__n33090 = ~new_new_n40644__ & ~new_new_n40791__;
  assign new_new_n40793__ = ~ys__n33091 & ys__n33090;
  assign new_new_n40794__ = ys__n33091 & ~ys__n33090;
  assign new_new_n40795__ = ~new_new_n40793__ & ~new_new_n40794__;
  assign new_new_n40796__ = new_new_n39848__ & new_new_n40627__;
  assign new_new_n40797__ = ys__n24768 & new_new_n40629__;
  assign new_new_n40798__ = new_new_n39848__ & new_new_n40631__;
  assign new_new_n40799__ = ~new_new_n40797__ & ~new_new_n40798__;
  assign new_new_n40800__ = ~new_new_n40796__ & new_new_n40799__;
  assign ys__n33089 = ~new_new_n40644__ & ~new_new_n40800__;
  assign new_new_n40802__ = ~ys__n33090 & ys__n33089;
  assign new_new_n40803__ = ys__n33090 & ~ys__n33089;
  assign new_new_n40804__ = ~new_new_n40802__ & ~new_new_n40803__;
  assign new_new_n40805__ = ~new_new_n40795__ & ~new_new_n40804__;
  assign new_new_n40806__ = new_new_n39822__ & new_new_n40627__;
  assign new_new_n40807__ = ys__n24765 & new_new_n40629__;
  assign new_new_n40808__ = new_new_n39822__ & new_new_n40631__;
  assign new_new_n40809__ = ~new_new_n40807__ & ~new_new_n40808__;
  assign new_new_n40810__ = ~new_new_n40806__ & new_new_n40809__;
  assign ys__n33088 = ~new_new_n40644__ & ~new_new_n40810__;
  assign new_new_n40812__ = ~ys__n33089 & ys__n33088;
  assign new_new_n40813__ = ys__n33089 & ~ys__n33088;
  assign new_new_n40814__ = ~new_new_n40812__ & ~new_new_n40813__;
  assign new_new_n40815__ = ys__n33087 & ~ys__n33088;
  assign new_new_n40816__ = ~ys__n33087 & ys__n33088;
  assign new_new_n40817__ = ~new_new_n40815__ & ~new_new_n40816__;
  assign new_new_n40818__ = ~new_new_n40814__ & ~new_new_n40817__;
  assign new_new_n40819__ = new_new_n40805__ & new_new_n40818__;
  assign new_new_n40820__ = new_new_n40786__ & new_new_n40819__;
  assign new_new_n40821__ = ~new_new_n40747__ & new_new_n40820__;
  assign new_new_n40822__ = ys__n33089 & ys__n33088;
  assign new_new_n40823__ = ys__n33087 & ys__n33088;
  assign new_new_n40824__ = ~new_new_n40814__ & new_new_n40823__;
  assign new_new_n40825__ = ~new_new_n40822__ & ~new_new_n40824__;
  assign new_new_n40826__ = new_new_n40805__ & ~new_new_n40825__;
  assign new_new_n40827__ = ys__n33091 & ys__n33090;
  assign new_new_n40828__ = ys__n33090 & ys__n33089;
  assign new_new_n40829__ = ~new_new_n40795__ & new_new_n40828__;
  assign new_new_n40830__ = ~new_new_n40827__ & ~new_new_n40829__;
  assign new_new_n40831__ = ~new_new_n40826__ & new_new_n40830__;
  assign new_new_n40832__ = new_new_n40786__ & ~new_new_n40831__;
  assign new_new_n40833__ = ys__n33093 & ys__n33092;
  assign new_new_n40834__ = ys__n33092 & ys__n33091;
  assign new_new_n40835__ = ~new_new_n40775__ & new_new_n40834__;
  assign new_new_n40836__ = ~new_new_n40833__ & ~new_new_n40835__;
  assign new_new_n40837__ = new_new_n40766__ & ~new_new_n40836__;
  assign new_new_n40838__ = ys__n33095 & ys__n33094;
  assign new_new_n40839__ = ys__n33094 & ys__n33093;
  assign new_new_n40840__ = ~new_new_n40756__ & new_new_n40839__;
  assign new_new_n40841__ = ~new_new_n40838__ & ~new_new_n40840__;
  assign new_new_n40842__ = ~new_new_n40837__ & new_new_n40841__;
  assign new_new_n40843__ = ~new_new_n40832__ & new_new_n40842__;
  assign new_new_n40844__ = ~new_new_n40821__ & new_new_n40843__;
  assign new_new_n40845__ = ~new_new_n40658__ & new_new_n40844__;
  assign new_new_n40846__ = new_new_n40658__ & ~new_new_n40844__;
  assign ys__n30616 = new_new_n40845__ | new_new_n40846__;
  assign new_new_n40848__ = ys__n24792 & new_new_n40629__;
  assign new_new_n40849__ = new_new_n40076__ & new_new_n40631__;
  assign new_new_n40850__ = ~new_new_n40848__ & ~new_new_n40849__;
  assign new_new_n40851__ = new_new_n39632__ & new_new_n40639__;
  assign new_new_n40852__ = new_new_n39632__ & new_new_n40641__;
  assign new_new_n40853__ = new_new_n40076__ & new_new_n40627__;
  assign new_new_n40854__ = ~new_new_n40852__ & ~new_new_n40853__;
  assign new_new_n40855__ = ~new_new_n40851__ & new_new_n40854__;
  assign new_new_n40856__ = new_new_n40850__ & new_new_n40855__;
  assign ys__n33097 = ~new_new_n40644__ & ~new_new_n40856__;
  assign new_new_n40858__ = ~ys__n33096 & ys__n33097;
  assign new_new_n40859__ = ys__n33096 & ~ys__n33097;
  assign new_new_n40860__ = ~new_new_n40858__ & ~new_new_n40859__;
  assign new_new_n40861__ = ys__n33095 & ys__n33096;
  assign new_new_n40862__ = new_new_n40860__ & new_new_n40861__;
  assign new_new_n40863__ = ~new_new_n40860__ & ~new_new_n40861__;
  assign new_new_n40864__ = ~new_new_n40862__ & ~new_new_n40863__;
  assign new_new_n40865__ = new_new_n40844__ & ~new_new_n40864__;
  assign new_new_n40866__ = ~new_new_n40658__ & new_new_n40864__;
  assign new_new_n40867__ = new_new_n40658__ & ~new_new_n40864__;
  assign new_new_n40868__ = ~new_new_n40866__ & ~new_new_n40867__;
  assign new_new_n40869__ = ~new_new_n40844__ & ~new_new_n40868__;
  assign ys__n30619 = new_new_n40865__ | new_new_n40869__;
  assign new_new_n40871__ = ys__n24795 & new_new_n40629__;
  assign new_new_n40872__ = new_new_n40108__ & new_new_n40631__;
  assign new_new_n40873__ = ~new_new_n40871__ & ~new_new_n40872__;
  assign new_new_n40874__ = new_new_n39659__ & new_new_n40639__;
  assign new_new_n40875__ = new_new_n39659__ & new_new_n40641__;
  assign new_new_n40876__ = new_new_n40108__ & new_new_n40627__;
  assign new_new_n40877__ = ~new_new_n40875__ & ~new_new_n40876__;
  assign new_new_n40878__ = ~new_new_n40874__ & new_new_n40877__;
  assign new_new_n40879__ = new_new_n40873__ & new_new_n40878__;
  assign ys__n33098 = ~new_new_n40644__ & ~new_new_n40879__;
  assign new_new_n40881__ = ~ys__n33097 & ys__n33098;
  assign new_new_n40882__ = ys__n33097 & ~ys__n33098;
  assign new_new_n40883__ = ~new_new_n40881__ & ~new_new_n40882__;
  assign new_new_n40884__ = ys__n33096 & ys__n33097;
  assign new_new_n40885__ = ~new_new_n40860__ & new_new_n40861__;
  assign new_new_n40886__ = ~new_new_n40884__ & ~new_new_n40885__;
  assign new_new_n40887__ = new_new_n40883__ & ~new_new_n40886__;
  assign new_new_n40888__ = ~new_new_n40883__ & new_new_n40886__;
  assign new_new_n40889__ = ~new_new_n40887__ & ~new_new_n40888__;
  assign new_new_n40890__ = new_new_n40844__ & ~new_new_n40889__;
  assign new_new_n40891__ = ~new_new_n40658__ & ~new_new_n40864__;
  assign new_new_n40892__ = new_new_n40889__ & new_new_n40891__;
  assign new_new_n40893__ = ~new_new_n40889__ & ~new_new_n40891__;
  assign new_new_n40894__ = ~new_new_n40892__ & ~new_new_n40893__;
  assign new_new_n40895__ = ~new_new_n40844__ & ~new_new_n40894__;
  assign ys__n30622 = new_new_n40890__ | new_new_n40895__;
  assign new_new_n40897__ = ys__n24798 & new_new_n40629__;
  assign new_new_n40898__ = new_new_n40143__ & new_new_n40631__;
  assign new_new_n40899__ = ~new_new_n40897__ & ~new_new_n40898__;
  assign new_new_n40900__ = new_new_n39685__ & new_new_n40639__;
  assign new_new_n40901__ = new_new_n39685__ & new_new_n40641__;
  assign new_new_n40902__ = new_new_n40143__ & new_new_n40627__;
  assign new_new_n40903__ = ~new_new_n40901__ & ~new_new_n40902__;
  assign new_new_n40904__ = ~new_new_n40900__ & new_new_n40903__;
  assign new_new_n40905__ = new_new_n40899__ & new_new_n40904__;
  assign ys__n33099 = ~new_new_n40644__ & ~new_new_n40905__;
  assign new_new_n40907__ = ~ys__n33098 & ys__n33099;
  assign new_new_n40908__ = ys__n33098 & ~ys__n33099;
  assign new_new_n40909__ = ~new_new_n40907__ & ~new_new_n40908__;
  assign new_new_n40910__ = ys__n33097 & ys__n33098;
  assign new_new_n40911__ = ~new_new_n40883__ & ~new_new_n40886__;
  assign new_new_n40912__ = ~new_new_n40910__ & ~new_new_n40911__;
  assign new_new_n40913__ = new_new_n40909__ & ~new_new_n40912__;
  assign new_new_n40914__ = ~new_new_n40909__ & new_new_n40912__;
  assign new_new_n40915__ = ~new_new_n40913__ & ~new_new_n40914__;
  assign new_new_n40916__ = new_new_n40844__ & ~new_new_n40915__;
  assign new_new_n40917__ = ~new_new_n40889__ & new_new_n40891__;
  assign new_new_n40918__ = new_new_n40915__ & new_new_n40917__;
  assign new_new_n40919__ = ~new_new_n40915__ & ~new_new_n40917__;
  assign new_new_n40920__ = ~new_new_n40918__ & ~new_new_n40919__;
  assign new_new_n40921__ = ~new_new_n40844__ & ~new_new_n40920__;
  assign ys__n30625 = new_new_n40916__ | new_new_n40921__;
  assign new_new_n40923__ = ys__n24801 & new_new_n40629__;
  assign new_new_n40924__ = new_new_n40178__ & new_new_n40631__;
  assign new_new_n40925__ = ~new_new_n40923__ & ~new_new_n40924__;
  assign new_new_n40926__ = new_new_n39711__ & new_new_n40639__;
  assign new_new_n40927__ = new_new_n39711__ & new_new_n40641__;
  assign new_new_n40928__ = new_new_n40178__ & new_new_n40627__;
  assign new_new_n40929__ = ~new_new_n40927__ & ~new_new_n40928__;
  assign new_new_n40930__ = ~new_new_n40926__ & new_new_n40929__;
  assign new_new_n40931__ = new_new_n40925__ & new_new_n40930__;
  assign ys__n33100 = ~new_new_n40644__ & ~new_new_n40931__;
  assign new_new_n40933__ = ~ys__n33099 & ys__n33100;
  assign new_new_n40934__ = ys__n33099 & ~ys__n33100;
  assign new_new_n40935__ = ~new_new_n40933__ & ~new_new_n40934__;
  assign new_new_n40936__ = ~new_new_n40883__ & ~new_new_n40909__;
  assign new_new_n40937__ = ~new_new_n40886__ & new_new_n40936__;
  assign new_new_n40938__ = ys__n33098 & ys__n33099;
  assign new_new_n40939__ = ~new_new_n40909__ & new_new_n40910__;
  assign new_new_n40940__ = ~new_new_n40938__ & ~new_new_n40939__;
  assign new_new_n40941__ = ~new_new_n40937__ & new_new_n40940__;
  assign new_new_n40942__ = new_new_n40935__ & ~new_new_n40941__;
  assign new_new_n40943__ = ~new_new_n40935__ & new_new_n40941__;
  assign new_new_n40944__ = ~new_new_n40942__ & ~new_new_n40943__;
  assign new_new_n40945__ = new_new_n40844__ & ~new_new_n40944__;
  assign new_new_n40946__ = ~new_new_n40915__ & new_new_n40917__;
  assign new_new_n40947__ = new_new_n40944__ & new_new_n40946__;
  assign new_new_n40948__ = ~new_new_n40944__ & ~new_new_n40946__;
  assign new_new_n40949__ = ~new_new_n40947__ & ~new_new_n40948__;
  assign new_new_n40950__ = ~new_new_n40844__ & ~new_new_n40949__;
  assign ys__n30628 = new_new_n40945__ | new_new_n40950__;
  assign new_new_n40952__ = ys__n24804 & new_new_n40629__;
  assign new_new_n40953__ = new_new_n40213__ & new_new_n40631__;
  assign new_new_n40954__ = ~new_new_n40952__ & ~new_new_n40953__;
  assign new_new_n40955__ = new_new_n39736__ & new_new_n40639__;
  assign new_new_n40956__ = new_new_n39736__ & new_new_n40641__;
  assign new_new_n40957__ = new_new_n40213__ & new_new_n40627__;
  assign new_new_n40958__ = ~new_new_n40956__ & ~new_new_n40957__;
  assign new_new_n40959__ = ~new_new_n40955__ & new_new_n40958__;
  assign new_new_n40960__ = new_new_n40954__ & new_new_n40959__;
  assign ys__n33101 = ~new_new_n40644__ & ~new_new_n40960__;
  assign new_new_n40962__ = ~ys__n33100 & ys__n33101;
  assign new_new_n40963__ = ys__n33100 & ~ys__n33101;
  assign new_new_n40964__ = ~new_new_n40962__ & ~new_new_n40963__;
  assign new_new_n40965__ = ys__n33099 & ys__n33100;
  assign new_new_n40966__ = ~new_new_n40935__ & ~new_new_n40941__;
  assign new_new_n40967__ = ~new_new_n40965__ & ~new_new_n40966__;
  assign new_new_n40968__ = new_new_n40964__ & ~new_new_n40967__;
  assign new_new_n40969__ = ~new_new_n40964__ & new_new_n40967__;
  assign new_new_n40970__ = ~new_new_n40968__ & ~new_new_n40969__;
  assign new_new_n40971__ = new_new_n40844__ & ~new_new_n40970__;
  assign new_new_n40972__ = ~new_new_n40944__ & new_new_n40946__;
  assign new_new_n40973__ = new_new_n40970__ & new_new_n40972__;
  assign new_new_n40974__ = ~new_new_n40970__ & ~new_new_n40972__;
  assign new_new_n40975__ = ~new_new_n40973__ & ~new_new_n40974__;
  assign new_new_n40976__ = ~new_new_n40844__ & ~new_new_n40975__;
  assign ys__n30631 = new_new_n40971__ | new_new_n40976__;
  assign new_new_n40978__ = ys__n24807 & new_new_n40629__;
  assign new_new_n40979__ = new_new_n40250__ & new_new_n40631__;
  assign new_new_n40980__ = ~new_new_n40978__ & ~new_new_n40979__;
  assign new_new_n40981__ = new_new_n39764__ & new_new_n40639__;
  assign new_new_n40982__ = new_new_n39764__ & new_new_n40641__;
  assign new_new_n40983__ = new_new_n40250__ & new_new_n40627__;
  assign new_new_n40984__ = ~new_new_n40982__ & ~new_new_n40983__;
  assign new_new_n40985__ = ~new_new_n40981__ & new_new_n40984__;
  assign new_new_n40986__ = new_new_n40980__ & new_new_n40985__;
  assign ys__n33102 = ~new_new_n40644__ & ~new_new_n40986__;
  assign new_new_n40988__ = ~ys__n33101 & ys__n33102;
  assign new_new_n40989__ = ys__n33101 & ~ys__n33102;
  assign new_new_n40990__ = ~new_new_n40988__ & ~new_new_n40989__;
  assign new_new_n40991__ = ys__n33100 & ys__n33101;
  assign new_new_n40992__ = ~new_new_n40964__ & new_new_n40965__;
  assign new_new_n40993__ = ~new_new_n40991__ & ~new_new_n40992__;
  assign new_new_n40994__ = ~new_new_n40935__ & ~new_new_n40964__;
  assign new_new_n40995__ = ~new_new_n40941__ & new_new_n40994__;
  assign new_new_n40996__ = new_new_n40993__ & ~new_new_n40995__;
  assign new_new_n40997__ = new_new_n40990__ & ~new_new_n40996__;
  assign new_new_n40998__ = ~new_new_n40990__ & new_new_n40996__;
  assign new_new_n40999__ = ~new_new_n40997__ & ~new_new_n40998__;
  assign new_new_n41000__ = new_new_n40844__ & ~new_new_n40999__;
  assign new_new_n41001__ = ~new_new_n40944__ & ~new_new_n40970__;
  assign new_new_n41002__ = new_new_n40946__ & new_new_n41001__;
  assign new_new_n41003__ = new_new_n40999__ & new_new_n41002__;
  assign new_new_n41004__ = ~new_new_n40999__ & ~new_new_n41002__;
  assign new_new_n41005__ = ~new_new_n41003__ & ~new_new_n41004__;
  assign new_new_n41006__ = ~new_new_n40844__ & ~new_new_n41005__;
  assign ys__n30634 = new_new_n41000__ | new_new_n41006__;
  assign new_new_n41008__ = ys__n24810 & new_new_n40629__;
  assign new_new_n41009__ = new_new_n40288__ & new_new_n40631__;
  assign new_new_n41010__ = ~new_new_n41008__ & ~new_new_n41009__;
  assign new_new_n41011__ = new_new_n39793__ & new_new_n40639__;
  assign new_new_n41012__ = new_new_n39793__ & new_new_n40641__;
  assign new_new_n41013__ = new_new_n40288__ & new_new_n40627__;
  assign new_new_n41014__ = ~new_new_n41012__ & ~new_new_n41013__;
  assign new_new_n41015__ = ~new_new_n41011__ & new_new_n41014__;
  assign new_new_n41016__ = new_new_n41010__ & new_new_n41015__;
  assign ys__n33103 = ~new_new_n40644__ & ~new_new_n41016__;
  assign new_new_n41018__ = ~ys__n33102 & ys__n33103;
  assign new_new_n41019__ = ys__n33102 & ~ys__n33103;
  assign new_new_n41020__ = ~new_new_n41018__ & ~new_new_n41019__;
  assign new_new_n41021__ = ys__n33101 & ys__n33102;
  assign new_new_n41022__ = ~new_new_n40990__ & ~new_new_n40996__;
  assign new_new_n41023__ = ~new_new_n41021__ & ~new_new_n41022__;
  assign new_new_n41024__ = new_new_n41020__ & ~new_new_n41023__;
  assign new_new_n41025__ = ~new_new_n41020__ & new_new_n41023__;
  assign new_new_n41026__ = ~new_new_n41024__ & ~new_new_n41025__;
  assign new_new_n41027__ = new_new_n40844__ & ~new_new_n41026__;
  assign new_new_n41028__ = ~new_new_n40999__ & new_new_n41002__;
  assign new_new_n41029__ = new_new_n41026__ & new_new_n41028__;
  assign new_new_n41030__ = ~new_new_n41026__ & ~new_new_n41028__;
  assign new_new_n41031__ = ~new_new_n41029__ & ~new_new_n41030__;
  assign new_new_n41032__ = ~new_new_n40844__ & ~new_new_n41031__;
  assign ys__n30637 = new_new_n41027__ | new_new_n41032__;
  assign new_new_n41034__ = ys__n24813 & new_new_n40629__;
  assign new_new_n41035__ = new_new_n40326__ & new_new_n40631__;
  assign new_new_n41036__ = ~new_new_n41034__ & ~new_new_n41035__;
  assign new_new_n41037__ = new_new_n39822__ & new_new_n40639__;
  assign new_new_n41038__ = new_new_n39822__ & new_new_n40641__;
  assign new_new_n41039__ = new_new_n40326__ & new_new_n40627__;
  assign new_new_n41040__ = ~new_new_n41038__ & ~new_new_n41039__;
  assign new_new_n41041__ = ~new_new_n41037__ & new_new_n41040__;
  assign new_new_n41042__ = new_new_n41036__ & new_new_n41041__;
  assign ys__n33104 = ~new_new_n40644__ & ~new_new_n41042__;
  assign new_new_n41044__ = ~ys__n33103 & ys__n33104;
  assign new_new_n41045__ = ys__n33103 & ~ys__n33104;
  assign new_new_n41046__ = ~new_new_n41044__ & ~new_new_n41045__;
  assign new_new_n41047__ = ~new_new_n40990__ & ~new_new_n41020__;
  assign new_new_n41048__ = new_new_n40994__ & new_new_n41047__;
  assign new_new_n41049__ = ~new_new_n40941__ & new_new_n41048__;
  assign new_new_n41050__ = ~new_new_n40993__ & new_new_n41047__;
  assign new_new_n41051__ = ys__n33102 & ys__n33103;
  assign new_new_n41052__ = ~new_new_n41020__ & new_new_n41021__;
  assign new_new_n41053__ = ~new_new_n41051__ & ~new_new_n41052__;
  assign new_new_n41054__ = ~new_new_n41050__ & new_new_n41053__;
  assign new_new_n41055__ = ~new_new_n41049__ & new_new_n41054__;
  assign new_new_n41056__ = new_new_n41046__ & ~new_new_n41055__;
  assign new_new_n41057__ = ~new_new_n41046__ & new_new_n41055__;
  assign new_new_n41058__ = ~new_new_n41056__ & ~new_new_n41057__;
  assign new_new_n41059__ = new_new_n40844__ & ~new_new_n41058__;
  assign new_new_n41060__ = new_new_n40946__ & ~new_new_n40999__;
  assign new_new_n41061__ = new_new_n41001__ & new_new_n41060__;
  assign new_new_n41062__ = ~new_new_n41026__ & new_new_n41061__;
  assign new_new_n41063__ = new_new_n41058__ & new_new_n41062__;
  assign new_new_n41064__ = ~new_new_n41058__ & ~new_new_n41062__;
  assign new_new_n41065__ = ~new_new_n41063__ & ~new_new_n41064__;
  assign new_new_n41066__ = ~new_new_n40844__ & ~new_new_n41065__;
  assign ys__n30640 = new_new_n41059__ | new_new_n41066__;
  assign new_new_n41068__ = ys__n24816 & new_new_n40629__;
  assign new_new_n41069__ = new_new_n40362__ & new_new_n40631__;
  assign new_new_n41070__ = ~new_new_n41068__ & ~new_new_n41069__;
  assign new_new_n41071__ = new_new_n39848__ & new_new_n40639__;
  assign new_new_n41072__ = new_new_n39848__ & new_new_n40641__;
  assign new_new_n41073__ = new_new_n40362__ & new_new_n40627__;
  assign new_new_n41074__ = ~new_new_n41072__ & ~new_new_n41073__;
  assign new_new_n41075__ = ~new_new_n41071__ & new_new_n41074__;
  assign new_new_n41076__ = new_new_n41070__ & new_new_n41075__;
  assign ys__n33105 = ~new_new_n40644__ & ~new_new_n41076__;
  assign new_new_n41078__ = ~ys__n33104 & ys__n33105;
  assign new_new_n41079__ = ys__n33104 & ~ys__n33105;
  assign new_new_n41080__ = ~new_new_n41078__ & ~new_new_n41079__;
  assign new_new_n41081__ = ys__n33103 & ys__n33104;
  assign new_new_n41082__ = ~new_new_n41046__ & ~new_new_n41055__;
  assign new_new_n41083__ = ~new_new_n41081__ & ~new_new_n41082__;
  assign new_new_n41084__ = new_new_n41080__ & ~new_new_n41083__;
  assign new_new_n41085__ = ~new_new_n41080__ & new_new_n41083__;
  assign new_new_n41086__ = ~new_new_n41084__ & ~new_new_n41085__;
  assign new_new_n41087__ = new_new_n40844__ & ~new_new_n41086__;
  assign new_new_n41088__ = ~new_new_n41058__ & new_new_n41062__;
  assign new_new_n41089__ = new_new_n41086__ & new_new_n41088__;
  assign new_new_n41090__ = ~new_new_n41086__ & ~new_new_n41088__;
  assign new_new_n41091__ = ~new_new_n41089__ & ~new_new_n41090__;
  assign new_new_n41092__ = ~new_new_n40844__ & ~new_new_n41091__;
  assign ys__n30643 = new_new_n41087__ | new_new_n41092__;
  assign new_new_n41094__ = ys__n24819 & new_new_n40629__;
  assign new_new_n41095__ = new_new_n40399__ & new_new_n40631__;
  assign new_new_n41096__ = ~new_new_n41094__ & ~new_new_n41095__;
  assign new_new_n41097__ = new_new_n39876__ & new_new_n40639__;
  assign new_new_n41098__ = new_new_n39876__ & new_new_n40641__;
  assign new_new_n41099__ = new_new_n40399__ & new_new_n40627__;
  assign new_new_n41100__ = ~new_new_n41098__ & ~new_new_n41099__;
  assign new_new_n41101__ = ~new_new_n41097__ & new_new_n41100__;
  assign new_new_n41102__ = new_new_n41096__ & new_new_n41101__;
  assign ys__n33106 = ~new_new_n40644__ & ~new_new_n41102__;
  assign new_new_n41104__ = ~ys__n33105 & ys__n33106;
  assign new_new_n41105__ = ys__n33105 & ~ys__n33106;
  assign new_new_n41106__ = ~new_new_n41104__ & ~new_new_n41105__;
  assign new_new_n41107__ = ys__n33104 & ys__n33105;
  assign new_new_n41108__ = ~new_new_n41080__ & new_new_n41081__;
  assign new_new_n41109__ = ~new_new_n41107__ & ~new_new_n41108__;
  assign new_new_n41110__ = ~new_new_n41046__ & ~new_new_n41080__;
  assign new_new_n41111__ = ~new_new_n41055__ & new_new_n41110__;
  assign new_new_n41112__ = new_new_n41109__ & ~new_new_n41111__;
  assign new_new_n41113__ = new_new_n41106__ & ~new_new_n41112__;
  assign new_new_n41114__ = ~new_new_n41106__ & new_new_n41112__;
  assign new_new_n41115__ = ~new_new_n41113__ & ~new_new_n41114__;
  assign new_new_n41116__ = new_new_n40844__ & ~new_new_n41115__;
  assign new_new_n41117__ = ~new_new_n41058__ & ~new_new_n41086__;
  assign new_new_n41118__ = new_new_n41062__ & new_new_n41117__;
  assign new_new_n41119__ = new_new_n41115__ & new_new_n41118__;
  assign new_new_n41120__ = ~new_new_n41115__ & ~new_new_n41118__;
  assign new_new_n41121__ = ~new_new_n41119__ & ~new_new_n41120__;
  assign new_new_n41122__ = ~new_new_n40844__ & ~new_new_n41121__;
  assign ys__n30646 = new_new_n41116__ | new_new_n41122__;
  assign new_new_n41124__ = ys__n24822 & new_new_n40629__;
  assign new_new_n41125__ = new_new_n40437__ & new_new_n40631__;
  assign new_new_n41126__ = ~new_new_n41124__ & ~new_new_n41125__;
  assign new_new_n41127__ = new_new_n39905__ & new_new_n40639__;
  assign new_new_n41128__ = new_new_n39905__ & new_new_n40641__;
  assign new_new_n41129__ = new_new_n40437__ & new_new_n40627__;
  assign new_new_n41130__ = ~new_new_n41128__ & ~new_new_n41129__;
  assign new_new_n41131__ = ~new_new_n41127__ & new_new_n41130__;
  assign new_new_n41132__ = new_new_n41126__ & new_new_n41131__;
  assign ys__n33107 = ~new_new_n40644__ & ~new_new_n41132__;
  assign new_new_n41134__ = ~ys__n33106 & ys__n33107;
  assign new_new_n41135__ = ys__n33106 & ~ys__n33107;
  assign new_new_n41136__ = ~new_new_n41134__ & ~new_new_n41135__;
  assign new_new_n41137__ = ys__n33105 & ys__n33106;
  assign new_new_n41138__ = ~new_new_n41106__ & ~new_new_n41112__;
  assign new_new_n41139__ = ~new_new_n41137__ & ~new_new_n41138__;
  assign new_new_n41140__ = new_new_n41136__ & ~new_new_n41139__;
  assign new_new_n41141__ = ~new_new_n41136__ & new_new_n41139__;
  assign new_new_n41142__ = ~new_new_n41140__ & ~new_new_n41141__;
  assign new_new_n41143__ = new_new_n40844__ & ~new_new_n41142__;
  assign new_new_n41144__ = ~new_new_n41115__ & new_new_n41118__;
  assign new_new_n41145__ = new_new_n41142__ & new_new_n41144__;
  assign new_new_n41146__ = ~new_new_n41142__ & ~new_new_n41144__;
  assign new_new_n41147__ = ~new_new_n41145__ & ~new_new_n41146__;
  assign new_new_n41148__ = ~new_new_n40844__ & ~new_new_n41147__;
  assign ys__n30649 = new_new_n41143__ | new_new_n41148__;
  assign new_new_n41150__ = ys__n24825 & new_new_n40629__;
  assign new_new_n41151__ = new_new_n40475__ & new_new_n40631__;
  assign new_new_n41152__ = ~new_new_n41150__ & ~new_new_n41151__;
  assign new_new_n41153__ = new_new_n39934__ & new_new_n40639__;
  assign new_new_n41154__ = new_new_n39934__ & new_new_n40641__;
  assign new_new_n41155__ = new_new_n40475__ & new_new_n40627__;
  assign new_new_n41156__ = ~new_new_n41154__ & ~new_new_n41155__;
  assign new_new_n41157__ = ~new_new_n41153__ & new_new_n41156__;
  assign new_new_n41158__ = new_new_n41152__ & new_new_n41157__;
  assign ys__n33108 = ~new_new_n40644__ & ~new_new_n41158__;
  assign new_new_n41160__ = ~ys__n33107 & ys__n33108;
  assign new_new_n41161__ = ys__n33107 & ~ys__n33108;
  assign new_new_n41162__ = ~new_new_n41160__ & ~new_new_n41161__;
  assign new_new_n41163__ = ~new_new_n41106__ & ~new_new_n41136__;
  assign new_new_n41164__ = ~new_new_n41109__ & new_new_n41163__;
  assign new_new_n41165__ = ys__n33106 & ys__n33107;
  assign new_new_n41166__ = ~new_new_n41136__ & new_new_n41137__;
  assign new_new_n41167__ = ~new_new_n41165__ & ~new_new_n41166__;
  assign new_new_n41168__ = ~new_new_n41164__ & new_new_n41167__;
  assign new_new_n41169__ = new_new_n41110__ & new_new_n41163__;
  assign new_new_n41170__ = ~new_new_n41055__ & new_new_n41169__;
  assign new_new_n41171__ = new_new_n41168__ & ~new_new_n41170__;
  assign new_new_n41172__ = new_new_n41162__ & ~new_new_n41171__;
  assign new_new_n41173__ = ~new_new_n41162__ & new_new_n41171__;
  assign new_new_n41174__ = ~new_new_n41172__ & ~new_new_n41173__;
  assign new_new_n41175__ = new_new_n40844__ & ~new_new_n41174__;
  assign new_new_n41176__ = ~new_new_n41115__ & new_new_n41117__;
  assign new_new_n41177__ = ~new_new_n41142__ & new_new_n41176__;
  assign new_new_n41178__ = new_new_n41062__ & new_new_n41177__;
  assign new_new_n41179__ = new_new_n41174__ & new_new_n41178__;
  assign new_new_n41180__ = ~new_new_n41174__ & ~new_new_n41178__;
  assign new_new_n41181__ = ~new_new_n41179__ & ~new_new_n41180__;
  assign new_new_n41182__ = ~new_new_n40844__ & ~new_new_n41181__;
  assign ys__n30652 = new_new_n41175__ | new_new_n41182__;
  assign new_new_n41184__ = ys__n24828 & new_new_n40629__;
  assign new_new_n41185__ = new_new_n40513__ & new_new_n40631__;
  assign new_new_n41186__ = ~new_new_n41184__ & ~new_new_n41185__;
  assign new_new_n41187__ = new_new_n39963__ & new_new_n40639__;
  assign new_new_n41188__ = new_new_n39963__ & new_new_n40641__;
  assign new_new_n41189__ = new_new_n40513__ & new_new_n40627__;
  assign new_new_n41190__ = ~new_new_n41188__ & ~new_new_n41189__;
  assign new_new_n41191__ = ~new_new_n41187__ & new_new_n41190__;
  assign new_new_n41192__ = new_new_n41186__ & new_new_n41191__;
  assign ys__n33109 = ~new_new_n40644__ & ~new_new_n41192__;
  assign new_new_n41194__ = ~ys__n33108 & ys__n33109;
  assign new_new_n41195__ = ys__n33108 & ~ys__n33109;
  assign new_new_n41196__ = ~new_new_n41194__ & ~new_new_n41195__;
  assign new_new_n41197__ = ys__n33107 & ys__n33108;
  assign new_new_n41198__ = ~new_new_n41162__ & ~new_new_n41171__;
  assign new_new_n41199__ = ~new_new_n41197__ & ~new_new_n41198__;
  assign new_new_n41200__ = new_new_n41196__ & ~new_new_n41199__;
  assign new_new_n41201__ = ~new_new_n41196__ & new_new_n41199__;
  assign new_new_n41202__ = ~new_new_n41200__ & ~new_new_n41201__;
  assign new_new_n41203__ = new_new_n40844__ & ~new_new_n41202__;
  assign new_new_n41204__ = ~new_new_n41174__ & new_new_n41178__;
  assign new_new_n41205__ = new_new_n41202__ & new_new_n41204__;
  assign new_new_n41206__ = ~new_new_n41202__ & ~new_new_n41204__;
  assign new_new_n41207__ = ~new_new_n41205__ & ~new_new_n41206__;
  assign new_new_n41208__ = ~new_new_n40844__ & ~new_new_n41207__;
  assign ys__n30655 = new_new_n41203__ | new_new_n41208__;
  assign new_new_n41210__ = ys__n24831 & new_new_n40629__;
  assign new_new_n41211__ = new_new_n40550__ & new_new_n40631__;
  assign new_new_n41212__ = ~new_new_n41210__ & ~new_new_n41211__;
  assign new_new_n41213__ = new_new_n39992__ & new_new_n40639__;
  assign new_new_n41214__ = new_new_n39992__ & new_new_n40641__;
  assign new_new_n41215__ = new_new_n40550__ & new_new_n40627__;
  assign new_new_n41216__ = ~new_new_n41214__ & ~new_new_n41215__;
  assign new_new_n41217__ = ~new_new_n41213__ & new_new_n41216__;
  assign new_new_n41218__ = new_new_n41212__ & new_new_n41217__;
  assign ys__n33110 = ~new_new_n40644__ & ~new_new_n41218__;
  assign new_new_n41220__ = ~ys__n33109 & ys__n33110;
  assign new_new_n41221__ = ys__n33109 & ~ys__n33110;
  assign new_new_n41222__ = ~new_new_n41220__ & ~new_new_n41221__;
  assign new_new_n41223__ = ys__n33108 & ys__n33109;
  assign new_new_n41224__ = ~new_new_n41196__ & new_new_n41197__;
  assign new_new_n41225__ = ~new_new_n41223__ & ~new_new_n41224__;
  assign new_new_n41226__ = ~new_new_n41162__ & ~new_new_n41196__;
  assign new_new_n41227__ = ~new_new_n41171__ & new_new_n41226__;
  assign new_new_n41228__ = new_new_n41225__ & ~new_new_n41227__;
  assign new_new_n41229__ = new_new_n41222__ & ~new_new_n41228__;
  assign new_new_n41230__ = ~new_new_n41222__ & new_new_n41228__;
  assign new_new_n41231__ = ~new_new_n41229__ & ~new_new_n41230__;
  assign new_new_n41232__ = new_new_n40844__ & ~new_new_n41231__;
  assign new_new_n41233__ = ~new_new_n41174__ & ~new_new_n41202__;
  assign new_new_n41234__ = new_new_n41178__ & new_new_n41233__;
  assign new_new_n41235__ = new_new_n41231__ & new_new_n41234__;
  assign new_new_n41236__ = ~new_new_n41231__ & ~new_new_n41234__;
  assign new_new_n41237__ = ~new_new_n41235__ & ~new_new_n41236__;
  assign new_new_n41238__ = ~new_new_n40844__ & ~new_new_n41237__;
  assign ys__n30658 = new_new_n41232__ | new_new_n41238__;
  assign new_new_n41240__ = new_new_n40588__ & new_new_n40631__;
  assign new_new_n41241__ = new_new_n40021__ & new_new_n40641__;
  assign new_new_n41242__ = ~new_new_n41240__ & ~new_new_n41241__;
  assign new_new_n41243__ = new_new_n40021__ & new_new_n40639__;
  assign new_new_n41244__ = ys__n24834 & new_new_n40629__;
  assign new_new_n41245__ = new_new_n40588__ & new_new_n40627__;
  assign new_new_n41246__ = ~new_new_n41244__ & ~new_new_n41245__;
  assign new_new_n41247__ = ~new_new_n41243__ & new_new_n41246__;
  assign new_new_n41248__ = new_new_n41242__ & new_new_n41247__;
  assign ys__n33111 = ~new_new_n40644__ & ~new_new_n41248__;
  assign new_new_n41250__ = ~ys__n33110 & ys__n33111;
  assign new_new_n41251__ = ys__n33110 & ~ys__n33111;
  assign new_new_n41252__ = ~new_new_n41250__ & ~new_new_n41251__;
  assign new_new_n41253__ = ys__n33109 & ys__n33110;
  assign new_new_n41254__ = ~new_new_n41222__ & ~new_new_n41228__;
  assign new_new_n41255__ = ~new_new_n41253__ & ~new_new_n41254__;
  assign new_new_n41256__ = new_new_n41252__ & ~new_new_n41255__;
  assign new_new_n41257__ = ~new_new_n41252__ & new_new_n41255__;
  assign new_new_n41258__ = ~new_new_n41256__ & ~new_new_n41257__;
  assign new_new_n41259__ = new_new_n40844__ & ~new_new_n41258__;
  assign new_new_n41260__ = ~new_new_n41231__ & new_new_n41234__;
  assign new_new_n41261__ = new_new_n41258__ & new_new_n41260__;
  assign new_new_n41262__ = ~new_new_n41258__ & ~new_new_n41260__;
  assign new_new_n41263__ = ~new_new_n41261__ & ~new_new_n41262__;
  assign new_new_n41264__ = ~new_new_n40844__ & ~new_new_n41263__;
  assign ys__n30661 = new_new_n41259__ | new_new_n41264__;
  assign new_new_n41266__ = ys__n39518 & new_new_n40629__;
  assign new_new_n41267__ = new_new_n41242__ & ~new_new_n41266__;
  assign ys__n30668 = ~new_new_n40644__ & ~new_new_n41267__;
  assign new_new_n41269__ = ~ys__n33111 & ys__n30668;
  assign new_new_n41270__ = ys__n33111 & ~ys__n30668;
  assign new_new_n41271__ = ~new_new_n41269__ & ~new_new_n41270__;
  assign new_new_n41272__ = ~new_new_n41222__ & ~new_new_n41252__;
  assign new_new_n41273__ = new_new_n41226__ & new_new_n41272__;
  assign new_new_n41274__ = new_new_n41169__ & new_new_n41273__;
  assign new_new_n41275__ = ~new_new_n41055__ & new_new_n41274__;
  assign new_new_n41276__ = ~new_new_n41168__ & new_new_n41273__;
  assign new_new_n41277__ = ~new_new_n41225__ & new_new_n41272__;
  assign new_new_n41278__ = ys__n33110 & ys__n33111;
  assign new_new_n41279__ = ~new_new_n41252__ & new_new_n41253__;
  assign new_new_n41280__ = ~new_new_n41278__ & ~new_new_n41279__;
  assign new_new_n41281__ = ~new_new_n41277__ & new_new_n41280__;
  assign new_new_n41282__ = ~new_new_n41276__ & new_new_n41281__;
  assign new_new_n41283__ = ~new_new_n41275__ & new_new_n41282__;
  assign new_new_n41284__ = new_new_n41271__ & ~new_new_n41283__;
  assign new_new_n41285__ = ~new_new_n41271__ & new_new_n41283__;
  assign new_new_n41286__ = ~new_new_n41284__ & ~new_new_n41285__;
  assign new_new_n41287__ = new_new_n40844__ & ~new_new_n41286__;
  assign new_new_n41288__ = new_new_n41062__ & ~new_new_n41231__;
  assign new_new_n41289__ = new_new_n41177__ & new_new_n41288__;
  assign new_new_n41290__ = new_new_n41233__ & new_new_n41289__;
  assign new_new_n41291__ = ~new_new_n41258__ & new_new_n41290__;
  assign new_new_n41292__ = new_new_n41286__ & new_new_n41291__;
  assign new_new_n41293__ = ~new_new_n41286__ & ~new_new_n41291__;
  assign new_new_n41294__ = ~new_new_n41292__ & ~new_new_n41293__;
  assign new_new_n41295__ = ~new_new_n40844__ & ~new_new_n41294__;
  assign ys__n30664 = new_new_n41287__ | new_new_n41295__;
  assign new_new_n41297__ = ys__n33111 & ys__n30668;
  assign new_new_n41298__ = ~new_new_n41271__ & ~new_new_n41283__;
  assign new_new_n41299__ = ~new_new_n41297__ & ~new_new_n41298__;
  assign new_new_n41300__ = new_new_n40844__ & ~new_new_n41299__;
  assign new_new_n41301__ = ~new_new_n41286__ & new_new_n41291__;
  assign new_new_n41302__ = new_new_n41299__ & new_new_n41301__;
  assign new_new_n41303__ = ~new_new_n41299__ & ~new_new_n41301__;
  assign new_new_n41304__ = ~new_new_n41302__ & ~new_new_n41303__;
  assign new_new_n41305__ = ~new_new_n40844__ & ~new_new_n41304__;
  assign ys__n30667 = new_new_n41300__ | new_new_n41305__;
  assign new_new_n41307__ = new_new_n40844__ & ys__n30668;
  assign new_new_n41308__ = ~new_new_n41286__ & ~new_new_n41299__;
  assign new_new_n41309__ = new_new_n41291__ & new_new_n41308__;
  assign new_new_n41310__ = ~ys__n30668 & new_new_n41309__;
  assign new_new_n41311__ = ys__n30668 & ~new_new_n41309__;
  assign new_new_n41312__ = ~new_new_n41310__ & ~new_new_n41311__;
  assign new_new_n41313__ = ~new_new_n40844__ & ~new_new_n41312__;
  assign ys__n30670 = new_new_n41307__ | new_new_n41313__;
  assign new_new_n41315__ = ~ys__n2535 & ~new_new_n24234__;
  assign new_new_n41316__ = ys__n2535 & ~new_new_n25508__;
  assign ys__n30797 = new_new_n41315__ | new_new_n41316__;
  assign new_new_n41318__ = ~ys__n2535 & ~new_new_n24312__;
  assign new_new_n41319__ = ys__n2535 & ~new_new_n25533__;
  assign ys__n30798 = new_new_n41318__ | new_new_n41319__;
  assign new_new_n41321__ = ~ys__n2535 & ~new_new_n24384__;
  assign new_new_n41322__ = ys__n2535 & ~new_new_n25560__;
  assign ys__n30799 = new_new_n41321__ | new_new_n41322__;
  assign new_new_n41324__ = ~ys__n2535 & ~new_new_n24459__;
  assign new_new_n41325__ = ys__n2535 & ~new_new_n25587__;
  assign ys__n30800 = new_new_n41324__ | new_new_n41325__;
  assign new_new_n41327__ = ~ys__n2535 & ~new_new_n24536__;
  assign new_new_n41328__ = ys__n2535 & ~new_new_n25617__;
  assign ys__n30801 = new_new_n41327__ | new_new_n41328__;
  assign new_new_n41330__ = ~ys__n2535 & ~new_new_n24611__;
  assign new_new_n41331__ = ys__n2535 & ~new_new_n25644__;
  assign ys__n30802 = new_new_n41330__ | new_new_n41331__;
  assign new_new_n41333__ = ~ys__n2535 & ~new_new_n24691__;
  assign new_new_n41334__ = ys__n2535 & ~new_new_n25674__;
  assign ys__n30803 = new_new_n41333__ | new_new_n41334__;
  assign new_new_n41336__ = ~ys__n2535 & ~new_new_n24767__;
  assign new_new_n41337__ = ys__n2535 & ~new_new_n25701__;
  assign ys__n30804 = new_new_n41336__ | new_new_n41337__;
  assign new_new_n41339__ = ~ys__n2535 & ~new_new_n24849__;
  assign new_new_n41340__ = ys__n2535 & ~new_new_n25734__;
  assign ys__n30805 = new_new_n41339__ | new_new_n41340__;
  assign new_new_n41342__ = ~ys__n2535 & ~new_new_n24924__;
  assign new_new_n41343__ = ys__n2535 & ~new_new_n25761__;
  assign ys__n30806 = new_new_n41342__ | new_new_n41343__;
  assign new_new_n41345__ = ~ys__n2535 & ~new_new_n25004__;
  assign new_new_n41346__ = ys__n2535 & ~new_new_n25791__;
  assign ys__n30807 = new_new_n41345__ | new_new_n41346__;
  assign new_new_n41348__ = ~ys__n2535 & ~new_new_n25080__;
  assign new_new_n41349__ = ys__n2535 & ~new_new_n25818__;
  assign ys__n30808 = new_new_n41348__ | new_new_n41349__;
  assign new_new_n41351__ = ~ys__n2535 & ~new_new_n25164__;
  assign new_new_n41352__ = ys__n2535 & ~new_new_n25851__;
  assign ys__n30809 = new_new_n41351__ | new_new_n41352__;
  assign new_new_n41354__ = ~ys__n2535 & ~new_new_n25240__;
  assign new_new_n41355__ = ys__n2535 & ~new_new_n25878__;
  assign ys__n30810 = new_new_n41354__ | new_new_n41355__;
  assign new_new_n41357__ = ~ys__n2535 & ~new_new_n25320__;
  assign new_new_n41358__ = ys__n2535 & ~new_new_n25908__;
  assign ys__n30811 = new_new_n41357__ | new_new_n41358__;
  assign new_new_n41360__ = ~ys__n2535 & ~new_new_n25394__;
  assign new_new_n41361__ = ys__n2535 & ~new_new_n25935__;
  assign ys__n30812 = new_new_n41360__ | new_new_n41361__;
  assign new_new_n41363__ = ~ys__n2535 & ~new_new_n24260__;
  assign new_new_n41364__ = ys__n2535 & new_new_n25961__;
  assign ys__n30813 = new_new_n41363__ | new_new_n41364__;
  assign new_new_n41366__ = ~ys__n152 & ys__n158;
  assign new_new_n41367__ = ~ys__n150 & ~ys__n156;
  assign new_new_n41368__ = new_new_n41366__ & new_new_n41367__;
  assign new_new_n41369__ = ys__n148 & new_new_n41368__;
  assign new_new_n41370__ = ys__n152 & ys__n158;
  assign new_new_n41371__ = ys__n148 & new_new_n41367__;
  assign new_new_n41372__ = new_new_n41370__ & new_new_n41371__;
  assign new_new_n41373__ = ~new_new_n41369__ & ~new_new_n41372__;
  assign new_new_n41374__ = ~ys__n150 & ys__n156;
  assign new_new_n41375__ = ~ys__n152 & ~ys__n158;
  assign new_new_n41376__ = ys__n148 & new_new_n41375__;
  assign new_new_n41377__ = new_new_n41374__ & new_new_n41376__;
  assign new_new_n41378__ = ys__n148 & new_new_n41366__;
  assign new_new_n41379__ = new_new_n41374__ & new_new_n41378__;
  assign new_new_n41380__ = ~new_new_n41377__ & ~new_new_n41379__;
  assign new_new_n41381__ = new_new_n41373__ & new_new_n41380__;
  assign new_new_n41382__ = ~ys__n30837 & ~new_new_n41381__;
  assign new_new_n41383__ = ys__n948 & new_new_n41382__;
  assign new_new_n41384__ = new_new_n12595__ & new_new_n12605__;
  assign new_new_n41385__ = ys__n352 & new_new_n12594__;
  assign new_new_n41386__ = new_new_n41384__ & new_new_n41385__;
  assign new_new_n41387__ = new_new_n12600__ & new_new_n12605__;
  assign new_new_n41388__ = new_new_n41385__ & new_new_n41387__;
  assign new_new_n41389__ = ~new_new_n41386__ & ~new_new_n41388__;
  assign new_new_n41390__ = new_new_n12604__ & new_new_n41389__;
  assign new_new_n41391__ = new_new_n12344__ & new_new_n12605__;
  assign new_new_n41392__ = new_new_n12607__ & new_new_n41391__;
  assign new_new_n41393__ = ~new_new_n12608__ & ~new_new_n41392__;
  assign new_new_n41394__ = new_new_n12342__ & new_new_n41387__;
  assign new_new_n41395__ = new_new_n12342__ & new_new_n12606__;
  assign new_new_n41396__ = ~new_new_n41394__ & ~new_new_n41395__;
  assign new_new_n41397__ = ys__n352 & new_new_n12336__;
  assign new_new_n41398__ = new_new_n12595__ & new_new_n41397__;
  assign new_new_n41399__ = new_new_n12341__ & new_new_n41398__;
  assign new_new_n41400__ = new_new_n12600__ & new_new_n41397__;
  assign new_new_n41401__ = new_new_n12341__ & new_new_n41400__;
  assign new_new_n41402__ = ~new_new_n41399__ & ~new_new_n41401__;
  assign new_new_n41403__ = new_new_n41396__ & new_new_n41402__;
  assign new_new_n41404__ = new_new_n41393__ & new_new_n41403__;
  assign new_new_n41405__ = new_new_n41390__ & new_new_n41404__;
  assign new_new_n41406__ = ys__n30832 & ~new_new_n41405__;
  assign ys__n30833 = new_new_n41383__ | new_new_n41406__;
  assign new_new_n41408__ = ~ys__n30837 & new_new_n41379__;
  assign new_new_n41409__ = ~ys__n4566 & new_new_n41408__;
  assign new_new_n41410__ = ~ys__n30832 & new_new_n41409__;
  assign new_new_n41411__ = ~new_new_n12603__ & ~new_new_n41401__;
  assign new_new_n41412__ = ~new_new_n41388__ & new_new_n41411__;
  assign new_new_n41413__ = ys__n30832 & ~new_new_n41412__;
  assign ys__n30835 = new_new_n41410__ | new_new_n41413__;
  assign new_new_n41415__ = ys__n30861 & ~ys__n30863;
  assign new_new_n41416__ = ys__n30862 & ys__n30863;
  assign ys__n30864 = new_new_n41415__ | new_new_n41416__;
  assign new_new_n41418__ = ys__n30865 & ~new_new_n13959__;
  assign new_new_n41419__ = new_new_n13962__ & new_new_n41418__;
  assign new_new_n41420__ = new_new_n13959__ & ys__n25842;
  assign ys__n30873 = new_new_n41419__ | new_new_n41420__;
  assign new_new_n41422__ = ys__n30867 & ~new_new_n13959__;
  assign new_new_n41423__ = new_new_n13962__ & new_new_n41422__;
  assign new_new_n41424__ = new_new_n13959__ & ys__n25844;
  assign ys__n30874 = new_new_n41423__ | new_new_n41424__;
  assign new_new_n41426__ = ys__n30869 & ~new_new_n13959__;
  assign new_new_n41427__ = new_new_n13962__ & new_new_n41426__;
  assign new_new_n41428__ = new_new_n13959__ & ys__n25846;
  assign ys__n30875 = new_new_n41427__ | new_new_n41428__;
  assign new_new_n41430__ = ys__n30871 & ~new_new_n13959__;
  assign new_new_n41431__ = new_new_n13962__ & new_new_n41430__;
  assign new_new_n41432__ = new_new_n13959__ & ys__n25852;
  assign ys__n30876 = new_new_n41431__ | new_new_n41432__;
  assign ys__n30942 = ys__n26425 & ~ys__n30941;
  assign ys__n30943 = ys__n26440 & ~ys__n30941;
  assign ys__n30944 = ys__n26446 & ~ys__n30941;
  assign new_new_n41437__ = ys__n26449 & ~ys__n30941;
  assign ys__n30945 = ys__n30941 | new_new_n41437__;
  assign ys__n30946 = ys__n26452 & ~ys__n30941;
  assign ys__n30947 = ys__n26466 & ~ys__n30941;
  assign ys__n30948 = ys__n26469 & ~ys__n30941;
  assign ys__n30949 = ys__n26472 & ~ys__n30941;
  assign new_new_n41443__ = ys__n26475 & ~ys__n30941;
  assign ys__n30950 = ys__n30941 | new_new_n41443__;
  assign new_new_n41445__ = ys__n26478 & ~ys__n30941;
  assign ys__n30951 = ys__n30941 | new_new_n41445__;
  assign ys__n30952 = ys__n26484 & ~ys__n30941;
  assign ys__n30953 = ys__n26496 & ~ys__n30941;
  assign ys__n30954 = ys__n26499 & ~ys__n30941;
  assign ys__n30955 = ys__n26502 & ~ys__n30941;
  assign ys__n30956 = ys__n26517 & ~ys__n30941;
  assign new_new_n41452__ = ~ys__n536 & ys__n538;
  assign new_new_n41453__ = new_new_n35345__ & new_new_n41452__;
  assign new_new_n41454__ = ys__n536 & ys__n538;
  assign new_new_n41455__ = new_new_n35343__ & new_new_n41454__;
  assign new_new_n41456__ = ~new_new_n41453__ & ~new_new_n41455__;
  assign new_new_n41457__ = new_new_n35345__ & new_new_n41454__;
  assign new_new_n41458__ = ys__n182 & ~ys__n536;
  assign new_new_n41459__ = ys__n538 & new_new_n41458__;
  assign new_new_n41460__ = ys__n182 & ys__n536;
  assign new_new_n41461__ = ys__n538 & new_new_n41460__;
  assign new_new_n41462__ = ~new_new_n41459__ & ~new_new_n41461__;
  assign new_new_n41463__ = ~new_new_n41457__ & new_new_n41462__;
  assign new_new_n41464__ = new_new_n35343__ & new_new_n41452__;
  assign new_new_n41465__ = ys__n538 & ~new_new_n41464__;
  assign new_new_n41466__ = new_new_n41456__ & new_new_n41465__;
  assign new_new_n41467__ = new_new_n41463__ & new_new_n41466__;
  assign new_new_n41468__ = ~new_new_n41456__ & ~new_new_n41467__;
  assign new_new_n41469__ = ~ys__n1386 & new_new_n12629__;
  assign new_new_n41470__ = new_new_n41468__ & new_new_n41469__;
  assign new_new_n41471__ = ys__n564 & new_new_n35343__;
  assign new_new_n41472__ = ys__n564 & ~new_new_n41471__;
  assign new_new_n41473__ = ys__n564 & new_new_n35345__;
  assign new_new_n41474__ = ys__n564 & ~new_new_n41473__;
  assign new_new_n41475__ = ys__n182 & ys__n564;
  assign new_new_n41476__ = ~new_new_n41471__ & ~new_new_n41475__;
  assign new_new_n41477__ = new_new_n41474__ & new_new_n41476__;
  assign new_new_n41478__ = ~new_new_n41472__ & ~new_new_n41477__;
  assign new_new_n41479__ = ys__n1386 & new_new_n41478__;
  assign new_new_n41480__ = ~new_new_n41470__ & ~new_new_n41479__;
  assign new_new_n41481__ = ~ys__n1386 & ~new_new_n41469__;
  assign ys__n31202 = ~new_new_n41480__ & ~new_new_n41481__;
  assign new_new_n41483__ = new_new_n41457__ & ~new_new_n41467__;
  assign new_new_n41484__ = new_new_n41469__ & new_new_n41483__;
  assign new_new_n41485__ = ~new_new_n41474__ & ~new_new_n41477__;
  assign new_new_n41486__ = ys__n1386 & new_new_n41485__;
  assign new_new_n41487__ = ~new_new_n41484__ & ~new_new_n41486__;
  assign ys__n31203 = ~new_new_n41481__ & ~new_new_n41487__;
  assign new_new_n41489__ = new_new_n39285__ & new_new_n39595__;
  assign new_new_n41490__ = ~new_new_n38879__ & ~new_new_n41489__;
  assign new_new_n41491__ = new_new_n39285__ & ~new_new_n39595__;
  assign new_new_n41492__ = ~new_new_n38879__ & ~new_new_n39620__;
  assign new_new_n41493__ = ~new_new_n41489__ & new_new_n41492__;
  assign new_new_n41494__ = ~new_new_n41491__ & new_new_n41493__;
  assign new_new_n41495__ = ~new_new_n41490__ & ~new_new_n41494__;
  assign new_new_n41496__ = ~ys__n30553 & ys__n30330;
  assign new_new_n41497__ = ys__n30553 & ~ys__n30330;
  assign new_new_n41498__ = ~new_new_n41496__ & ~new_new_n41497__;
  assign new_new_n41499__ = ~new_new_n41495__ & ~new_new_n41498__;
  assign new_new_n41500__ = new_new_n41495__ & new_new_n41498__;
  assign new_new_n41501__ = ~new_new_n41499__ & ~new_new_n41500__;
  assign new_new_n41502__ = ys__n39167 & ~new_new_n41501__;
  assign new_new_n41503__ = ys__n562 & ys__n47010;
  assign new_new_n41504__ = ys__n398 & ~ys__n33614;
  assign new_new_n41505__ = new_new_n41503__ & new_new_n41504__;
  assign new_new_n41506__ = ys__n2652 & ys__n17803;
  assign new_new_n41507__ = ys__n398 & ys__n33614;
  assign new_new_n41508__ = ~new_new_n41503__ & new_new_n41507__;
  assign new_new_n41509__ = ~new_new_n41506__ & ~new_new_n41508__;
  assign new_new_n41510__ = ~new_new_n41505__ & new_new_n41509__;
  assign new_new_n41511__ = ~new_new_n41502__ & new_new_n41510__;
  assign new_new_n41512__ = new_new_n12219__ & ~new_new_n41511__;
  assign new_new_n41513__ = ys__n30820 & ~new_new_n23477__;
  assign new_new_n41514__ = ys__n30819 & ~new_new_n23477__;
  assign new_new_n41515__ = ~new_new_n41513__ & ~new_new_n41514__;
  assign new_new_n41516__ = ys__n314 & new_new_n41515__;
  assign new_new_n41517__ = ~new_new_n24260__ & ~new_new_n41515__;
  assign new_new_n41518__ = ~new_new_n41516__ & ~new_new_n41517__;
  assign new_new_n41519__ = ~new_new_n12216__ & ~new_new_n41518__;
  assign new_new_n41520__ = ys__n314 & new_new_n12216__;
  assign new_new_n41521__ = ~new_new_n41519__ & ~new_new_n41520__;
  assign new_new_n41522__ = new_new_n12218__ & ~new_new_n41521__;
  assign new_new_n41523__ = ~new_new_n41512__ & ~new_new_n41522__;
  assign ys__n31207 = ys__n888 & ~new_new_n41523__;
  assign new_new_n41525__ = ~new_new_n41492__ & ~new_new_n41494__;
  assign new_new_n41526__ = ~new_new_n41498__ & ~new_new_n41525__;
  assign new_new_n41527__ = new_new_n41498__ & new_new_n41525__;
  assign new_new_n41528__ = ~new_new_n41526__ & ~new_new_n41527__;
  assign new_new_n41529__ = ys__n39167 & ~new_new_n41528__;
  assign new_new_n41530__ = ys__n562 & ys__n47011;
  assign new_new_n41531__ = new_new_n41503__ & ~new_new_n41530__;
  assign new_new_n41532__ = ~new_new_n41503__ & new_new_n41530__;
  assign new_new_n41533__ = ~new_new_n41531__ & ~new_new_n41532__;
  assign new_new_n41534__ = new_new_n41507__ & ~new_new_n41533__;
  assign new_new_n41535__ = ys__n2652 & ys__n17804;
  assign new_new_n41536__ = new_new_n41504__ & new_new_n41530__;
  assign new_new_n41537__ = ~new_new_n41535__ & ~new_new_n41536__;
  assign new_new_n41538__ = ~new_new_n41534__ & new_new_n41537__;
  assign new_new_n41539__ = ~new_new_n41529__ & new_new_n41538__;
  assign new_new_n41540__ = new_new_n12219__ & ~new_new_n41539__;
  assign new_new_n41541__ = ys__n170 & new_new_n41515__;
  assign new_new_n41542__ = ~new_new_n24329__ & ~new_new_n41515__;
  assign new_new_n41543__ = ~new_new_n41541__ & ~new_new_n41542__;
  assign new_new_n41544__ = ~new_new_n12216__ & ~new_new_n41543__;
  assign new_new_n41545__ = ys__n170 & new_new_n12216__;
  assign new_new_n41546__ = ~new_new_n41544__ & ~new_new_n41545__;
  assign new_new_n41547__ = new_new_n12218__ & ~new_new_n41546__;
  assign new_new_n41548__ = ~new_new_n41540__ & ~new_new_n41547__;
  assign ys__n31208 = ys__n888 & ~new_new_n41548__;
  assign new_new_n41550__ = ys__n562 & ys__n47012;
  assign new_new_n41551__ = new_new_n41503__ & new_new_n41530__;
  assign new_new_n41552__ = ~new_new_n41550__ & new_new_n41551__;
  assign new_new_n41553__ = new_new_n41550__ & ~new_new_n41551__;
  assign new_new_n41554__ = ~new_new_n41552__ & ~new_new_n41553__;
  assign new_new_n41555__ = new_new_n41507__ & ~new_new_n41554__;
  assign new_new_n41556__ = new_new_n41504__ & new_new_n41550__;
  assign new_new_n41557__ = ys__n2652 & ys__n17806;
  assign new_new_n41558__ = ys__n39167 & new_new_n41503__;
  assign new_new_n41559__ = ~new_new_n41557__ & ~new_new_n41558__;
  assign new_new_n41560__ = ~new_new_n41556__ & new_new_n41559__;
  assign new_new_n41561__ = ~new_new_n41555__ & new_new_n41560__;
  assign new_new_n41562__ = new_new_n12219__ & ~new_new_n41561__;
  assign new_new_n41563__ = ys__n380 & new_new_n41515__;
  assign new_new_n41564__ = ~new_new_n24401__ & ~new_new_n41515__;
  assign new_new_n41565__ = ~new_new_n41563__ & ~new_new_n41564__;
  assign new_new_n41566__ = ~new_new_n12216__ & ~new_new_n41565__;
  assign new_new_n41567__ = ys__n380 & new_new_n12216__;
  assign new_new_n41568__ = ~new_new_n41566__ & ~new_new_n41567__;
  assign new_new_n41569__ = new_new_n12218__ & ~new_new_n41568__;
  assign new_new_n41570__ = ~new_new_n41562__ & ~new_new_n41569__;
  assign ys__n31209 = ys__n888 & ~new_new_n41570__;
  assign new_new_n41572__ = ys__n562 & ys__n47013;
  assign new_new_n41573__ = new_new_n41550__ & new_new_n41551__;
  assign new_new_n41574__ = ~new_new_n41572__ & new_new_n41573__;
  assign new_new_n41575__ = new_new_n41572__ & ~new_new_n41573__;
  assign new_new_n41576__ = ~new_new_n41574__ & ~new_new_n41575__;
  assign new_new_n41577__ = new_new_n41507__ & ~new_new_n41576__;
  assign new_new_n41578__ = new_new_n41504__ & new_new_n41572__;
  assign new_new_n41579__ = ys__n2652 & ys__n17807;
  assign new_new_n41580__ = ys__n39167 & new_new_n41530__;
  assign new_new_n41581__ = ~new_new_n41579__ & ~new_new_n41580__;
  assign new_new_n41582__ = ~new_new_n41578__ & new_new_n41581__;
  assign new_new_n41583__ = ~new_new_n41577__ & new_new_n41582__;
  assign new_new_n41584__ = new_new_n12219__ & ~new_new_n41583__;
  assign new_new_n41585__ = ys__n378 & new_new_n41515__;
  assign new_new_n41586__ = ~new_new_n24476__ & ~new_new_n41515__;
  assign new_new_n41587__ = ~new_new_n41585__ & ~new_new_n41586__;
  assign new_new_n41588__ = ~new_new_n12216__ & ~new_new_n41587__;
  assign new_new_n41589__ = ys__n378 & new_new_n12216__;
  assign new_new_n41590__ = ~new_new_n41588__ & ~new_new_n41589__;
  assign new_new_n41591__ = new_new_n12218__ & ~new_new_n41590__;
  assign new_new_n41592__ = ~new_new_n41584__ & ~new_new_n41591__;
  assign ys__n31210 = ys__n888 & ~new_new_n41592__;
  assign new_new_n41594__ = ys__n562 & ys__n47014;
  assign new_new_n41595__ = new_new_n41550__ & new_new_n41572__;
  assign new_new_n41596__ = new_new_n41551__ & new_new_n41595__;
  assign new_new_n41597__ = ~new_new_n41594__ & new_new_n41596__;
  assign new_new_n41598__ = new_new_n41594__ & ~new_new_n41596__;
  assign new_new_n41599__ = ~new_new_n41597__ & ~new_new_n41598__;
  assign new_new_n41600__ = new_new_n41507__ & ~new_new_n41599__;
  assign new_new_n41601__ = new_new_n41504__ & new_new_n41594__;
  assign new_new_n41602__ = ys__n2652 & ys__n17809;
  assign new_new_n41603__ = ys__n39167 & new_new_n41550__;
  assign new_new_n41604__ = ~new_new_n41602__ & ~new_new_n41603__;
  assign new_new_n41605__ = ~new_new_n41601__ & new_new_n41604__;
  assign new_new_n41606__ = ~new_new_n41600__ & new_new_n41605__;
  assign new_new_n41607__ = new_new_n12219__ & ~new_new_n41606__;
  assign new_new_n41608__ = ys__n382 & new_new_n41515__;
  assign new_new_n41609__ = ~new_new_n24553__ & ~new_new_n41515__;
  assign new_new_n41610__ = ~new_new_n41608__ & ~new_new_n41609__;
  assign new_new_n41611__ = ~new_new_n12216__ & ~new_new_n41610__;
  assign new_new_n41612__ = ys__n382 & new_new_n12216__;
  assign new_new_n41613__ = ~new_new_n41611__ & ~new_new_n41612__;
  assign new_new_n41614__ = new_new_n12218__ & ~new_new_n41613__;
  assign new_new_n41615__ = ~new_new_n41607__ & ~new_new_n41614__;
  assign ys__n31211 = ys__n888 & ~new_new_n41615__;
  assign new_new_n41617__ = ys__n562 & ys__n47015;
  assign new_new_n41618__ = new_new_n41594__ & new_new_n41596__;
  assign new_new_n41619__ = ~new_new_n41617__ & new_new_n41618__;
  assign new_new_n41620__ = new_new_n41617__ & ~new_new_n41618__;
  assign new_new_n41621__ = ~new_new_n41619__ & ~new_new_n41620__;
  assign new_new_n41622__ = new_new_n41507__ & ~new_new_n41621__;
  assign new_new_n41623__ = new_new_n41504__ & new_new_n41617__;
  assign new_new_n41624__ = ys__n2652 & ys__n17810;
  assign new_new_n41625__ = ys__n39167 & new_new_n41572__;
  assign new_new_n41626__ = ~new_new_n41624__ & ~new_new_n41625__;
  assign new_new_n41627__ = ~new_new_n41623__ & new_new_n41626__;
  assign new_new_n41628__ = ~new_new_n41622__ & new_new_n41627__;
  assign new_new_n41629__ = new_new_n12219__ & ~new_new_n41628__;
  assign new_new_n41630__ = ys__n374 & new_new_n41515__;
  assign new_new_n41631__ = ~new_new_n24629__ & ~new_new_n41515__;
  assign new_new_n41632__ = ~new_new_n41630__ & ~new_new_n41631__;
  assign new_new_n41633__ = ~new_new_n12216__ & ~new_new_n41632__;
  assign new_new_n41634__ = ys__n374 & new_new_n12216__;
  assign new_new_n41635__ = ~new_new_n41633__ & ~new_new_n41634__;
  assign new_new_n41636__ = new_new_n12218__ & ~new_new_n41635__;
  assign new_new_n41637__ = ~new_new_n41629__ & ~new_new_n41636__;
  assign ys__n31212 = ys__n888 & ~new_new_n41637__;
  assign new_new_n41639__ = ys__n562 & ys__n47016;
  assign new_new_n41640__ = new_new_n41594__ & new_new_n41617__;
  assign new_new_n41641__ = new_new_n41596__ & new_new_n41640__;
  assign new_new_n41642__ = ~new_new_n41639__ & new_new_n41641__;
  assign new_new_n41643__ = new_new_n41639__ & ~new_new_n41641__;
  assign new_new_n41644__ = ~new_new_n41642__ & ~new_new_n41643__;
  assign new_new_n41645__ = new_new_n41507__ & ~new_new_n41644__;
  assign new_new_n41646__ = new_new_n41504__ & new_new_n41639__;
  assign new_new_n41647__ = ys__n2652 & ys__n17812;
  assign new_new_n41648__ = ys__n39167 & new_new_n41594__;
  assign new_new_n41649__ = ~new_new_n41647__ & ~new_new_n41648__;
  assign new_new_n41650__ = ~new_new_n41646__ & new_new_n41649__;
  assign new_new_n41651__ = ~new_new_n41645__ & new_new_n41650__;
  assign new_new_n41652__ = new_new_n12219__ & ~new_new_n41651__;
  assign new_new_n41653__ = ys__n376 & new_new_n41515__;
  assign new_new_n41654__ = ~new_new_n24709__ & ~new_new_n41515__;
  assign new_new_n41655__ = ~new_new_n41653__ & ~new_new_n41654__;
  assign new_new_n41656__ = ~new_new_n12216__ & ~new_new_n41655__;
  assign new_new_n41657__ = ys__n376 & new_new_n12216__;
  assign new_new_n41658__ = ~new_new_n41656__ & ~new_new_n41657__;
  assign new_new_n41659__ = new_new_n12218__ & ~new_new_n41658__;
  assign new_new_n41660__ = ~new_new_n41652__ & ~new_new_n41659__;
  assign ys__n31213 = ys__n888 & ~new_new_n41660__;
  assign new_new_n41662__ = ys__n562 & ys__n47017;
  assign new_new_n41663__ = new_new_n41639__ & new_new_n41641__;
  assign new_new_n41664__ = ~new_new_n41662__ & new_new_n41663__;
  assign new_new_n41665__ = new_new_n41662__ & ~new_new_n41663__;
  assign new_new_n41666__ = ~new_new_n41664__ & ~new_new_n41665__;
  assign new_new_n41667__ = new_new_n41507__ & ~new_new_n41666__;
  assign new_new_n41668__ = new_new_n41504__ & new_new_n41662__;
  assign new_new_n41669__ = ys__n2652 & ys__n17813;
  assign new_new_n41670__ = ys__n39167 & new_new_n41617__;
  assign new_new_n41671__ = ~new_new_n41669__ & ~new_new_n41670__;
  assign new_new_n41672__ = ~new_new_n41668__ & new_new_n41671__;
  assign new_new_n41673__ = ~new_new_n41667__ & new_new_n41672__;
  assign new_new_n41674__ = new_new_n12219__ & ~new_new_n41673__;
  assign new_new_n41675__ = ys__n372 & new_new_n41515__;
  assign new_new_n41676__ = ~new_new_n24785__ & ~new_new_n41515__;
  assign new_new_n41677__ = ~new_new_n41675__ & ~new_new_n41676__;
  assign new_new_n41678__ = ~new_new_n12216__ & ~new_new_n41677__;
  assign new_new_n41679__ = ys__n372 & new_new_n12216__;
  assign new_new_n41680__ = ~new_new_n41678__ & ~new_new_n41679__;
  assign new_new_n41681__ = new_new_n12218__ & ~new_new_n41680__;
  assign new_new_n41682__ = ~new_new_n41674__ & ~new_new_n41681__;
  assign ys__n31214 = ys__n888 & ~new_new_n41682__;
  assign new_new_n41684__ = ys__n562 & ys__n47018;
  assign new_new_n41685__ = new_new_n41639__ & new_new_n41662__;
  assign new_new_n41686__ = new_new_n41640__ & new_new_n41685__;
  assign new_new_n41687__ = new_new_n41596__ & new_new_n41686__;
  assign new_new_n41688__ = ~new_new_n41684__ & new_new_n41687__;
  assign new_new_n41689__ = new_new_n41684__ & ~new_new_n41687__;
  assign new_new_n41690__ = ~new_new_n41688__ & ~new_new_n41689__;
  assign new_new_n41691__ = new_new_n41507__ & ~new_new_n41690__;
  assign new_new_n41692__ = new_new_n41504__ & new_new_n41684__;
  assign new_new_n41693__ = ys__n2652 & ys__n17815;
  assign new_new_n41694__ = ys__n39167 & new_new_n41639__;
  assign new_new_n41695__ = ~new_new_n41693__ & ~new_new_n41694__;
  assign new_new_n41696__ = ~new_new_n41692__ & new_new_n41695__;
  assign new_new_n41697__ = ~new_new_n41691__ & new_new_n41696__;
  assign new_new_n41698__ = new_new_n12219__ & ~new_new_n41697__;
  assign new_new_n41699__ = ys__n384 & new_new_n41515__;
  assign new_new_n41700__ = ~new_new_n24866__ & ~new_new_n41515__;
  assign new_new_n41701__ = ~new_new_n41699__ & ~new_new_n41700__;
  assign new_new_n41702__ = ~new_new_n12216__ & ~new_new_n41701__;
  assign new_new_n41703__ = ys__n384 & new_new_n12216__;
  assign new_new_n41704__ = ~new_new_n41702__ & ~new_new_n41703__;
  assign new_new_n41705__ = new_new_n12218__ & ~new_new_n41704__;
  assign new_new_n41706__ = ~new_new_n41698__ & ~new_new_n41705__;
  assign ys__n31215 = ys__n888 & ~new_new_n41706__;
  assign new_new_n41708__ = ys__n562 & ys__n47019;
  assign new_new_n41709__ = new_new_n41684__ & new_new_n41687__;
  assign new_new_n41710__ = ~new_new_n41708__ & new_new_n41709__;
  assign new_new_n41711__ = new_new_n41708__ & ~new_new_n41709__;
  assign new_new_n41712__ = ~new_new_n41710__ & ~new_new_n41711__;
  assign new_new_n41713__ = new_new_n41507__ & ~new_new_n41712__;
  assign new_new_n41714__ = new_new_n41504__ & new_new_n41708__;
  assign new_new_n41715__ = ys__n2652 & ys__n17816;
  assign new_new_n41716__ = ys__n39167 & new_new_n41662__;
  assign new_new_n41717__ = ~new_new_n41715__ & ~new_new_n41716__;
  assign new_new_n41718__ = ~new_new_n41714__ & new_new_n41717__;
  assign new_new_n41719__ = ~new_new_n41713__ & new_new_n41718__;
  assign new_new_n41720__ = new_new_n12219__ & ~new_new_n41719__;
  assign new_new_n41721__ = ys__n366 & new_new_n41515__;
  assign new_new_n41722__ = ~new_new_n24942__ & ~new_new_n41515__;
  assign new_new_n41723__ = ~new_new_n41721__ & ~new_new_n41722__;
  assign new_new_n41724__ = ~new_new_n12216__ & ~new_new_n41723__;
  assign new_new_n41725__ = ys__n366 & new_new_n12216__;
  assign new_new_n41726__ = ~new_new_n41724__ & ~new_new_n41725__;
  assign new_new_n41727__ = new_new_n12218__ & ~new_new_n41726__;
  assign new_new_n41728__ = ~new_new_n41720__ & ~new_new_n41727__;
  assign ys__n31216 = ys__n888 & ~new_new_n41728__;
  assign new_new_n41730__ = ys__n562 & ys__n47020;
  assign new_new_n41731__ = new_new_n41684__ & new_new_n41708__;
  assign new_new_n41732__ = new_new_n41687__ & new_new_n41731__;
  assign new_new_n41733__ = ~new_new_n41730__ & new_new_n41732__;
  assign new_new_n41734__ = new_new_n41730__ & ~new_new_n41732__;
  assign new_new_n41735__ = ~new_new_n41733__ & ~new_new_n41734__;
  assign new_new_n41736__ = new_new_n41507__ & ~new_new_n41735__;
  assign new_new_n41737__ = new_new_n41504__ & new_new_n41730__;
  assign new_new_n41738__ = ys__n2652 & ys__n17818;
  assign new_new_n41739__ = ys__n39167 & new_new_n41684__;
  assign new_new_n41740__ = ~new_new_n41738__ & ~new_new_n41739__;
  assign new_new_n41741__ = ~new_new_n41737__ & new_new_n41740__;
  assign new_new_n41742__ = ~new_new_n41736__ & new_new_n41741__;
  assign new_new_n41743__ = new_new_n12219__ & ~new_new_n41742__;
  assign new_new_n41744__ = ys__n368 & new_new_n41515__;
  assign new_new_n41745__ = ~new_new_n25022__ & ~new_new_n41515__;
  assign new_new_n41746__ = ~new_new_n41744__ & ~new_new_n41745__;
  assign new_new_n41747__ = ~new_new_n12216__ & ~new_new_n41746__;
  assign new_new_n41748__ = ys__n368 & new_new_n12216__;
  assign new_new_n41749__ = ~new_new_n41747__ & ~new_new_n41748__;
  assign new_new_n41750__ = new_new_n12218__ & ~new_new_n41749__;
  assign new_new_n41751__ = ~new_new_n41743__ & ~new_new_n41750__;
  assign ys__n31217 = ys__n888 & ~new_new_n41751__;
  assign new_new_n41753__ = ys__n562 & ys__n47021;
  assign new_new_n41754__ = new_new_n41730__ & new_new_n41732__;
  assign new_new_n41755__ = ~new_new_n41753__ & new_new_n41754__;
  assign new_new_n41756__ = new_new_n41753__ & ~new_new_n41754__;
  assign new_new_n41757__ = ~new_new_n41755__ & ~new_new_n41756__;
  assign new_new_n41758__ = new_new_n41507__ & ~new_new_n41757__;
  assign new_new_n41759__ = new_new_n41504__ & new_new_n41753__;
  assign new_new_n41760__ = ys__n2652 & ys__n17819;
  assign new_new_n41761__ = ys__n39167 & new_new_n41708__;
  assign new_new_n41762__ = ~new_new_n41760__ & ~new_new_n41761__;
  assign new_new_n41763__ = ~new_new_n41759__ & new_new_n41762__;
  assign new_new_n41764__ = ~new_new_n41758__ & new_new_n41763__;
  assign new_new_n41765__ = new_new_n12219__ & ~new_new_n41764__;
  assign new_new_n41766__ = ys__n364 & new_new_n41515__;
  assign new_new_n41767__ = ~new_new_n25098__ & ~new_new_n41515__;
  assign new_new_n41768__ = ~new_new_n41766__ & ~new_new_n41767__;
  assign new_new_n41769__ = ~new_new_n12216__ & ~new_new_n41768__;
  assign new_new_n41770__ = ys__n364 & new_new_n12216__;
  assign new_new_n41771__ = ~new_new_n41769__ & ~new_new_n41770__;
  assign new_new_n41772__ = new_new_n12218__ & ~new_new_n41771__;
  assign new_new_n41773__ = ~new_new_n41765__ & ~new_new_n41772__;
  assign ys__n31218 = ys__n888 & ~new_new_n41773__;
  assign new_new_n41775__ = ys__n562 & ys__n47022;
  assign new_new_n41776__ = new_new_n41730__ & new_new_n41753__;
  assign new_new_n41777__ = new_new_n41731__ & new_new_n41776__;
  assign new_new_n41778__ = new_new_n41687__ & new_new_n41777__;
  assign new_new_n41779__ = ~new_new_n41775__ & new_new_n41778__;
  assign new_new_n41780__ = new_new_n41775__ & ~new_new_n41778__;
  assign new_new_n41781__ = ~new_new_n41779__ & ~new_new_n41780__;
  assign new_new_n41782__ = new_new_n41507__ & ~new_new_n41781__;
  assign new_new_n41783__ = new_new_n41504__ & new_new_n41775__;
  assign new_new_n41784__ = ys__n2652 & ys__n17821;
  assign new_new_n41785__ = ys__n39167 & new_new_n41730__;
  assign new_new_n41786__ = ~new_new_n41784__ & ~new_new_n41785__;
  assign new_new_n41787__ = ~new_new_n41783__ & new_new_n41786__;
  assign new_new_n41788__ = ~new_new_n41782__ & new_new_n41787__;
  assign new_new_n41789__ = new_new_n12219__ & ~new_new_n41788__;
  assign new_new_n41790__ = ys__n370 & new_new_n41515__;
  assign new_new_n41791__ = ~new_new_n25182__ & ~new_new_n41515__;
  assign new_new_n41792__ = ~new_new_n41790__ & ~new_new_n41791__;
  assign new_new_n41793__ = ~new_new_n12216__ & ~new_new_n41792__;
  assign new_new_n41794__ = ys__n370 & new_new_n12216__;
  assign new_new_n41795__ = ~new_new_n41793__ & ~new_new_n41794__;
  assign new_new_n41796__ = new_new_n12218__ & ~new_new_n41795__;
  assign new_new_n41797__ = ~new_new_n41789__ & ~new_new_n41796__;
  assign ys__n31219 = ys__n888 & ~new_new_n41797__;
  assign new_new_n41799__ = ys__n562 & ys__n47023;
  assign new_new_n41800__ = new_new_n41775__ & new_new_n41778__;
  assign new_new_n41801__ = ~new_new_n41799__ & new_new_n41800__;
  assign new_new_n41802__ = new_new_n41799__ & ~new_new_n41800__;
  assign new_new_n41803__ = ~new_new_n41801__ & ~new_new_n41802__;
  assign new_new_n41804__ = new_new_n41507__ & ~new_new_n41803__;
  assign new_new_n41805__ = new_new_n41504__ & new_new_n41799__;
  assign new_new_n41806__ = ys__n2652 & ys__n17822;
  assign new_new_n41807__ = ys__n39167 & new_new_n41753__;
  assign new_new_n41808__ = ~new_new_n41806__ & ~new_new_n41807__;
  assign new_new_n41809__ = ~new_new_n41805__ & new_new_n41808__;
  assign new_new_n41810__ = ~new_new_n41804__ & new_new_n41809__;
  assign new_new_n41811__ = new_new_n12219__ & ~new_new_n41810__;
  assign new_new_n41812__ = ys__n360 & new_new_n41515__;
  assign new_new_n41813__ = ~new_new_n25258__ & ~new_new_n41515__;
  assign new_new_n41814__ = ~new_new_n41812__ & ~new_new_n41813__;
  assign new_new_n41815__ = ~new_new_n12216__ & ~new_new_n41814__;
  assign new_new_n41816__ = ys__n360 & new_new_n12216__;
  assign new_new_n41817__ = ~new_new_n41815__ & ~new_new_n41816__;
  assign new_new_n41818__ = new_new_n12218__ & ~new_new_n41817__;
  assign new_new_n41819__ = ~new_new_n41811__ & ~new_new_n41818__;
  assign ys__n31220 = ys__n888 & ~new_new_n41819__;
  assign new_new_n41821__ = ys__n562 & ys__n47024;
  assign new_new_n41822__ = new_new_n41775__ & new_new_n41799__;
  assign new_new_n41823__ = new_new_n41778__ & new_new_n41822__;
  assign new_new_n41824__ = ~new_new_n41821__ & new_new_n41823__;
  assign new_new_n41825__ = new_new_n41821__ & ~new_new_n41823__;
  assign new_new_n41826__ = ~new_new_n41824__ & ~new_new_n41825__;
  assign new_new_n41827__ = new_new_n41507__ & ~new_new_n41826__;
  assign new_new_n41828__ = new_new_n41504__ & new_new_n41821__;
  assign new_new_n41829__ = ys__n2652 & ys__n17824;
  assign new_new_n41830__ = ys__n39167 & new_new_n41775__;
  assign new_new_n41831__ = ~new_new_n41829__ & ~new_new_n41830__;
  assign new_new_n41832__ = ~new_new_n41828__ & new_new_n41831__;
  assign new_new_n41833__ = ~new_new_n41827__ & new_new_n41832__;
  assign new_new_n41834__ = new_new_n12219__ & ~new_new_n41833__;
  assign new_new_n41835__ = ys__n362 & new_new_n41515__;
  assign new_new_n41836__ = ~new_new_n25338__ & ~new_new_n41515__;
  assign new_new_n41837__ = ~new_new_n41835__ & ~new_new_n41836__;
  assign new_new_n41838__ = ~new_new_n12216__ & ~new_new_n41837__;
  assign new_new_n41839__ = ys__n362 & new_new_n12216__;
  assign new_new_n41840__ = ~new_new_n41838__ & ~new_new_n41839__;
  assign new_new_n41841__ = new_new_n12218__ & ~new_new_n41840__;
  assign new_new_n41842__ = ~new_new_n41834__ & ~new_new_n41841__;
  assign ys__n31221 = ys__n888 & ~new_new_n41842__;
  assign new_new_n41844__ = ys__n562 & ys__n47025;
  assign new_new_n41845__ = new_new_n41821__ & new_new_n41823__;
  assign new_new_n41846__ = ~new_new_n41844__ & new_new_n41845__;
  assign new_new_n41847__ = new_new_n41844__ & ~new_new_n41845__;
  assign new_new_n41848__ = ~new_new_n41846__ & ~new_new_n41847__;
  assign new_new_n41849__ = new_new_n41507__ & ~new_new_n41848__;
  assign new_new_n41850__ = new_new_n41504__ & new_new_n41844__;
  assign new_new_n41851__ = ys__n2652 & ys__n17825;
  assign new_new_n41852__ = ys__n39167 & new_new_n41799__;
  assign new_new_n41853__ = ~new_new_n41851__ & ~new_new_n41852__;
  assign new_new_n41854__ = ~new_new_n41850__ & new_new_n41853__;
  assign new_new_n41855__ = ~new_new_n41849__ & new_new_n41854__;
  assign new_new_n41856__ = new_new_n12219__ & ~new_new_n41855__;
  assign new_new_n41857__ = ys__n358 & new_new_n41515__;
  assign new_new_n41858__ = ~new_new_n25412__ & ~new_new_n41515__;
  assign new_new_n41859__ = ~new_new_n41857__ & ~new_new_n41858__;
  assign new_new_n41860__ = ~new_new_n12216__ & ~new_new_n41859__;
  assign new_new_n41861__ = ys__n358 & new_new_n12216__;
  assign new_new_n41862__ = ~new_new_n41860__ & ~new_new_n41861__;
  assign new_new_n41863__ = new_new_n12218__ & ~new_new_n41862__;
  assign new_new_n41864__ = ~new_new_n41856__ & ~new_new_n41863__;
  assign ys__n31222 = ys__n888 & ~new_new_n41864__;
  assign new_new_n41866__ = ys__n562 & ys__n47026;
  assign new_new_n41867__ = new_new_n41821__ & new_new_n41844__;
  assign new_new_n41868__ = new_new_n41822__ & new_new_n41867__;
  assign new_new_n41869__ = new_new_n41777__ & new_new_n41868__;
  assign new_new_n41870__ = new_new_n41687__ & new_new_n41869__;
  assign new_new_n41871__ = ~new_new_n41866__ & new_new_n41870__;
  assign new_new_n41872__ = new_new_n41866__ & ~new_new_n41870__;
  assign new_new_n41873__ = ~new_new_n41871__ & ~new_new_n41872__;
  assign new_new_n41874__ = new_new_n41507__ & ~new_new_n41873__;
  assign new_new_n41875__ = new_new_n41504__ & new_new_n41866__;
  assign new_new_n41876__ = ys__n2652 & ys__n17827;
  assign new_new_n41877__ = ys__n39167 & new_new_n41821__;
  assign new_new_n41878__ = ~new_new_n41876__ & ~new_new_n41877__;
  assign new_new_n41879__ = ~new_new_n41875__ & new_new_n41878__;
  assign new_new_n41880__ = ~new_new_n41874__ & new_new_n41879__;
  assign new_new_n41881__ = new_new_n12219__ & ~new_new_n41880__;
  assign new_new_n41882__ = ~new_new_n24234__ & new_new_n41515__;
  assign new_new_n41883__ = ~new_new_n24227__ & ~new_new_n41515__;
  assign new_new_n41884__ = ~new_new_n41882__ & ~new_new_n41883__;
  assign new_new_n41885__ = ~new_new_n12216__ & ~new_new_n41884__;
  assign new_new_n41886__ = new_new_n12216__ & ~new_new_n24234__;
  assign new_new_n41887__ = ~new_new_n41885__ & ~new_new_n41886__;
  assign new_new_n41888__ = new_new_n12218__ & ~new_new_n41887__;
  assign new_new_n41889__ = ~new_new_n41881__ & ~new_new_n41888__;
  assign ys__n31223 = ys__n888 & ~new_new_n41889__;
  assign new_new_n41891__ = ys__n562 & ys__n47027;
  assign new_new_n41892__ = new_new_n41866__ & new_new_n41870__;
  assign new_new_n41893__ = ~new_new_n41891__ & new_new_n41892__;
  assign new_new_n41894__ = new_new_n41891__ & ~new_new_n41892__;
  assign new_new_n41895__ = ~new_new_n41893__ & ~new_new_n41894__;
  assign new_new_n41896__ = new_new_n41507__ & ~new_new_n41895__;
  assign new_new_n41897__ = new_new_n41504__ & new_new_n41891__;
  assign new_new_n41898__ = ys__n2652 & ys__n17828;
  assign new_new_n41899__ = ys__n39167 & new_new_n41844__;
  assign new_new_n41900__ = ~new_new_n41898__ & ~new_new_n41899__;
  assign new_new_n41901__ = ~new_new_n41897__ & new_new_n41900__;
  assign new_new_n41902__ = ~new_new_n41896__ & new_new_n41901__;
  assign new_new_n41903__ = new_new_n12219__ & ~new_new_n41902__;
  assign new_new_n41904__ = ~new_new_n24312__ & new_new_n41515__;
  assign new_new_n41905__ = ~new_new_n24306__ & ~new_new_n41515__;
  assign new_new_n41906__ = ~new_new_n41904__ & ~new_new_n41905__;
  assign new_new_n41907__ = ~new_new_n12216__ & ~new_new_n41906__;
  assign new_new_n41908__ = new_new_n12216__ & ~new_new_n24312__;
  assign new_new_n41909__ = ~new_new_n41907__ & ~new_new_n41908__;
  assign new_new_n41910__ = new_new_n12218__ & ~new_new_n41909__;
  assign new_new_n41911__ = ~new_new_n41903__ & ~new_new_n41910__;
  assign ys__n31224 = ys__n888 & ~new_new_n41911__;
  assign new_new_n41913__ = ys__n562 & ys__n47028;
  assign new_new_n41914__ = new_new_n41866__ & new_new_n41891__;
  assign new_new_n41915__ = new_new_n41870__ & new_new_n41914__;
  assign new_new_n41916__ = ~new_new_n41913__ & new_new_n41915__;
  assign new_new_n41917__ = new_new_n41913__ & ~new_new_n41915__;
  assign new_new_n41918__ = ~new_new_n41916__ & ~new_new_n41917__;
  assign new_new_n41919__ = new_new_n41507__ & ~new_new_n41918__;
  assign new_new_n41920__ = new_new_n41504__ & new_new_n41913__;
  assign new_new_n41921__ = ys__n2652 & ys__n17830;
  assign new_new_n41922__ = ys__n39167 & new_new_n41866__;
  assign new_new_n41923__ = ~new_new_n41921__ & ~new_new_n41922__;
  assign new_new_n41924__ = ~new_new_n41920__ & new_new_n41923__;
  assign new_new_n41925__ = ~new_new_n41919__ & new_new_n41924__;
  assign new_new_n41926__ = new_new_n12219__ & ~new_new_n41925__;
  assign new_new_n41927__ = ~new_new_n24384__ & new_new_n41515__;
  assign new_new_n41928__ = ~new_new_n24378__ & ~new_new_n41515__;
  assign new_new_n41929__ = ~new_new_n41927__ & ~new_new_n41928__;
  assign new_new_n41930__ = ~new_new_n12216__ & ~new_new_n41929__;
  assign new_new_n41931__ = new_new_n12216__ & ~new_new_n24384__;
  assign new_new_n41932__ = ~new_new_n41930__ & ~new_new_n41931__;
  assign new_new_n41933__ = new_new_n12218__ & ~new_new_n41932__;
  assign new_new_n41934__ = ~new_new_n41926__ & ~new_new_n41933__;
  assign ys__n31225 = ys__n888 & ~new_new_n41934__;
  assign new_new_n41936__ = ys__n562 & ys__n47029;
  assign new_new_n41937__ = new_new_n41913__ & new_new_n41915__;
  assign new_new_n41938__ = ~new_new_n41936__ & new_new_n41937__;
  assign new_new_n41939__ = new_new_n41936__ & ~new_new_n41937__;
  assign new_new_n41940__ = ~new_new_n41938__ & ~new_new_n41939__;
  assign new_new_n41941__ = new_new_n41507__ & ~new_new_n41940__;
  assign new_new_n41942__ = new_new_n41504__ & new_new_n41936__;
  assign new_new_n41943__ = ys__n2652 & ys__n17831;
  assign new_new_n41944__ = ys__n39167 & new_new_n41891__;
  assign new_new_n41945__ = ~new_new_n41943__ & ~new_new_n41944__;
  assign new_new_n41946__ = ~new_new_n41942__ & new_new_n41945__;
  assign new_new_n41947__ = ~new_new_n41941__ & new_new_n41946__;
  assign new_new_n41948__ = new_new_n12219__ & ~new_new_n41947__;
  assign new_new_n41949__ = ~new_new_n24459__ & new_new_n41515__;
  assign new_new_n41950__ = ~new_new_n24451__ & ~new_new_n41515__;
  assign new_new_n41951__ = ~new_new_n41949__ & ~new_new_n41950__;
  assign new_new_n41952__ = ~new_new_n12216__ & ~new_new_n41951__;
  assign new_new_n41953__ = new_new_n12216__ & ~new_new_n24459__;
  assign new_new_n41954__ = ~new_new_n41952__ & ~new_new_n41953__;
  assign new_new_n41955__ = new_new_n12218__ & ~new_new_n41954__;
  assign new_new_n41956__ = ~new_new_n41948__ & ~new_new_n41955__;
  assign ys__n31226 = ys__n888 & ~new_new_n41956__;
  assign new_new_n41958__ = ys__n562 & ys__n47030;
  assign new_new_n41959__ = new_new_n41913__ & new_new_n41936__;
  assign new_new_n41960__ = new_new_n41914__ & new_new_n41959__;
  assign new_new_n41961__ = new_new_n41870__ & new_new_n41960__;
  assign new_new_n41962__ = ~new_new_n41958__ & new_new_n41961__;
  assign new_new_n41963__ = new_new_n41958__ & ~new_new_n41961__;
  assign new_new_n41964__ = ~new_new_n41962__ & ~new_new_n41963__;
  assign new_new_n41965__ = new_new_n41507__ & ~new_new_n41964__;
  assign new_new_n41966__ = new_new_n41504__ & new_new_n41958__;
  assign new_new_n41967__ = ys__n2652 & ys__n17833;
  assign new_new_n41968__ = ys__n39167 & new_new_n41913__;
  assign new_new_n41969__ = ~new_new_n41967__ & ~new_new_n41968__;
  assign new_new_n41970__ = ~new_new_n41966__ & new_new_n41969__;
  assign new_new_n41971__ = ~new_new_n41965__ & new_new_n41970__;
  assign new_new_n41972__ = new_new_n12219__ & ~new_new_n41971__;
  assign new_new_n41973__ = ~new_new_n24536__ & new_new_n41515__;
  assign new_new_n41974__ = ~new_new_n24530__ & ~new_new_n41515__;
  assign new_new_n41975__ = ~new_new_n41973__ & ~new_new_n41974__;
  assign new_new_n41976__ = ~new_new_n12216__ & ~new_new_n41975__;
  assign new_new_n41977__ = new_new_n12216__ & ~new_new_n24536__;
  assign new_new_n41978__ = ~new_new_n41976__ & ~new_new_n41977__;
  assign new_new_n41979__ = new_new_n12218__ & ~new_new_n41978__;
  assign new_new_n41980__ = ~new_new_n41972__ & ~new_new_n41979__;
  assign ys__n31227 = ys__n888 & ~new_new_n41980__;
  assign new_new_n41982__ = ys__n562 & ys__n47031;
  assign new_new_n41983__ = new_new_n41958__ & new_new_n41961__;
  assign new_new_n41984__ = ~new_new_n41982__ & new_new_n41983__;
  assign new_new_n41985__ = new_new_n41982__ & ~new_new_n41983__;
  assign new_new_n41986__ = ~new_new_n41984__ & ~new_new_n41985__;
  assign new_new_n41987__ = new_new_n41507__ & ~new_new_n41986__;
  assign new_new_n41988__ = new_new_n41504__ & new_new_n41982__;
  assign new_new_n41989__ = ys__n2652 & ys__n17834;
  assign new_new_n41990__ = ys__n39167 & new_new_n41936__;
  assign new_new_n41991__ = ~new_new_n41989__ & ~new_new_n41990__;
  assign new_new_n41992__ = ~new_new_n41988__ & new_new_n41991__;
  assign new_new_n41993__ = ~new_new_n41987__ & new_new_n41992__;
  assign new_new_n41994__ = new_new_n12219__ & ~new_new_n41993__;
  assign new_new_n41995__ = ~new_new_n24611__ & new_new_n41515__;
  assign new_new_n41996__ = ~new_new_n24603__ & ~new_new_n41515__;
  assign new_new_n41997__ = ~new_new_n41995__ & ~new_new_n41996__;
  assign new_new_n41998__ = ~new_new_n12216__ & ~new_new_n41997__;
  assign new_new_n41999__ = new_new_n12216__ & ~new_new_n24611__;
  assign new_new_n42000__ = ~new_new_n41998__ & ~new_new_n41999__;
  assign new_new_n42001__ = new_new_n12218__ & ~new_new_n42000__;
  assign new_new_n42002__ = ~new_new_n41994__ & ~new_new_n42001__;
  assign ys__n31228 = ys__n888 & ~new_new_n42002__;
  assign new_new_n42004__ = ys__n562 & ys__n47032;
  assign new_new_n42005__ = new_new_n41958__ & new_new_n41982__;
  assign new_new_n42006__ = new_new_n41961__ & new_new_n42005__;
  assign new_new_n42007__ = ~new_new_n42004__ & new_new_n42006__;
  assign new_new_n42008__ = new_new_n42004__ & ~new_new_n42006__;
  assign new_new_n42009__ = ~new_new_n42007__ & ~new_new_n42008__;
  assign new_new_n42010__ = new_new_n41507__ & ~new_new_n42009__;
  assign new_new_n42011__ = new_new_n41504__ & new_new_n42004__;
  assign new_new_n42012__ = ys__n2652 & ys__n17836;
  assign new_new_n42013__ = ys__n39167 & new_new_n41958__;
  assign new_new_n42014__ = ~new_new_n42012__ & ~new_new_n42013__;
  assign new_new_n42015__ = ~new_new_n42011__ & new_new_n42014__;
  assign new_new_n42016__ = ~new_new_n42010__ & new_new_n42015__;
  assign new_new_n42017__ = new_new_n12219__ & ~new_new_n42016__;
  assign new_new_n42018__ = ~new_new_n24691__ & new_new_n41515__;
  assign new_new_n42019__ = ~new_new_n24683__ & ~new_new_n41515__;
  assign new_new_n42020__ = ~new_new_n42018__ & ~new_new_n42019__;
  assign new_new_n42021__ = ~new_new_n12216__ & ~new_new_n42020__;
  assign new_new_n42022__ = new_new_n12216__ & ~new_new_n24691__;
  assign new_new_n42023__ = ~new_new_n42021__ & ~new_new_n42022__;
  assign new_new_n42024__ = new_new_n12218__ & ~new_new_n42023__;
  assign new_new_n42025__ = ~new_new_n42017__ & ~new_new_n42024__;
  assign ys__n31229 = ys__n888 & ~new_new_n42025__;
  assign new_new_n42027__ = ys__n562 & ys__n47033;
  assign new_new_n42028__ = new_new_n42004__ & new_new_n42006__;
  assign new_new_n42029__ = ~new_new_n42027__ & new_new_n42028__;
  assign new_new_n42030__ = new_new_n42027__ & ~new_new_n42028__;
  assign new_new_n42031__ = ~new_new_n42029__ & ~new_new_n42030__;
  assign new_new_n42032__ = new_new_n41507__ & ~new_new_n42031__;
  assign new_new_n42033__ = new_new_n41504__ & new_new_n42027__;
  assign new_new_n42034__ = ys__n2652 & ys__n17837;
  assign new_new_n42035__ = ys__n39167 & new_new_n41982__;
  assign new_new_n42036__ = ~new_new_n42034__ & ~new_new_n42035__;
  assign new_new_n42037__ = ~new_new_n42033__ & new_new_n42036__;
  assign new_new_n42038__ = ~new_new_n42032__ & new_new_n42037__;
  assign new_new_n42039__ = new_new_n12219__ & ~new_new_n42038__;
  assign new_new_n42040__ = ~new_new_n24767__ & new_new_n41515__;
  assign new_new_n42041__ = ~new_new_n24759__ & ~new_new_n41515__;
  assign new_new_n42042__ = ~new_new_n42040__ & ~new_new_n42041__;
  assign new_new_n42043__ = ~new_new_n12216__ & ~new_new_n42042__;
  assign new_new_n42044__ = new_new_n12216__ & ~new_new_n24767__;
  assign new_new_n42045__ = ~new_new_n42043__ & ~new_new_n42044__;
  assign new_new_n42046__ = new_new_n12218__ & ~new_new_n42045__;
  assign new_new_n42047__ = ~new_new_n42039__ & ~new_new_n42046__;
  assign ys__n31230 = ys__n888 & ~new_new_n42047__;
  assign new_new_n42049__ = ys__n562 & ys__n47034;
  assign new_new_n42050__ = new_new_n42004__ & new_new_n42027__;
  assign new_new_n42051__ = new_new_n42005__ & new_new_n42050__;
  assign new_new_n42052__ = new_new_n41960__ & new_new_n42051__;
  assign new_new_n42053__ = new_new_n41870__ & new_new_n42052__;
  assign new_new_n42054__ = ~new_new_n42049__ & new_new_n42053__;
  assign new_new_n42055__ = new_new_n42049__ & ~new_new_n42053__;
  assign new_new_n42056__ = ~new_new_n42054__ & ~new_new_n42055__;
  assign new_new_n42057__ = new_new_n41507__ & ~new_new_n42056__;
  assign new_new_n42058__ = new_new_n41504__ & new_new_n42049__;
  assign new_new_n42059__ = ys__n2652 & ys__n17839;
  assign new_new_n42060__ = ys__n39167 & new_new_n42004__;
  assign new_new_n42061__ = ~new_new_n42059__ & ~new_new_n42060__;
  assign new_new_n42062__ = ~new_new_n42058__ & new_new_n42061__;
  assign new_new_n42063__ = ~new_new_n42057__ & new_new_n42062__;
  assign new_new_n42064__ = new_new_n12219__ & ~new_new_n42063__;
  assign new_new_n42065__ = ~new_new_n24849__ & new_new_n41515__;
  assign new_new_n42066__ = ~new_new_n24843__ & ~new_new_n41515__;
  assign new_new_n42067__ = ~new_new_n42065__ & ~new_new_n42066__;
  assign new_new_n42068__ = ~new_new_n12216__ & ~new_new_n42067__;
  assign new_new_n42069__ = new_new_n12216__ & ~new_new_n24849__;
  assign new_new_n42070__ = ~new_new_n42068__ & ~new_new_n42069__;
  assign new_new_n42071__ = new_new_n12218__ & ~new_new_n42070__;
  assign new_new_n42072__ = ~new_new_n42064__ & ~new_new_n42071__;
  assign ys__n31231 = ys__n888 & ~new_new_n42072__;
  assign new_new_n42074__ = ys__n562 & ys__n47035;
  assign new_new_n42075__ = new_new_n42049__ & new_new_n42053__;
  assign new_new_n42076__ = ~new_new_n42074__ & new_new_n42075__;
  assign new_new_n42077__ = new_new_n42074__ & ~new_new_n42075__;
  assign new_new_n42078__ = ~new_new_n42076__ & ~new_new_n42077__;
  assign new_new_n42079__ = new_new_n41507__ & ~new_new_n42078__;
  assign new_new_n42080__ = new_new_n41504__ & new_new_n42074__;
  assign new_new_n42081__ = ys__n2652 & ys__n17840;
  assign new_new_n42082__ = ys__n39167 & new_new_n42027__;
  assign new_new_n42083__ = ~new_new_n42081__ & ~new_new_n42082__;
  assign new_new_n42084__ = ~new_new_n42080__ & new_new_n42083__;
  assign new_new_n42085__ = ~new_new_n42079__ & new_new_n42084__;
  assign new_new_n42086__ = new_new_n12219__ & ~new_new_n42085__;
  assign new_new_n42087__ = ~new_new_n24924__ & new_new_n41515__;
  assign new_new_n42088__ = ~new_new_n24916__ & ~new_new_n41515__;
  assign new_new_n42089__ = ~new_new_n42087__ & ~new_new_n42088__;
  assign new_new_n42090__ = ~new_new_n12216__ & ~new_new_n42089__;
  assign new_new_n42091__ = new_new_n12216__ & ~new_new_n24924__;
  assign new_new_n42092__ = ~new_new_n42090__ & ~new_new_n42091__;
  assign new_new_n42093__ = new_new_n12218__ & ~new_new_n42092__;
  assign new_new_n42094__ = ~new_new_n42086__ & ~new_new_n42093__;
  assign ys__n31232 = ys__n888 & ~new_new_n42094__;
  assign new_new_n42096__ = ys__n562 & ys__n47036;
  assign new_new_n42097__ = new_new_n42049__ & new_new_n42074__;
  assign new_new_n42098__ = new_new_n42053__ & new_new_n42097__;
  assign new_new_n42099__ = ~new_new_n42096__ & new_new_n42098__;
  assign new_new_n42100__ = new_new_n42096__ & ~new_new_n42098__;
  assign new_new_n42101__ = ~new_new_n42099__ & ~new_new_n42100__;
  assign new_new_n42102__ = new_new_n41507__ & ~new_new_n42101__;
  assign new_new_n42103__ = new_new_n41504__ & new_new_n42096__;
  assign new_new_n42104__ = ys__n2652 & ys__n17842;
  assign new_new_n42105__ = ys__n39167 & new_new_n42049__;
  assign new_new_n42106__ = ~new_new_n42104__ & ~new_new_n42105__;
  assign new_new_n42107__ = ~new_new_n42103__ & new_new_n42106__;
  assign new_new_n42108__ = ~new_new_n42102__ & new_new_n42107__;
  assign new_new_n42109__ = new_new_n12219__ & ~new_new_n42108__;
  assign new_new_n42110__ = ~new_new_n25004__ & new_new_n41515__;
  assign new_new_n42111__ = ~new_new_n24996__ & ~new_new_n41515__;
  assign new_new_n42112__ = ~new_new_n42110__ & ~new_new_n42111__;
  assign new_new_n42113__ = ~new_new_n12216__ & ~new_new_n42112__;
  assign new_new_n42114__ = new_new_n12216__ & ~new_new_n25004__;
  assign new_new_n42115__ = ~new_new_n42113__ & ~new_new_n42114__;
  assign new_new_n42116__ = new_new_n12218__ & ~new_new_n42115__;
  assign new_new_n42117__ = ~new_new_n42109__ & ~new_new_n42116__;
  assign ys__n31233 = ys__n888 & ~new_new_n42117__;
  assign new_new_n42119__ = ys__n562 & ys__n47037;
  assign new_new_n42120__ = new_new_n42096__ & new_new_n42098__;
  assign new_new_n42121__ = ~new_new_n42119__ & new_new_n42120__;
  assign new_new_n42122__ = new_new_n42119__ & ~new_new_n42120__;
  assign new_new_n42123__ = ~new_new_n42121__ & ~new_new_n42122__;
  assign new_new_n42124__ = new_new_n41507__ & ~new_new_n42123__;
  assign new_new_n42125__ = new_new_n41504__ & new_new_n42119__;
  assign new_new_n42126__ = ys__n2652 & ys__n17843;
  assign new_new_n42127__ = ys__n39167 & new_new_n42074__;
  assign new_new_n42128__ = ~new_new_n42126__ & ~new_new_n42127__;
  assign new_new_n42129__ = ~new_new_n42125__ & new_new_n42128__;
  assign new_new_n42130__ = ~new_new_n42124__ & new_new_n42129__;
  assign new_new_n42131__ = new_new_n12219__ & ~new_new_n42130__;
  assign new_new_n42132__ = ~new_new_n25080__ & new_new_n41515__;
  assign new_new_n42133__ = ~new_new_n25072__ & ~new_new_n41515__;
  assign new_new_n42134__ = ~new_new_n42132__ & ~new_new_n42133__;
  assign new_new_n42135__ = ~new_new_n12216__ & ~new_new_n42134__;
  assign new_new_n42136__ = new_new_n12216__ & ~new_new_n25080__;
  assign new_new_n42137__ = ~new_new_n42135__ & ~new_new_n42136__;
  assign new_new_n42138__ = new_new_n12218__ & ~new_new_n42137__;
  assign new_new_n42139__ = ~new_new_n42131__ & ~new_new_n42138__;
  assign ys__n31234 = ys__n888 & ~new_new_n42139__;
  assign new_new_n42141__ = ys__n562 & ys__n47038;
  assign new_new_n42142__ = new_new_n42096__ & new_new_n42119__;
  assign new_new_n42143__ = new_new_n42097__ & new_new_n42142__;
  assign new_new_n42144__ = new_new_n42053__ & new_new_n42143__;
  assign new_new_n42145__ = ~new_new_n42141__ & new_new_n42144__;
  assign new_new_n42146__ = new_new_n42141__ & ~new_new_n42144__;
  assign new_new_n42147__ = ~new_new_n42145__ & ~new_new_n42146__;
  assign new_new_n42148__ = new_new_n41507__ & ~new_new_n42147__;
  assign new_new_n42149__ = new_new_n41504__ & new_new_n42141__;
  assign new_new_n42150__ = ys__n2652 & ys__n17845;
  assign new_new_n42151__ = ys__n39167 & new_new_n42096__;
  assign new_new_n42152__ = ~new_new_n42150__ & ~new_new_n42151__;
  assign new_new_n42153__ = ~new_new_n42149__ & new_new_n42152__;
  assign new_new_n42154__ = ~new_new_n42148__ & new_new_n42153__;
  assign new_new_n42155__ = new_new_n12219__ & ~new_new_n42154__;
  assign new_new_n42156__ = ~new_new_n25164__ & new_new_n41515__;
  assign new_new_n42157__ = ~new_new_n25156__ & ~new_new_n41515__;
  assign new_new_n42158__ = ~new_new_n42156__ & ~new_new_n42157__;
  assign new_new_n42159__ = ~new_new_n12216__ & ~new_new_n42158__;
  assign new_new_n42160__ = new_new_n12216__ & ~new_new_n25164__;
  assign new_new_n42161__ = ~new_new_n42159__ & ~new_new_n42160__;
  assign new_new_n42162__ = new_new_n12218__ & ~new_new_n42161__;
  assign new_new_n42163__ = ~new_new_n42155__ & ~new_new_n42162__;
  assign ys__n31235 = ys__n888 & ~new_new_n42163__;
  assign new_new_n42165__ = ys__n562 & ys__n47039;
  assign new_new_n42166__ = new_new_n42141__ & new_new_n42144__;
  assign new_new_n42167__ = ~new_new_n42165__ & new_new_n42166__;
  assign new_new_n42168__ = new_new_n42165__ & ~new_new_n42166__;
  assign new_new_n42169__ = ~new_new_n42167__ & ~new_new_n42168__;
  assign new_new_n42170__ = new_new_n41507__ & ~new_new_n42169__;
  assign new_new_n42171__ = new_new_n41504__ & new_new_n42165__;
  assign new_new_n42172__ = ys__n2652 & ys__n17846;
  assign new_new_n42173__ = ys__n39167 & new_new_n42119__;
  assign new_new_n42174__ = ~new_new_n42172__ & ~new_new_n42173__;
  assign new_new_n42175__ = ~new_new_n42171__ & new_new_n42174__;
  assign new_new_n42176__ = ~new_new_n42170__ & new_new_n42175__;
  assign new_new_n42177__ = new_new_n12219__ & ~new_new_n42176__;
  assign new_new_n42178__ = ~new_new_n25240__ & new_new_n41515__;
  assign new_new_n42179__ = ~new_new_n25232__ & ~new_new_n41515__;
  assign new_new_n42180__ = ~new_new_n42178__ & ~new_new_n42179__;
  assign new_new_n42181__ = ~new_new_n12216__ & ~new_new_n42180__;
  assign new_new_n42182__ = new_new_n12216__ & ~new_new_n25240__;
  assign new_new_n42183__ = ~new_new_n42181__ & ~new_new_n42182__;
  assign new_new_n42184__ = new_new_n12218__ & ~new_new_n42183__;
  assign new_new_n42185__ = ~new_new_n42177__ & ~new_new_n42184__;
  assign ys__n31236 = ys__n888 & ~new_new_n42185__;
  assign new_new_n42187__ = ys__n562 & ys__n47040;
  assign new_new_n42188__ = new_new_n42141__ & new_new_n42165__;
  assign new_new_n42189__ = new_new_n42144__ & new_new_n42188__;
  assign new_new_n42190__ = ~new_new_n42187__ & new_new_n42189__;
  assign new_new_n42191__ = new_new_n42187__ & ~new_new_n42189__;
  assign new_new_n42192__ = ~new_new_n42190__ & ~new_new_n42191__;
  assign new_new_n42193__ = new_new_n41507__ & ~new_new_n42192__;
  assign new_new_n42194__ = new_new_n41504__ & new_new_n42187__;
  assign new_new_n42195__ = ys__n2652 & ys__n17848;
  assign new_new_n42196__ = ys__n39167 & new_new_n42141__;
  assign new_new_n42197__ = ~new_new_n42195__ & ~new_new_n42196__;
  assign new_new_n42198__ = ~new_new_n42194__ & new_new_n42197__;
  assign ys__n39392 = new_new_n42193__ | ~new_new_n42198__;
  assign new_new_n42200__ = new_new_n12219__ & ys__n39392;
  assign new_new_n42201__ = ~new_new_n25320__ & new_new_n41515__;
  assign new_new_n42202__ = ~new_new_n25312__ & ~new_new_n41515__;
  assign new_new_n42203__ = ~new_new_n42201__ & ~new_new_n42202__;
  assign new_new_n42204__ = ~new_new_n12216__ & ~new_new_n42203__;
  assign new_new_n42205__ = new_new_n12216__ & ~new_new_n25320__;
  assign new_new_n42206__ = ~new_new_n42204__ & ~new_new_n42205__;
  assign new_new_n42207__ = new_new_n12218__ & ~new_new_n42206__;
  assign new_new_n42208__ = ~new_new_n42200__ & ~new_new_n42207__;
  assign ys__n31237 = ys__n888 & ~new_new_n42208__;
  assign new_new_n42210__ = ys__n562 & ys__n47041;
  assign new_new_n42211__ = new_new_n42187__ & new_new_n42189__;
  assign new_new_n42212__ = ~new_new_n42210__ & new_new_n42211__;
  assign new_new_n42213__ = new_new_n42210__ & ~new_new_n42211__;
  assign new_new_n42214__ = ~new_new_n42212__ & ~new_new_n42213__;
  assign new_new_n42215__ = new_new_n41507__ & ~new_new_n42214__;
  assign new_new_n42216__ = new_new_n41504__ & new_new_n42210__;
  assign new_new_n42217__ = ys__n2652 & ys__n17849;
  assign new_new_n42218__ = ys__n39167 & new_new_n42165__;
  assign new_new_n42219__ = ~new_new_n42217__ & ~new_new_n42218__;
  assign new_new_n42220__ = ~new_new_n42216__ & new_new_n42219__;
  assign ys__n39393 = new_new_n42215__ | ~new_new_n42220__;
  assign new_new_n42222__ = new_new_n12219__ & ys__n39393;
  assign new_new_n42223__ = ~new_new_n25394__ & new_new_n41515__;
  assign new_new_n42224__ = ~new_new_n25386__ & ~new_new_n41515__;
  assign new_new_n42225__ = ~new_new_n42223__ & ~new_new_n42224__;
  assign new_new_n42226__ = ~new_new_n12216__ & ~new_new_n42225__;
  assign new_new_n42227__ = new_new_n12216__ & ~new_new_n25394__;
  assign new_new_n42228__ = ~new_new_n42226__ & ~new_new_n42227__;
  assign new_new_n42229__ = new_new_n12218__ & ~new_new_n42228__;
  assign new_new_n42230__ = ~new_new_n42222__ & ~new_new_n42229__;
  assign ys__n31238 = ys__n888 & ~new_new_n42230__;
  assign new_new_n42232__ = ys__n842 & new_new_n12106__;
  assign new_new_n42233__ = ys__n47234 & new_new_n42232__;
  assign new_new_n42234__ = ~ys__n844 & ~new_new_n12106__;
  assign new_new_n42235__ = ~ys__n842 & new_new_n12106__;
  assign new_new_n42236__ = ~new_new_n42234__ & ~new_new_n42235__;
  assign new_new_n42237__ = ys__n47202 & ~new_new_n42236__;
  assign new_new_n42238__ = ~new_new_n42233__ & ~new_new_n42237__;
  assign new_new_n42239__ = ~new_new_n42232__ & new_new_n42236__;
  assign ys__n31326 = ~new_new_n42238__ & ~new_new_n42239__;
  assign new_new_n42241__ = ys__n47235 & new_new_n42232__;
  assign new_new_n42242__ = ys__n47203 & ~new_new_n42236__;
  assign new_new_n42243__ = ~new_new_n42241__ & ~new_new_n42242__;
  assign ys__n31327 = ~new_new_n42239__ & ~new_new_n42243__;
  assign new_new_n42245__ = ys__n47236 & new_new_n42232__;
  assign new_new_n42246__ = ys__n47204 & ~new_new_n42236__;
  assign new_new_n42247__ = ~new_new_n42245__ & ~new_new_n42246__;
  assign ys__n31328 = ~new_new_n42239__ & ~new_new_n42247__;
  assign new_new_n42249__ = ys__n47237 & new_new_n42232__;
  assign new_new_n42250__ = ys__n47205 & ~new_new_n42236__;
  assign new_new_n42251__ = ~new_new_n42249__ & ~new_new_n42250__;
  assign ys__n31329 = ~new_new_n42239__ & ~new_new_n42251__;
  assign new_new_n42253__ = ys__n47238 & new_new_n42232__;
  assign new_new_n42254__ = ys__n47206 & ~new_new_n42236__;
  assign new_new_n42255__ = ~new_new_n42253__ & ~new_new_n42254__;
  assign ys__n31330 = ~new_new_n42239__ & ~new_new_n42255__;
  assign new_new_n42257__ = ys__n47239 & new_new_n42232__;
  assign new_new_n42258__ = ys__n47207 & ~new_new_n42236__;
  assign new_new_n42259__ = ~new_new_n42257__ & ~new_new_n42258__;
  assign ys__n31331 = ~new_new_n42239__ & ~new_new_n42259__;
  assign new_new_n42261__ = ys__n47240 & new_new_n42232__;
  assign new_new_n42262__ = ys__n47208 & ~new_new_n42236__;
  assign new_new_n42263__ = ~new_new_n42261__ & ~new_new_n42262__;
  assign ys__n31332 = ~new_new_n42239__ & ~new_new_n42263__;
  assign new_new_n42265__ = ys__n47241 & new_new_n42232__;
  assign new_new_n42266__ = ys__n47209 & ~new_new_n42236__;
  assign new_new_n42267__ = ~new_new_n42265__ & ~new_new_n42266__;
  assign ys__n31333 = ~new_new_n42239__ & ~new_new_n42267__;
  assign new_new_n42269__ = ys__n47242 & new_new_n42232__;
  assign new_new_n42270__ = ys__n47210 & ~new_new_n42236__;
  assign new_new_n42271__ = ~new_new_n42269__ & ~new_new_n42270__;
  assign ys__n31334 = ~new_new_n42239__ & ~new_new_n42271__;
  assign new_new_n42273__ = ys__n47243 & new_new_n42232__;
  assign new_new_n42274__ = ys__n47211 & ~new_new_n42236__;
  assign new_new_n42275__ = ~new_new_n42273__ & ~new_new_n42274__;
  assign ys__n31335 = ~new_new_n42239__ & ~new_new_n42275__;
  assign new_new_n42277__ = ys__n47244 & new_new_n42232__;
  assign new_new_n42278__ = ys__n47212 & ~new_new_n42236__;
  assign new_new_n42279__ = ~new_new_n42277__ & ~new_new_n42278__;
  assign ys__n31336 = ~new_new_n42239__ & ~new_new_n42279__;
  assign new_new_n42281__ = ys__n47245 & new_new_n42232__;
  assign new_new_n42282__ = ys__n47213 & ~new_new_n42236__;
  assign new_new_n42283__ = ~new_new_n42281__ & ~new_new_n42282__;
  assign ys__n31337 = ~new_new_n42239__ & ~new_new_n42283__;
  assign new_new_n42285__ = ys__n47246 & new_new_n42232__;
  assign new_new_n42286__ = ys__n47214 & ~new_new_n42236__;
  assign new_new_n42287__ = ~new_new_n42285__ & ~new_new_n42286__;
  assign ys__n31338 = ~new_new_n42239__ & ~new_new_n42287__;
  assign new_new_n42289__ = ys__n47247 & new_new_n42232__;
  assign new_new_n42290__ = ys__n47215 & ~new_new_n42236__;
  assign new_new_n42291__ = ~new_new_n42289__ & ~new_new_n42290__;
  assign ys__n31339 = ~new_new_n42239__ & ~new_new_n42291__;
  assign new_new_n42293__ = ys__n47248 & new_new_n42232__;
  assign new_new_n42294__ = ys__n47216 & ~new_new_n42236__;
  assign new_new_n42295__ = ~new_new_n42293__ & ~new_new_n42294__;
  assign ys__n31340 = ~new_new_n42239__ & ~new_new_n42295__;
  assign new_new_n42297__ = ys__n47249 & new_new_n42232__;
  assign new_new_n42298__ = ys__n47217 & ~new_new_n42236__;
  assign new_new_n42299__ = ~new_new_n42297__ & ~new_new_n42298__;
  assign ys__n31341 = ~new_new_n42239__ & ~new_new_n42299__;
  assign new_new_n42301__ = ys__n47250 & new_new_n42232__;
  assign new_new_n42302__ = ys__n47218 & ~new_new_n42236__;
  assign new_new_n42303__ = ~new_new_n42301__ & ~new_new_n42302__;
  assign ys__n31342 = ~new_new_n42239__ & ~new_new_n42303__;
  assign new_new_n42305__ = ys__n47251 & new_new_n42232__;
  assign new_new_n42306__ = ys__n47219 & ~new_new_n42236__;
  assign new_new_n42307__ = ~new_new_n42305__ & ~new_new_n42306__;
  assign ys__n31343 = ~new_new_n42239__ & ~new_new_n42307__;
  assign new_new_n42309__ = ys__n47252 & new_new_n42232__;
  assign new_new_n42310__ = ys__n47220 & ~new_new_n42236__;
  assign new_new_n42311__ = ~new_new_n42309__ & ~new_new_n42310__;
  assign ys__n31344 = ~new_new_n42239__ & ~new_new_n42311__;
  assign new_new_n42313__ = ys__n47253 & new_new_n42232__;
  assign new_new_n42314__ = ys__n47221 & ~new_new_n42236__;
  assign new_new_n42315__ = ~new_new_n42313__ & ~new_new_n42314__;
  assign ys__n31345 = ~new_new_n42239__ & ~new_new_n42315__;
  assign new_new_n42317__ = ys__n47254 & new_new_n42232__;
  assign new_new_n42318__ = ys__n47222 & ~new_new_n42236__;
  assign new_new_n42319__ = ~new_new_n42317__ & ~new_new_n42318__;
  assign ys__n31346 = ~new_new_n42239__ & ~new_new_n42319__;
  assign new_new_n42321__ = ys__n47255 & new_new_n42232__;
  assign new_new_n42322__ = ys__n47223 & ~new_new_n42236__;
  assign new_new_n42323__ = ~new_new_n42321__ & ~new_new_n42322__;
  assign ys__n31347 = ~new_new_n42239__ & ~new_new_n42323__;
  assign new_new_n42325__ = ys__n47256 & new_new_n42232__;
  assign new_new_n42326__ = ys__n47224 & ~new_new_n42236__;
  assign new_new_n42327__ = ~new_new_n42325__ & ~new_new_n42326__;
  assign ys__n31348 = ~new_new_n42239__ & ~new_new_n42327__;
  assign new_new_n42329__ = ys__n47257 & new_new_n42232__;
  assign new_new_n42330__ = ys__n47225 & ~new_new_n42236__;
  assign new_new_n42331__ = ~new_new_n42329__ & ~new_new_n42330__;
  assign ys__n31349 = ~new_new_n42239__ & ~new_new_n42331__;
  assign new_new_n42333__ = ys__n47258 & new_new_n42232__;
  assign new_new_n42334__ = ys__n47226 & ~new_new_n42236__;
  assign new_new_n42335__ = ~new_new_n42333__ & ~new_new_n42334__;
  assign ys__n31350 = ~new_new_n42239__ & ~new_new_n42335__;
  assign new_new_n42337__ = ys__n47259 & new_new_n42232__;
  assign new_new_n42338__ = ys__n47227 & ~new_new_n42236__;
  assign new_new_n42339__ = ~new_new_n42337__ & ~new_new_n42338__;
  assign ys__n31351 = ~new_new_n42239__ & ~new_new_n42339__;
  assign new_new_n42341__ = ys__n47260 & new_new_n42232__;
  assign new_new_n42342__ = ys__n47228 & ~new_new_n42236__;
  assign new_new_n42343__ = ~new_new_n42341__ & ~new_new_n42342__;
  assign ys__n31352 = ~new_new_n42239__ & ~new_new_n42343__;
  assign new_new_n42345__ = ys__n47261 & new_new_n42232__;
  assign new_new_n42346__ = ys__n47229 & ~new_new_n42236__;
  assign new_new_n42347__ = ~new_new_n42345__ & ~new_new_n42346__;
  assign ys__n31353 = ~new_new_n42239__ & ~new_new_n42347__;
  assign new_new_n42349__ = ys__n47262 & new_new_n42232__;
  assign new_new_n42350__ = ys__n47230 & ~new_new_n42236__;
  assign new_new_n42351__ = ~new_new_n42349__ & ~new_new_n42350__;
  assign ys__n31354 = ~new_new_n42239__ & ~new_new_n42351__;
  assign new_new_n42353__ = ys__n47263 & new_new_n42232__;
  assign new_new_n42354__ = ys__n47231 & ~new_new_n42236__;
  assign new_new_n42355__ = ~new_new_n42353__ & ~new_new_n42354__;
  assign ys__n31355 = ~new_new_n42239__ & ~new_new_n42355__;
  assign new_new_n42357__ = ys__n47264 & new_new_n42232__;
  assign new_new_n42358__ = ys__n47232 & ~new_new_n42236__;
  assign new_new_n42359__ = ~new_new_n42357__ & ~new_new_n42358__;
  assign ys__n31356 = ~new_new_n42239__ & ~new_new_n42359__;
  assign new_new_n42361__ = ys__n47265 & new_new_n42232__;
  assign new_new_n42362__ = ys__n47233 & ~new_new_n42236__;
  assign new_new_n42363__ = ~new_new_n42361__ & ~new_new_n42362__;
  assign ys__n31357 = ~new_new_n42239__ & ~new_new_n42363__;
  assign new_new_n42365__ = ys__n47266 & new_new_n42232__;
  assign new_new_n42366__ = ys__n18762 & ~new_new_n42236__;
  assign new_new_n42367__ = ~new_new_n42365__ & ~new_new_n42366__;
  assign ys__n31358 = ~new_new_n42239__ & ~new_new_n42367__;
  assign new_new_n42369__ = ys__n47267 & new_new_n42232__;
  assign new_new_n42370__ = ys__n18750 & ~new_new_n42236__;
  assign new_new_n42371__ = ~new_new_n42369__ & ~new_new_n42370__;
  assign ys__n31359 = ~new_new_n42239__ & ~new_new_n42371__;
  assign new_new_n42373__ = ys__n47268 & new_new_n42232__;
  assign new_new_n42374__ = ys__n18753 & ~new_new_n42236__;
  assign new_new_n42375__ = ~new_new_n42373__ & ~new_new_n42374__;
  assign ys__n31360 = ~new_new_n42239__ & ~new_new_n42375__;
  assign new_new_n42377__ = ys__n840 & new_new_n12106__;
  assign new_new_n42378__ = ys__n47269 & new_new_n42377__;
  assign new_new_n42379__ = ~ys__n842 & ~new_new_n12106__;
  assign new_new_n42380__ = ~ys__n840 & new_new_n12106__;
  assign new_new_n42381__ = ~new_new_n42379__ & ~new_new_n42380__;
  assign new_new_n42382__ = ys__n47202 & ~new_new_n42381__;
  assign new_new_n42383__ = ~new_new_n42378__ & ~new_new_n42382__;
  assign new_new_n42384__ = ~new_new_n42377__ & new_new_n42381__;
  assign ys__n31361 = ~new_new_n42383__ & ~new_new_n42384__;
  assign new_new_n42386__ = ys__n47270 & new_new_n42377__;
  assign new_new_n42387__ = ys__n47203 & ~new_new_n42381__;
  assign new_new_n42388__ = ~new_new_n42386__ & ~new_new_n42387__;
  assign ys__n31362 = ~new_new_n42384__ & ~new_new_n42388__;
  assign new_new_n42390__ = ys__n47271 & new_new_n42377__;
  assign new_new_n42391__ = ys__n47204 & ~new_new_n42381__;
  assign new_new_n42392__ = ~new_new_n42390__ & ~new_new_n42391__;
  assign ys__n31363 = ~new_new_n42384__ & ~new_new_n42392__;
  assign new_new_n42394__ = ys__n47272 & new_new_n42377__;
  assign new_new_n42395__ = ys__n47205 & ~new_new_n42381__;
  assign new_new_n42396__ = ~new_new_n42394__ & ~new_new_n42395__;
  assign ys__n31364 = ~new_new_n42384__ & ~new_new_n42396__;
  assign new_new_n42398__ = ys__n47273 & new_new_n42377__;
  assign new_new_n42399__ = ys__n47206 & ~new_new_n42381__;
  assign new_new_n42400__ = ~new_new_n42398__ & ~new_new_n42399__;
  assign ys__n31365 = ~new_new_n42384__ & ~new_new_n42400__;
  assign new_new_n42402__ = ys__n47274 & new_new_n42377__;
  assign new_new_n42403__ = ys__n47207 & ~new_new_n42381__;
  assign new_new_n42404__ = ~new_new_n42402__ & ~new_new_n42403__;
  assign ys__n31366 = ~new_new_n42384__ & ~new_new_n42404__;
  assign new_new_n42406__ = ys__n47275 & new_new_n42377__;
  assign new_new_n42407__ = ys__n47208 & ~new_new_n42381__;
  assign new_new_n42408__ = ~new_new_n42406__ & ~new_new_n42407__;
  assign ys__n31367 = ~new_new_n42384__ & ~new_new_n42408__;
  assign new_new_n42410__ = ys__n47276 & new_new_n42377__;
  assign new_new_n42411__ = ys__n47209 & ~new_new_n42381__;
  assign new_new_n42412__ = ~new_new_n42410__ & ~new_new_n42411__;
  assign ys__n31368 = ~new_new_n42384__ & ~new_new_n42412__;
  assign new_new_n42414__ = ys__n47277 & new_new_n42377__;
  assign new_new_n42415__ = ys__n47210 & ~new_new_n42381__;
  assign new_new_n42416__ = ~new_new_n42414__ & ~new_new_n42415__;
  assign ys__n31369 = ~new_new_n42384__ & ~new_new_n42416__;
  assign new_new_n42418__ = ys__n47278 & new_new_n42377__;
  assign new_new_n42419__ = ys__n47211 & ~new_new_n42381__;
  assign new_new_n42420__ = ~new_new_n42418__ & ~new_new_n42419__;
  assign ys__n31370 = ~new_new_n42384__ & ~new_new_n42420__;
  assign new_new_n42422__ = ys__n47279 & new_new_n42377__;
  assign new_new_n42423__ = ys__n47212 & ~new_new_n42381__;
  assign new_new_n42424__ = ~new_new_n42422__ & ~new_new_n42423__;
  assign ys__n31371 = ~new_new_n42384__ & ~new_new_n42424__;
  assign new_new_n42426__ = ys__n47280 & new_new_n42377__;
  assign new_new_n42427__ = ys__n47213 & ~new_new_n42381__;
  assign new_new_n42428__ = ~new_new_n42426__ & ~new_new_n42427__;
  assign ys__n31372 = ~new_new_n42384__ & ~new_new_n42428__;
  assign new_new_n42430__ = ys__n47281 & new_new_n42377__;
  assign new_new_n42431__ = ys__n47214 & ~new_new_n42381__;
  assign new_new_n42432__ = ~new_new_n42430__ & ~new_new_n42431__;
  assign ys__n31373 = ~new_new_n42384__ & ~new_new_n42432__;
  assign new_new_n42434__ = ys__n47282 & new_new_n42377__;
  assign new_new_n42435__ = ys__n47215 & ~new_new_n42381__;
  assign new_new_n42436__ = ~new_new_n42434__ & ~new_new_n42435__;
  assign ys__n31374 = ~new_new_n42384__ & ~new_new_n42436__;
  assign new_new_n42438__ = ys__n47283 & new_new_n42377__;
  assign new_new_n42439__ = ys__n47216 & ~new_new_n42381__;
  assign new_new_n42440__ = ~new_new_n42438__ & ~new_new_n42439__;
  assign ys__n31375 = ~new_new_n42384__ & ~new_new_n42440__;
  assign new_new_n42442__ = ys__n47284 & new_new_n42377__;
  assign new_new_n42443__ = ys__n47217 & ~new_new_n42381__;
  assign new_new_n42444__ = ~new_new_n42442__ & ~new_new_n42443__;
  assign ys__n31376 = ~new_new_n42384__ & ~new_new_n42444__;
  assign new_new_n42446__ = ys__n47285 & new_new_n42377__;
  assign new_new_n42447__ = ys__n47218 & ~new_new_n42381__;
  assign new_new_n42448__ = ~new_new_n42446__ & ~new_new_n42447__;
  assign ys__n31377 = ~new_new_n42384__ & ~new_new_n42448__;
  assign new_new_n42450__ = ys__n47286 & new_new_n42377__;
  assign new_new_n42451__ = ys__n47219 & ~new_new_n42381__;
  assign new_new_n42452__ = ~new_new_n42450__ & ~new_new_n42451__;
  assign ys__n31378 = ~new_new_n42384__ & ~new_new_n42452__;
  assign new_new_n42454__ = ys__n47287 & new_new_n42377__;
  assign new_new_n42455__ = ys__n47220 & ~new_new_n42381__;
  assign new_new_n42456__ = ~new_new_n42454__ & ~new_new_n42455__;
  assign ys__n31379 = ~new_new_n42384__ & ~new_new_n42456__;
  assign new_new_n42458__ = ys__n47288 & new_new_n42377__;
  assign new_new_n42459__ = ys__n47221 & ~new_new_n42381__;
  assign new_new_n42460__ = ~new_new_n42458__ & ~new_new_n42459__;
  assign ys__n31380 = ~new_new_n42384__ & ~new_new_n42460__;
  assign new_new_n42462__ = ys__n47289 & new_new_n42377__;
  assign new_new_n42463__ = ys__n47222 & ~new_new_n42381__;
  assign new_new_n42464__ = ~new_new_n42462__ & ~new_new_n42463__;
  assign ys__n31381 = ~new_new_n42384__ & ~new_new_n42464__;
  assign new_new_n42466__ = ys__n47290 & new_new_n42377__;
  assign new_new_n42467__ = ys__n47223 & ~new_new_n42381__;
  assign new_new_n42468__ = ~new_new_n42466__ & ~new_new_n42467__;
  assign ys__n31382 = ~new_new_n42384__ & ~new_new_n42468__;
  assign new_new_n42470__ = ys__n47291 & new_new_n42377__;
  assign new_new_n42471__ = ys__n47224 & ~new_new_n42381__;
  assign new_new_n42472__ = ~new_new_n42470__ & ~new_new_n42471__;
  assign ys__n31383 = ~new_new_n42384__ & ~new_new_n42472__;
  assign new_new_n42474__ = ys__n47292 & new_new_n42377__;
  assign new_new_n42475__ = ys__n47225 & ~new_new_n42381__;
  assign new_new_n42476__ = ~new_new_n42474__ & ~new_new_n42475__;
  assign ys__n31384 = ~new_new_n42384__ & ~new_new_n42476__;
  assign new_new_n42478__ = ys__n47293 & new_new_n42377__;
  assign new_new_n42479__ = ys__n47226 & ~new_new_n42381__;
  assign new_new_n42480__ = ~new_new_n42478__ & ~new_new_n42479__;
  assign ys__n31385 = ~new_new_n42384__ & ~new_new_n42480__;
  assign new_new_n42482__ = ys__n47294 & new_new_n42377__;
  assign new_new_n42483__ = ys__n47227 & ~new_new_n42381__;
  assign new_new_n42484__ = ~new_new_n42482__ & ~new_new_n42483__;
  assign ys__n31386 = ~new_new_n42384__ & ~new_new_n42484__;
  assign new_new_n42486__ = ys__n47295 & new_new_n42377__;
  assign new_new_n42487__ = ys__n47228 & ~new_new_n42381__;
  assign new_new_n42488__ = ~new_new_n42486__ & ~new_new_n42487__;
  assign ys__n31387 = ~new_new_n42384__ & ~new_new_n42488__;
  assign new_new_n42490__ = ys__n47296 & new_new_n42377__;
  assign new_new_n42491__ = ys__n47229 & ~new_new_n42381__;
  assign new_new_n42492__ = ~new_new_n42490__ & ~new_new_n42491__;
  assign ys__n31388 = ~new_new_n42384__ & ~new_new_n42492__;
  assign new_new_n42494__ = ys__n47297 & new_new_n42377__;
  assign new_new_n42495__ = ys__n47230 & ~new_new_n42381__;
  assign new_new_n42496__ = ~new_new_n42494__ & ~new_new_n42495__;
  assign ys__n31389 = ~new_new_n42384__ & ~new_new_n42496__;
  assign new_new_n42498__ = ys__n47298 & new_new_n42377__;
  assign new_new_n42499__ = ys__n47231 & ~new_new_n42381__;
  assign new_new_n42500__ = ~new_new_n42498__ & ~new_new_n42499__;
  assign ys__n31390 = ~new_new_n42384__ & ~new_new_n42500__;
  assign new_new_n42502__ = ys__n47299 & new_new_n42377__;
  assign new_new_n42503__ = ys__n47232 & ~new_new_n42381__;
  assign new_new_n42504__ = ~new_new_n42502__ & ~new_new_n42503__;
  assign ys__n31391 = ~new_new_n42384__ & ~new_new_n42504__;
  assign new_new_n42506__ = ys__n47300 & new_new_n42377__;
  assign new_new_n42507__ = ys__n47233 & ~new_new_n42381__;
  assign new_new_n42508__ = ~new_new_n42506__ & ~new_new_n42507__;
  assign ys__n31392 = ~new_new_n42384__ & ~new_new_n42508__;
  assign new_new_n42510__ = ys__n47301 & new_new_n42377__;
  assign new_new_n42511__ = ys__n18762 & ~new_new_n42381__;
  assign new_new_n42512__ = ~new_new_n42510__ & ~new_new_n42511__;
  assign ys__n31393 = ~new_new_n42384__ & ~new_new_n42512__;
  assign new_new_n42514__ = ys__n47302 & new_new_n42377__;
  assign new_new_n42515__ = ys__n18750 & ~new_new_n42381__;
  assign new_new_n42516__ = ~new_new_n42514__ & ~new_new_n42515__;
  assign ys__n31394 = ~new_new_n42384__ & ~new_new_n42516__;
  assign new_new_n42518__ = ys__n47303 & new_new_n42377__;
  assign new_new_n42519__ = ys__n18753 & ~new_new_n42381__;
  assign new_new_n42520__ = ~new_new_n42518__ & ~new_new_n42519__;
  assign ys__n31395 = ~new_new_n42384__ & ~new_new_n42520__;
  assign new_new_n42522__ = ys__n838 & new_new_n12106__;
  assign new_new_n42523__ = ys__n47305 & new_new_n42522__;
  assign new_new_n42524__ = ~ys__n840 & ~new_new_n12106__;
  assign new_new_n42525__ = ~ys__n838 & new_new_n12106__;
  assign new_new_n42526__ = ~new_new_n42524__ & ~new_new_n42525__;
  assign new_new_n42527__ = ys__n47202 & ~new_new_n42526__;
  assign new_new_n42528__ = ~new_new_n42523__ & ~new_new_n42527__;
  assign new_new_n42529__ = ~new_new_n42522__ & new_new_n42526__;
  assign ys__n31397 = ~new_new_n42528__ & ~new_new_n42529__;
  assign new_new_n42531__ = ys__n47306 & new_new_n42522__;
  assign new_new_n42532__ = ys__n47203 & ~new_new_n42526__;
  assign new_new_n42533__ = ~new_new_n42531__ & ~new_new_n42532__;
  assign ys__n31398 = ~new_new_n42529__ & ~new_new_n42533__;
  assign new_new_n42535__ = ys__n47307 & new_new_n42522__;
  assign new_new_n42536__ = ys__n47204 & ~new_new_n42526__;
  assign new_new_n42537__ = ~new_new_n42535__ & ~new_new_n42536__;
  assign ys__n31399 = ~new_new_n42529__ & ~new_new_n42537__;
  assign new_new_n42539__ = ys__n47308 & new_new_n42522__;
  assign new_new_n42540__ = ys__n47205 & ~new_new_n42526__;
  assign new_new_n42541__ = ~new_new_n42539__ & ~new_new_n42540__;
  assign ys__n31400 = ~new_new_n42529__ & ~new_new_n42541__;
  assign new_new_n42543__ = ys__n47309 & new_new_n42522__;
  assign new_new_n42544__ = ys__n47206 & ~new_new_n42526__;
  assign new_new_n42545__ = ~new_new_n42543__ & ~new_new_n42544__;
  assign ys__n31401 = ~new_new_n42529__ & ~new_new_n42545__;
  assign new_new_n42547__ = ys__n47310 & new_new_n42522__;
  assign new_new_n42548__ = ys__n47207 & ~new_new_n42526__;
  assign new_new_n42549__ = ~new_new_n42547__ & ~new_new_n42548__;
  assign ys__n31402 = ~new_new_n42529__ & ~new_new_n42549__;
  assign new_new_n42551__ = ys__n47311 & new_new_n42522__;
  assign new_new_n42552__ = ys__n47208 & ~new_new_n42526__;
  assign new_new_n42553__ = ~new_new_n42551__ & ~new_new_n42552__;
  assign ys__n31403 = ~new_new_n42529__ & ~new_new_n42553__;
  assign new_new_n42555__ = ys__n47312 & new_new_n42522__;
  assign new_new_n42556__ = ys__n47209 & ~new_new_n42526__;
  assign new_new_n42557__ = ~new_new_n42555__ & ~new_new_n42556__;
  assign ys__n31404 = ~new_new_n42529__ & ~new_new_n42557__;
  assign new_new_n42559__ = ys__n47313 & new_new_n42522__;
  assign new_new_n42560__ = ys__n47210 & ~new_new_n42526__;
  assign new_new_n42561__ = ~new_new_n42559__ & ~new_new_n42560__;
  assign ys__n31405 = ~new_new_n42529__ & ~new_new_n42561__;
  assign new_new_n42563__ = ys__n47314 & new_new_n42522__;
  assign new_new_n42564__ = ys__n47211 & ~new_new_n42526__;
  assign new_new_n42565__ = ~new_new_n42563__ & ~new_new_n42564__;
  assign ys__n31406 = ~new_new_n42529__ & ~new_new_n42565__;
  assign new_new_n42567__ = ys__n47315 & new_new_n42522__;
  assign new_new_n42568__ = ys__n47212 & ~new_new_n42526__;
  assign new_new_n42569__ = ~new_new_n42567__ & ~new_new_n42568__;
  assign ys__n31407 = ~new_new_n42529__ & ~new_new_n42569__;
  assign new_new_n42571__ = ys__n47316 & new_new_n42522__;
  assign new_new_n42572__ = ys__n47213 & ~new_new_n42526__;
  assign new_new_n42573__ = ~new_new_n42571__ & ~new_new_n42572__;
  assign ys__n31408 = ~new_new_n42529__ & ~new_new_n42573__;
  assign new_new_n42575__ = ys__n47317 & new_new_n42522__;
  assign new_new_n42576__ = ys__n47214 & ~new_new_n42526__;
  assign new_new_n42577__ = ~new_new_n42575__ & ~new_new_n42576__;
  assign ys__n31409 = ~new_new_n42529__ & ~new_new_n42577__;
  assign new_new_n42579__ = ys__n47318 & new_new_n42522__;
  assign new_new_n42580__ = ys__n47215 & ~new_new_n42526__;
  assign new_new_n42581__ = ~new_new_n42579__ & ~new_new_n42580__;
  assign ys__n31410 = ~new_new_n42529__ & ~new_new_n42581__;
  assign new_new_n42583__ = ys__n47319 & new_new_n42522__;
  assign new_new_n42584__ = ys__n47216 & ~new_new_n42526__;
  assign new_new_n42585__ = ~new_new_n42583__ & ~new_new_n42584__;
  assign ys__n31411 = ~new_new_n42529__ & ~new_new_n42585__;
  assign new_new_n42587__ = ys__n47320 & new_new_n42522__;
  assign new_new_n42588__ = ys__n47217 & ~new_new_n42526__;
  assign new_new_n42589__ = ~new_new_n42587__ & ~new_new_n42588__;
  assign ys__n31412 = ~new_new_n42529__ & ~new_new_n42589__;
  assign new_new_n42591__ = ys__n47321 & new_new_n42522__;
  assign new_new_n42592__ = ys__n47218 & ~new_new_n42526__;
  assign new_new_n42593__ = ~new_new_n42591__ & ~new_new_n42592__;
  assign ys__n31413 = ~new_new_n42529__ & ~new_new_n42593__;
  assign new_new_n42595__ = ys__n47322 & new_new_n42522__;
  assign new_new_n42596__ = ys__n47219 & ~new_new_n42526__;
  assign new_new_n42597__ = ~new_new_n42595__ & ~new_new_n42596__;
  assign ys__n31414 = ~new_new_n42529__ & ~new_new_n42597__;
  assign new_new_n42599__ = ys__n47323 & new_new_n42522__;
  assign new_new_n42600__ = ys__n47220 & ~new_new_n42526__;
  assign new_new_n42601__ = ~new_new_n42599__ & ~new_new_n42600__;
  assign ys__n31415 = ~new_new_n42529__ & ~new_new_n42601__;
  assign new_new_n42603__ = ys__n47324 & new_new_n42522__;
  assign new_new_n42604__ = ys__n47221 & ~new_new_n42526__;
  assign new_new_n42605__ = ~new_new_n42603__ & ~new_new_n42604__;
  assign ys__n31416 = ~new_new_n42529__ & ~new_new_n42605__;
  assign new_new_n42607__ = ys__n47325 & new_new_n42522__;
  assign new_new_n42608__ = ys__n47222 & ~new_new_n42526__;
  assign new_new_n42609__ = ~new_new_n42607__ & ~new_new_n42608__;
  assign ys__n31417 = ~new_new_n42529__ & ~new_new_n42609__;
  assign new_new_n42611__ = ys__n47326 & new_new_n42522__;
  assign new_new_n42612__ = ys__n47223 & ~new_new_n42526__;
  assign new_new_n42613__ = ~new_new_n42611__ & ~new_new_n42612__;
  assign ys__n31418 = ~new_new_n42529__ & ~new_new_n42613__;
  assign new_new_n42615__ = ys__n47327 & new_new_n42522__;
  assign new_new_n42616__ = ys__n47224 & ~new_new_n42526__;
  assign new_new_n42617__ = ~new_new_n42615__ & ~new_new_n42616__;
  assign ys__n31419 = ~new_new_n42529__ & ~new_new_n42617__;
  assign new_new_n42619__ = ys__n47328 & new_new_n42522__;
  assign new_new_n42620__ = ys__n47225 & ~new_new_n42526__;
  assign new_new_n42621__ = ~new_new_n42619__ & ~new_new_n42620__;
  assign ys__n31420 = ~new_new_n42529__ & ~new_new_n42621__;
  assign new_new_n42623__ = ys__n47329 & new_new_n42522__;
  assign new_new_n42624__ = ys__n47226 & ~new_new_n42526__;
  assign new_new_n42625__ = ~new_new_n42623__ & ~new_new_n42624__;
  assign ys__n31421 = ~new_new_n42529__ & ~new_new_n42625__;
  assign new_new_n42627__ = ys__n47330 & new_new_n42522__;
  assign new_new_n42628__ = ys__n47227 & ~new_new_n42526__;
  assign new_new_n42629__ = ~new_new_n42627__ & ~new_new_n42628__;
  assign ys__n31422 = ~new_new_n42529__ & ~new_new_n42629__;
  assign new_new_n42631__ = ys__n47331 & new_new_n42522__;
  assign new_new_n42632__ = ys__n47228 & ~new_new_n42526__;
  assign new_new_n42633__ = ~new_new_n42631__ & ~new_new_n42632__;
  assign ys__n31423 = ~new_new_n42529__ & ~new_new_n42633__;
  assign new_new_n42635__ = ys__n47332 & new_new_n42522__;
  assign new_new_n42636__ = ys__n47229 & ~new_new_n42526__;
  assign new_new_n42637__ = ~new_new_n42635__ & ~new_new_n42636__;
  assign ys__n31424 = ~new_new_n42529__ & ~new_new_n42637__;
  assign new_new_n42639__ = ys__n47333 & new_new_n42522__;
  assign new_new_n42640__ = ys__n47230 & ~new_new_n42526__;
  assign new_new_n42641__ = ~new_new_n42639__ & ~new_new_n42640__;
  assign ys__n31425 = ~new_new_n42529__ & ~new_new_n42641__;
  assign new_new_n42643__ = ys__n47334 & new_new_n42522__;
  assign new_new_n42644__ = ys__n47231 & ~new_new_n42526__;
  assign new_new_n42645__ = ~new_new_n42643__ & ~new_new_n42644__;
  assign ys__n31426 = ~new_new_n42529__ & ~new_new_n42645__;
  assign new_new_n42647__ = ys__n47335 & new_new_n42522__;
  assign new_new_n42648__ = ys__n47232 & ~new_new_n42526__;
  assign new_new_n42649__ = ~new_new_n42647__ & ~new_new_n42648__;
  assign ys__n31427 = ~new_new_n42529__ & ~new_new_n42649__;
  assign new_new_n42651__ = ys__n47336 & new_new_n42522__;
  assign new_new_n42652__ = ys__n47233 & ~new_new_n42526__;
  assign new_new_n42653__ = ~new_new_n42651__ & ~new_new_n42652__;
  assign ys__n31428 = ~new_new_n42529__ & ~new_new_n42653__;
  assign new_new_n42655__ = ys__n47337 & new_new_n42522__;
  assign new_new_n42656__ = ys__n18762 & ~new_new_n42526__;
  assign new_new_n42657__ = ~new_new_n42655__ & ~new_new_n42656__;
  assign ys__n31429 = ~new_new_n42529__ & ~new_new_n42657__;
  assign new_new_n42659__ = ys__n47338 & new_new_n42522__;
  assign new_new_n42660__ = ys__n18750 & ~new_new_n42526__;
  assign new_new_n42661__ = ~new_new_n42659__ & ~new_new_n42660__;
  assign ys__n31430 = ~new_new_n42529__ & ~new_new_n42661__;
  assign new_new_n42663__ = ys__n47339 & new_new_n42522__;
  assign new_new_n42664__ = ys__n18753 & ~new_new_n42526__;
  assign new_new_n42665__ = ~new_new_n42663__ & ~new_new_n42664__;
  assign ys__n31431 = ~new_new_n42529__ & ~new_new_n42665__;
  assign new_new_n42667__ = ys__n1386 & ys__n24188;
  assign new_new_n42668__ = ys__n47340 & ~ys__n2152;
  assign new_new_n42669__ = ys__n47342 & new_new_n35343__;
  assign new_new_n42670__ = ys__n47341 & new_new_n35345__;
  assign new_new_n42671__ = ~new_new_n42669__ & ~new_new_n42670__;
  assign new_new_n42672__ = ~ys__n182 & ~new_new_n35343__;
  assign new_new_n42673__ = ~new_new_n35345__ & new_new_n42672__;
  assign new_new_n42674__ = ~new_new_n42671__ & ~new_new_n42673__;
  assign new_new_n42675__ = new_new_n41469__ & new_new_n42674__;
  assign new_new_n42676__ = ~new_new_n42668__ & ~new_new_n42675__;
  assign new_new_n42677__ = ~new_new_n42667__ & new_new_n42676__;
  assign new_new_n42678__ = ys__n2152 & new_new_n41481__;
  assign ys__n33007 = ~new_new_n42677__ & ~new_new_n42678__;
  assign new_new_n42680__ = ~ys__n500 & new_new_n12629__;
  assign new_new_n42681__ = ~ys__n1386 & new_new_n42680__;
  assign new_new_n42682__ = ~ys__n1386 & ~new_new_n42681__;
  assign new_new_n42683__ = ys__n33007 & ~new_new_n42682__;
  assign new_new_n42684__ = ys__n502 & ~ys__n2152;
  assign new_new_n42685__ = ~ys__n504 & ~ys__n2152;
  assign new_new_n42686__ = ~ys__n502 & new_new_n42685__;
  assign new_new_n42687__ = ~new_new_n42684__ & ~new_new_n42686__;
  assign new_new_n42688__ = ys__n28787 & ~new_new_n42687__;
  assign new_new_n42689__ = ys__n504 & ~ys__n2152;
  assign new_new_n42690__ = ~ys__n502 & new_new_n42689__;
  assign new_new_n42691__ = ys__n47185 & new_new_n42690__;
  assign new_new_n42692__ = ys__n500 & new_new_n12629__;
  assign new_new_n42693__ = ~ys__n1386 & new_new_n42692__;
  assign new_new_n42694__ = ys__n47340 & new_new_n42693__;
  assign new_new_n42695__ = ~new_new_n42691__ & ~new_new_n42694__;
  assign new_new_n42696__ = ~new_new_n42688__ & new_new_n42695__;
  assign new_new_n42697__ = ~new_new_n42683__ & new_new_n42696__;
  assign new_new_n42698__ = new_new_n42682__ & ~new_new_n42693__;
  assign new_new_n42699__ = ~new_new_n42690__ & new_new_n42698__;
  assign new_new_n42700__ = new_new_n42687__ & new_new_n42699__;
  assign ys__n31432 = ~new_new_n42697__ & ~new_new_n42700__;
  assign new_new_n42702__ = ys__n1386 & ys__n24191;
  assign new_new_n42703__ = ys__n47341 & ~ys__n2152;
  assign new_new_n42704__ = ys__n47342 & new_new_n35345__;
  assign new_new_n42705__ = ~new_new_n42673__ & new_new_n42704__;
  assign new_new_n42706__ = new_new_n41469__ & new_new_n42705__;
  assign new_new_n42707__ = ~new_new_n42703__ & ~new_new_n42706__;
  assign new_new_n42708__ = ~new_new_n42702__ & new_new_n42707__;
  assign ys__n33008 = ~new_new_n42678__ & ~new_new_n42708__;
  assign new_new_n42710__ = ~new_new_n42682__ & ys__n33008;
  assign new_new_n42711__ = ys__n28788 & ~new_new_n42687__;
  assign new_new_n42712__ = ys__n47184 & new_new_n42690__;
  assign new_new_n42713__ = ys__n47341 & new_new_n42693__;
  assign new_new_n42714__ = ~new_new_n42712__ & ~new_new_n42713__;
  assign new_new_n42715__ = ~new_new_n42711__ & new_new_n42714__;
  assign new_new_n42716__ = ~new_new_n42710__ & new_new_n42715__;
  assign ys__n31433 = ~new_new_n42700__ & ~new_new_n42716__;
  assign new_new_n42718__ = ys__n47342 & ~ys__n2152;
  assign new_new_n42719__ = ys__n714 & ys__n1386;
  assign new_new_n42720__ = ~new_new_n42718__ & ~new_new_n42719__;
  assign ys__n33009 = ~new_new_n42678__ & ~new_new_n42720__;
  assign new_new_n42722__ = ~new_new_n42682__ & ys__n33009;
  assign new_new_n42723__ = ys__n28789 & ~new_new_n42687__;
  assign new_new_n42724__ = ys__n46956 & new_new_n42690__;
  assign new_new_n42725__ = ys__n47342 & new_new_n42693__;
  assign new_new_n42726__ = ~new_new_n42724__ & ~new_new_n42725__;
  assign new_new_n42727__ = ~new_new_n42723__ & new_new_n42726__;
  assign new_new_n42728__ = ~new_new_n42722__ & new_new_n42727__;
  assign ys__n31434 = ~new_new_n42700__ & ~new_new_n42728__;
  assign new_new_n42730__ = ys__n46957 & new_new_n42690__;
  assign new_new_n42731__ = ys__n28790 & ~new_new_n42687__;
  assign new_new_n42732__ = ~new_new_n42730__ & ~new_new_n42731__;
  assign ys__n31435 = ~new_new_n42700__ & ~new_new_n42732__;
  assign new_new_n42734__ = ys__n46958 & new_new_n42690__;
  assign new_new_n42735__ = ys__n28791 & ~new_new_n42687__;
  assign new_new_n42736__ = ~new_new_n42734__ & ~new_new_n42735__;
  assign ys__n31436 = ~new_new_n42700__ & ~new_new_n42736__;
  assign new_new_n42738__ = ys__n46959 & new_new_n42690__;
  assign new_new_n42739__ = ys__n28792 & ~new_new_n42687__;
  assign new_new_n42740__ = ~new_new_n42738__ & ~new_new_n42739__;
  assign ys__n31437 = ~new_new_n42700__ & ~new_new_n42740__;
  assign new_new_n42742__ = ys__n46960 & new_new_n42690__;
  assign new_new_n42743__ = ys__n28793 & ~new_new_n42687__;
  assign new_new_n42744__ = ~new_new_n42742__ & ~new_new_n42743__;
  assign ys__n31438 = ~new_new_n42700__ & ~new_new_n42744__;
  assign new_new_n42746__ = ys__n46961 & new_new_n42690__;
  assign new_new_n42747__ = ys__n28794 & ~new_new_n42687__;
  assign new_new_n42748__ = ~new_new_n42746__ & ~new_new_n42747__;
  assign ys__n31439 = ~new_new_n42700__ & ~new_new_n42748__;
  assign new_new_n42750__ = ys__n836 & new_new_n12106__;
  assign new_new_n42751__ = ys__n47343 & new_new_n42750__;
  assign new_new_n42752__ = ~ys__n838 & ~new_new_n12106__;
  assign new_new_n42753__ = ~ys__n836 & new_new_n12106__;
  assign new_new_n42754__ = ~new_new_n42752__ & ~new_new_n42753__;
  assign new_new_n42755__ = ys__n47202 & ~new_new_n42754__;
  assign new_new_n42756__ = ~new_new_n42751__ & ~new_new_n42755__;
  assign new_new_n42757__ = ~new_new_n42750__ & new_new_n42754__;
  assign ys__n31440 = ~new_new_n42756__ & ~new_new_n42757__;
  assign new_new_n42759__ = ys__n47344 & new_new_n42750__;
  assign new_new_n42760__ = ys__n47203 & ~new_new_n42754__;
  assign new_new_n42761__ = ~new_new_n42759__ & ~new_new_n42760__;
  assign ys__n31441 = ~new_new_n42757__ & ~new_new_n42761__;
  assign new_new_n42763__ = ys__n47345 & new_new_n42750__;
  assign new_new_n42764__ = ys__n47204 & ~new_new_n42754__;
  assign new_new_n42765__ = ~new_new_n42763__ & ~new_new_n42764__;
  assign ys__n31442 = ~new_new_n42757__ & ~new_new_n42765__;
  assign new_new_n42767__ = ys__n47346 & new_new_n42750__;
  assign new_new_n42768__ = ys__n47205 & ~new_new_n42754__;
  assign new_new_n42769__ = ~new_new_n42767__ & ~new_new_n42768__;
  assign ys__n31443 = ~new_new_n42757__ & ~new_new_n42769__;
  assign new_new_n42771__ = ys__n47347 & new_new_n42750__;
  assign new_new_n42772__ = ys__n47206 & ~new_new_n42754__;
  assign new_new_n42773__ = ~new_new_n42771__ & ~new_new_n42772__;
  assign ys__n31444 = ~new_new_n42757__ & ~new_new_n42773__;
  assign new_new_n42775__ = ys__n47348 & new_new_n42750__;
  assign new_new_n42776__ = ys__n47207 & ~new_new_n42754__;
  assign new_new_n42777__ = ~new_new_n42775__ & ~new_new_n42776__;
  assign ys__n31445 = ~new_new_n42757__ & ~new_new_n42777__;
  assign new_new_n42779__ = ys__n47349 & new_new_n42750__;
  assign new_new_n42780__ = ys__n47208 & ~new_new_n42754__;
  assign new_new_n42781__ = ~new_new_n42779__ & ~new_new_n42780__;
  assign ys__n31446 = ~new_new_n42757__ & ~new_new_n42781__;
  assign new_new_n42783__ = ys__n47350 & new_new_n42750__;
  assign new_new_n42784__ = ys__n47209 & ~new_new_n42754__;
  assign new_new_n42785__ = ~new_new_n42783__ & ~new_new_n42784__;
  assign ys__n31447 = ~new_new_n42757__ & ~new_new_n42785__;
  assign new_new_n42787__ = ys__n47351 & new_new_n42750__;
  assign new_new_n42788__ = ys__n47210 & ~new_new_n42754__;
  assign new_new_n42789__ = ~new_new_n42787__ & ~new_new_n42788__;
  assign ys__n31448 = ~new_new_n42757__ & ~new_new_n42789__;
  assign new_new_n42791__ = ys__n47352 & new_new_n42750__;
  assign new_new_n42792__ = ys__n47211 & ~new_new_n42754__;
  assign new_new_n42793__ = ~new_new_n42791__ & ~new_new_n42792__;
  assign ys__n31449 = ~new_new_n42757__ & ~new_new_n42793__;
  assign new_new_n42795__ = ys__n47353 & new_new_n42750__;
  assign new_new_n42796__ = ys__n47212 & ~new_new_n42754__;
  assign new_new_n42797__ = ~new_new_n42795__ & ~new_new_n42796__;
  assign ys__n31450 = ~new_new_n42757__ & ~new_new_n42797__;
  assign new_new_n42799__ = ys__n47354 & new_new_n42750__;
  assign new_new_n42800__ = ys__n47213 & ~new_new_n42754__;
  assign new_new_n42801__ = ~new_new_n42799__ & ~new_new_n42800__;
  assign ys__n31451 = ~new_new_n42757__ & ~new_new_n42801__;
  assign new_new_n42803__ = ys__n47355 & new_new_n42750__;
  assign new_new_n42804__ = ys__n47214 & ~new_new_n42754__;
  assign new_new_n42805__ = ~new_new_n42803__ & ~new_new_n42804__;
  assign ys__n31452 = ~new_new_n42757__ & ~new_new_n42805__;
  assign new_new_n42807__ = ys__n47356 & new_new_n42750__;
  assign new_new_n42808__ = ys__n47215 & ~new_new_n42754__;
  assign new_new_n42809__ = ~new_new_n42807__ & ~new_new_n42808__;
  assign ys__n31453 = ~new_new_n42757__ & ~new_new_n42809__;
  assign new_new_n42811__ = ys__n47357 & new_new_n42750__;
  assign new_new_n42812__ = ys__n47216 & ~new_new_n42754__;
  assign new_new_n42813__ = ~new_new_n42811__ & ~new_new_n42812__;
  assign ys__n31454 = ~new_new_n42757__ & ~new_new_n42813__;
  assign new_new_n42815__ = ys__n47358 & new_new_n42750__;
  assign new_new_n42816__ = ys__n47217 & ~new_new_n42754__;
  assign new_new_n42817__ = ~new_new_n42815__ & ~new_new_n42816__;
  assign ys__n31455 = ~new_new_n42757__ & ~new_new_n42817__;
  assign new_new_n42819__ = ys__n47359 & new_new_n42750__;
  assign new_new_n42820__ = ys__n47218 & ~new_new_n42754__;
  assign new_new_n42821__ = ~new_new_n42819__ & ~new_new_n42820__;
  assign ys__n31456 = ~new_new_n42757__ & ~new_new_n42821__;
  assign new_new_n42823__ = ys__n47360 & new_new_n42750__;
  assign new_new_n42824__ = ys__n47219 & ~new_new_n42754__;
  assign new_new_n42825__ = ~new_new_n42823__ & ~new_new_n42824__;
  assign ys__n31457 = ~new_new_n42757__ & ~new_new_n42825__;
  assign new_new_n42827__ = ys__n47361 & new_new_n42750__;
  assign new_new_n42828__ = ys__n47220 & ~new_new_n42754__;
  assign new_new_n42829__ = ~new_new_n42827__ & ~new_new_n42828__;
  assign ys__n31458 = ~new_new_n42757__ & ~new_new_n42829__;
  assign new_new_n42831__ = ys__n47362 & new_new_n42750__;
  assign new_new_n42832__ = ys__n47221 & ~new_new_n42754__;
  assign new_new_n42833__ = ~new_new_n42831__ & ~new_new_n42832__;
  assign ys__n31459 = ~new_new_n42757__ & ~new_new_n42833__;
  assign new_new_n42835__ = ys__n47363 & new_new_n42750__;
  assign new_new_n42836__ = ys__n47222 & ~new_new_n42754__;
  assign new_new_n42837__ = ~new_new_n42835__ & ~new_new_n42836__;
  assign ys__n31460 = ~new_new_n42757__ & ~new_new_n42837__;
  assign new_new_n42839__ = ys__n47364 & new_new_n42750__;
  assign new_new_n42840__ = ys__n47223 & ~new_new_n42754__;
  assign new_new_n42841__ = ~new_new_n42839__ & ~new_new_n42840__;
  assign ys__n31461 = ~new_new_n42757__ & ~new_new_n42841__;
  assign new_new_n42843__ = ys__n47365 & new_new_n42750__;
  assign new_new_n42844__ = ys__n47224 & ~new_new_n42754__;
  assign new_new_n42845__ = ~new_new_n42843__ & ~new_new_n42844__;
  assign ys__n31462 = ~new_new_n42757__ & ~new_new_n42845__;
  assign new_new_n42847__ = ys__n47366 & new_new_n42750__;
  assign new_new_n42848__ = ys__n47225 & ~new_new_n42754__;
  assign new_new_n42849__ = ~new_new_n42847__ & ~new_new_n42848__;
  assign ys__n31463 = ~new_new_n42757__ & ~new_new_n42849__;
  assign new_new_n42851__ = ys__n47367 & new_new_n42750__;
  assign new_new_n42852__ = ys__n47226 & ~new_new_n42754__;
  assign new_new_n42853__ = ~new_new_n42851__ & ~new_new_n42852__;
  assign ys__n31464 = ~new_new_n42757__ & ~new_new_n42853__;
  assign new_new_n42855__ = ys__n47368 & new_new_n42750__;
  assign new_new_n42856__ = ys__n47227 & ~new_new_n42754__;
  assign new_new_n42857__ = ~new_new_n42855__ & ~new_new_n42856__;
  assign ys__n31465 = ~new_new_n42757__ & ~new_new_n42857__;
  assign new_new_n42859__ = ys__n47369 & new_new_n42750__;
  assign new_new_n42860__ = ys__n47228 & ~new_new_n42754__;
  assign new_new_n42861__ = ~new_new_n42859__ & ~new_new_n42860__;
  assign ys__n31466 = ~new_new_n42757__ & ~new_new_n42861__;
  assign new_new_n42863__ = ys__n47370 & new_new_n42750__;
  assign new_new_n42864__ = ys__n47229 & ~new_new_n42754__;
  assign new_new_n42865__ = ~new_new_n42863__ & ~new_new_n42864__;
  assign ys__n31467 = ~new_new_n42757__ & ~new_new_n42865__;
  assign new_new_n42867__ = ys__n47371 & new_new_n42750__;
  assign new_new_n42868__ = ys__n47230 & ~new_new_n42754__;
  assign new_new_n42869__ = ~new_new_n42867__ & ~new_new_n42868__;
  assign ys__n31468 = ~new_new_n42757__ & ~new_new_n42869__;
  assign new_new_n42871__ = ys__n47372 & new_new_n42750__;
  assign new_new_n42872__ = ys__n47231 & ~new_new_n42754__;
  assign new_new_n42873__ = ~new_new_n42871__ & ~new_new_n42872__;
  assign ys__n31469 = ~new_new_n42757__ & ~new_new_n42873__;
  assign new_new_n42875__ = ys__n47373 & new_new_n42750__;
  assign new_new_n42876__ = ys__n47232 & ~new_new_n42754__;
  assign new_new_n42877__ = ~new_new_n42875__ & ~new_new_n42876__;
  assign ys__n31470 = ~new_new_n42757__ & ~new_new_n42877__;
  assign new_new_n42879__ = ys__n47374 & new_new_n42750__;
  assign new_new_n42880__ = ys__n47233 & ~new_new_n42754__;
  assign new_new_n42881__ = ~new_new_n42879__ & ~new_new_n42880__;
  assign ys__n31471 = ~new_new_n42757__ & ~new_new_n42881__;
  assign new_new_n42883__ = ys__n47375 & new_new_n42750__;
  assign new_new_n42884__ = ys__n18762 & ~new_new_n42754__;
  assign new_new_n42885__ = ~new_new_n42883__ & ~new_new_n42884__;
  assign ys__n31472 = ~new_new_n42757__ & ~new_new_n42885__;
  assign new_new_n42887__ = ys__n47376 & new_new_n42750__;
  assign new_new_n42888__ = ys__n18750 & ~new_new_n42754__;
  assign new_new_n42889__ = ~new_new_n42887__ & ~new_new_n42888__;
  assign ys__n31473 = ~new_new_n42757__ & ~new_new_n42889__;
  assign new_new_n42891__ = ys__n47377 & new_new_n42750__;
  assign new_new_n42892__ = ys__n18753 & ~new_new_n42754__;
  assign new_new_n42893__ = ~new_new_n42891__ & ~new_new_n42892__;
  assign ys__n31474 = ~new_new_n42757__ & ~new_new_n42893__;
  assign new_new_n42895__ = ys__n832 & new_new_n12106__;
  assign new_new_n42896__ = ys__n47378 & new_new_n42895__;
  assign new_new_n42897__ = ~ys__n834 & ~new_new_n12106__;
  assign new_new_n42898__ = ~ys__n832 & new_new_n12106__;
  assign new_new_n42899__ = ~new_new_n42897__ & ~new_new_n42898__;
  assign new_new_n42900__ = ys__n47202 & ~new_new_n42899__;
  assign new_new_n42901__ = ~new_new_n42896__ & ~new_new_n42900__;
  assign new_new_n42902__ = ~new_new_n42895__ & new_new_n42899__;
  assign ys__n31475 = ~new_new_n42901__ & ~new_new_n42902__;
  assign new_new_n42904__ = ys__n47379 & new_new_n42895__;
  assign new_new_n42905__ = ys__n47203 & ~new_new_n42899__;
  assign new_new_n42906__ = ~new_new_n42904__ & ~new_new_n42905__;
  assign ys__n31476 = ~new_new_n42902__ & ~new_new_n42906__;
  assign new_new_n42908__ = ys__n47380 & new_new_n42895__;
  assign new_new_n42909__ = ys__n47204 & ~new_new_n42899__;
  assign new_new_n42910__ = ~new_new_n42908__ & ~new_new_n42909__;
  assign ys__n31477 = ~new_new_n42902__ & ~new_new_n42910__;
  assign new_new_n42912__ = ys__n47381 & new_new_n42895__;
  assign new_new_n42913__ = ys__n47205 & ~new_new_n42899__;
  assign new_new_n42914__ = ~new_new_n42912__ & ~new_new_n42913__;
  assign ys__n31478 = ~new_new_n42902__ & ~new_new_n42914__;
  assign new_new_n42916__ = ys__n47382 & new_new_n42895__;
  assign new_new_n42917__ = ys__n47206 & ~new_new_n42899__;
  assign new_new_n42918__ = ~new_new_n42916__ & ~new_new_n42917__;
  assign ys__n31479 = ~new_new_n42902__ & ~new_new_n42918__;
  assign new_new_n42920__ = ys__n47383 & new_new_n42895__;
  assign new_new_n42921__ = ys__n47207 & ~new_new_n42899__;
  assign new_new_n42922__ = ~new_new_n42920__ & ~new_new_n42921__;
  assign ys__n31480 = ~new_new_n42902__ & ~new_new_n42922__;
  assign new_new_n42924__ = ys__n47384 & new_new_n42895__;
  assign new_new_n42925__ = ys__n47208 & ~new_new_n42899__;
  assign new_new_n42926__ = ~new_new_n42924__ & ~new_new_n42925__;
  assign ys__n31481 = ~new_new_n42902__ & ~new_new_n42926__;
  assign new_new_n42928__ = ys__n47385 & new_new_n42895__;
  assign new_new_n42929__ = ys__n47209 & ~new_new_n42899__;
  assign new_new_n42930__ = ~new_new_n42928__ & ~new_new_n42929__;
  assign ys__n31482 = ~new_new_n42902__ & ~new_new_n42930__;
  assign new_new_n42932__ = ys__n47386 & new_new_n42895__;
  assign new_new_n42933__ = ys__n47210 & ~new_new_n42899__;
  assign new_new_n42934__ = ~new_new_n42932__ & ~new_new_n42933__;
  assign ys__n31483 = ~new_new_n42902__ & ~new_new_n42934__;
  assign new_new_n42936__ = ys__n47387 & new_new_n42895__;
  assign new_new_n42937__ = ys__n47211 & ~new_new_n42899__;
  assign new_new_n42938__ = ~new_new_n42936__ & ~new_new_n42937__;
  assign ys__n31484 = ~new_new_n42902__ & ~new_new_n42938__;
  assign new_new_n42940__ = ys__n47388 & new_new_n42895__;
  assign new_new_n42941__ = ys__n47212 & ~new_new_n42899__;
  assign new_new_n42942__ = ~new_new_n42940__ & ~new_new_n42941__;
  assign ys__n31485 = ~new_new_n42902__ & ~new_new_n42942__;
  assign new_new_n42944__ = ys__n47389 & new_new_n42895__;
  assign new_new_n42945__ = ys__n47213 & ~new_new_n42899__;
  assign new_new_n42946__ = ~new_new_n42944__ & ~new_new_n42945__;
  assign ys__n31486 = ~new_new_n42902__ & ~new_new_n42946__;
  assign new_new_n42948__ = ys__n47390 & new_new_n42895__;
  assign new_new_n42949__ = ys__n47214 & ~new_new_n42899__;
  assign new_new_n42950__ = ~new_new_n42948__ & ~new_new_n42949__;
  assign ys__n31487 = ~new_new_n42902__ & ~new_new_n42950__;
  assign new_new_n42952__ = ys__n47391 & new_new_n42895__;
  assign new_new_n42953__ = ys__n47215 & ~new_new_n42899__;
  assign new_new_n42954__ = ~new_new_n42952__ & ~new_new_n42953__;
  assign ys__n31488 = ~new_new_n42902__ & ~new_new_n42954__;
  assign new_new_n42956__ = ys__n47392 & new_new_n42895__;
  assign new_new_n42957__ = ys__n47216 & ~new_new_n42899__;
  assign new_new_n42958__ = ~new_new_n42956__ & ~new_new_n42957__;
  assign ys__n31489 = ~new_new_n42902__ & ~new_new_n42958__;
  assign new_new_n42960__ = ys__n47393 & new_new_n42895__;
  assign new_new_n42961__ = ys__n47217 & ~new_new_n42899__;
  assign new_new_n42962__ = ~new_new_n42960__ & ~new_new_n42961__;
  assign ys__n31490 = ~new_new_n42902__ & ~new_new_n42962__;
  assign new_new_n42964__ = ys__n47394 & new_new_n42895__;
  assign new_new_n42965__ = ys__n47218 & ~new_new_n42899__;
  assign new_new_n42966__ = ~new_new_n42964__ & ~new_new_n42965__;
  assign ys__n31491 = ~new_new_n42902__ & ~new_new_n42966__;
  assign new_new_n42968__ = ys__n47395 & new_new_n42895__;
  assign new_new_n42969__ = ys__n47219 & ~new_new_n42899__;
  assign new_new_n42970__ = ~new_new_n42968__ & ~new_new_n42969__;
  assign ys__n31492 = ~new_new_n42902__ & ~new_new_n42970__;
  assign new_new_n42972__ = ys__n47396 & new_new_n42895__;
  assign new_new_n42973__ = ys__n47220 & ~new_new_n42899__;
  assign new_new_n42974__ = ~new_new_n42972__ & ~new_new_n42973__;
  assign ys__n31493 = ~new_new_n42902__ & ~new_new_n42974__;
  assign new_new_n42976__ = ys__n47397 & new_new_n42895__;
  assign new_new_n42977__ = ys__n47221 & ~new_new_n42899__;
  assign new_new_n42978__ = ~new_new_n42976__ & ~new_new_n42977__;
  assign ys__n31494 = ~new_new_n42902__ & ~new_new_n42978__;
  assign new_new_n42980__ = ys__n47398 & new_new_n42895__;
  assign new_new_n42981__ = ys__n47222 & ~new_new_n42899__;
  assign new_new_n42982__ = ~new_new_n42980__ & ~new_new_n42981__;
  assign ys__n31495 = ~new_new_n42902__ & ~new_new_n42982__;
  assign new_new_n42984__ = ys__n47399 & new_new_n42895__;
  assign new_new_n42985__ = ys__n47223 & ~new_new_n42899__;
  assign new_new_n42986__ = ~new_new_n42984__ & ~new_new_n42985__;
  assign ys__n31496 = ~new_new_n42902__ & ~new_new_n42986__;
  assign new_new_n42988__ = ys__n47400 & new_new_n42895__;
  assign new_new_n42989__ = ys__n47224 & ~new_new_n42899__;
  assign new_new_n42990__ = ~new_new_n42988__ & ~new_new_n42989__;
  assign ys__n31497 = ~new_new_n42902__ & ~new_new_n42990__;
  assign new_new_n42992__ = ys__n47401 & new_new_n42895__;
  assign new_new_n42993__ = ys__n47225 & ~new_new_n42899__;
  assign new_new_n42994__ = ~new_new_n42992__ & ~new_new_n42993__;
  assign ys__n31498 = ~new_new_n42902__ & ~new_new_n42994__;
  assign new_new_n42996__ = ys__n47402 & new_new_n42895__;
  assign new_new_n42997__ = ys__n47226 & ~new_new_n42899__;
  assign new_new_n42998__ = ~new_new_n42996__ & ~new_new_n42997__;
  assign ys__n31499 = ~new_new_n42902__ & ~new_new_n42998__;
  assign new_new_n43000__ = ys__n47403 & new_new_n42895__;
  assign new_new_n43001__ = ys__n47227 & ~new_new_n42899__;
  assign new_new_n43002__ = ~new_new_n43000__ & ~new_new_n43001__;
  assign ys__n31500 = ~new_new_n42902__ & ~new_new_n43002__;
  assign new_new_n43004__ = ys__n47404 & new_new_n42895__;
  assign new_new_n43005__ = ys__n47228 & ~new_new_n42899__;
  assign new_new_n43006__ = ~new_new_n43004__ & ~new_new_n43005__;
  assign ys__n31501 = ~new_new_n42902__ & ~new_new_n43006__;
  assign new_new_n43008__ = ys__n47405 & new_new_n42895__;
  assign new_new_n43009__ = ys__n47229 & ~new_new_n42899__;
  assign new_new_n43010__ = ~new_new_n43008__ & ~new_new_n43009__;
  assign ys__n31502 = ~new_new_n42902__ & ~new_new_n43010__;
  assign new_new_n43012__ = ys__n47406 & new_new_n42895__;
  assign new_new_n43013__ = ys__n47230 & ~new_new_n42899__;
  assign new_new_n43014__ = ~new_new_n43012__ & ~new_new_n43013__;
  assign ys__n31503 = ~new_new_n42902__ & ~new_new_n43014__;
  assign new_new_n43016__ = ys__n47407 & new_new_n42895__;
  assign new_new_n43017__ = ys__n47231 & ~new_new_n42899__;
  assign new_new_n43018__ = ~new_new_n43016__ & ~new_new_n43017__;
  assign ys__n31504 = ~new_new_n42902__ & ~new_new_n43018__;
  assign new_new_n43020__ = ys__n47408 & new_new_n42895__;
  assign new_new_n43021__ = ys__n47232 & ~new_new_n42899__;
  assign new_new_n43022__ = ~new_new_n43020__ & ~new_new_n43021__;
  assign ys__n31505 = ~new_new_n42902__ & ~new_new_n43022__;
  assign new_new_n43024__ = ys__n47409 & new_new_n42895__;
  assign new_new_n43025__ = ys__n47233 & ~new_new_n42899__;
  assign new_new_n43026__ = ~new_new_n43024__ & ~new_new_n43025__;
  assign ys__n31506 = ~new_new_n42902__ & ~new_new_n43026__;
  assign new_new_n43028__ = ys__n47410 & new_new_n42895__;
  assign new_new_n43029__ = ys__n18762 & ~new_new_n42899__;
  assign new_new_n43030__ = ~new_new_n43028__ & ~new_new_n43029__;
  assign ys__n31507 = ~new_new_n42902__ & ~new_new_n43030__;
  assign new_new_n43032__ = ys__n47411 & new_new_n42895__;
  assign new_new_n43033__ = ys__n18750 & ~new_new_n42899__;
  assign new_new_n43034__ = ~new_new_n43032__ & ~new_new_n43033__;
  assign ys__n31508 = ~new_new_n42902__ & ~new_new_n43034__;
  assign new_new_n43036__ = ys__n47412 & new_new_n42895__;
  assign new_new_n43037__ = ys__n18753 & ~new_new_n42899__;
  assign new_new_n43038__ = ~new_new_n43036__ & ~new_new_n43037__;
  assign ys__n31509 = ~new_new_n42902__ & ~new_new_n43038__;
  assign new_new_n43040__ = ys__n834 & new_new_n12106__;
  assign new_new_n43041__ = ys__n47413 & new_new_n43040__;
  assign new_new_n43042__ = ~ys__n836 & ~new_new_n12106__;
  assign new_new_n43043__ = ~ys__n834 & new_new_n12106__;
  assign new_new_n43044__ = ~new_new_n43042__ & ~new_new_n43043__;
  assign new_new_n43045__ = ys__n47202 & ~new_new_n43044__;
  assign new_new_n43046__ = ~new_new_n43041__ & ~new_new_n43045__;
  assign new_new_n43047__ = ~new_new_n43040__ & new_new_n43044__;
  assign ys__n31510 = ~new_new_n43046__ & ~new_new_n43047__;
  assign new_new_n43049__ = ys__n47414 & new_new_n43040__;
  assign new_new_n43050__ = ys__n47203 & ~new_new_n43044__;
  assign new_new_n43051__ = ~new_new_n43049__ & ~new_new_n43050__;
  assign ys__n31511 = ~new_new_n43047__ & ~new_new_n43051__;
  assign new_new_n43053__ = ys__n47415 & new_new_n43040__;
  assign new_new_n43054__ = ys__n47204 & ~new_new_n43044__;
  assign new_new_n43055__ = ~new_new_n43053__ & ~new_new_n43054__;
  assign ys__n31512 = ~new_new_n43047__ & ~new_new_n43055__;
  assign new_new_n43057__ = ys__n47416 & new_new_n43040__;
  assign new_new_n43058__ = ys__n47205 & ~new_new_n43044__;
  assign new_new_n43059__ = ~new_new_n43057__ & ~new_new_n43058__;
  assign ys__n31513 = ~new_new_n43047__ & ~new_new_n43059__;
  assign new_new_n43061__ = ys__n47417 & new_new_n43040__;
  assign new_new_n43062__ = ys__n47206 & ~new_new_n43044__;
  assign new_new_n43063__ = ~new_new_n43061__ & ~new_new_n43062__;
  assign ys__n31514 = ~new_new_n43047__ & ~new_new_n43063__;
  assign new_new_n43065__ = ys__n47418 & new_new_n43040__;
  assign new_new_n43066__ = ys__n47207 & ~new_new_n43044__;
  assign new_new_n43067__ = ~new_new_n43065__ & ~new_new_n43066__;
  assign ys__n31515 = ~new_new_n43047__ & ~new_new_n43067__;
  assign new_new_n43069__ = ys__n47419 & new_new_n43040__;
  assign new_new_n43070__ = ys__n47208 & ~new_new_n43044__;
  assign new_new_n43071__ = ~new_new_n43069__ & ~new_new_n43070__;
  assign ys__n31516 = ~new_new_n43047__ & ~new_new_n43071__;
  assign new_new_n43073__ = ys__n47420 & new_new_n43040__;
  assign new_new_n43074__ = ys__n47209 & ~new_new_n43044__;
  assign new_new_n43075__ = ~new_new_n43073__ & ~new_new_n43074__;
  assign ys__n31517 = ~new_new_n43047__ & ~new_new_n43075__;
  assign new_new_n43077__ = ys__n47421 & new_new_n43040__;
  assign new_new_n43078__ = ys__n47210 & ~new_new_n43044__;
  assign new_new_n43079__ = ~new_new_n43077__ & ~new_new_n43078__;
  assign ys__n31518 = ~new_new_n43047__ & ~new_new_n43079__;
  assign new_new_n43081__ = ys__n47422 & new_new_n43040__;
  assign new_new_n43082__ = ys__n47211 & ~new_new_n43044__;
  assign new_new_n43083__ = ~new_new_n43081__ & ~new_new_n43082__;
  assign ys__n31519 = ~new_new_n43047__ & ~new_new_n43083__;
  assign new_new_n43085__ = ys__n47423 & new_new_n43040__;
  assign new_new_n43086__ = ys__n47212 & ~new_new_n43044__;
  assign new_new_n43087__ = ~new_new_n43085__ & ~new_new_n43086__;
  assign ys__n31520 = ~new_new_n43047__ & ~new_new_n43087__;
  assign new_new_n43089__ = ys__n47424 & new_new_n43040__;
  assign new_new_n43090__ = ys__n47213 & ~new_new_n43044__;
  assign new_new_n43091__ = ~new_new_n43089__ & ~new_new_n43090__;
  assign ys__n31521 = ~new_new_n43047__ & ~new_new_n43091__;
  assign new_new_n43093__ = ys__n47425 & new_new_n43040__;
  assign new_new_n43094__ = ys__n47214 & ~new_new_n43044__;
  assign new_new_n43095__ = ~new_new_n43093__ & ~new_new_n43094__;
  assign ys__n31522 = ~new_new_n43047__ & ~new_new_n43095__;
  assign new_new_n43097__ = ys__n47426 & new_new_n43040__;
  assign new_new_n43098__ = ys__n47215 & ~new_new_n43044__;
  assign new_new_n43099__ = ~new_new_n43097__ & ~new_new_n43098__;
  assign ys__n31523 = ~new_new_n43047__ & ~new_new_n43099__;
  assign new_new_n43101__ = ys__n47427 & new_new_n43040__;
  assign new_new_n43102__ = ys__n47216 & ~new_new_n43044__;
  assign new_new_n43103__ = ~new_new_n43101__ & ~new_new_n43102__;
  assign ys__n31524 = ~new_new_n43047__ & ~new_new_n43103__;
  assign new_new_n43105__ = ys__n47428 & new_new_n43040__;
  assign new_new_n43106__ = ys__n47217 & ~new_new_n43044__;
  assign new_new_n43107__ = ~new_new_n43105__ & ~new_new_n43106__;
  assign ys__n31525 = ~new_new_n43047__ & ~new_new_n43107__;
  assign new_new_n43109__ = ys__n47429 & new_new_n43040__;
  assign new_new_n43110__ = ys__n47218 & ~new_new_n43044__;
  assign new_new_n43111__ = ~new_new_n43109__ & ~new_new_n43110__;
  assign ys__n31526 = ~new_new_n43047__ & ~new_new_n43111__;
  assign new_new_n43113__ = ys__n47430 & new_new_n43040__;
  assign new_new_n43114__ = ys__n47219 & ~new_new_n43044__;
  assign new_new_n43115__ = ~new_new_n43113__ & ~new_new_n43114__;
  assign ys__n31527 = ~new_new_n43047__ & ~new_new_n43115__;
  assign new_new_n43117__ = ys__n47431 & new_new_n43040__;
  assign new_new_n43118__ = ys__n47220 & ~new_new_n43044__;
  assign new_new_n43119__ = ~new_new_n43117__ & ~new_new_n43118__;
  assign ys__n31528 = ~new_new_n43047__ & ~new_new_n43119__;
  assign new_new_n43121__ = ys__n47432 & new_new_n43040__;
  assign new_new_n43122__ = ys__n47221 & ~new_new_n43044__;
  assign new_new_n43123__ = ~new_new_n43121__ & ~new_new_n43122__;
  assign ys__n31529 = ~new_new_n43047__ & ~new_new_n43123__;
  assign new_new_n43125__ = ys__n47433 & new_new_n43040__;
  assign new_new_n43126__ = ys__n47222 & ~new_new_n43044__;
  assign new_new_n43127__ = ~new_new_n43125__ & ~new_new_n43126__;
  assign ys__n31530 = ~new_new_n43047__ & ~new_new_n43127__;
  assign new_new_n43129__ = ys__n47434 & new_new_n43040__;
  assign new_new_n43130__ = ys__n47223 & ~new_new_n43044__;
  assign new_new_n43131__ = ~new_new_n43129__ & ~new_new_n43130__;
  assign ys__n31531 = ~new_new_n43047__ & ~new_new_n43131__;
  assign new_new_n43133__ = ys__n47435 & new_new_n43040__;
  assign new_new_n43134__ = ys__n47224 & ~new_new_n43044__;
  assign new_new_n43135__ = ~new_new_n43133__ & ~new_new_n43134__;
  assign ys__n31532 = ~new_new_n43047__ & ~new_new_n43135__;
  assign new_new_n43137__ = ys__n47436 & new_new_n43040__;
  assign new_new_n43138__ = ys__n47225 & ~new_new_n43044__;
  assign new_new_n43139__ = ~new_new_n43137__ & ~new_new_n43138__;
  assign ys__n31533 = ~new_new_n43047__ & ~new_new_n43139__;
  assign new_new_n43141__ = ys__n47437 & new_new_n43040__;
  assign new_new_n43142__ = ys__n47226 & ~new_new_n43044__;
  assign new_new_n43143__ = ~new_new_n43141__ & ~new_new_n43142__;
  assign ys__n31534 = ~new_new_n43047__ & ~new_new_n43143__;
  assign new_new_n43145__ = ys__n47438 & new_new_n43040__;
  assign new_new_n43146__ = ys__n47227 & ~new_new_n43044__;
  assign new_new_n43147__ = ~new_new_n43145__ & ~new_new_n43146__;
  assign ys__n31535 = ~new_new_n43047__ & ~new_new_n43147__;
  assign new_new_n43149__ = ys__n47439 & new_new_n43040__;
  assign new_new_n43150__ = ys__n47228 & ~new_new_n43044__;
  assign new_new_n43151__ = ~new_new_n43149__ & ~new_new_n43150__;
  assign ys__n31536 = ~new_new_n43047__ & ~new_new_n43151__;
  assign new_new_n43153__ = ys__n47440 & new_new_n43040__;
  assign new_new_n43154__ = ys__n47229 & ~new_new_n43044__;
  assign new_new_n43155__ = ~new_new_n43153__ & ~new_new_n43154__;
  assign ys__n31537 = ~new_new_n43047__ & ~new_new_n43155__;
  assign new_new_n43157__ = ys__n47441 & new_new_n43040__;
  assign new_new_n43158__ = ys__n47230 & ~new_new_n43044__;
  assign new_new_n43159__ = ~new_new_n43157__ & ~new_new_n43158__;
  assign ys__n31538 = ~new_new_n43047__ & ~new_new_n43159__;
  assign new_new_n43161__ = ys__n47442 & new_new_n43040__;
  assign new_new_n43162__ = ys__n47231 & ~new_new_n43044__;
  assign new_new_n43163__ = ~new_new_n43161__ & ~new_new_n43162__;
  assign ys__n31539 = ~new_new_n43047__ & ~new_new_n43163__;
  assign new_new_n43165__ = ys__n47443 & new_new_n43040__;
  assign new_new_n43166__ = ys__n47232 & ~new_new_n43044__;
  assign new_new_n43167__ = ~new_new_n43165__ & ~new_new_n43166__;
  assign ys__n31540 = ~new_new_n43047__ & ~new_new_n43167__;
  assign new_new_n43169__ = ys__n47444 & new_new_n43040__;
  assign new_new_n43170__ = ys__n47233 & ~new_new_n43044__;
  assign new_new_n43171__ = ~new_new_n43169__ & ~new_new_n43170__;
  assign ys__n31541 = ~new_new_n43047__ & ~new_new_n43171__;
  assign new_new_n43173__ = ys__n47445 & new_new_n43040__;
  assign new_new_n43174__ = ys__n18762 & ~new_new_n43044__;
  assign new_new_n43175__ = ~new_new_n43173__ & ~new_new_n43174__;
  assign ys__n31542 = ~new_new_n43047__ & ~new_new_n43175__;
  assign new_new_n43177__ = ys__n47446 & new_new_n43040__;
  assign new_new_n43178__ = ys__n18750 & ~new_new_n43044__;
  assign new_new_n43179__ = ~new_new_n43177__ & ~new_new_n43178__;
  assign ys__n31543 = ~new_new_n43047__ & ~new_new_n43179__;
  assign new_new_n43181__ = ys__n47447 & new_new_n43040__;
  assign new_new_n43182__ = ys__n18753 & ~new_new_n43044__;
  assign new_new_n43183__ = ~new_new_n43181__ & ~new_new_n43182__;
  assign ys__n31544 = ~new_new_n43047__ & ~new_new_n43183__;
  assign new_new_n43185__ = ys__n35057 & ~ys__n35059;
  assign new_new_n43186__ = ~ys__n488 & ys__n490;
  assign new_new_n43187__ = ~new_new_n43185__ & new_new_n43186__;
  assign new_new_n43188__ = ~ys__n35057 & ~ys__n35059;
  assign new_new_n43189__ = ~ys__n488 & ~ys__n490;
  assign new_new_n43190__ = ~new_new_n43188__ & new_new_n43189__;
  assign new_new_n43191__ = ~new_new_n43187__ & ~new_new_n43190__;
  assign new_new_n43192__ = ys__n488 & ys__n490;
  assign new_new_n43193__ = ~new_new_n43186__ & ~new_new_n43192__;
  assign new_new_n43194__ = ys__n488 & ~ys__n490;
  assign new_new_n43195__ = ~new_new_n43189__ & ~new_new_n43194__;
  assign new_new_n43196__ = new_new_n43193__ & new_new_n43195__;
  assign ys__n31559 = ~new_new_n43191__ & ~new_new_n43196__;
  assign new_new_n43198__ = ~ys__n35057 & ys__n35059;
  assign new_new_n43199__ = new_new_n43194__ & ~new_new_n43198__;
  assign new_new_n43200__ = ~new_new_n43187__ & ~new_new_n43199__;
  assign ys__n31560 = ~new_new_n43196__ & ~new_new_n43200__;
  assign new_new_n43202__ = ~new_new_n43188__ & ~new_new_n43198__;
  assign new_new_n43203__ = new_new_n43189__ & ~new_new_n43202__;
  assign new_new_n43204__ = ys__n35057 & ys__n35059;
  assign new_new_n43205__ = new_new_n43186__ & new_new_n43204__;
  assign new_new_n43206__ = new_new_n43185__ & new_new_n43194__;
  assign new_new_n43207__ = ~new_new_n43205__ & ~new_new_n43206__;
  assign new_new_n43208__ = ~new_new_n43203__ & new_new_n43207__;
  assign ys__n31562 = ~new_new_n43196__ & ~new_new_n43208__;
  assign new_new_n43210__ = new_new_n43194__ & new_new_n43198__;
  assign ys__n31564 = ~new_new_n43196__ & new_new_n43210__;
  assign new_new_n43212__ = new_new_n43185__ & new_new_n43186__;
  assign ys__n31567 = ~new_new_n43196__ & new_new_n43212__;
  assign new_new_n43214__ = ~new_new_n43189__ & ~new_new_n43192__;
  assign new_new_n43215__ = ~new_new_n43186__ & ~new_new_n43194__;
  assign new_new_n43216__ = new_new_n43214__ & new_new_n43215__;
  assign new_new_n43217__ = new_new_n43204__ & ~new_new_n43214__;
  assign ys__n31571 = ~new_new_n43216__ & new_new_n43217__;
  assign new_new_n43219__ = ys__n830 & new_new_n12106__;
  assign new_new_n43220__ = ys__n47449 & new_new_n43219__;
  assign new_new_n43221__ = ~ys__n832 & ~new_new_n12106__;
  assign new_new_n43222__ = ~ys__n830 & new_new_n12106__;
  assign new_new_n43223__ = ~new_new_n43221__ & ~new_new_n43222__;
  assign new_new_n43224__ = ys__n47202 & ~new_new_n43223__;
  assign new_new_n43225__ = ~new_new_n43220__ & ~new_new_n43224__;
  assign new_new_n43226__ = ~new_new_n43219__ & new_new_n43223__;
  assign ys__n31740 = ~new_new_n43225__ & ~new_new_n43226__;
  assign new_new_n43228__ = ys__n47450 & new_new_n43219__;
  assign new_new_n43229__ = ys__n47203 & ~new_new_n43223__;
  assign new_new_n43230__ = ~new_new_n43228__ & ~new_new_n43229__;
  assign ys__n31741 = ~new_new_n43226__ & ~new_new_n43230__;
  assign new_new_n43232__ = ys__n47451 & new_new_n43219__;
  assign new_new_n43233__ = ys__n47204 & ~new_new_n43223__;
  assign new_new_n43234__ = ~new_new_n43232__ & ~new_new_n43233__;
  assign ys__n31742 = ~new_new_n43226__ & ~new_new_n43234__;
  assign new_new_n43236__ = ys__n47452 & new_new_n43219__;
  assign new_new_n43237__ = ys__n47205 & ~new_new_n43223__;
  assign new_new_n43238__ = ~new_new_n43236__ & ~new_new_n43237__;
  assign ys__n31743 = ~new_new_n43226__ & ~new_new_n43238__;
  assign new_new_n43240__ = ys__n47453 & new_new_n43219__;
  assign new_new_n43241__ = ys__n47206 & ~new_new_n43223__;
  assign new_new_n43242__ = ~new_new_n43240__ & ~new_new_n43241__;
  assign ys__n31744 = ~new_new_n43226__ & ~new_new_n43242__;
  assign new_new_n43244__ = ys__n47454 & new_new_n43219__;
  assign new_new_n43245__ = ys__n47207 & ~new_new_n43223__;
  assign new_new_n43246__ = ~new_new_n43244__ & ~new_new_n43245__;
  assign ys__n31745 = ~new_new_n43226__ & ~new_new_n43246__;
  assign new_new_n43248__ = ys__n47455 & new_new_n43219__;
  assign new_new_n43249__ = ys__n47208 & ~new_new_n43223__;
  assign new_new_n43250__ = ~new_new_n43248__ & ~new_new_n43249__;
  assign ys__n31746 = ~new_new_n43226__ & ~new_new_n43250__;
  assign new_new_n43252__ = ys__n47456 & new_new_n43219__;
  assign new_new_n43253__ = ys__n47209 & ~new_new_n43223__;
  assign new_new_n43254__ = ~new_new_n43252__ & ~new_new_n43253__;
  assign ys__n31747 = ~new_new_n43226__ & ~new_new_n43254__;
  assign new_new_n43256__ = ys__n47457 & new_new_n43219__;
  assign new_new_n43257__ = ys__n47210 & ~new_new_n43223__;
  assign new_new_n43258__ = ~new_new_n43256__ & ~new_new_n43257__;
  assign ys__n31748 = ~new_new_n43226__ & ~new_new_n43258__;
  assign new_new_n43260__ = ys__n47458 & new_new_n43219__;
  assign new_new_n43261__ = ys__n47211 & ~new_new_n43223__;
  assign new_new_n43262__ = ~new_new_n43260__ & ~new_new_n43261__;
  assign ys__n31749 = ~new_new_n43226__ & ~new_new_n43262__;
  assign new_new_n43264__ = ys__n47459 & new_new_n43219__;
  assign new_new_n43265__ = ys__n47212 & ~new_new_n43223__;
  assign new_new_n43266__ = ~new_new_n43264__ & ~new_new_n43265__;
  assign ys__n31750 = ~new_new_n43226__ & ~new_new_n43266__;
  assign new_new_n43268__ = ys__n47460 & new_new_n43219__;
  assign new_new_n43269__ = ys__n47213 & ~new_new_n43223__;
  assign new_new_n43270__ = ~new_new_n43268__ & ~new_new_n43269__;
  assign ys__n31751 = ~new_new_n43226__ & ~new_new_n43270__;
  assign new_new_n43272__ = ys__n47461 & new_new_n43219__;
  assign new_new_n43273__ = ys__n47214 & ~new_new_n43223__;
  assign new_new_n43274__ = ~new_new_n43272__ & ~new_new_n43273__;
  assign ys__n31752 = ~new_new_n43226__ & ~new_new_n43274__;
  assign new_new_n43276__ = ys__n47462 & new_new_n43219__;
  assign new_new_n43277__ = ys__n47215 & ~new_new_n43223__;
  assign new_new_n43278__ = ~new_new_n43276__ & ~new_new_n43277__;
  assign ys__n31753 = ~new_new_n43226__ & ~new_new_n43278__;
  assign new_new_n43280__ = ys__n47463 & new_new_n43219__;
  assign new_new_n43281__ = ys__n47216 & ~new_new_n43223__;
  assign new_new_n43282__ = ~new_new_n43280__ & ~new_new_n43281__;
  assign ys__n31754 = ~new_new_n43226__ & ~new_new_n43282__;
  assign new_new_n43284__ = ys__n47464 & new_new_n43219__;
  assign new_new_n43285__ = ys__n47217 & ~new_new_n43223__;
  assign new_new_n43286__ = ~new_new_n43284__ & ~new_new_n43285__;
  assign ys__n31755 = ~new_new_n43226__ & ~new_new_n43286__;
  assign new_new_n43288__ = ys__n47465 & new_new_n43219__;
  assign new_new_n43289__ = ys__n47218 & ~new_new_n43223__;
  assign new_new_n43290__ = ~new_new_n43288__ & ~new_new_n43289__;
  assign ys__n31756 = ~new_new_n43226__ & ~new_new_n43290__;
  assign new_new_n43292__ = ys__n47466 & new_new_n43219__;
  assign new_new_n43293__ = ys__n47219 & ~new_new_n43223__;
  assign new_new_n43294__ = ~new_new_n43292__ & ~new_new_n43293__;
  assign ys__n31757 = ~new_new_n43226__ & ~new_new_n43294__;
  assign new_new_n43296__ = ys__n47467 & new_new_n43219__;
  assign new_new_n43297__ = ys__n47220 & ~new_new_n43223__;
  assign new_new_n43298__ = ~new_new_n43296__ & ~new_new_n43297__;
  assign ys__n31758 = ~new_new_n43226__ & ~new_new_n43298__;
  assign new_new_n43300__ = ys__n47468 & new_new_n43219__;
  assign new_new_n43301__ = ys__n47221 & ~new_new_n43223__;
  assign new_new_n43302__ = ~new_new_n43300__ & ~new_new_n43301__;
  assign ys__n31759 = ~new_new_n43226__ & ~new_new_n43302__;
  assign new_new_n43304__ = ys__n47469 & new_new_n43219__;
  assign new_new_n43305__ = ys__n47222 & ~new_new_n43223__;
  assign new_new_n43306__ = ~new_new_n43304__ & ~new_new_n43305__;
  assign ys__n31760 = ~new_new_n43226__ & ~new_new_n43306__;
  assign new_new_n43308__ = ys__n47470 & new_new_n43219__;
  assign new_new_n43309__ = ys__n47223 & ~new_new_n43223__;
  assign new_new_n43310__ = ~new_new_n43308__ & ~new_new_n43309__;
  assign ys__n31761 = ~new_new_n43226__ & ~new_new_n43310__;
  assign new_new_n43312__ = ys__n47471 & new_new_n43219__;
  assign new_new_n43313__ = ys__n47224 & ~new_new_n43223__;
  assign new_new_n43314__ = ~new_new_n43312__ & ~new_new_n43313__;
  assign ys__n31762 = ~new_new_n43226__ & ~new_new_n43314__;
  assign new_new_n43316__ = ys__n47472 & new_new_n43219__;
  assign new_new_n43317__ = ys__n47225 & ~new_new_n43223__;
  assign new_new_n43318__ = ~new_new_n43316__ & ~new_new_n43317__;
  assign ys__n31763 = ~new_new_n43226__ & ~new_new_n43318__;
  assign new_new_n43320__ = ys__n47473 & new_new_n43219__;
  assign new_new_n43321__ = ys__n47226 & ~new_new_n43223__;
  assign new_new_n43322__ = ~new_new_n43320__ & ~new_new_n43321__;
  assign ys__n31764 = ~new_new_n43226__ & ~new_new_n43322__;
  assign new_new_n43324__ = ys__n47474 & new_new_n43219__;
  assign new_new_n43325__ = ys__n47227 & ~new_new_n43223__;
  assign new_new_n43326__ = ~new_new_n43324__ & ~new_new_n43325__;
  assign ys__n31765 = ~new_new_n43226__ & ~new_new_n43326__;
  assign new_new_n43328__ = ys__n47475 & new_new_n43219__;
  assign new_new_n43329__ = ys__n47228 & ~new_new_n43223__;
  assign new_new_n43330__ = ~new_new_n43328__ & ~new_new_n43329__;
  assign ys__n31766 = ~new_new_n43226__ & ~new_new_n43330__;
  assign new_new_n43332__ = ys__n47476 & new_new_n43219__;
  assign new_new_n43333__ = ys__n47229 & ~new_new_n43223__;
  assign new_new_n43334__ = ~new_new_n43332__ & ~new_new_n43333__;
  assign ys__n31767 = ~new_new_n43226__ & ~new_new_n43334__;
  assign new_new_n43336__ = ys__n47477 & new_new_n43219__;
  assign new_new_n43337__ = ys__n47230 & ~new_new_n43223__;
  assign new_new_n43338__ = ~new_new_n43336__ & ~new_new_n43337__;
  assign ys__n31768 = ~new_new_n43226__ & ~new_new_n43338__;
  assign new_new_n43340__ = ys__n47478 & new_new_n43219__;
  assign new_new_n43341__ = ys__n47231 & ~new_new_n43223__;
  assign new_new_n43342__ = ~new_new_n43340__ & ~new_new_n43341__;
  assign ys__n31769 = ~new_new_n43226__ & ~new_new_n43342__;
  assign new_new_n43344__ = ys__n47479 & new_new_n43219__;
  assign new_new_n43345__ = ys__n47232 & ~new_new_n43223__;
  assign new_new_n43346__ = ~new_new_n43344__ & ~new_new_n43345__;
  assign ys__n31770 = ~new_new_n43226__ & ~new_new_n43346__;
  assign new_new_n43348__ = ys__n47480 & new_new_n43219__;
  assign new_new_n43349__ = ys__n47233 & ~new_new_n43223__;
  assign new_new_n43350__ = ~new_new_n43348__ & ~new_new_n43349__;
  assign ys__n31771 = ~new_new_n43226__ & ~new_new_n43350__;
  assign new_new_n43352__ = ys__n47481 & new_new_n43219__;
  assign new_new_n43353__ = ys__n18762 & ~new_new_n43223__;
  assign new_new_n43354__ = ~new_new_n43352__ & ~new_new_n43353__;
  assign ys__n31772 = ~new_new_n43226__ & ~new_new_n43354__;
  assign new_new_n43356__ = ys__n47482 & new_new_n43219__;
  assign new_new_n43357__ = ys__n18750 & ~new_new_n43223__;
  assign new_new_n43358__ = ~new_new_n43356__ & ~new_new_n43357__;
  assign ys__n31773 = ~new_new_n43226__ & ~new_new_n43358__;
  assign new_new_n43360__ = ys__n47483 & new_new_n43219__;
  assign new_new_n43361__ = ys__n18753 & ~new_new_n43223__;
  assign new_new_n43362__ = ~new_new_n43360__ & ~new_new_n43361__;
  assign ys__n31774 = ~new_new_n43226__ & ~new_new_n43362__;
  assign new_new_n43364__ = ys__n858 & new_new_n12106__;
  assign new_new_n43365__ = ys__n47484 & new_new_n43364__;
  assign new_new_n43366__ = ~ys__n830 & ~new_new_n12106__;
  assign new_new_n43367__ = ~ys__n858 & new_new_n12106__;
  assign new_new_n43368__ = ~new_new_n43366__ & ~new_new_n43367__;
  assign new_new_n43369__ = ys__n47202 & ~new_new_n43368__;
  assign new_new_n43370__ = ~new_new_n43365__ & ~new_new_n43369__;
  assign new_new_n43371__ = ~new_new_n43364__ & new_new_n43368__;
  assign ys__n31775 = ~new_new_n43370__ & ~new_new_n43371__;
  assign new_new_n43373__ = ys__n47485 & new_new_n43364__;
  assign new_new_n43374__ = ys__n47203 & ~new_new_n43368__;
  assign new_new_n43375__ = ~new_new_n43373__ & ~new_new_n43374__;
  assign ys__n31776 = ~new_new_n43371__ & ~new_new_n43375__;
  assign new_new_n43377__ = ys__n47486 & new_new_n43364__;
  assign new_new_n43378__ = ys__n47204 & ~new_new_n43368__;
  assign new_new_n43379__ = ~new_new_n43377__ & ~new_new_n43378__;
  assign ys__n31777 = ~new_new_n43371__ & ~new_new_n43379__;
  assign new_new_n43381__ = ys__n47487 & new_new_n43364__;
  assign new_new_n43382__ = ys__n47205 & ~new_new_n43368__;
  assign new_new_n43383__ = ~new_new_n43381__ & ~new_new_n43382__;
  assign ys__n31778 = ~new_new_n43371__ & ~new_new_n43383__;
  assign new_new_n43385__ = ys__n47488 & new_new_n43364__;
  assign new_new_n43386__ = ys__n47206 & ~new_new_n43368__;
  assign new_new_n43387__ = ~new_new_n43385__ & ~new_new_n43386__;
  assign ys__n31779 = ~new_new_n43371__ & ~new_new_n43387__;
  assign new_new_n43389__ = ys__n47489 & new_new_n43364__;
  assign new_new_n43390__ = ys__n47207 & ~new_new_n43368__;
  assign new_new_n43391__ = ~new_new_n43389__ & ~new_new_n43390__;
  assign ys__n31780 = ~new_new_n43371__ & ~new_new_n43391__;
  assign new_new_n43393__ = ys__n47490 & new_new_n43364__;
  assign new_new_n43394__ = ys__n47208 & ~new_new_n43368__;
  assign new_new_n43395__ = ~new_new_n43393__ & ~new_new_n43394__;
  assign ys__n31781 = ~new_new_n43371__ & ~new_new_n43395__;
  assign new_new_n43397__ = ys__n47491 & new_new_n43364__;
  assign new_new_n43398__ = ys__n47209 & ~new_new_n43368__;
  assign new_new_n43399__ = ~new_new_n43397__ & ~new_new_n43398__;
  assign ys__n31782 = ~new_new_n43371__ & ~new_new_n43399__;
  assign new_new_n43401__ = ys__n47492 & new_new_n43364__;
  assign new_new_n43402__ = ys__n47210 & ~new_new_n43368__;
  assign new_new_n43403__ = ~new_new_n43401__ & ~new_new_n43402__;
  assign ys__n31783 = ~new_new_n43371__ & ~new_new_n43403__;
  assign new_new_n43405__ = ys__n47493 & new_new_n43364__;
  assign new_new_n43406__ = ys__n47211 & ~new_new_n43368__;
  assign new_new_n43407__ = ~new_new_n43405__ & ~new_new_n43406__;
  assign ys__n31784 = ~new_new_n43371__ & ~new_new_n43407__;
  assign new_new_n43409__ = ys__n47494 & new_new_n43364__;
  assign new_new_n43410__ = ys__n47212 & ~new_new_n43368__;
  assign new_new_n43411__ = ~new_new_n43409__ & ~new_new_n43410__;
  assign ys__n31785 = ~new_new_n43371__ & ~new_new_n43411__;
  assign new_new_n43413__ = ys__n47495 & new_new_n43364__;
  assign new_new_n43414__ = ys__n47213 & ~new_new_n43368__;
  assign new_new_n43415__ = ~new_new_n43413__ & ~new_new_n43414__;
  assign ys__n31786 = ~new_new_n43371__ & ~new_new_n43415__;
  assign new_new_n43417__ = ys__n47496 & new_new_n43364__;
  assign new_new_n43418__ = ys__n47214 & ~new_new_n43368__;
  assign new_new_n43419__ = ~new_new_n43417__ & ~new_new_n43418__;
  assign ys__n31787 = ~new_new_n43371__ & ~new_new_n43419__;
  assign new_new_n43421__ = ys__n47497 & new_new_n43364__;
  assign new_new_n43422__ = ys__n47215 & ~new_new_n43368__;
  assign new_new_n43423__ = ~new_new_n43421__ & ~new_new_n43422__;
  assign ys__n31788 = ~new_new_n43371__ & ~new_new_n43423__;
  assign new_new_n43425__ = ys__n47498 & new_new_n43364__;
  assign new_new_n43426__ = ys__n47216 & ~new_new_n43368__;
  assign new_new_n43427__ = ~new_new_n43425__ & ~new_new_n43426__;
  assign ys__n31789 = ~new_new_n43371__ & ~new_new_n43427__;
  assign new_new_n43429__ = ys__n47499 & new_new_n43364__;
  assign new_new_n43430__ = ys__n47217 & ~new_new_n43368__;
  assign new_new_n43431__ = ~new_new_n43429__ & ~new_new_n43430__;
  assign ys__n31790 = ~new_new_n43371__ & ~new_new_n43431__;
  assign new_new_n43433__ = ys__n47500 & new_new_n43364__;
  assign new_new_n43434__ = ys__n47218 & ~new_new_n43368__;
  assign new_new_n43435__ = ~new_new_n43433__ & ~new_new_n43434__;
  assign ys__n31791 = ~new_new_n43371__ & ~new_new_n43435__;
  assign new_new_n43437__ = ys__n47501 & new_new_n43364__;
  assign new_new_n43438__ = ys__n47219 & ~new_new_n43368__;
  assign new_new_n43439__ = ~new_new_n43437__ & ~new_new_n43438__;
  assign ys__n31792 = ~new_new_n43371__ & ~new_new_n43439__;
  assign new_new_n43441__ = ys__n47502 & new_new_n43364__;
  assign new_new_n43442__ = ys__n47220 & ~new_new_n43368__;
  assign new_new_n43443__ = ~new_new_n43441__ & ~new_new_n43442__;
  assign ys__n31793 = ~new_new_n43371__ & ~new_new_n43443__;
  assign new_new_n43445__ = ys__n47503 & new_new_n43364__;
  assign new_new_n43446__ = ys__n47221 & ~new_new_n43368__;
  assign new_new_n43447__ = ~new_new_n43445__ & ~new_new_n43446__;
  assign ys__n31794 = ~new_new_n43371__ & ~new_new_n43447__;
  assign new_new_n43449__ = ys__n47504 & new_new_n43364__;
  assign new_new_n43450__ = ys__n47222 & ~new_new_n43368__;
  assign new_new_n43451__ = ~new_new_n43449__ & ~new_new_n43450__;
  assign ys__n31795 = ~new_new_n43371__ & ~new_new_n43451__;
  assign new_new_n43453__ = ys__n47505 & new_new_n43364__;
  assign new_new_n43454__ = ys__n47223 & ~new_new_n43368__;
  assign new_new_n43455__ = ~new_new_n43453__ & ~new_new_n43454__;
  assign ys__n31796 = ~new_new_n43371__ & ~new_new_n43455__;
  assign new_new_n43457__ = ys__n47506 & new_new_n43364__;
  assign new_new_n43458__ = ys__n47224 & ~new_new_n43368__;
  assign new_new_n43459__ = ~new_new_n43457__ & ~new_new_n43458__;
  assign ys__n31797 = ~new_new_n43371__ & ~new_new_n43459__;
  assign new_new_n43461__ = ys__n47507 & new_new_n43364__;
  assign new_new_n43462__ = ys__n47225 & ~new_new_n43368__;
  assign new_new_n43463__ = ~new_new_n43461__ & ~new_new_n43462__;
  assign ys__n31798 = ~new_new_n43371__ & ~new_new_n43463__;
  assign new_new_n43465__ = ys__n47508 & new_new_n43364__;
  assign new_new_n43466__ = ys__n47226 & ~new_new_n43368__;
  assign new_new_n43467__ = ~new_new_n43465__ & ~new_new_n43466__;
  assign ys__n31799 = ~new_new_n43371__ & ~new_new_n43467__;
  assign new_new_n43469__ = ys__n47509 & new_new_n43364__;
  assign new_new_n43470__ = ys__n47227 & ~new_new_n43368__;
  assign new_new_n43471__ = ~new_new_n43469__ & ~new_new_n43470__;
  assign ys__n31800 = ~new_new_n43371__ & ~new_new_n43471__;
  assign new_new_n43473__ = ys__n47510 & new_new_n43364__;
  assign new_new_n43474__ = ys__n47228 & ~new_new_n43368__;
  assign new_new_n43475__ = ~new_new_n43473__ & ~new_new_n43474__;
  assign ys__n31801 = ~new_new_n43371__ & ~new_new_n43475__;
  assign new_new_n43477__ = ys__n47511 & new_new_n43364__;
  assign new_new_n43478__ = ys__n47229 & ~new_new_n43368__;
  assign new_new_n43479__ = ~new_new_n43477__ & ~new_new_n43478__;
  assign ys__n31802 = ~new_new_n43371__ & ~new_new_n43479__;
  assign new_new_n43481__ = ys__n47512 & new_new_n43364__;
  assign new_new_n43482__ = ys__n47230 & ~new_new_n43368__;
  assign new_new_n43483__ = ~new_new_n43481__ & ~new_new_n43482__;
  assign ys__n31803 = ~new_new_n43371__ & ~new_new_n43483__;
  assign new_new_n43485__ = ys__n47513 & new_new_n43364__;
  assign new_new_n43486__ = ys__n47231 & ~new_new_n43368__;
  assign new_new_n43487__ = ~new_new_n43485__ & ~new_new_n43486__;
  assign ys__n31804 = ~new_new_n43371__ & ~new_new_n43487__;
  assign new_new_n43489__ = ys__n47514 & new_new_n43364__;
  assign new_new_n43490__ = ys__n47232 & ~new_new_n43368__;
  assign new_new_n43491__ = ~new_new_n43489__ & ~new_new_n43490__;
  assign ys__n31805 = ~new_new_n43371__ & ~new_new_n43491__;
  assign new_new_n43493__ = ys__n47515 & new_new_n43364__;
  assign new_new_n43494__ = ys__n47233 & ~new_new_n43368__;
  assign new_new_n43495__ = ~new_new_n43493__ & ~new_new_n43494__;
  assign ys__n31806 = ~new_new_n43371__ & ~new_new_n43495__;
  assign new_new_n43497__ = ys__n47516 & new_new_n43364__;
  assign new_new_n43498__ = ys__n18762 & ~new_new_n43368__;
  assign new_new_n43499__ = ~new_new_n43497__ & ~new_new_n43498__;
  assign ys__n31807 = ~new_new_n43371__ & ~new_new_n43499__;
  assign new_new_n43501__ = ys__n47517 & new_new_n43364__;
  assign new_new_n43502__ = ys__n18750 & ~new_new_n43368__;
  assign new_new_n43503__ = ~new_new_n43501__ & ~new_new_n43502__;
  assign ys__n31808 = ~new_new_n43371__ & ~new_new_n43503__;
  assign new_new_n43505__ = ys__n47518 & new_new_n43364__;
  assign new_new_n43506__ = ys__n18753 & ~new_new_n43368__;
  assign new_new_n43507__ = ~new_new_n43505__ & ~new_new_n43506__;
  assign ys__n31809 = ~new_new_n43371__ & ~new_new_n43507__;
  assign new_new_n43509__ = ys__n856 & new_new_n12106__;
  assign new_new_n43510__ = ys__n47519 & new_new_n43509__;
  assign new_new_n43511__ = ~ys__n858 & ~new_new_n12106__;
  assign new_new_n43512__ = ~ys__n856 & new_new_n12106__;
  assign new_new_n43513__ = ~new_new_n43511__ & ~new_new_n43512__;
  assign new_new_n43514__ = ys__n47202 & ~new_new_n43513__;
  assign new_new_n43515__ = ~new_new_n43510__ & ~new_new_n43514__;
  assign new_new_n43516__ = ~new_new_n43509__ & new_new_n43513__;
  assign ys__n31810 = ~new_new_n43515__ & ~new_new_n43516__;
  assign new_new_n43518__ = ys__n47520 & new_new_n43509__;
  assign new_new_n43519__ = ys__n47203 & ~new_new_n43513__;
  assign new_new_n43520__ = ~new_new_n43518__ & ~new_new_n43519__;
  assign ys__n31811 = ~new_new_n43516__ & ~new_new_n43520__;
  assign new_new_n43522__ = ys__n47521 & new_new_n43509__;
  assign new_new_n43523__ = ys__n47204 & ~new_new_n43513__;
  assign new_new_n43524__ = ~new_new_n43522__ & ~new_new_n43523__;
  assign ys__n31812 = ~new_new_n43516__ & ~new_new_n43524__;
  assign new_new_n43526__ = ys__n47522 & new_new_n43509__;
  assign new_new_n43527__ = ys__n47205 & ~new_new_n43513__;
  assign new_new_n43528__ = ~new_new_n43526__ & ~new_new_n43527__;
  assign ys__n31813 = ~new_new_n43516__ & ~new_new_n43528__;
  assign new_new_n43530__ = ys__n47523 & new_new_n43509__;
  assign new_new_n43531__ = ys__n47206 & ~new_new_n43513__;
  assign new_new_n43532__ = ~new_new_n43530__ & ~new_new_n43531__;
  assign ys__n31814 = ~new_new_n43516__ & ~new_new_n43532__;
  assign new_new_n43534__ = ys__n47524 & new_new_n43509__;
  assign new_new_n43535__ = ys__n47207 & ~new_new_n43513__;
  assign new_new_n43536__ = ~new_new_n43534__ & ~new_new_n43535__;
  assign ys__n31815 = ~new_new_n43516__ & ~new_new_n43536__;
  assign new_new_n43538__ = ys__n47525 & new_new_n43509__;
  assign new_new_n43539__ = ys__n47208 & ~new_new_n43513__;
  assign new_new_n43540__ = ~new_new_n43538__ & ~new_new_n43539__;
  assign ys__n31816 = ~new_new_n43516__ & ~new_new_n43540__;
  assign new_new_n43542__ = ys__n47526 & new_new_n43509__;
  assign new_new_n43543__ = ys__n47209 & ~new_new_n43513__;
  assign new_new_n43544__ = ~new_new_n43542__ & ~new_new_n43543__;
  assign ys__n31817 = ~new_new_n43516__ & ~new_new_n43544__;
  assign new_new_n43546__ = ys__n47527 & new_new_n43509__;
  assign new_new_n43547__ = ys__n47210 & ~new_new_n43513__;
  assign new_new_n43548__ = ~new_new_n43546__ & ~new_new_n43547__;
  assign ys__n31818 = ~new_new_n43516__ & ~new_new_n43548__;
  assign new_new_n43550__ = ys__n47528 & new_new_n43509__;
  assign new_new_n43551__ = ys__n47211 & ~new_new_n43513__;
  assign new_new_n43552__ = ~new_new_n43550__ & ~new_new_n43551__;
  assign ys__n31819 = ~new_new_n43516__ & ~new_new_n43552__;
  assign new_new_n43554__ = ys__n47529 & new_new_n43509__;
  assign new_new_n43555__ = ys__n47212 & ~new_new_n43513__;
  assign new_new_n43556__ = ~new_new_n43554__ & ~new_new_n43555__;
  assign ys__n31820 = ~new_new_n43516__ & ~new_new_n43556__;
  assign new_new_n43558__ = ys__n47530 & new_new_n43509__;
  assign new_new_n43559__ = ys__n47213 & ~new_new_n43513__;
  assign new_new_n43560__ = ~new_new_n43558__ & ~new_new_n43559__;
  assign ys__n31821 = ~new_new_n43516__ & ~new_new_n43560__;
  assign new_new_n43562__ = ys__n47531 & new_new_n43509__;
  assign new_new_n43563__ = ys__n47214 & ~new_new_n43513__;
  assign new_new_n43564__ = ~new_new_n43562__ & ~new_new_n43563__;
  assign ys__n31822 = ~new_new_n43516__ & ~new_new_n43564__;
  assign new_new_n43566__ = ys__n47532 & new_new_n43509__;
  assign new_new_n43567__ = ys__n47215 & ~new_new_n43513__;
  assign new_new_n43568__ = ~new_new_n43566__ & ~new_new_n43567__;
  assign ys__n31823 = ~new_new_n43516__ & ~new_new_n43568__;
  assign new_new_n43570__ = ys__n47533 & new_new_n43509__;
  assign new_new_n43571__ = ys__n47216 & ~new_new_n43513__;
  assign new_new_n43572__ = ~new_new_n43570__ & ~new_new_n43571__;
  assign ys__n31824 = ~new_new_n43516__ & ~new_new_n43572__;
  assign new_new_n43574__ = ys__n47534 & new_new_n43509__;
  assign new_new_n43575__ = ys__n47217 & ~new_new_n43513__;
  assign new_new_n43576__ = ~new_new_n43574__ & ~new_new_n43575__;
  assign ys__n31825 = ~new_new_n43516__ & ~new_new_n43576__;
  assign new_new_n43578__ = ys__n47535 & new_new_n43509__;
  assign new_new_n43579__ = ys__n47218 & ~new_new_n43513__;
  assign new_new_n43580__ = ~new_new_n43578__ & ~new_new_n43579__;
  assign ys__n31826 = ~new_new_n43516__ & ~new_new_n43580__;
  assign new_new_n43582__ = ys__n47536 & new_new_n43509__;
  assign new_new_n43583__ = ys__n47219 & ~new_new_n43513__;
  assign new_new_n43584__ = ~new_new_n43582__ & ~new_new_n43583__;
  assign ys__n31827 = ~new_new_n43516__ & ~new_new_n43584__;
  assign new_new_n43586__ = ys__n47537 & new_new_n43509__;
  assign new_new_n43587__ = ys__n47220 & ~new_new_n43513__;
  assign new_new_n43588__ = ~new_new_n43586__ & ~new_new_n43587__;
  assign ys__n31828 = ~new_new_n43516__ & ~new_new_n43588__;
  assign new_new_n43590__ = ys__n47538 & new_new_n43509__;
  assign new_new_n43591__ = ys__n47221 & ~new_new_n43513__;
  assign new_new_n43592__ = ~new_new_n43590__ & ~new_new_n43591__;
  assign ys__n31829 = ~new_new_n43516__ & ~new_new_n43592__;
  assign new_new_n43594__ = ys__n47539 & new_new_n43509__;
  assign new_new_n43595__ = ys__n47222 & ~new_new_n43513__;
  assign new_new_n43596__ = ~new_new_n43594__ & ~new_new_n43595__;
  assign ys__n31830 = ~new_new_n43516__ & ~new_new_n43596__;
  assign new_new_n43598__ = ys__n47540 & new_new_n43509__;
  assign new_new_n43599__ = ys__n47223 & ~new_new_n43513__;
  assign new_new_n43600__ = ~new_new_n43598__ & ~new_new_n43599__;
  assign ys__n31831 = ~new_new_n43516__ & ~new_new_n43600__;
  assign new_new_n43602__ = ys__n47541 & new_new_n43509__;
  assign new_new_n43603__ = ys__n47224 & ~new_new_n43513__;
  assign new_new_n43604__ = ~new_new_n43602__ & ~new_new_n43603__;
  assign ys__n31832 = ~new_new_n43516__ & ~new_new_n43604__;
  assign new_new_n43606__ = ys__n47542 & new_new_n43509__;
  assign new_new_n43607__ = ys__n47225 & ~new_new_n43513__;
  assign new_new_n43608__ = ~new_new_n43606__ & ~new_new_n43607__;
  assign ys__n31833 = ~new_new_n43516__ & ~new_new_n43608__;
  assign new_new_n43610__ = ys__n47543 & new_new_n43509__;
  assign new_new_n43611__ = ys__n47226 & ~new_new_n43513__;
  assign new_new_n43612__ = ~new_new_n43610__ & ~new_new_n43611__;
  assign ys__n31834 = ~new_new_n43516__ & ~new_new_n43612__;
  assign new_new_n43614__ = ys__n47544 & new_new_n43509__;
  assign new_new_n43615__ = ys__n47227 & ~new_new_n43513__;
  assign new_new_n43616__ = ~new_new_n43614__ & ~new_new_n43615__;
  assign ys__n31835 = ~new_new_n43516__ & ~new_new_n43616__;
  assign new_new_n43618__ = ys__n47545 & new_new_n43509__;
  assign new_new_n43619__ = ys__n47228 & ~new_new_n43513__;
  assign new_new_n43620__ = ~new_new_n43618__ & ~new_new_n43619__;
  assign ys__n31836 = ~new_new_n43516__ & ~new_new_n43620__;
  assign new_new_n43622__ = ys__n47546 & new_new_n43509__;
  assign new_new_n43623__ = ys__n47229 & ~new_new_n43513__;
  assign new_new_n43624__ = ~new_new_n43622__ & ~new_new_n43623__;
  assign ys__n31837 = ~new_new_n43516__ & ~new_new_n43624__;
  assign new_new_n43626__ = ys__n47547 & new_new_n43509__;
  assign new_new_n43627__ = ys__n47230 & ~new_new_n43513__;
  assign new_new_n43628__ = ~new_new_n43626__ & ~new_new_n43627__;
  assign ys__n31838 = ~new_new_n43516__ & ~new_new_n43628__;
  assign new_new_n43630__ = ys__n47548 & new_new_n43509__;
  assign new_new_n43631__ = ys__n47231 & ~new_new_n43513__;
  assign new_new_n43632__ = ~new_new_n43630__ & ~new_new_n43631__;
  assign ys__n31839 = ~new_new_n43516__ & ~new_new_n43632__;
  assign new_new_n43634__ = ys__n47549 & new_new_n43509__;
  assign new_new_n43635__ = ys__n47232 & ~new_new_n43513__;
  assign new_new_n43636__ = ~new_new_n43634__ & ~new_new_n43635__;
  assign ys__n31840 = ~new_new_n43516__ & ~new_new_n43636__;
  assign new_new_n43638__ = ys__n47550 & new_new_n43509__;
  assign new_new_n43639__ = ys__n47233 & ~new_new_n43513__;
  assign new_new_n43640__ = ~new_new_n43638__ & ~new_new_n43639__;
  assign ys__n31841 = ~new_new_n43516__ & ~new_new_n43640__;
  assign new_new_n43642__ = ys__n47551 & new_new_n43509__;
  assign new_new_n43643__ = ys__n18762 & ~new_new_n43513__;
  assign new_new_n43644__ = ~new_new_n43642__ & ~new_new_n43643__;
  assign ys__n31842 = ~new_new_n43516__ & ~new_new_n43644__;
  assign new_new_n43646__ = ys__n47552 & new_new_n43509__;
  assign new_new_n43647__ = ys__n18750 & ~new_new_n43513__;
  assign new_new_n43648__ = ~new_new_n43646__ & ~new_new_n43647__;
  assign ys__n31843 = ~new_new_n43516__ & ~new_new_n43648__;
  assign new_new_n43650__ = ys__n47553 & new_new_n43509__;
  assign new_new_n43651__ = ys__n18753 & ~new_new_n43513__;
  assign new_new_n43652__ = ~new_new_n43650__ & ~new_new_n43651__;
  assign ys__n31844 = ~new_new_n43516__ & ~new_new_n43652__;
  assign new_new_n43654__ = ys__n854 & new_new_n12106__;
  assign new_new_n43655__ = ys__n47554 & new_new_n43654__;
  assign new_new_n43656__ = ~ys__n856 & ~new_new_n12106__;
  assign new_new_n43657__ = ~ys__n854 & new_new_n12106__;
  assign new_new_n43658__ = ~new_new_n43656__ & ~new_new_n43657__;
  assign new_new_n43659__ = ys__n47202 & ~new_new_n43658__;
  assign new_new_n43660__ = ~new_new_n43655__ & ~new_new_n43659__;
  assign new_new_n43661__ = ~new_new_n43654__ & new_new_n43658__;
  assign ys__n31845 = ~new_new_n43660__ & ~new_new_n43661__;
  assign new_new_n43663__ = ys__n47555 & new_new_n43654__;
  assign new_new_n43664__ = ys__n47203 & ~new_new_n43658__;
  assign new_new_n43665__ = ~new_new_n43663__ & ~new_new_n43664__;
  assign ys__n31846 = ~new_new_n43661__ & ~new_new_n43665__;
  assign new_new_n43667__ = ys__n47556 & new_new_n43654__;
  assign new_new_n43668__ = ys__n47204 & ~new_new_n43658__;
  assign new_new_n43669__ = ~new_new_n43667__ & ~new_new_n43668__;
  assign ys__n31847 = ~new_new_n43661__ & ~new_new_n43669__;
  assign new_new_n43671__ = ys__n47557 & new_new_n43654__;
  assign new_new_n43672__ = ys__n47205 & ~new_new_n43658__;
  assign new_new_n43673__ = ~new_new_n43671__ & ~new_new_n43672__;
  assign ys__n31848 = ~new_new_n43661__ & ~new_new_n43673__;
  assign new_new_n43675__ = ys__n47558 & new_new_n43654__;
  assign new_new_n43676__ = ys__n47206 & ~new_new_n43658__;
  assign new_new_n43677__ = ~new_new_n43675__ & ~new_new_n43676__;
  assign ys__n31849 = ~new_new_n43661__ & ~new_new_n43677__;
  assign new_new_n43679__ = ys__n47559 & new_new_n43654__;
  assign new_new_n43680__ = ys__n47207 & ~new_new_n43658__;
  assign new_new_n43681__ = ~new_new_n43679__ & ~new_new_n43680__;
  assign ys__n31850 = ~new_new_n43661__ & ~new_new_n43681__;
  assign new_new_n43683__ = ys__n47560 & new_new_n43654__;
  assign new_new_n43684__ = ys__n47208 & ~new_new_n43658__;
  assign new_new_n43685__ = ~new_new_n43683__ & ~new_new_n43684__;
  assign ys__n31851 = ~new_new_n43661__ & ~new_new_n43685__;
  assign new_new_n43687__ = ys__n47561 & new_new_n43654__;
  assign new_new_n43688__ = ys__n47209 & ~new_new_n43658__;
  assign new_new_n43689__ = ~new_new_n43687__ & ~new_new_n43688__;
  assign ys__n31852 = ~new_new_n43661__ & ~new_new_n43689__;
  assign new_new_n43691__ = ys__n47562 & new_new_n43654__;
  assign new_new_n43692__ = ys__n47210 & ~new_new_n43658__;
  assign new_new_n43693__ = ~new_new_n43691__ & ~new_new_n43692__;
  assign ys__n31853 = ~new_new_n43661__ & ~new_new_n43693__;
  assign new_new_n43695__ = ys__n47563 & new_new_n43654__;
  assign new_new_n43696__ = ys__n47211 & ~new_new_n43658__;
  assign new_new_n43697__ = ~new_new_n43695__ & ~new_new_n43696__;
  assign ys__n31854 = ~new_new_n43661__ & ~new_new_n43697__;
  assign new_new_n43699__ = ys__n47564 & new_new_n43654__;
  assign new_new_n43700__ = ys__n47212 & ~new_new_n43658__;
  assign new_new_n43701__ = ~new_new_n43699__ & ~new_new_n43700__;
  assign ys__n31855 = ~new_new_n43661__ & ~new_new_n43701__;
  assign new_new_n43703__ = ys__n47565 & new_new_n43654__;
  assign new_new_n43704__ = ys__n47213 & ~new_new_n43658__;
  assign new_new_n43705__ = ~new_new_n43703__ & ~new_new_n43704__;
  assign ys__n31856 = ~new_new_n43661__ & ~new_new_n43705__;
  assign new_new_n43707__ = ys__n47566 & new_new_n43654__;
  assign new_new_n43708__ = ys__n47214 & ~new_new_n43658__;
  assign new_new_n43709__ = ~new_new_n43707__ & ~new_new_n43708__;
  assign ys__n31857 = ~new_new_n43661__ & ~new_new_n43709__;
  assign new_new_n43711__ = ys__n47567 & new_new_n43654__;
  assign new_new_n43712__ = ys__n47215 & ~new_new_n43658__;
  assign new_new_n43713__ = ~new_new_n43711__ & ~new_new_n43712__;
  assign ys__n31858 = ~new_new_n43661__ & ~new_new_n43713__;
  assign new_new_n43715__ = ys__n47568 & new_new_n43654__;
  assign new_new_n43716__ = ys__n47216 & ~new_new_n43658__;
  assign new_new_n43717__ = ~new_new_n43715__ & ~new_new_n43716__;
  assign ys__n31859 = ~new_new_n43661__ & ~new_new_n43717__;
  assign new_new_n43719__ = ys__n47569 & new_new_n43654__;
  assign new_new_n43720__ = ys__n47217 & ~new_new_n43658__;
  assign new_new_n43721__ = ~new_new_n43719__ & ~new_new_n43720__;
  assign ys__n31860 = ~new_new_n43661__ & ~new_new_n43721__;
  assign new_new_n43723__ = ys__n47570 & new_new_n43654__;
  assign new_new_n43724__ = ys__n47218 & ~new_new_n43658__;
  assign new_new_n43725__ = ~new_new_n43723__ & ~new_new_n43724__;
  assign ys__n31861 = ~new_new_n43661__ & ~new_new_n43725__;
  assign new_new_n43727__ = ys__n47571 & new_new_n43654__;
  assign new_new_n43728__ = ys__n47219 & ~new_new_n43658__;
  assign new_new_n43729__ = ~new_new_n43727__ & ~new_new_n43728__;
  assign ys__n31862 = ~new_new_n43661__ & ~new_new_n43729__;
  assign new_new_n43731__ = ys__n47572 & new_new_n43654__;
  assign new_new_n43732__ = ys__n47220 & ~new_new_n43658__;
  assign new_new_n43733__ = ~new_new_n43731__ & ~new_new_n43732__;
  assign ys__n31863 = ~new_new_n43661__ & ~new_new_n43733__;
  assign new_new_n43735__ = ys__n47573 & new_new_n43654__;
  assign new_new_n43736__ = ys__n47221 & ~new_new_n43658__;
  assign new_new_n43737__ = ~new_new_n43735__ & ~new_new_n43736__;
  assign ys__n31864 = ~new_new_n43661__ & ~new_new_n43737__;
  assign new_new_n43739__ = ys__n47574 & new_new_n43654__;
  assign new_new_n43740__ = ys__n47222 & ~new_new_n43658__;
  assign new_new_n43741__ = ~new_new_n43739__ & ~new_new_n43740__;
  assign ys__n31865 = ~new_new_n43661__ & ~new_new_n43741__;
  assign new_new_n43743__ = ys__n47575 & new_new_n43654__;
  assign new_new_n43744__ = ys__n47223 & ~new_new_n43658__;
  assign new_new_n43745__ = ~new_new_n43743__ & ~new_new_n43744__;
  assign ys__n31866 = ~new_new_n43661__ & ~new_new_n43745__;
  assign new_new_n43747__ = ys__n47576 & new_new_n43654__;
  assign new_new_n43748__ = ys__n47224 & ~new_new_n43658__;
  assign new_new_n43749__ = ~new_new_n43747__ & ~new_new_n43748__;
  assign ys__n31867 = ~new_new_n43661__ & ~new_new_n43749__;
  assign new_new_n43751__ = ys__n47577 & new_new_n43654__;
  assign new_new_n43752__ = ys__n47225 & ~new_new_n43658__;
  assign new_new_n43753__ = ~new_new_n43751__ & ~new_new_n43752__;
  assign ys__n31868 = ~new_new_n43661__ & ~new_new_n43753__;
  assign new_new_n43755__ = ys__n47578 & new_new_n43654__;
  assign new_new_n43756__ = ys__n47226 & ~new_new_n43658__;
  assign new_new_n43757__ = ~new_new_n43755__ & ~new_new_n43756__;
  assign ys__n31869 = ~new_new_n43661__ & ~new_new_n43757__;
  assign new_new_n43759__ = ys__n47579 & new_new_n43654__;
  assign new_new_n43760__ = ys__n47227 & ~new_new_n43658__;
  assign new_new_n43761__ = ~new_new_n43759__ & ~new_new_n43760__;
  assign ys__n31870 = ~new_new_n43661__ & ~new_new_n43761__;
  assign new_new_n43763__ = ys__n47580 & new_new_n43654__;
  assign new_new_n43764__ = ys__n47228 & ~new_new_n43658__;
  assign new_new_n43765__ = ~new_new_n43763__ & ~new_new_n43764__;
  assign ys__n31871 = ~new_new_n43661__ & ~new_new_n43765__;
  assign new_new_n43767__ = ys__n47581 & new_new_n43654__;
  assign new_new_n43768__ = ys__n47229 & ~new_new_n43658__;
  assign new_new_n43769__ = ~new_new_n43767__ & ~new_new_n43768__;
  assign ys__n31872 = ~new_new_n43661__ & ~new_new_n43769__;
  assign new_new_n43771__ = ys__n47582 & new_new_n43654__;
  assign new_new_n43772__ = ys__n47230 & ~new_new_n43658__;
  assign new_new_n43773__ = ~new_new_n43771__ & ~new_new_n43772__;
  assign ys__n31873 = ~new_new_n43661__ & ~new_new_n43773__;
  assign new_new_n43775__ = ys__n47583 & new_new_n43654__;
  assign new_new_n43776__ = ys__n47231 & ~new_new_n43658__;
  assign new_new_n43777__ = ~new_new_n43775__ & ~new_new_n43776__;
  assign ys__n31874 = ~new_new_n43661__ & ~new_new_n43777__;
  assign new_new_n43779__ = ys__n47584 & new_new_n43654__;
  assign new_new_n43780__ = ys__n47232 & ~new_new_n43658__;
  assign new_new_n43781__ = ~new_new_n43779__ & ~new_new_n43780__;
  assign ys__n31875 = ~new_new_n43661__ & ~new_new_n43781__;
  assign new_new_n43783__ = ys__n47585 & new_new_n43654__;
  assign new_new_n43784__ = ys__n47233 & ~new_new_n43658__;
  assign new_new_n43785__ = ~new_new_n43783__ & ~new_new_n43784__;
  assign ys__n31876 = ~new_new_n43661__ & ~new_new_n43785__;
  assign new_new_n43787__ = ys__n47586 & new_new_n43654__;
  assign new_new_n43788__ = ys__n18762 & ~new_new_n43658__;
  assign new_new_n43789__ = ~new_new_n43787__ & ~new_new_n43788__;
  assign ys__n31877 = ~new_new_n43661__ & ~new_new_n43789__;
  assign new_new_n43791__ = ys__n47587 & new_new_n43654__;
  assign new_new_n43792__ = ys__n18750 & ~new_new_n43658__;
  assign new_new_n43793__ = ~new_new_n43791__ & ~new_new_n43792__;
  assign ys__n31878 = ~new_new_n43661__ & ~new_new_n43793__;
  assign new_new_n43795__ = ys__n47588 & new_new_n43654__;
  assign new_new_n43796__ = ys__n18753 & ~new_new_n43658__;
  assign new_new_n43797__ = ~new_new_n43795__ & ~new_new_n43796__;
  assign ys__n31879 = ~new_new_n43661__ & ~new_new_n43797__;
  assign new_new_n43799__ = ys__n852 & new_new_n12106__;
  assign new_new_n43800__ = ys__n47589 & new_new_n43799__;
  assign new_new_n43801__ = ~ys__n854 & ~new_new_n12106__;
  assign new_new_n43802__ = ~ys__n852 & new_new_n12106__;
  assign new_new_n43803__ = ~new_new_n43801__ & ~new_new_n43802__;
  assign new_new_n43804__ = ys__n47202 & ~new_new_n43803__;
  assign new_new_n43805__ = ~new_new_n43800__ & ~new_new_n43804__;
  assign new_new_n43806__ = ~new_new_n43799__ & new_new_n43803__;
  assign ys__n31880 = ~new_new_n43805__ & ~new_new_n43806__;
  assign new_new_n43808__ = ys__n47590 & new_new_n43799__;
  assign new_new_n43809__ = ys__n47203 & ~new_new_n43803__;
  assign new_new_n43810__ = ~new_new_n43808__ & ~new_new_n43809__;
  assign ys__n31881 = ~new_new_n43806__ & ~new_new_n43810__;
  assign new_new_n43812__ = ys__n47591 & new_new_n43799__;
  assign new_new_n43813__ = ys__n47204 & ~new_new_n43803__;
  assign new_new_n43814__ = ~new_new_n43812__ & ~new_new_n43813__;
  assign ys__n31882 = ~new_new_n43806__ & ~new_new_n43814__;
  assign new_new_n43816__ = ys__n47592 & new_new_n43799__;
  assign new_new_n43817__ = ys__n47205 & ~new_new_n43803__;
  assign new_new_n43818__ = ~new_new_n43816__ & ~new_new_n43817__;
  assign ys__n31883 = ~new_new_n43806__ & ~new_new_n43818__;
  assign new_new_n43820__ = ys__n47593 & new_new_n43799__;
  assign new_new_n43821__ = ys__n47206 & ~new_new_n43803__;
  assign new_new_n43822__ = ~new_new_n43820__ & ~new_new_n43821__;
  assign ys__n31884 = ~new_new_n43806__ & ~new_new_n43822__;
  assign new_new_n43824__ = ys__n47594 & new_new_n43799__;
  assign new_new_n43825__ = ys__n47207 & ~new_new_n43803__;
  assign new_new_n43826__ = ~new_new_n43824__ & ~new_new_n43825__;
  assign ys__n31885 = ~new_new_n43806__ & ~new_new_n43826__;
  assign new_new_n43828__ = ys__n47595 & new_new_n43799__;
  assign new_new_n43829__ = ys__n47208 & ~new_new_n43803__;
  assign new_new_n43830__ = ~new_new_n43828__ & ~new_new_n43829__;
  assign ys__n31886 = ~new_new_n43806__ & ~new_new_n43830__;
  assign new_new_n43832__ = ys__n47596 & new_new_n43799__;
  assign new_new_n43833__ = ys__n47209 & ~new_new_n43803__;
  assign new_new_n43834__ = ~new_new_n43832__ & ~new_new_n43833__;
  assign ys__n31887 = ~new_new_n43806__ & ~new_new_n43834__;
  assign new_new_n43836__ = ys__n47597 & new_new_n43799__;
  assign new_new_n43837__ = ys__n47210 & ~new_new_n43803__;
  assign new_new_n43838__ = ~new_new_n43836__ & ~new_new_n43837__;
  assign ys__n31888 = ~new_new_n43806__ & ~new_new_n43838__;
  assign new_new_n43840__ = ys__n47598 & new_new_n43799__;
  assign new_new_n43841__ = ys__n47211 & ~new_new_n43803__;
  assign new_new_n43842__ = ~new_new_n43840__ & ~new_new_n43841__;
  assign ys__n31889 = ~new_new_n43806__ & ~new_new_n43842__;
  assign new_new_n43844__ = ys__n47599 & new_new_n43799__;
  assign new_new_n43845__ = ys__n47212 & ~new_new_n43803__;
  assign new_new_n43846__ = ~new_new_n43844__ & ~new_new_n43845__;
  assign ys__n31890 = ~new_new_n43806__ & ~new_new_n43846__;
  assign new_new_n43848__ = ys__n47600 & new_new_n43799__;
  assign new_new_n43849__ = ys__n47213 & ~new_new_n43803__;
  assign new_new_n43850__ = ~new_new_n43848__ & ~new_new_n43849__;
  assign ys__n31891 = ~new_new_n43806__ & ~new_new_n43850__;
  assign new_new_n43852__ = ys__n47601 & new_new_n43799__;
  assign new_new_n43853__ = ys__n47214 & ~new_new_n43803__;
  assign new_new_n43854__ = ~new_new_n43852__ & ~new_new_n43853__;
  assign ys__n31892 = ~new_new_n43806__ & ~new_new_n43854__;
  assign new_new_n43856__ = ys__n47602 & new_new_n43799__;
  assign new_new_n43857__ = ys__n47215 & ~new_new_n43803__;
  assign new_new_n43858__ = ~new_new_n43856__ & ~new_new_n43857__;
  assign ys__n31893 = ~new_new_n43806__ & ~new_new_n43858__;
  assign new_new_n43860__ = ys__n47603 & new_new_n43799__;
  assign new_new_n43861__ = ys__n47216 & ~new_new_n43803__;
  assign new_new_n43862__ = ~new_new_n43860__ & ~new_new_n43861__;
  assign ys__n31894 = ~new_new_n43806__ & ~new_new_n43862__;
  assign new_new_n43864__ = ys__n47604 & new_new_n43799__;
  assign new_new_n43865__ = ys__n47217 & ~new_new_n43803__;
  assign new_new_n43866__ = ~new_new_n43864__ & ~new_new_n43865__;
  assign ys__n31895 = ~new_new_n43806__ & ~new_new_n43866__;
  assign new_new_n43868__ = ys__n47605 & new_new_n43799__;
  assign new_new_n43869__ = ys__n47218 & ~new_new_n43803__;
  assign new_new_n43870__ = ~new_new_n43868__ & ~new_new_n43869__;
  assign ys__n31896 = ~new_new_n43806__ & ~new_new_n43870__;
  assign new_new_n43872__ = ys__n47606 & new_new_n43799__;
  assign new_new_n43873__ = ys__n47219 & ~new_new_n43803__;
  assign new_new_n43874__ = ~new_new_n43872__ & ~new_new_n43873__;
  assign ys__n31897 = ~new_new_n43806__ & ~new_new_n43874__;
  assign new_new_n43876__ = ys__n47607 & new_new_n43799__;
  assign new_new_n43877__ = ys__n47220 & ~new_new_n43803__;
  assign new_new_n43878__ = ~new_new_n43876__ & ~new_new_n43877__;
  assign ys__n31898 = ~new_new_n43806__ & ~new_new_n43878__;
  assign new_new_n43880__ = ys__n47608 & new_new_n43799__;
  assign new_new_n43881__ = ys__n47221 & ~new_new_n43803__;
  assign new_new_n43882__ = ~new_new_n43880__ & ~new_new_n43881__;
  assign ys__n31899 = ~new_new_n43806__ & ~new_new_n43882__;
  assign new_new_n43884__ = ys__n47609 & new_new_n43799__;
  assign new_new_n43885__ = ys__n47222 & ~new_new_n43803__;
  assign new_new_n43886__ = ~new_new_n43884__ & ~new_new_n43885__;
  assign ys__n31900 = ~new_new_n43806__ & ~new_new_n43886__;
  assign new_new_n43888__ = ys__n47610 & new_new_n43799__;
  assign new_new_n43889__ = ys__n47223 & ~new_new_n43803__;
  assign new_new_n43890__ = ~new_new_n43888__ & ~new_new_n43889__;
  assign ys__n31901 = ~new_new_n43806__ & ~new_new_n43890__;
  assign new_new_n43892__ = ys__n47611 & new_new_n43799__;
  assign new_new_n43893__ = ys__n47224 & ~new_new_n43803__;
  assign new_new_n43894__ = ~new_new_n43892__ & ~new_new_n43893__;
  assign ys__n31902 = ~new_new_n43806__ & ~new_new_n43894__;
  assign new_new_n43896__ = ys__n47612 & new_new_n43799__;
  assign new_new_n43897__ = ys__n47225 & ~new_new_n43803__;
  assign new_new_n43898__ = ~new_new_n43896__ & ~new_new_n43897__;
  assign ys__n31903 = ~new_new_n43806__ & ~new_new_n43898__;
  assign new_new_n43900__ = ys__n47613 & new_new_n43799__;
  assign new_new_n43901__ = ys__n47226 & ~new_new_n43803__;
  assign new_new_n43902__ = ~new_new_n43900__ & ~new_new_n43901__;
  assign ys__n31904 = ~new_new_n43806__ & ~new_new_n43902__;
  assign new_new_n43904__ = ys__n47614 & new_new_n43799__;
  assign new_new_n43905__ = ys__n47227 & ~new_new_n43803__;
  assign new_new_n43906__ = ~new_new_n43904__ & ~new_new_n43905__;
  assign ys__n31905 = ~new_new_n43806__ & ~new_new_n43906__;
  assign new_new_n43908__ = ys__n47615 & new_new_n43799__;
  assign new_new_n43909__ = ys__n47228 & ~new_new_n43803__;
  assign new_new_n43910__ = ~new_new_n43908__ & ~new_new_n43909__;
  assign ys__n31906 = ~new_new_n43806__ & ~new_new_n43910__;
  assign new_new_n43912__ = ys__n47616 & new_new_n43799__;
  assign new_new_n43913__ = ys__n47229 & ~new_new_n43803__;
  assign new_new_n43914__ = ~new_new_n43912__ & ~new_new_n43913__;
  assign ys__n31907 = ~new_new_n43806__ & ~new_new_n43914__;
  assign new_new_n43916__ = ys__n47617 & new_new_n43799__;
  assign new_new_n43917__ = ys__n47230 & ~new_new_n43803__;
  assign new_new_n43918__ = ~new_new_n43916__ & ~new_new_n43917__;
  assign ys__n31908 = ~new_new_n43806__ & ~new_new_n43918__;
  assign new_new_n43920__ = ys__n47618 & new_new_n43799__;
  assign new_new_n43921__ = ys__n47231 & ~new_new_n43803__;
  assign new_new_n43922__ = ~new_new_n43920__ & ~new_new_n43921__;
  assign ys__n31909 = ~new_new_n43806__ & ~new_new_n43922__;
  assign new_new_n43924__ = ys__n47619 & new_new_n43799__;
  assign new_new_n43925__ = ys__n47232 & ~new_new_n43803__;
  assign new_new_n43926__ = ~new_new_n43924__ & ~new_new_n43925__;
  assign ys__n31910 = ~new_new_n43806__ & ~new_new_n43926__;
  assign new_new_n43928__ = ys__n47620 & new_new_n43799__;
  assign new_new_n43929__ = ys__n47233 & ~new_new_n43803__;
  assign new_new_n43930__ = ~new_new_n43928__ & ~new_new_n43929__;
  assign ys__n31911 = ~new_new_n43806__ & ~new_new_n43930__;
  assign new_new_n43932__ = ys__n47621 & new_new_n43799__;
  assign new_new_n43933__ = ys__n18762 & ~new_new_n43803__;
  assign new_new_n43934__ = ~new_new_n43932__ & ~new_new_n43933__;
  assign ys__n31912 = ~new_new_n43806__ & ~new_new_n43934__;
  assign new_new_n43936__ = ys__n47622 & new_new_n43799__;
  assign new_new_n43937__ = ys__n18750 & ~new_new_n43803__;
  assign new_new_n43938__ = ~new_new_n43936__ & ~new_new_n43937__;
  assign ys__n31913 = ~new_new_n43806__ & ~new_new_n43938__;
  assign new_new_n43940__ = ys__n47623 & new_new_n43799__;
  assign new_new_n43941__ = ys__n18753 & ~new_new_n43803__;
  assign new_new_n43942__ = ~new_new_n43940__ & ~new_new_n43941__;
  assign ys__n31914 = ~new_new_n43806__ & ~new_new_n43942__;
  assign new_new_n43944__ = ys__n850 & new_new_n12106__;
  assign new_new_n43945__ = ys__n47624 & new_new_n43944__;
  assign new_new_n43946__ = ~ys__n852 & ~new_new_n12106__;
  assign new_new_n43947__ = ~ys__n850 & new_new_n12106__;
  assign new_new_n43948__ = ~new_new_n43946__ & ~new_new_n43947__;
  assign new_new_n43949__ = ys__n47202 & ~new_new_n43948__;
  assign new_new_n43950__ = ~new_new_n43945__ & ~new_new_n43949__;
  assign new_new_n43951__ = ~new_new_n43944__ & new_new_n43948__;
  assign ys__n31915 = ~new_new_n43950__ & ~new_new_n43951__;
  assign new_new_n43953__ = ys__n47625 & new_new_n43944__;
  assign new_new_n43954__ = ys__n47203 & ~new_new_n43948__;
  assign new_new_n43955__ = ~new_new_n43953__ & ~new_new_n43954__;
  assign ys__n31916 = ~new_new_n43951__ & ~new_new_n43955__;
  assign new_new_n43957__ = ys__n47626 & new_new_n43944__;
  assign new_new_n43958__ = ys__n47204 & ~new_new_n43948__;
  assign new_new_n43959__ = ~new_new_n43957__ & ~new_new_n43958__;
  assign ys__n31917 = ~new_new_n43951__ & ~new_new_n43959__;
  assign new_new_n43961__ = ys__n47627 & new_new_n43944__;
  assign new_new_n43962__ = ys__n47205 & ~new_new_n43948__;
  assign new_new_n43963__ = ~new_new_n43961__ & ~new_new_n43962__;
  assign ys__n31918 = ~new_new_n43951__ & ~new_new_n43963__;
  assign new_new_n43965__ = ys__n47628 & new_new_n43944__;
  assign new_new_n43966__ = ys__n47206 & ~new_new_n43948__;
  assign new_new_n43967__ = ~new_new_n43965__ & ~new_new_n43966__;
  assign ys__n31919 = ~new_new_n43951__ & ~new_new_n43967__;
  assign new_new_n43969__ = ys__n47629 & new_new_n43944__;
  assign new_new_n43970__ = ys__n47207 & ~new_new_n43948__;
  assign new_new_n43971__ = ~new_new_n43969__ & ~new_new_n43970__;
  assign ys__n31920 = ~new_new_n43951__ & ~new_new_n43971__;
  assign new_new_n43973__ = ys__n47630 & new_new_n43944__;
  assign new_new_n43974__ = ys__n47208 & ~new_new_n43948__;
  assign new_new_n43975__ = ~new_new_n43973__ & ~new_new_n43974__;
  assign ys__n31921 = ~new_new_n43951__ & ~new_new_n43975__;
  assign new_new_n43977__ = ys__n47631 & new_new_n43944__;
  assign new_new_n43978__ = ys__n47209 & ~new_new_n43948__;
  assign new_new_n43979__ = ~new_new_n43977__ & ~new_new_n43978__;
  assign ys__n31922 = ~new_new_n43951__ & ~new_new_n43979__;
  assign new_new_n43981__ = ys__n47632 & new_new_n43944__;
  assign new_new_n43982__ = ys__n47210 & ~new_new_n43948__;
  assign new_new_n43983__ = ~new_new_n43981__ & ~new_new_n43982__;
  assign ys__n31923 = ~new_new_n43951__ & ~new_new_n43983__;
  assign new_new_n43985__ = ys__n47633 & new_new_n43944__;
  assign new_new_n43986__ = ys__n47211 & ~new_new_n43948__;
  assign new_new_n43987__ = ~new_new_n43985__ & ~new_new_n43986__;
  assign ys__n31924 = ~new_new_n43951__ & ~new_new_n43987__;
  assign new_new_n43989__ = ys__n47634 & new_new_n43944__;
  assign new_new_n43990__ = ys__n47212 & ~new_new_n43948__;
  assign new_new_n43991__ = ~new_new_n43989__ & ~new_new_n43990__;
  assign ys__n31925 = ~new_new_n43951__ & ~new_new_n43991__;
  assign new_new_n43993__ = ys__n47635 & new_new_n43944__;
  assign new_new_n43994__ = ys__n47213 & ~new_new_n43948__;
  assign new_new_n43995__ = ~new_new_n43993__ & ~new_new_n43994__;
  assign ys__n31926 = ~new_new_n43951__ & ~new_new_n43995__;
  assign new_new_n43997__ = ys__n47636 & new_new_n43944__;
  assign new_new_n43998__ = ys__n47214 & ~new_new_n43948__;
  assign new_new_n43999__ = ~new_new_n43997__ & ~new_new_n43998__;
  assign ys__n31927 = ~new_new_n43951__ & ~new_new_n43999__;
  assign new_new_n44001__ = ys__n47637 & new_new_n43944__;
  assign new_new_n44002__ = ys__n47215 & ~new_new_n43948__;
  assign new_new_n44003__ = ~new_new_n44001__ & ~new_new_n44002__;
  assign ys__n31928 = ~new_new_n43951__ & ~new_new_n44003__;
  assign new_new_n44005__ = ys__n47638 & new_new_n43944__;
  assign new_new_n44006__ = ys__n47216 & ~new_new_n43948__;
  assign new_new_n44007__ = ~new_new_n44005__ & ~new_new_n44006__;
  assign ys__n31929 = ~new_new_n43951__ & ~new_new_n44007__;
  assign new_new_n44009__ = ys__n47639 & new_new_n43944__;
  assign new_new_n44010__ = ys__n47217 & ~new_new_n43948__;
  assign new_new_n44011__ = ~new_new_n44009__ & ~new_new_n44010__;
  assign ys__n31930 = ~new_new_n43951__ & ~new_new_n44011__;
  assign new_new_n44013__ = ys__n47640 & new_new_n43944__;
  assign new_new_n44014__ = ys__n47218 & ~new_new_n43948__;
  assign new_new_n44015__ = ~new_new_n44013__ & ~new_new_n44014__;
  assign ys__n31931 = ~new_new_n43951__ & ~new_new_n44015__;
  assign new_new_n44017__ = ys__n47641 & new_new_n43944__;
  assign new_new_n44018__ = ys__n47219 & ~new_new_n43948__;
  assign new_new_n44019__ = ~new_new_n44017__ & ~new_new_n44018__;
  assign ys__n31932 = ~new_new_n43951__ & ~new_new_n44019__;
  assign new_new_n44021__ = ys__n47642 & new_new_n43944__;
  assign new_new_n44022__ = ys__n47220 & ~new_new_n43948__;
  assign new_new_n44023__ = ~new_new_n44021__ & ~new_new_n44022__;
  assign ys__n31933 = ~new_new_n43951__ & ~new_new_n44023__;
  assign new_new_n44025__ = ys__n47643 & new_new_n43944__;
  assign new_new_n44026__ = ys__n47221 & ~new_new_n43948__;
  assign new_new_n44027__ = ~new_new_n44025__ & ~new_new_n44026__;
  assign ys__n31934 = ~new_new_n43951__ & ~new_new_n44027__;
  assign new_new_n44029__ = ys__n47644 & new_new_n43944__;
  assign new_new_n44030__ = ys__n47222 & ~new_new_n43948__;
  assign new_new_n44031__ = ~new_new_n44029__ & ~new_new_n44030__;
  assign ys__n31935 = ~new_new_n43951__ & ~new_new_n44031__;
  assign new_new_n44033__ = ys__n47645 & new_new_n43944__;
  assign new_new_n44034__ = ys__n47223 & ~new_new_n43948__;
  assign new_new_n44035__ = ~new_new_n44033__ & ~new_new_n44034__;
  assign ys__n31936 = ~new_new_n43951__ & ~new_new_n44035__;
  assign new_new_n44037__ = ys__n47646 & new_new_n43944__;
  assign new_new_n44038__ = ys__n47224 & ~new_new_n43948__;
  assign new_new_n44039__ = ~new_new_n44037__ & ~new_new_n44038__;
  assign ys__n31937 = ~new_new_n43951__ & ~new_new_n44039__;
  assign new_new_n44041__ = ys__n47647 & new_new_n43944__;
  assign new_new_n44042__ = ys__n47225 & ~new_new_n43948__;
  assign new_new_n44043__ = ~new_new_n44041__ & ~new_new_n44042__;
  assign ys__n31938 = ~new_new_n43951__ & ~new_new_n44043__;
  assign new_new_n44045__ = ys__n47648 & new_new_n43944__;
  assign new_new_n44046__ = ys__n47226 & ~new_new_n43948__;
  assign new_new_n44047__ = ~new_new_n44045__ & ~new_new_n44046__;
  assign ys__n31939 = ~new_new_n43951__ & ~new_new_n44047__;
  assign new_new_n44049__ = ys__n47649 & new_new_n43944__;
  assign new_new_n44050__ = ys__n47227 & ~new_new_n43948__;
  assign new_new_n44051__ = ~new_new_n44049__ & ~new_new_n44050__;
  assign ys__n31940 = ~new_new_n43951__ & ~new_new_n44051__;
  assign new_new_n44053__ = ys__n47650 & new_new_n43944__;
  assign new_new_n44054__ = ys__n47228 & ~new_new_n43948__;
  assign new_new_n44055__ = ~new_new_n44053__ & ~new_new_n44054__;
  assign ys__n31941 = ~new_new_n43951__ & ~new_new_n44055__;
  assign new_new_n44057__ = ys__n47651 & new_new_n43944__;
  assign new_new_n44058__ = ys__n47229 & ~new_new_n43948__;
  assign new_new_n44059__ = ~new_new_n44057__ & ~new_new_n44058__;
  assign ys__n31942 = ~new_new_n43951__ & ~new_new_n44059__;
  assign new_new_n44061__ = ys__n47652 & new_new_n43944__;
  assign new_new_n44062__ = ys__n47230 & ~new_new_n43948__;
  assign new_new_n44063__ = ~new_new_n44061__ & ~new_new_n44062__;
  assign ys__n31943 = ~new_new_n43951__ & ~new_new_n44063__;
  assign new_new_n44065__ = ys__n47653 & new_new_n43944__;
  assign new_new_n44066__ = ys__n47231 & ~new_new_n43948__;
  assign new_new_n44067__ = ~new_new_n44065__ & ~new_new_n44066__;
  assign ys__n31944 = ~new_new_n43951__ & ~new_new_n44067__;
  assign new_new_n44069__ = ys__n47654 & new_new_n43944__;
  assign new_new_n44070__ = ys__n47232 & ~new_new_n43948__;
  assign new_new_n44071__ = ~new_new_n44069__ & ~new_new_n44070__;
  assign ys__n31945 = ~new_new_n43951__ & ~new_new_n44071__;
  assign new_new_n44073__ = ys__n47655 & new_new_n43944__;
  assign new_new_n44074__ = ys__n47233 & ~new_new_n43948__;
  assign new_new_n44075__ = ~new_new_n44073__ & ~new_new_n44074__;
  assign ys__n31946 = ~new_new_n43951__ & ~new_new_n44075__;
  assign new_new_n44077__ = ys__n47656 & new_new_n43944__;
  assign new_new_n44078__ = ys__n18762 & ~new_new_n43948__;
  assign new_new_n44079__ = ~new_new_n44077__ & ~new_new_n44078__;
  assign ys__n31947 = ~new_new_n43951__ & ~new_new_n44079__;
  assign new_new_n44081__ = ys__n47657 & new_new_n43944__;
  assign new_new_n44082__ = ys__n18750 & ~new_new_n43948__;
  assign new_new_n44083__ = ~new_new_n44081__ & ~new_new_n44082__;
  assign ys__n31948 = ~new_new_n43951__ & ~new_new_n44083__;
  assign new_new_n44085__ = ys__n47658 & new_new_n43944__;
  assign new_new_n44086__ = ys__n18753 & ~new_new_n43948__;
  assign new_new_n44087__ = ~new_new_n44085__ & ~new_new_n44086__;
  assign ys__n31949 = ~new_new_n43951__ & ~new_new_n44087__;
  assign new_new_n44089__ = ~ys__n556 & ys__n558;
  assign new_new_n44090__ = ~ys__n935 & ~ys__n1802;
  assign new_new_n44091__ = new_new_n44089__ & new_new_n44090__;
  assign new_new_n44092__ = ys__n556 & ~ys__n935;
  assign new_new_n44093__ = ~ys__n1802 & new_new_n44092__;
  assign new_new_n44094__ = ~new_new_n44091__ & ~new_new_n44093__;
  assign new_new_n44095__ = ~ys__n556 & ~ys__n558;
  assign new_new_n44096__ = ys__n935 & ~ys__n1802;
  assign new_new_n44097__ = new_new_n44095__ & new_new_n44096__;
  assign new_new_n44098__ = ys__n556 & ys__n935;
  assign new_new_n44099__ = ~ys__n1802 & new_new_n44098__;
  assign new_new_n44100__ = ~ys__n1802 & ~new_new_n44099__;
  assign new_new_n44101__ = ~new_new_n44097__ & new_new_n44100__;
  assign new_new_n44102__ = new_new_n44089__ & new_new_n44096__;
  assign new_new_n44103__ = new_new_n44090__ & new_new_n44095__;
  assign new_new_n44104__ = ~new_new_n44102__ & ~new_new_n44103__;
  assign new_new_n44105__ = new_new_n44101__ & new_new_n44104__;
  assign new_new_n44106__ = new_new_n44094__ & new_new_n44105__;
  assign new_new_n44107__ = new_new_n12583__ & ~new_new_n44094__;
  assign new_new_n44108__ = ~new_new_n44106__ & new_new_n44107__;
  assign new_new_n44109__ = ys__n556 & ~ys__n1802;
  assign new_new_n44110__ = ys__n178 & new_new_n10990__;
  assign new_new_n44111__ = ~ys__n176 & ~ys__n558;
  assign new_new_n44112__ = new_new_n44110__ & new_new_n44111__;
  assign new_new_n44113__ = new_new_n44109__ & new_new_n44112__;
  assign new_new_n44114__ = ys__n178 & ~new_new_n10990__;
  assign new_new_n44115__ = new_new_n44111__ & new_new_n44114__;
  assign new_new_n44116__ = new_new_n44109__ & new_new_n44115__;
  assign new_new_n44117__ = ~new_new_n44113__ & ~new_new_n44116__;
  assign new_new_n44118__ = ~ys__n176 & ys__n558;
  assign new_new_n44119__ = new_new_n44110__ & new_new_n44118__;
  assign new_new_n44120__ = new_new_n44109__ & new_new_n44119__;
  assign new_new_n44121__ = new_new_n44114__ & new_new_n44118__;
  assign new_new_n44122__ = new_new_n44109__ & new_new_n44121__;
  assign new_new_n44123__ = ~new_new_n44120__ & ~new_new_n44122__;
  assign new_new_n44124__ = new_new_n44117__ & new_new_n44123__;
  assign new_new_n44125__ = new_new_n10993__ & new_new_n44089__;
  assign new_new_n44126__ = ~ys__n1802 & new_new_n44125__;
  assign new_new_n44127__ = ys__n556 & ~ys__n558;
  assign new_new_n44128__ = new_new_n10993__ & new_new_n44127__;
  assign new_new_n44129__ = ~ys__n1802 & new_new_n44128__;
  assign new_new_n44130__ = ~new_new_n44126__ & ~new_new_n44129__;
  assign new_new_n44131__ = ys__n556 & ys__n558;
  assign new_new_n44132__ = new_new_n11001__ & new_new_n44131__;
  assign new_new_n44133__ = ~ys__n1802 & new_new_n44132__;
  assign new_new_n44134__ = new_new_n11000__ & new_new_n44131__;
  assign new_new_n44135__ = ~ys__n1802 & new_new_n44134__;
  assign new_new_n44136__ = new_new_n10993__ & new_new_n44131__;
  assign new_new_n44137__ = ~ys__n1802 & new_new_n44136__;
  assign new_new_n44138__ = ~new_new_n44135__ & ~new_new_n44137__;
  assign new_new_n44139__ = ~new_new_n44133__ & new_new_n44138__;
  assign new_new_n44140__ = new_new_n44130__ & new_new_n44139__;
  assign new_new_n44141__ = ~ys__n556 & ~ys__n1802;
  assign new_new_n44142__ = new_new_n44119__ & new_new_n44141__;
  assign new_new_n44143__ = new_new_n44121__ & new_new_n44141__;
  assign new_new_n44144__ = ~new_new_n44142__ & ~new_new_n44143__;
  assign new_new_n44145__ = new_new_n44140__ & new_new_n44144__;
  assign new_new_n44146__ = new_new_n44124__ & new_new_n44145__;
  assign new_new_n44147__ = new_new_n11000__ & new_new_n44089__;
  assign new_new_n44148__ = ~ys__n1802 & new_new_n44147__;
  assign new_new_n44149__ = new_new_n11001__ & new_new_n44089__;
  assign new_new_n44150__ = ~ys__n1802 & new_new_n44149__;
  assign new_new_n44151__ = ~new_new_n44148__ & ~new_new_n44150__;
  assign new_new_n44152__ = new_new_n11000__ & new_new_n44127__;
  assign new_new_n44153__ = ~ys__n1802 & new_new_n44152__;
  assign new_new_n44154__ = new_new_n11001__ & new_new_n44127__;
  assign new_new_n44155__ = ~ys__n1802 & new_new_n44154__;
  assign new_new_n44156__ = ~new_new_n44153__ & ~new_new_n44155__;
  assign new_new_n44157__ = new_new_n44151__ & new_new_n44156__;
  assign new_new_n44158__ = new_new_n11000__ & new_new_n44095__;
  assign new_new_n44159__ = ~ys__n1802 & new_new_n44158__;
  assign new_new_n44160__ = ~ys__n1802 & ~new_new_n44159__;
  assign new_new_n44161__ = new_new_n10993__ & new_new_n44095__;
  assign new_new_n44162__ = ~ys__n1802 & new_new_n44161__;
  assign new_new_n44163__ = new_new_n11001__ & new_new_n44095__;
  assign new_new_n44164__ = ~ys__n1802 & new_new_n44163__;
  assign new_new_n44165__ = ~new_new_n44162__ & ~new_new_n44164__;
  assign new_new_n44166__ = new_new_n44160__ & new_new_n44165__;
  assign new_new_n44167__ = new_new_n44157__ & new_new_n44166__;
  assign new_new_n44168__ = new_new_n44112__ & new_new_n44141__;
  assign new_new_n44169__ = new_new_n44115__ & new_new_n44141__;
  assign new_new_n44170__ = ~new_new_n44168__ & ~new_new_n44169__;
  assign new_new_n44171__ = new_new_n44167__ & new_new_n44170__;
  assign new_new_n44172__ = new_new_n44146__ & new_new_n44171__;
  assign new_new_n44173__ = new_new_n11006__ & ~new_new_n44146__;
  assign new_new_n44174__ = ~new_new_n44172__ & new_new_n44173__;
  assign new_new_n44175__ = ~new_new_n44108__ & ~new_new_n44174__;
  assign new_new_n44176__ = ~ys__n738 & ~new_new_n11006__;
  assign new_new_n44177__ = ~new_new_n12583__ & new_new_n44176__;
  assign ys__n31950 = ~new_new_n44175__ & ~new_new_n44177__;
  assign new_new_n44179__ = ~new_new_n44137__ & ~new_new_n44162__;
  assign new_new_n44180__ = new_new_n44130__ & new_new_n44179__;
  assign new_new_n44181__ = ~new_new_n44142__ & new_new_n44180__;
  assign new_new_n44182__ = ~new_new_n44113__ & ~new_new_n44120__;
  assign new_new_n44183__ = ~new_new_n44168__ & new_new_n44182__;
  assign new_new_n44184__ = new_new_n44181__ & new_new_n44183__;
  assign new_new_n44185__ = ~new_new_n44133__ & ~new_new_n44150__;
  assign new_new_n44186__ = ~new_new_n44155__ & new_new_n44185__;
  assign new_new_n44187__ = new_new_n44184__ & new_new_n44186__;
  assign new_new_n44188__ = ~new_new_n44116__ & ~new_new_n44143__;
  assign new_new_n44189__ = ~new_new_n44122__ & ~new_new_n44169__;
  assign new_new_n44190__ = new_new_n44188__ & new_new_n44189__;
  assign new_new_n44191__ = ~new_new_n44135__ & ~new_new_n44148__;
  assign new_new_n44192__ = ~new_new_n44153__ & new_new_n44191__;
  assign new_new_n44193__ = new_new_n44190__ & new_new_n44192__;
  assign new_new_n44194__ = ~new_new_n44159__ & ~new_new_n44164__;
  assign new_new_n44195__ = ~ys__n1802 & new_new_n44194__;
  assign new_new_n44196__ = new_new_n44193__ & new_new_n44195__;
  assign new_new_n44197__ = new_new_n44187__ & new_new_n44196__;
  assign new_new_n44198__ = new_new_n44193__ & new_new_n44194__;
  assign new_new_n44199__ = new_new_n11006__ & ~new_new_n44198__;
  assign new_new_n44200__ = ~new_new_n44197__ & new_new_n44199__;
  assign new_new_n44201__ = ~new_new_n44109__ & ~new_new_n44141__;
  assign new_new_n44202__ = ~ys__n1802 & new_new_n44201__;
  assign new_new_n44203__ = ys__n738 & new_new_n44141__;
  assign new_new_n44204__ = ~new_new_n44202__ & new_new_n44203__;
  assign new_new_n44205__ = new_new_n44094__ & ~new_new_n44103__;
  assign new_new_n44206__ = ~new_new_n44099__ & ~new_new_n44102__;
  assign new_new_n44207__ = ~ys__n1802 & ~new_new_n44097__;
  assign new_new_n44208__ = new_new_n44206__ & new_new_n44207__;
  assign new_new_n44209__ = new_new_n44205__ & new_new_n44208__;
  assign new_new_n44210__ = new_new_n12583__ & new_new_n44097__;
  assign new_new_n44211__ = ~new_new_n44209__ & new_new_n44210__;
  assign new_new_n44212__ = ~new_new_n44204__ & ~new_new_n44211__;
  assign new_new_n44213__ = ~new_new_n44200__ & new_new_n44212__;
  assign ys__n31953 = ~new_new_n44177__ & ~new_new_n44213__;
  assign new_new_n44215__ = new_new_n44187__ & new_new_n44194__;
  assign new_new_n44216__ = new_new_n11006__ & ~new_new_n44197__;
  assign new_new_n44217__ = ~new_new_n44215__ & new_new_n44216__;
  assign new_new_n44218__ = ys__n738 & ~new_new_n44201__;
  assign new_new_n44219__ = ~new_new_n44202__ & new_new_n44218__;
  assign new_new_n44220__ = ~new_new_n44097__ & new_new_n44206__;
  assign new_new_n44221__ = new_new_n12583__ & ~new_new_n44220__;
  assign new_new_n44222__ = ~new_new_n44209__ & new_new_n44221__;
  assign new_new_n44223__ = ~new_new_n44219__ & ~new_new_n44222__;
  assign new_new_n44224__ = ~new_new_n44217__ & new_new_n44223__;
  assign ys__n31954 = ~new_new_n44177__ & ~new_new_n44224__;
  assign new_new_n44226__ = ~new_new_n44164__ & new_new_n44190__;
  assign new_new_n44227__ = new_new_n44184__ & new_new_n44226__;
  assign new_new_n44228__ = new_new_n11006__ & ~new_new_n44227__;
  assign new_new_n44229__ = ~new_new_n44197__ & new_new_n44228__;
  assign new_new_n44230__ = ~new_new_n44097__ & new_new_n44205__;
  assign new_new_n44231__ = new_new_n12583__ & ~new_new_n44209__;
  assign new_new_n44232__ = ~new_new_n44230__ & new_new_n44231__;
  assign new_new_n44233__ = ~new_new_n44204__ & ~new_new_n44232__;
  assign new_new_n44234__ = ~new_new_n44229__ & new_new_n44233__;
  assign ys__n31955 = ~new_new_n44177__ & ~new_new_n44234__;
  assign new_new_n44236__ = ys__n29846 & new_new_n10601__;
  assign new_new_n44237__ = ~new_new_n10601__ & ys__n29847;
  assign new_new_n44238__ = ~new_new_n44236__ & ~new_new_n44237__;
  assign new_new_n44239__ = ~ys__n23764 & ~new_new_n44238__;
  assign new_new_n44240__ = ys__n29898 & ~new_new_n10603__;
  assign new_new_n44241__ = ~new_new_n10601__ & new_new_n44240__;
  assign new_new_n44242__ = ~ys__n22466 & new_new_n44241__;
  assign new_new_n44243__ = ys__n22466 & ~new_new_n44238__;
  assign new_new_n44244__ = ~new_new_n44242__ & ~new_new_n44243__;
  assign new_new_n44245__ = ys__n23764 & ~new_new_n44244__;
  assign new_new_n44246__ = ~new_new_n44239__ & ~new_new_n44245__;
  assign ys__n31965 = new_new_n10866__ & ~new_new_n44246__;
  assign new_new_n44248__ = ys__n29887 & ~new_new_n10603__;
  assign new_new_n44249__ = ~new_new_n10601__ & new_new_n44248__;
  assign new_new_n44250__ = ~ys__n23764 & new_new_n44249__;
  assign new_new_n44251__ = ys__n29903 & ~new_new_n10603__;
  assign new_new_n44252__ = ~new_new_n10601__ & new_new_n44251__;
  assign new_new_n44253__ = ~ys__n22466 & new_new_n44252__;
  assign new_new_n44254__ = ys__n22466 & new_new_n44249__;
  assign new_new_n44255__ = ~new_new_n44253__ & ~new_new_n44254__;
  assign new_new_n44256__ = ys__n23764 & ~new_new_n44255__;
  assign new_new_n44257__ = ~new_new_n44250__ & ~new_new_n44256__;
  assign ys__n31971 = new_new_n10866__ & ~new_new_n44257__;
  assign new_new_n44259__ = ys__n29888 & ~new_new_n10603__;
  assign new_new_n44260__ = ~new_new_n10601__ & new_new_n44259__;
  assign new_new_n44261__ = ~ys__n23764 & new_new_n44260__;
  assign new_new_n44262__ = ys__n29904 & ~new_new_n10603__;
  assign new_new_n44263__ = ~new_new_n10601__ & new_new_n44262__;
  assign new_new_n44264__ = ~ys__n22466 & new_new_n44263__;
  assign new_new_n44265__ = ys__n22466 & new_new_n44260__;
  assign new_new_n44266__ = ~new_new_n44264__ & ~new_new_n44265__;
  assign new_new_n44267__ = ys__n23764 & ~new_new_n44266__;
  assign new_new_n44268__ = ~new_new_n44261__ & ~new_new_n44267__;
  assign ys__n31973 = new_new_n10866__ & ~new_new_n44268__;
  assign new_new_n44270__ = ys__n29889 & ~new_new_n10603__;
  assign new_new_n44271__ = ~new_new_n10601__ & new_new_n44270__;
  assign new_new_n44272__ = ~ys__n23764 & new_new_n44271__;
  assign new_new_n44273__ = ys__n29905 & ~new_new_n10603__;
  assign new_new_n44274__ = ~new_new_n10601__ & new_new_n44273__;
  assign new_new_n44275__ = ~ys__n22466 & new_new_n44274__;
  assign new_new_n44276__ = ys__n22466 & new_new_n44271__;
  assign new_new_n44277__ = ~new_new_n44275__ & ~new_new_n44276__;
  assign new_new_n44278__ = ys__n23764 & ~new_new_n44277__;
  assign new_new_n44279__ = ~new_new_n44272__ & ~new_new_n44278__;
  assign ys__n31975 = new_new_n10866__ & ~new_new_n44279__;
  assign new_new_n44281__ = ys__n29890 & ~new_new_n10603__;
  assign new_new_n44282__ = ~new_new_n10601__ & new_new_n44281__;
  assign new_new_n44283__ = ~ys__n23764 & new_new_n44282__;
  assign new_new_n44284__ = ys__n29906 & ~new_new_n10603__;
  assign new_new_n44285__ = ~new_new_n10601__ & new_new_n44284__;
  assign new_new_n44286__ = ~ys__n22466 & new_new_n44285__;
  assign new_new_n44287__ = ys__n22466 & new_new_n44282__;
  assign new_new_n44288__ = ~new_new_n44286__ & ~new_new_n44287__;
  assign new_new_n44289__ = ys__n23764 & ~new_new_n44288__;
  assign new_new_n44290__ = ~new_new_n44283__ & ~new_new_n44289__;
  assign new_new_n44291__ = ~new_new_n10859__ & ~new_new_n44290__;
  assign new_new_n44292__ = ~new_new_n12064__ & ~new_new_n44291__;
  assign ys__n31976 = ~new_new_n10865__ & ~new_new_n44292__;
  assign new_new_n44294__ = ys__n29891 & ~new_new_n10603__;
  assign new_new_n44295__ = ~new_new_n10601__ & new_new_n44294__;
  assign new_new_n44296__ = ~ys__n23764 & new_new_n44295__;
  assign new_new_n44297__ = ys__n29907 & ~new_new_n10603__;
  assign new_new_n44298__ = ~new_new_n10601__ & new_new_n44297__;
  assign new_new_n44299__ = ~ys__n22466 & new_new_n44298__;
  assign new_new_n44300__ = ys__n22466 & new_new_n44295__;
  assign new_new_n44301__ = ~new_new_n44299__ & ~new_new_n44300__;
  assign new_new_n44302__ = ys__n23764 & ~new_new_n44301__;
  assign new_new_n44303__ = ~new_new_n44296__ & ~new_new_n44302__;
  assign ys__n31978 = new_new_n10866__ & ~new_new_n44303__;
  assign new_new_n44305__ = ys__n29892 & ~new_new_n10603__;
  assign new_new_n44306__ = ~new_new_n10601__ & new_new_n44305__;
  assign new_new_n44307__ = ~ys__n23764 & new_new_n44306__;
  assign new_new_n44308__ = ys__n29908 & ~new_new_n10603__;
  assign new_new_n44309__ = ~new_new_n10601__ & new_new_n44308__;
  assign new_new_n44310__ = ~ys__n22466 & new_new_n44309__;
  assign new_new_n44311__ = ys__n22466 & new_new_n44306__;
  assign new_new_n44312__ = ~new_new_n44310__ & ~new_new_n44311__;
  assign new_new_n44313__ = ys__n23764 & ~new_new_n44312__;
  assign new_new_n44314__ = ~new_new_n44307__ & ~new_new_n44313__;
  assign new_new_n44315__ = ~new_new_n10859__ & ~new_new_n44314__;
  assign new_new_n44316__ = ~new_new_n12064__ & ~new_new_n44315__;
  assign ys__n31979 = ~new_new_n10865__ & ~new_new_n44316__;
  assign new_new_n44318__ = ~ys__n23764 & ~new_new_n10859__;
  assign new_new_n44319__ = ~new_new_n10865__ & new_new_n44318__;
  assign ys__n31984 = new_new_n44241__ & new_new_n44319__;
  assign ys__n31986 = new_new_n26170__ & new_new_n44319__;
  assign ys__n31988 = new_new_n26181__ & new_new_n44319__;
  assign ys__n31990 = new_new_n26192__ & new_new_n44319__;
  assign ys__n31992 = new_new_n16892__ & new_new_n44319__;
  assign ys__n31994 = new_new_n44252__ & new_new_n44319__;
  assign ys__n31996 = new_new_n44263__ & new_new_n44319__;
  assign ys__n31998 = new_new_n44274__ & new_new_n44319__;
  assign ys__n32000 = new_new_n44285__ & new_new_n44319__;
  assign ys__n32002 = new_new_n44298__ & new_new_n44319__;
  assign new_new_n44330__ = ~ys__n23764 & new_new_n44309__;
  assign new_new_n44331__ = ~new_new_n16911__ & ~new_new_n44330__;
  assign ys__n32004 = new_new_n10866__ & ~new_new_n44331__;
  assign new_new_n44333__ = ~ys__n23764 & new_new_n16907__;
  assign new_new_n44334__ = ~new_new_n12137__ & ~new_new_n44333__;
  assign ys__n32006 = new_new_n10866__ & ~new_new_n44334__;
  assign new_new_n44336__ = ~ys__n23764 & new_new_n12133__;
  assign new_new_n44337__ = ~new_new_n12119__ & ~new_new_n44336__;
  assign new_new_n44338__ = ~new_new_n10859__ & ~new_new_n44337__;
  assign new_new_n44339__ = ~new_new_n12064__ & ~new_new_n44338__;
  assign ys__n32007 = ~new_new_n10865__ & ~new_new_n44339__;
  assign new_new_n44341__ = ~ys__n23764 & new_new_n12115__;
  assign new_new_n44342__ = ~new_new_n12061__ & ~new_new_n44341__;
  assign new_new_n44343__ = ~new_new_n10859__ & ~new_new_n44342__;
  assign new_new_n44344__ = ~new_new_n12064__ & ~new_new_n44343__;
  assign ys__n32008 = ~new_new_n10865__ & ~new_new_n44344__;
  assign ys__n32010 = new_new_n12057__ & new_new_n44319__;
  assign new_new_n44347__ = ~ys__n23764 & new_new_n10620__;
  assign new_new_n44348__ = ~new_new_n10627__ & ~new_new_n44347__;
  assign ys__n32012 = new_new_n10866__ & ~new_new_n44348__;
  assign new_new_n44350__ = new_new_n11323__ & new_new_n21497__;
  assign ys__n32014 = ~new_new_n21499__ & new_new_n44350__;
  assign new_new_n44352__ = new_new_n11343__ & new_new_n21497__;
  assign ys__n32016 = ~new_new_n21499__ & new_new_n44352__;
  assign new_new_n44354__ = new_new_n11319__ & new_new_n21497__;
  assign ys__n32018 = ~new_new_n21499__ & new_new_n44354__;
  assign new_new_n44356__ = ~ys__n23661 & ys__n23663;
  assign new_new_n44357__ = ~ys__n28459 & new_new_n44356__;
  assign new_new_n44358__ = ys__n23661 & ~ys__n28457;
  assign new_new_n44359__ = ~new_new_n44357__ & ~new_new_n44358__;
  assign new_new_n44360__ = ~ys__n23658 & ~new_new_n44359__;
  assign new_new_n44361__ = ys__n23658 & ~ys__n28455;
  assign new_new_n44362__ = ~new_new_n44360__ & ~new_new_n44361__;
  assign new_new_n44363__ = ~ys__n23655 & ~new_new_n44362__;
  assign new_new_n44364__ = ys__n23655 & ~ys__n28453;
  assign new_new_n44365__ = ys__n38315 & new_new_n44364__;
  assign new_new_n44366__ = ~new_new_n44363__ & ~new_new_n44365__;
  assign new_new_n44367__ = ~ys__n352 & ~ys__n19973;
  assign new_new_n44368__ = ys__n38424 & new_new_n44367__;
  assign new_new_n44369__ = new_new_n44366__ & ~new_new_n44368__;
  assign new_new_n44370__ = ys__n544 & ~ys__n546;
  assign new_new_n44371__ = new_new_n44369__ & new_new_n44370__;
  assign new_new_n44372__ = ~ys__n544 & ~ys__n546;
  assign new_new_n44373__ = ~new_new_n44368__ & new_new_n44372__;
  assign new_new_n44374__ = ~new_new_n44366__ & new_new_n44373__;
  assign new_new_n44375__ = ~new_new_n44371__ & ~new_new_n44374__;
  assign new_new_n44376__ = new_new_n44368__ & new_new_n44372__;
  assign new_new_n44377__ = new_new_n44366__ & new_new_n44376__;
  assign new_new_n44378__ = ~new_new_n44374__ & ~new_new_n44377__;
  assign new_new_n44379__ = ~ys__n544 & ys__n546;
  assign new_new_n44380__ = new_new_n44369__ & new_new_n44379__;
  assign new_new_n44381__ = ~new_new_n44371__ & ~new_new_n44380__;
  assign ys__n32024 = ~new_new_n44378__ | ~new_new_n44381__;
  assign ys__n32022 = ~new_new_n44375__ & ys__n32024;
  assign ys__n32023 = ~new_new_n44378__ & ys__n32024;
  assign new_new_n44385__ = ys__n47692 & ~new_new_n12625__;
  assign new_new_n44386__ = ys__n47723 & new_new_n12626__;
  assign new_new_n44387__ = ~new_new_n44385__ & ~new_new_n44386__;
  assign ys__n32025 = ~new_new_n12627__ & ~new_new_n44387__;
  assign new_new_n44389__ = ys__n47693 & ~new_new_n12625__;
  assign new_new_n44390__ = ys__n47724 & new_new_n12626__;
  assign new_new_n44391__ = ~new_new_n44389__ & ~new_new_n44390__;
  assign ys__n32026 = ~new_new_n12627__ & ~new_new_n44391__;
  assign new_new_n44393__ = ys__n47694 & ~new_new_n12625__;
  assign new_new_n44394__ = ys__n47725 & new_new_n12626__;
  assign new_new_n44395__ = ~new_new_n44393__ & ~new_new_n44394__;
  assign ys__n32027 = ~new_new_n12627__ & ~new_new_n44395__;
  assign new_new_n44397__ = ys__n47695 & ~new_new_n12625__;
  assign new_new_n44398__ = ys__n47726 & new_new_n12626__;
  assign new_new_n44399__ = ~new_new_n44397__ & ~new_new_n44398__;
  assign ys__n32028 = ~new_new_n12627__ & ~new_new_n44399__;
  assign new_new_n44401__ = ys__n47696 & ~new_new_n12625__;
  assign new_new_n44402__ = ys__n47727 & new_new_n12626__;
  assign new_new_n44403__ = ~new_new_n44401__ & ~new_new_n44402__;
  assign ys__n32029 = ~new_new_n12627__ & ~new_new_n44403__;
  assign new_new_n44405__ = ys__n47697 & ~new_new_n12625__;
  assign new_new_n44406__ = ys__n47728 & new_new_n12626__;
  assign new_new_n44407__ = ~new_new_n44405__ & ~new_new_n44406__;
  assign ys__n32030 = ~new_new_n12627__ & ~new_new_n44407__;
  assign new_new_n44409__ = ys__n47698 & ~new_new_n12625__;
  assign new_new_n44410__ = ys__n47729 & new_new_n12626__;
  assign new_new_n44411__ = ~new_new_n44409__ & ~new_new_n44410__;
  assign ys__n32031 = ~new_new_n12627__ & ~new_new_n44411__;
  assign new_new_n44413__ = ys__n47699 & ~new_new_n12625__;
  assign new_new_n44414__ = ys__n47730 & new_new_n12626__;
  assign new_new_n44415__ = ~new_new_n44413__ & ~new_new_n44414__;
  assign ys__n32032 = ~new_new_n12627__ & ~new_new_n44415__;
  assign new_new_n44417__ = ys__n47700 & ~new_new_n12625__;
  assign new_new_n44418__ = ys__n47731 & new_new_n12626__;
  assign new_new_n44419__ = ~new_new_n44417__ & ~new_new_n44418__;
  assign ys__n32033 = ~new_new_n12627__ & ~new_new_n44419__;
  assign new_new_n44421__ = ys__n47701 & ~new_new_n12625__;
  assign new_new_n44422__ = ys__n47732 & new_new_n12626__;
  assign new_new_n44423__ = ~new_new_n44421__ & ~new_new_n44422__;
  assign ys__n32034 = ~new_new_n12627__ & ~new_new_n44423__;
  assign new_new_n44425__ = ys__n47702 & ~new_new_n12625__;
  assign new_new_n44426__ = ys__n47733 & new_new_n12626__;
  assign new_new_n44427__ = ~new_new_n44425__ & ~new_new_n44426__;
  assign ys__n32035 = ~new_new_n12627__ & ~new_new_n44427__;
  assign new_new_n44429__ = ys__n47703 & ~new_new_n12625__;
  assign new_new_n44430__ = ys__n47734 & new_new_n12626__;
  assign new_new_n44431__ = ~new_new_n44429__ & ~new_new_n44430__;
  assign ys__n32036 = ~new_new_n12627__ & ~new_new_n44431__;
  assign new_new_n44433__ = ys__n47704 & ~new_new_n12625__;
  assign new_new_n44434__ = ys__n47735 & new_new_n12626__;
  assign new_new_n44435__ = ~new_new_n44433__ & ~new_new_n44434__;
  assign ys__n32037 = ~new_new_n12627__ & ~new_new_n44435__;
  assign new_new_n44437__ = ys__n47705 & ~new_new_n12625__;
  assign new_new_n44438__ = ys__n47736 & new_new_n12626__;
  assign new_new_n44439__ = ~new_new_n44437__ & ~new_new_n44438__;
  assign ys__n32038 = ~new_new_n12627__ & ~new_new_n44439__;
  assign new_new_n44441__ = ys__n47706 & ~new_new_n12625__;
  assign new_new_n44442__ = ys__n47737 & new_new_n12626__;
  assign new_new_n44443__ = ~new_new_n44441__ & ~new_new_n44442__;
  assign ys__n32039 = ~new_new_n12627__ & ~new_new_n44443__;
  assign new_new_n44445__ = ys__n47707 & ~new_new_n12625__;
  assign new_new_n44446__ = ys__n47738 & new_new_n12626__;
  assign new_new_n44447__ = ~new_new_n44445__ & ~new_new_n44446__;
  assign ys__n32040 = ~new_new_n12627__ & ~new_new_n44447__;
  assign new_new_n44449__ = ys__n47708 & ~new_new_n12625__;
  assign new_new_n44450__ = ys__n47739 & new_new_n12626__;
  assign new_new_n44451__ = ~new_new_n44449__ & ~new_new_n44450__;
  assign ys__n32041 = ~new_new_n12627__ & ~new_new_n44451__;
  assign new_new_n44453__ = ys__n47709 & ~new_new_n12625__;
  assign new_new_n44454__ = ys__n47740 & new_new_n12626__;
  assign new_new_n44455__ = ~new_new_n44453__ & ~new_new_n44454__;
  assign ys__n32042 = ~new_new_n12627__ & ~new_new_n44455__;
  assign new_new_n44457__ = ys__n47710 & ~new_new_n12625__;
  assign new_new_n44458__ = ys__n47741 & new_new_n12626__;
  assign new_new_n44459__ = ~new_new_n44457__ & ~new_new_n44458__;
  assign ys__n32043 = ~new_new_n12627__ & ~new_new_n44459__;
  assign new_new_n44461__ = ys__n47711 & ~new_new_n12625__;
  assign new_new_n44462__ = ys__n47742 & new_new_n12626__;
  assign new_new_n44463__ = ~new_new_n44461__ & ~new_new_n44462__;
  assign ys__n32044 = ~new_new_n12627__ & ~new_new_n44463__;
  assign new_new_n44465__ = ys__n47712 & ~new_new_n12625__;
  assign new_new_n44466__ = ys__n47743 & new_new_n12626__;
  assign new_new_n44467__ = ~new_new_n44465__ & ~new_new_n44466__;
  assign ys__n32045 = ~new_new_n12627__ & ~new_new_n44467__;
  assign new_new_n44469__ = ys__n47713 & ~new_new_n12625__;
  assign new_new_n44470__ = ys__n47744 & new_new_n12626__;
  assign new_new_n44471__ = ~new_new_n44469__ & ~new_new_n44470__;
  assign ys__n32046 = ~new_new_n12627__ & ~new_new_n44471__;
  assign new_new_n44473__ = ys__n47714 & ~new_new_n12625__;
  assign new_new_n44474__ = ys__n47745 & new_new_n12626__;
  assign new_new_n44475__ = ~new_new_n44473__ & ~new_new_n44474__;
  assign ys__n32047 = ~new_new_n12627__ & ~new_new_n44475__;
  assign new_new_n44477__ = ys__n47715 & ~new_new_n12625__;
  assign new_new_n44478__ = ys__n47746 & new_new_n12626__;
  assign new_new_n44479__ = ~new_new_n44477__ & ~new_new_n44478__;
  assign ys__n32048 = ~new_new_n12627__ & ~new_new_n44479__;
  assign new_new_n44481__ = ys__n47716 & ~new_new_n12625__;
  assign new_new_n44482__ = ys__n47747 & new_new_n12626__;
  assign new_new_n44483__ = ~new_new_n44481__ & ~new_new_n44482__;
  assign ys__n32049 = ~new_new_n12627__ & ~new_new_n44483__;
  assign new_new_n44485__ = ys__n47717 & ~new_new_n12625__;
  assign new_new_n44486__ = ys__n47748 & new_new_n12626__;
  assign new_new_n44487__ = ~new_new_n44485__ & ~new_new_n44486__;
  assign ys__n32050 = ~new_new_n12627__ & ~new_new_n44487__;
  assign new_new_n44489__ = ys__n47718 & ~new_new_n12625__;
  assign new_new_n44490__ = ys__n47749 & new_new_n12626__;
  assign new_new_n44491__ = ~new_new_n44489__ & ~new_new_n44490__;
  assign ys__n32051 = ~new_new_n12627__ & ~new_new_n44491__;
  assign new_new_n44493__ = ys__n47719 & ~new_new_n12625__;
  assign new_new_n44494__ = ys__n47750 & new_new_n12626__;
  assign new_new_n44495__ = ~new_new_n44493__ & ~new_new_n44494__;
  assign ys__n32052 = ~new_new_n12627__ & ~new_new_n44495__;
  assign new_new_n44497__ = ys__n47720 & ~new_new_n12625__;
  assign new_new_n44498__ = ys__n47751 & new_new_n12626__;
  assign new_new_n44499__ = ~new_new_n44497__ & ~new_new_n44498__;
  assign ys__n32053 = ~new_new_n12627__ & ~new_new_n44499__;
  assign new_new_n44501__ = ys__n47721 & ~new_new_n12625__;
  assign new_new_n44502__ = ys__n47752 & new_new_n12626__;
  assign new_new_n44503__ = ~new_new_n44501__ & ~new_new_n44502__;
  assign ys__n32054 = ~new_new_n12627__ & ~new_new_n44503__;
  assign new_new_n44505__ = ys__n47722 & ~new_new_n12625__;
  assign new_new_n44506__ = ys__n47753 & new_new_n12626__;
  assign new_new_n44507__ = ~new_new_n44505__ & ~new_new_n44506__;
  assign ys__n32055 = ~new_new_n12627__ & ~new_new_n44507__;
  assign new_new_n44509__ = ys__n38323 & ~new_new_n12625__;
  assign new_new_n44510__ = ys__n47754 & new_new_n12626__;
  assign new_new_n44511__ = ~new_new_n44509__ & ~new_new_n44510__;
  assign ys__n32056 = ~new_new_n12627__ & ~new_new_n44511__;
  assign new_new_n44513__ = ~ys__n935 & new_new_n12297__;
  assign new_new_n44514__ = ys__n28462 & new_new_n44513__;
  assign new_new_n44515__ = ~ys__n226 & ys__n935;
  assign new_new_n44516__ = new_new_n12303__ & new_new_n44515__;
  assign new_new_n44517__ = ys__n23077 & new_new_n44516__;
  assign new_new_n44518__ = ys__n226 & ys__n935;
  assign new_new_n44519__ = ys__n22918 & new_new_n44518__;
  assign new_new_n44520__ = ~new_new_n12303__ & new_new_n44515__;
  assign new_new_n44521__ = ys__n23014 & new_new_n44520__;
  assign new_new_n44522__ = ~new_new_n44519__ & ~new_new_n44521__;
  assign new_new_n44523__ = ~new_new_n44517__ & new_new_n44522__;
  assign new_new_n44524__ = ~new_new_n44514__ & new_new_n44523__;
  assign new_new_n44525__ = ~new_new_n44518__ & ~new_new_n44520__;
  assign new_new_n44526__ = ~new_new_n44516__ & new_new_n44525__;
  assign new_new_n44527__ = ~new_new_n44513__ & new_new_n44526__;
  assign ys__n32057 = ~new_new_n44524__ & ~new_new_n44527__;
  assign new_new_n44529__ = ys__n28464 & new_new_n44513__;
  assign new_new_n44530__ = ys__n23078 & new_new_n44516__;
  assign new_new_n44531__ = ys__n22921 & new_new_n44518__;
  assign new_new_n44532__ = ys__n23016 & new_new_n44520__;
  assign new_new_n44533__ = ~new_new_n44531__ & ~new_new_n44532__;
  assign new_new_n44534__ = ~new_new_n44530__ & new_new_n44533__;
  assign new_new_n44535__ = ~new_new_n44529__ & new_new_n44534__;
  assign ys__n32058 = ~new_new_n44527__ & ~new_new_n44535__;
  assign new_new_n44537__ = ys__n28466 & new_new_n44513__;
  assign new_new_n44538__ = ys__n23079 & new_new_n44516__;
  assign new_new_n44539__ = ys__n22924 & new_new_n44518__;
  assign new_new_n44540__ = ys__n23018 & new_new_n44520__;
  assign new_new_n44541__ = ~new_new_n44539__ & ~new_new_n44540__;
  assign new_new_n44542__ = ~new_new_n44538__ & new_new_n44541__;
  assign new_new_n44543__ = ~new_new_n44537__ & new_new_n44542__;
  assign ys__n32059 = ~new_new_n44527__ & ~new_new_n44543__;
  assign new_new_n44545__ = ys__n28468 & new_new_n44513__;
  assign new_new_n44546__ = ys__n23080 & new_new_n44516__;
  assign new_new_n44547__ = ys__n22927 & new_new_n44518__;
  assign new_new_n44548__ = ys__n23020 & new_new_n44520__;
  assign new_new_n44549__ = ~new_new_n44547__ & ~new_new_n44548__;
  assign new_new_n44550__ = ~new_new_n44546__ & new_new_n44549__;
  assign new_new_n44551__ = ~new_new_n44545__ & new_new_n44550__;
  assign ys__n32060 = ~new_new_n44527__ & ~new_new_n44551__;
  assign new_new_n44553__ = ys__n28470 & new_new_n44513__;
  assign new_new_n44554__ = ys__n23081 & new_new_n44516__;
  assign new_new_n44555__ = ys__n22930 & new_new_n44518__;
  assign new_new_n44556__ = ys__n23022 & new_new_n44520__;
  assign new_new_n44557__ = ~new_new_n44555__ & ~new_new_n44556__;
  assign new_new_n44558__ = ~new_new_n44554__ & new_new_n44557__;
  assign new_new_n44559__ = ~new_new_n44553__ & new_new_n44558__;
  assign ys__n32061 = ~new_new_n44527__ & ~new_new_n44559__;
  assign new_new_n44561__ = ys__n28472 & new_new_n44513__;
  assign new_new_n44562__ = ys__n23082 & new_new_n44516__;
  assign new_new_n44563__ = ys__n22933 & new_new_n44518__;
  assign new_new_n44564__ = ys__n23024 & new_new_n44520__;
  assign new_new_n44565__ = ~new_new_n44563__ & ~new_new_n44564__;
  assign new_new_n44566__ = ~new_new_n44562__ & new_new_n44565__;
  assign new_new_n44567__ = ~new_new_n44561__ & new_new_n44566__;
  assign ys__n32062 = ~new_new_n44527__ & ~new_new_n44567__;
  assign new_new_n44569__ = ys__n29558 & new_new_n44513__;
  assign new_new_n44570__ = ys__n23083 & new_new_n44516__;
  assign new_new_n44571__ = ys__n22936 & new_new_n44518__;
  assign new_new_n44572__ = ys__n23026 & new_new_n44520__;
  assign new_new_n44573__ = ~new_new_n44571__ & ~new_new_n44572__;
  assign new_new_n44574__ = ~new_new_n44570__ & new_new_n44573__;
  assign new_new_n44575__ = ~new_new_n44569__ & new_new_n44574__;
  assign ys__n32063 = ~new_new_n44527__ & ~new_new_n44575__;
  assign new_new_n44577__ = ys__n29560 & new_new_n44513__;
  assign new_new_n44578__ = ys__n23084 & new_new_n44516__;
  assign new_new_n44579__ = ys__n22939 & new_new_n44518__;
  assign new_new_n44580__ = ys__n23028 & new_new_n44520__;
  assign new_new_n44581__ = ~new_new_n44579__ & ~new_new_n44580__;
  assign new_new_n44582__ = ~new_new_n44578__ & new_new_n44581__;
  assign new_new_n44583__ = ~new_new_n44577__ & new_new_n44582__;
  assign ys__n32064 = ~new_new_n44527__ & ~new_new_n44583__;
  assign new_new_n44585__ = ys__n29562 & new_new_n44513__;
  assign new_new_n44586__ = ys__n23085 & new_new_n44516__;
  assign new_new_n44587__ = ys__n22942 & new_new_n44518__;
  assign new_new_n44588__ = ys__n23030 & new_new_n44520__;
  assign new_new_n44589__ = ~new_new_n44587__ & ~new_new_n44588__;
  assign new_new_n44590__ = ~new_new_n44586__ & new_new_n44589__;
  assign new_new_n44591__ = ~new_new_n44585__ & new_new_n44590__;
  assign ys__n32065 = ~new_new_n44527__ & ~new_new_n44591__;
  assign new_new_n44593__ = ys__n29564 & new_new_n44513__;
  assign new_new_n44594__ = ys__n23086 & new_new_n44516__;
  assign new_new_n44595__ = ys__n22945 & new_new_n44518__;
  assign new_new_n44596__ = ys__n23032 & new_new_n44520__;
  assign new_new_n44597__ = ~new_new_n44595__ & ~new_new_n44596__;
  assign new_new_n44598__ = ~new_new_n44594__ & new_new_n44597__;
  assign new_new_n44599__ = ~new_new_n44593__ & new_new_n44598__;
  assign ys__n32066 = ~new_new_n44527__ & ~new_new_n44599__;
  assign new_new_n44601__ = ys__n29566 & new_new_n44513__;
  assign new_new_n44602__ = ys__n23087 & new_new_n44516__;
  assign new_new_n44603__ = ys__n22948 & new_new_n44518__;
  assign new_new_n44604__ = ys__n23034 & new_new_n44520__;
  assign new_new_n44605__ = ~new_new_n44603__ & ~new_new_n44604__;
  assign new_new_n44606__ = ~new_new_n44602__ & new_new_n44605__;
  assign new_new_n44607__ = ~new_new_n44601__ & new_new_n44606__;
  assign ys__n32067 = ~new_new_n44527__ & ~new_new_n44607__;
  assign new_new_n44609__ = ys__n29568 & new_new_n44513__;
  assign new_new_n44610__ = ys__n23088 & new_new_n44516__;
  assign new_new_n44611__ = ys__n22951 & new_new_n44518__;
  assign new_new_n44612__ = ys__n23036 & new_new_n44520__;
  assign new_new_n44613__ = ~new_new_n44611__ & ~new_new_n44612__;
  assign new_new_n44614__ = ~new_new_n44610__ & new_new_n44613__;
  assign new_new_n44615__ = ~new_new_n44609__ & new_new_n44614__;
  assign ys__n32068 = ~new_new_n44527__ & ~new_new_n44615__;
  assign new_new_n44617__ = ys__n29570 & new_new_n44513__;
  assign new_new_n44618__ = ys__n23089 & new_new_n44516__;
  assign new_new_n44619__ = ys__n22954 & new_new_n44518__;
  assign new_new_n44620__ = ys__n23038 & new_new_n44520__;
  assign new_new_n44621__ = ~new_new_n44619__ & ~new_new_n44620__;
  assign new_new_n44622__ = ~new_new_n44618__ & new_new_n44621__;
  assign new_new_n44623__ = ~new_new_n44617__ & new_new_n44622__;
  assign ys__n32069 = ~new_new_n44527__ & ~new_new_n44623__;
  assign new_new_n44625__ = ys__n29572 & new_new_n44513__;
  assign new_new_n44626__ = ys__n23090 & new_new_n44516__;
  assign new_new_n44627__ = ys__n22957 & new_new_n44518__;
  assign new_new_n44628__ = ys__n23040 & new_new_n44520__;
  assign new_new_n44629__ = ~new_new_n44627__ & ~new_new_n44628__;
  assign new_new_n44630__ = ~new_new_n44626__ & new_new_n44629__;
  assign new_new_n44631__ = ~new_new_n44625__ & new_new_n44630__;
  assign ys__n32070 = ~new_new_n44527__ & ~new_new_n44631__;
  assign new_new_n44633__ = ys__n29574 & new_new_n44513__;
  assign new_new_n44634__ = ys__n23091 & new_new_n44516__;
  assign new_new_n44635__ = ys__n22960 & new_new_n44518__;
  assign new_new_n44636__ = ys__n23042 & new_new_n44520__;
  assign new_new_n44637__ = ~new_new_n44635__ & ~new_new_n44636__;
  assign new_new_n44638__ = ~new_new_n44634__ & new_new_n44637__;
  assign new_new_n44639__ = ~new_new_n44633__ & new_new_n44638__;
  assign ys__n32071 = ~new_new_n44527__ & ~new_new_n44639__;
  assign new_new_n44641__ = ys__n29576 & new_new_n44513__;
  assign new_new_n44642__ = ys__n23092 & new_new_n44516__;
  assign new_new_n44643__ = ys__n22963 & new_new_n44518__;
  assign new_new_n44644__ = ys__n23044 & new_new_n44520__;
  assign new_new_n44645__ = ~new_new_n44643__ & ~new_new_n44644__;
  assign new_new_n44646__ = ~new_new_n44642__ & new_new_n44645__;
  assign new_new_n44647__ = ~new_new_n44641__ & new_new_n44646__;
  assign ys__n32072 = ~new_new_n44527__ & ~new_new_n44647__;
  assign new_new_n44649__ = ys__n29578 & new_new_n44513__;
  assign new_new_n44650__ = ys__n23093 & new_new_n44516__;
  assign new_new_n44651__ = ys__n22966 & new_new_n44518__;
  assign new_new_n44652__ = ys__n23046 & new_new_n44520__;
  assign new_new_n44653__ = ~new_new_n44651__ & ~new_new_n44652__;
  assign new_new_n44654__ = ~new_new_n44650__ & new_new_n44653__;
  assign new_new_n44655__ = ~new_new_n44649__ & new_new_n44654__;
  assign ys__n32073 = ~new_new_n44527__ & ~new_new_n44655__;
  assign new_new_n44657__ = ys__n29580 & new_new_n44513__;
  assign new_new_n44658__ = ys__n23094 & new_new_n44516__;
  assign new_new_n44659__ = ys__n22969 & new_new_n44518__;
  assign new_new_n44660__ = ys__n23048 & new_new_n44520__;
  assign new_new_n44661__ = ~new_new_n44659__ & ~new_new_n44660__;
  assign new_new_n44662__ = ~new_new_n44658__ & new_new_n44661__;
  assign new_new_n44663__ = ~new_new_n44657__ & new_new_n44662__;
  assign ys__n32074 = ~new_new_n44527__ & ~new_new_n44663__;
  assign new_new_n44665__ = ys__n29582 & new_new_n44513__;
  assign new_new_n44666__ = ys__n23095 & new_new_n44516__;
  assign new_new_n44667__ = ys__n22972 & new_new_n44518__;
  assign new_new_n44668__ = ys__n23050 & new_new_n44520__;
  assign new_new_n44669__ = ~new_new_n44667__ & ~new_new_n44668__;
  assign new_new_n44670__ = ~new_new_n44666__ & new_new_n44669__;
  assign new_new_n44671__ = ~new_new_n44665__ & new_new_n44670__;
  assign ys__n32075 = ~new_new_n44527__ & ~new_new_n44671__;
  assign new_new_n44673__ = ys__n29584 & new_new_n44513__;
  assign new_new_n44674__ = ys__n23096 & new_new_n44516__;
  assign new_new_n44675__ = ys__n22975 & new_new_n44518__;
  assign new_new_n44676__ = ys__n23052 & new_new_n44520__;
  assign new_new_n44677__ = ~new_new_n44675__ & ~new_new_n44676__;
  assign new_new_n44678__ = ~new_new_n44674__ & new_new_n44677__;
  assign new_new_n44679__ = ~new_new_n44673__ & new_new_n44678__;
  assign ys__n32076 = ~new_new_n44527__ & ~new_new_n44679__;
  assign new_new_n44681__ = ys__n29586 & new_new_n44513__;
  assign new_new_n44682__ = ys__n23097 & new_new_n44516__;
  assign new_new_n44683__ = ys__n22978 & new_new_n44518__;
  assign new_new_n44684__ = ys__n23054 & new_new_n44520__;
  assign new_new_n44685__ = ~new_new_n44683__ & ~new_new_n44684__;
  assign new_new_n44686__ = ~new_new_n44682__ & new_new_n44685__;
  assign new_new_n44687__ = ~new_new_n44681__ & new_new_n44686__;
  assign ys__n32077 = ~new_new_n44527__ & ~new_new_n44687__;
  assign new_new_n44689__ = ys__n29588 & new_new_n44513__;
  assign new_new_n44690__ = ys__n23098 & new_new_n44516__;
  assign new_new_n44691__ = ys__n22981 & new_new_n44518__;
  assign new_new_n44692__ = ys__n23056 & new_new_n44520__;
  assign new_new_n44693__ = ~new_new_n44691__ & ~new_new_n44692__;
  assign new_new_n44694__ = ~new_new_n44690__ & new_new_n44693__;
  assign new_new_n44695__ = ~new_new_n44689__ & new_new_n44694__;
  assign ys__n32078 = ~new_new_n44527__ & ~new_new_n44695__;
  assign new_new_n44697__ = ys__n29590 & new_new_n44513__;
  assign new_new_n44698__ = ys__n23099 & new_new_n44516__;
  assign new_new_n44699__ = ys__n22984 & new_new_n44518__;
  assign new_new_n44700__ = ys__n23058 & new_new_n44520__;
  assign new_new_n44701__ = ~new_new_n44699__ & ~new_new_n44700__;
  assign new_new_n44702__ = ~new_new_n44698__ & new_new_n44701__;
  assign new_new_n44703__ = ~new_new_n44697__ & new_new_n44702__;
  assign ys__n32079 = ~new_new_n44527__ & ~new_new_n44703__;
  assign new_new_n44705__ = ys__n29592 & new_new_n44513__;
  assign new_new_n44706__ = ys__n23100 & new_new_n44516__;
  assign new_new_n44707__ = ys__n22987 & new_new_n44518__;
  assign new_new_n44708__ = ys__n23060 & new_new_n44520__;
  assign new_new_n44709__ = ~new_new_n44707__ & ~new_new_n44708__;
  assign new_new_n44710__ = ~new_new_n44706__ & new_new_n44709__;
  assign new_new_n44711__ = ~new_new_n44705__ & new_new_n44710__;
  assign ys__n32080 = ~new_new_n44527__ & ~new_new_n44711__;
  assign new_new_n44713__ = ys__n29594 & new_new_n44513__;
  assign new_new_n44714__ = ys__n23101 & new_new_n44516__;
  assign new_new_n44715__ = ys__n22990 & new_new_n44518__;
  assign new_new_n44716__ = ys__n23062 & new_new_n44520__;
  assign new_new_n44717__ = ~new_new_n44715__ & ~new_new_n44716__;
  assign new_new_n44718__ = ~new_new_n44714__ & new_new_n44717__;
  assign new_new_n44719__ = ~new_new_n44713__ & new_new_n44718__;
  assign ys__n32081 = ~new_new_n44527__ & ~new_new_n44719__;
  assign new_new_n44721__ = ys__n29596 & new_new_n44513__;
  assign new_new_n44722__ = ys__n23102 & new_new_n44516__;
  assign new_new_n44723__ = ys__n22993 & new_new_n44518__;
  assign new_new_n44724__ = ys__n23064 & new_new_n44520__;
  assign new_new_n44725__ = ~new_new_n44723__ & ~new_new_n44724__;
  assign new_new_n44726__ = ~new_new_n44722__ & new_new_n44725__;
  assign new_new_n44727__ = ~new_new_n44721__ & new_new_n44726__;
  assign ys__n32082 = ~new_new_n44527__ & ~new_new_n44727__;
  assign new_new_n44729__ = ys__n29598 & new_new_n44513__;
  assign new_new_n44730__ = ys__n23103 & new_new_n44516__;
  assign new_new_n44731__ = ys__n22996 & new_new_n44518__;
  assign new_new_n44732__ = ys__n23066 & new_new_n44520__;
  assign new_new_n44733__ = ~new_new_n44731__ & ~new_new_n44732__;
  assign new_new_n44734__ = ~new_new_n44730__ & new_new_n44733__;
  assign new_new_n44735__ = ~new_new_n44729__ & new_new_n44734__;
  assign ys__n32083 = ~new_new_n44527__ & ~new_new_n44735__;
  assign new_new_n44737__ = ys__n29600 & new_new_n44513__;
  assign new_new_n44738__ = ys__n23104 & new_new_n44516__;
  assign new_new_n44739__ = ys__n22999 & new_new_n44518__;
  assign new_new_n44740__ = ys__n23068 & new_new_n44520__;
  assign new_new_n44741__ = ~new_new_n44739__ & ~new_new_n44740__;
  assign new_new_n44742__ = ~new_new_n44738__ & new_new_n44741__;
  assign new_new_n44743__ = ~new_new_n44737__ & new_new_n44742__;
  assign ys__n32084 = ~new_new_n44527__ & ~new_new_n44743__;
  assign new_new_n44745__ = ys__n29602 & new_new_n44513__;
  assign new_new_n44746__ = ys__n23105 & new_new_n44516__;
  assign new_new_n44747__ = ys__n23002 & new_new_n44518__;
  assign new_new_n44748__ = ys__n23070 & new_new_n44520__;
  assign new_new_n44749__ = ~new_new_n44747__ & ~new_new_n44748__;
  assign new_new_n44750__ = ~new_new_n44746__ & new_new_n44749__;
  assign new_new_n44751__ = ~new_new_n44745__ & new_new_n44750__;
  assign ys__n32085 = ~new_new_n44527__ & ~new_new_n44751__;
  assign new_new_n44753__ = ys__n29604 & new_new_n44513__;
  assign new_new_n44754__ = ys__n23106 & new_new_n44516__;
  assign new_new_n44755__ = ys__n23005 & new_new_n44518__;
  assign new_new_n44756__ = ys__n23072 & new_new_n44520__;
  assign new_new_n44757__ = ~new_new_n44755__ & ~new_new_n44756__;
  assign new_new_n44758__ = ~new_new_n44754__ & new_new_n44757__;
  assign new_new_n44759__ = ~new_new_n44753__ & new_new_n44758__;
  assign ys__n32086 = ~new_new_n44527__ & ~new_new_n44759__;
  assign new_new_n44761__ = ys__n29606 & new_new_n44513__;
  assign new_new_n44762__ = ys__n23107 & new_new_n44516__;
  assign new_new_n44763__ = ys__n23008 & new_new_n44518__;
  assign new_new_n44764__ = ys__n23074 & new_new_n44520__;
  assign new_new_n44765__ = ~new_new_n44763__ & ~new_new_n44764__;
  assign new_new_n44766__ = ~new_new_n44762__ & new_new_n44765__;
  assign new_new_n44767__ = ~new_new_n44761__ & new_new_n44766__;
  assign ys__n32087 = ~new_new_n44527__ & ~new_new_n44767__;
  assign new_new_n44769__ = ys__n29608 & new_new_n44513__;
  assign new_new_n44770__ = ys__n23108 & new_new_n44516__;
  assign new_new_n44771__ = ys__n23011 & new_new_n44518__;
  assign new_new_n44772__ = ys__n23076 & new_new_n44520__;
  assign new_new_n44773__ = ~new_new_n44771__ & ~new_new_n44772__;
  assign new_new_n44774__ = ~new_new_n44770__ & new_new_n44773__;
  assign new_new_n44775__ = ~new_new_n44769__ & new_new_n44774__;
  assign ys__n32088 = ~new_new_n44527__ & ~new_new_n44775__;
  assign new_new_n44777__ = ~new_new_n22623__ & ~new_new_n37452__;
  assign new_new_n44778__ = ~new_new_n23118__ & ~new_new_n44777__;
  assign new_new_n44779__ = ys__n38486 & new_new_n22618__;
  assign new_new_n44780__ = ~new_new_n44778__ & ~new_new_n44779__;
  assign new_new_n44781__ = ys__n27743 & new_new_n44779__;
  assign new_new_n44782__ = ~new_new_n44780__ & ~new_new_n44781__;
  assign new_new_n44783__ = ~ys__n278 & ~ys__n814;
  assign new_new_n44784__ = new_new_n12566__ & new_new_n44783__;
  assign new_new_n44785__ = ys__n20273 & ~ys__n250;
  assign new_new_n44786__ = ~ys__n252 & new_new_n44785__;
  assign new_new_n44787__ = new_new_n44784__ & new_new_n44786__;
  assign new_new_n44788__ = ys__n254 & new_new_n44787__;
  assign new_new_n44789__ = ~new_new_n44782__ & new_new_n44788__;
  assign new_new_n44790__ = ys__n20273 & ys__n250;
  assign new_new_n44791__ = new_new_n44784__ & new_new_n44790__;
  assign new_new_n44792__ = new_new_n12564__ & new_new_n44791__;
  assign new_new_n44793__ = ys__n19878 & new_new_n44792__;
  assign new_new_n44794__ = ys__n20956 & ~ys__n28243;
  assign new_new_n44795__ = ys__n21276 & ys__n28243;
  assign new_new_n44796__ = ~new_new_n44794__ & ~new_new_n44795__;
  assign new_new_n44797__ = ys__n28243 & ~new_new_n44796__;
  assign new_new_n44798__ = ~ys__n28243 & new_new_n44797__;
  assign new_new_n44799__ = ys__n21500 & ~ys__n28243;
  assign new_new_n44800__ = ys__n21820 & ys__n28243;
  assign new_new_n44801__ = ~new_new_n44799__ & ~new_new_n44800__;
  assign new_new_n44802__ = ~ys__n28243 & ~new_new_n44801__;
  assign new_new_n44803__ = ys__n21980 & ~ys__n28243;
  assign new_new_n44804__ = ys__n22300 & ys__n28243;
  assign new_new_n44805__ = ~new_new_n44803__ & ~new_new_n44804__;
  assign new_new_n44806__ = ys__n28243 & ~new_new_n44805__;
  assign new_new_n44807__ = ~new_new_n44802__ & ~new_new_n44806__;
  assign new_new_n44808__ = ys__n28243 & ~new_new_n44807__;
  assign new_new_n44809__ = ~new_new_n44798__ & ~new_new_n44808__;
  assign new_new_n44810__ = ys__n20273 & ~ys__n814;
  assign new_new_n44811__ = ys__n278 & new_new_n44810__;
  assign new_new_n44812__ = new_new_n12566__ & new_new_n44811__;
  assign new_new_n44813__ = new_new_n12565__ & new_new_n44812__;
  assign new_new_n44814__ = ~new_new_n44809__ & new_new_n44813__;
  assign new_new_n44815__ = ys__n252 & new_new_n44785__;
  assign new_new_n44816__ = new_new_n44784__ & new_new_n44815__;
  assign new_new_n44817__ = ~ys__n254 & new_new_n44816__;
  assign new_new_n44818__ = ys__n47791 & new_new_n44817__;
  assign new_new_n44819__ = ~new_new_n44814__ & ~new_new_n44818__;
  assign new_new_n44820__ = ys__n20273 & ~ys__n246;
  assign new_new_n44821__ = ys__n270 & new_new_n44820__;
  assign new_new_n44822__ = new_new_n44783__ & new_new_n44821__;
  assign new_new_n44823__ = new_new_n12565__ & new_new_n44822__;
  assign new_new_n44824__ = ys__n47759 & new_new_n44823__;
  assign new_new_n44825__ = ys__n464 & ~ys__n28243;
  assign new_new_n44826__ = ys__n28288 & ys__n28296;
  assign new_new_n44827__ = ys__n28243 & new_new_n44826__;
  assign new_new_n44828__ = ~new_new_n44825__ & ~new_new_n44827__;
  assign new_new_n44829__ = ys__n20273 & ys__n246;
  assign new_new_n44830__ = ~ys__n270 & new_new_n44829__;
  assign new_new_n44831__ = new_new_n44783__ & new_new_n44830__;
  assign new_new_n44832__ = new_new_n12565__ & new_new_n44831__;
  assign new_new_n44833__ = ~new_new_n44828__ & new_new_n44832__;
  assign new_new_n44834__ = ~new_new_n44824__ & ~new_new_n44833__;
  assign new_new_n44835__ = new_new_n44819__ & new_new_n44834__;
  assign new_new_n44836__ = ~new_new_n44793__ & new_new_n44835__;
  assign new_new_n44837__ = ~new_new_n44789__ & new_new_n44836__;
  assign new_new_n44838__ = ~new_new_n44788__ & ~new_new_n44817__;
  assign new_new_n44839__ = ~new_new_n44792__ & new_new_n44838__;
  assign new_new_n44840__ = ~new_new_n44813__ & new_new_n44839__;
  assign new_new_n44841__ = ~ys__n20273 & new_new_n44784__;
  assign new_new_n44842__ = new_new_n12565__ & new_new_n44841__;
  assign new_new_n44843__ = ~new_new_n44823__ & ~new_new_n44832__;
  assign new_new_n44844__ = ~new_new_n44842__ & new_new_n44843__;
  assign new_new_n44845__ = new_new_n44840__ & new_new_n44844__;
  assign ys__n32124 = ~new_new_n44837__ & ~new_new_n44845__;
  assign new_new_n44847__ = ~new_new_n22623__ & ~new_new_n37461__;
  assign new_new_n44848__ = ~new_new_n23137__ & ~new_new_n44847__;
  assign new_new_n44849__ = ~new_new_n44779__ & ~new_new_n44848__;
  assign new_new_n44850__ = ys__n27747 & new_new_n44779__;
  assign new_new_n44851__ = ~new_new_n44849__ & ~new_new_n44850__;
  assign new_new_n44852__ = new_new_n44788__ & ~new_new_n44851__;
  assign new_new_n44853__ = ys__n19881 & new_new_n44792__;
  assign new_new_n44854__ = ys__n20958 & ~ys__n28243;
  assign new_new_n44855__ = ys__n21278 & ys__n28243;
  assign new_new_n44856__ = ~new_new_n44854__ & ~new_new_n44855__;
  assign new_new_n44857__ = ys__n28243 & ~new_new_n44856__;
  assign new_new_n44858__ = ~ys__n28243 & new_new_n44857__;
  assign new_new_n44859__ = ys__n21502 & ~ys__n28243;
  assign new_new_n44860__ = ys__n21822 & ys__n28243;
  assign new_new_n44861__ = ~new_new_n44859__ & ~new_new_n44860__;
  assign new_new_n44862__ = ~ys__n28243 & ~new_new_n44861__;
  assign new_new_n44863__ = ys__n21982 & ~ys__n28243;
  assign new_new_n44864__ = ys__n22302 & ys__n28243;
  assign new_new_n44865__ = ~new_new_n44863__ & ~new_new_n44864__;
  assign new_new_n44866__ = ys__n28243 & ~new_new_n44865__;
  assign new_new_n44867__ = ~new_new_n44862__ & ~new_new_n44866__;
  assign new_new_n44868__ = ys__n28243 & ~new_new_n44867__;
  assign new_new_n44869__ = ~new_new_n44858__ & ~new_new_n44868__;
  assign new_new_n44870__ = new_new_n44813__ & ~new_new_n44869__;
  assign new_new_n44871__ = ys__n47792 & new_new_n44817__;
  assign new_new_n44872__ = ~new_new_n44870__ & ~new_new_n44871__;
  assign new_new_n44873__ = ys__n47760 & new_new_n44823__;
  assign new_new_n44874__ = ys__n4340 & ~ys__n28243;
  assign new_new_n44875__ = ys__n28287 & ys__n28288;
  assign new_new_n44876__ = ys__n28243 & new_new_n44875__;
  assign new_new_n44877__ = ~new_new_n44874__ & ~new_new_n44876__;
  assign new_new_n44878__ = new_new_n44832__ & ~new_new_n44877__;
  assign new_new_n44879__ = ~new_new_n44873__ & ~new_new_n44878__;
  assign new_new_n44880__ = new_new_n44872__ & new_new_n44879__;
  assign new_new_n44881__ = ~new_new_n44853__ & new_new_n44880__;
  assign new_new_n44882__ = ~new_new_n44852__ & new_new_n44881__;
  assign ys__n32125 = ~new_new_n44845__ & ~new_new_n44882__;
  assign new_new_n44884__ = ~new_new_n22623__ & ~new_new_n37469__;
  assign new_new_n44885__ = ~new_new_n23156__ & ~new_new_n44884__;
  assign new_new_n44886__ = ~new_new_n44779__ & ~new_new_n44885__;
  assign new_new_n44887__ = ys__n27750 & new_new_n44779__;
  assign new_new_n44888__ = ~new_new_n44886__ & ~new_new_n44887__;
  assign new_new_n44889__ = new_new_n44788__ & ~new_new_n44888__;
  assign new_new_n44890__ = ys__n19884 & new_new_n44792__;
  assign new_new_n44891__ = ys__n20960 & ~ys__n28243;
  assign new_new_n44892__ = ys__n21280 & ys__n28243;
  assign new_new_n44893__ = ~new_new_n44891__ & ~new_new_n44892__;
  assign new_new_n44894__ = ys__n28243 & ~new_new_n44893__;
  assign new_new_n44895__ = ~ys__n28243 & new_new_n44894__;
  assign new_new_n44896__ = ys__n21504 & ~ys__n28243;
  assign new_new_n44897__ = ys__n21824 & ys__n28243;
  assign new_new_n44898__ = ~new_new_n44896__ & ~new_new_n44897__;
  assign new_new_n44899__ = ~ys__n28243 & ~new_new_n44898__;
  assign new_new_n44900__ = ys__n21984 & ~ys__n28243;
  assign new_new_n44901__ = ys__n22304 & ys__n28243;
  assign new_new_n44902__ = ~new_new_n44900__ & ~new_new_n44901__;
  assign new_new_n44903__ = ys__n28243 & ~new_new_n44902__;
  assign new_new_n44904__ = ~new_new_n44899__ & ~new_new_n44903__;
  assign new_new_n44905__ = ys__n28243 & ~new_new_n44904__;
  assign new_new_n44906__ = ~new_new_n44895__ & ~new_new_n44905__;
  assign new_new_n44907__ = new_new_n44813__ & ~new_new_n44906__;
  assign new_new_n44908__ = ys__n47793 & new_new_n44817__;
  assign new_new_n44909__ = ~new_new_n44907__ & ~new_new_n44908__;
  assign new_new_n44910__ = ys__n47761 & new_new_n44823__;
  assign new_new_n44911__ = ys__n240 & ~ys__n28243;
  assign new_new_n44912__ = ys__n464 & ~ys__n28288;
  assign new_new_n44913__ = ys__n28288 & ys__n28290;
  assign new_new_n44914__ = ~new_new_n44912__ & ~new_new_n44913__;
  assign new_new_n44915__ = ys__n28243 & ~new_new_n44914__;
  assign new_new_n44916__ = ~new_new_n44911__ & ~new_new_n44915__;
  assign new_new_n44917__ = new_new_n44832__ & ~new_new_n44916__;
  assign new_new_n44918__ = ~new_new_n44910__ & ~new_new_n44917__;
  assign new_new_n44919__ = new_new_n44909__ & new_new_n44918__;
  assign new_new_n44920__ = ~new_new_n44890__ & new_new_n44919__;
  assign new_new_n44921__ = ~new_new_n44889__ & new_new_n44920__;
  assign ys__n32126 = ~new_new_n44845__ & ~new_new_n44921__;
  assign new_new_n44923__ = ~new_new_n22623__ & ~new_new_n37477__;
  assign new_new_n44924__ = ~new_new_n23175__ & ~new_new_n44923__;
  assign new_new_n44925__ = ~new_new_n44779__ & ~new_new_n44924__;
  assign new_new_n44926__ = ys__n27753 & new_new_n44779__;
  assign new_new_n44927__ = ~new_new_n44925__ & ~new_new_n44926__;
  assign new_new_n44928__ = new_new_n44788__ & ~new_new_n44927__;
  assign new_new_n44929__ = ys__n19887 & new_new_n44792__;
  assign new_new_n44930__ = ys__n20962 & ~ys__n28243;
  assign new_new_n44931__ = ys__n21282 & ys__n28243;
  assign new_new_n44932__ = ~new_new_n44930__ & ~new_new_n44931__;
  assign new_new_n44933__ = ys__n28243 & ~new_new_n44932__;
  assign new_new_n44934__ = ~ys__n28243 & new_new_n44933__;
  assign new_new_n44935__ = ys__n21506 & ~ys__n28243;
  assign new_new_n44936__ = ys__n21826 & ys__n28243;
  assign new_new_n44937__ = ~new_new_n44935__ & ~new_new_n44936__;
  assign new_new_n44938__ = ~ys__n28243 & ~new_new_n44937__;
  assign new_new_n44939__ = ys__n21986 & ~ys__n28243;
  assign new_new_n44940__ = ys__n22306 & ys__n28243;
  assign new_new_n44941__ = ~new_new_n44939__ & ~new_new_n44940__;
  assign new_new_n44942__ = ys__n28243 & ~new_new_n44941__;
  assign new_new_n44943__ = ~new_new_n44938__ & ~new_new_n44942__;
  assign new_new_n44944__ = ys__n28243 & ~new_new_n44943__;
  assign new_new_n44945__ = ~new_new_n44934__ & ~new_new_n44944__;
  assign new_new_n44946__ = new_new_n44813__ & ~new_new_n44945__;
  assign new_new_n44947__ = ys__n47794 & new_new_n44817__;
  assign new_new_n44948__ = ~new_new_n44946__ & ~new_new_n44947__;
  assign new_new_n44949__ = ys__n47762 & new_new_n44823__;
  assign new_new_n44950__ = ys__n238 & ~ys__n28243;
  assign new_new_n44951__ = ys__n4340 & ~ys__n28288;
  assign new_new_n44952__ = ys__n28288 & ys__n28292;
  assign new_new_n44953__ = ~new_new_n44951__ & ~new_new_n44952__;
  assign new_new_n44954__ = ys__n28243 & ~new_new_n44953__;
  assign new_new_n44955__ = ~new_new_n44950__ & ~new_new_n44954__;
  assign new_new_n44956__ = new_new_n44832__ & ~new_new_n44955__;
  assign new_new_n44957__ = ~new_new_n44949__ & ~new_new_n44956__;
  assign new_new_n44958__ = new_new_n44948__ & new_new_n44957__;
  assign new_new_n44959__ = ~new_new_n44929__ & new_new_n44958__;
  assign new_new_n44960__ = ~new_new_n44928__ & new_new_n44959__;
  assign ys__n32127 = ~new_new_n44845__ & ~new_new_n44960__;
  assign new_new_n44962__ = ~new_new_n22623__ & ~new_new_n37485__;
  assign new_new_n44963__ = ~new_new_n23194__ & ~new_new_n44962__;
  assign new_new_n44964__ = ~new_new_n44779__ & ~new_new_n44963__;
  assign new_new_n44965__ = ys__n27756 & new_new_n44779__;
  assign new_new_n44966__ = ~new_new_n44964__ & ~new_new_n44965__;
  assign new_new_n44967__ = new_new_n44788__ & ~new_new_n44966__;
  assign new_new_n44968__ = ys__n19890 & new_new_n44792__;
  assign new_new_n44969__ = ys__n20964 & ~ys__n28243;
  assign new_new_n44970__ = ys__n21284 & ys__n28243;
  assign new_new_n44971__ = ~new_new_n44969__ & ~new_new_n44970__;
  assign new_new_n44972__ = ys__n28243 & ~new_new_n44971__;
  assign new_new_n44973__ = ~ys__n28243 & new_new_n44972__;
  assign new_new_n44974__ = ys__n21508 & ~ys__n28243;
  assign new_new_n44975__ = ys__n21828 & ys__n28243;
  assign new_new_n44976__ = ~new_new_n44974__ & ~new_new_n44975__;
  assign new_new_n44977__ = ~ys__n28243 & ~new_new_n44976__;
  assign new_new_n44978__ = ys__n21988 & ~ys__n28243;
  assign new_new_n44979__ = ys__n22308 & ys__n28243;
  assign new_new_n44980__ = ~new_new_n44978__ & ~new_new_n44979__;
  assign new_new_n44981__ = ys__n28243 & ~new_new_n44980__;
  assign new_new_n44982__ = ~new_new_n44977__ & ~new_new_n44981__;
  assign new_new_n44983__ = ys__n28243 & ~new_new_n44982__;
  assign new_new_n44984__ = ~new_new_n44973__ & ~new_new_n44983__;
  assign new_new_n44985__ = new_new_n44813__ & ~new_new_n44984__;
  assign new_new_n44986__ = ys__n47795 & new_new_n44817__;
  assign new_new_n44987__ = ~new_new_n44985__ & ~new_new_n44986__;
  assign new_new_n44988__ = ys__n47763 & new_new_n44823__;
  assign new_new_n44989__ = ys__n242 & ~ys__n28243;
  assign new_new_n44990__ = ys__n28288 & ys__n28294;
  assign new_new_n44991__ = ys__n28243 & new_new_n44990__;
  assign new_new_n44992__ = ~new_new_n44989__ & ~new_new_n44991__;
  assign new_new_n44993__ = new_new_n44832__ & ~new_new_n44992__;
  assign new_new_n44994__ = ~new_new_n44988__ & ~new_new_n44993__;
  assign new_new_n44995__ = new_new_n44987__ & new_new_n44994__;
  assign new_new_n44996__ = ~new_new_n44968__ & new_new_n44995__;
  assign new_new_n44997__ = ~new_new_n44967__ & new_new_n44996__;
  assign ys__n32128 = ~new_new_n44845__ & ~new_new_n44997__;
  assign new_new_n44999__ = ~new_new_n22623__ & ~new_new_n37493__;
  assign new_new_n45000__ = ~new_new_n23213__ & ~new_new_n44999__;
  assign new_new_n45001__ = ~new_new_n44779__ & ~new_new_n45000__;
  assign new_new_n45002__ = ys__n27759 & new_new_n44779__;
  assign new_new_n45003__ = ~new_new_n45001__ & ~new_new_n45002__;
  assign new_new_n45004__ = new_new_n44788__ & ~new_new_n45003__;
  assign new_new_n45005__ = ys__n19893 & new_new_n44792__;
  assign new_new_n45006__ = ys__n47764 & new_new_n44823__;
  assign new_new_n45007__ = ys__n20966 & ~ys__n28243;
  assign new_new_n45008__ = ys__n21286 & ys__n28243;
  assign new_new_n45009__ = ~new_new_n45007__ & ~new_new_n45008__;
  assign new_new_n45010__ = ys__n28243 & ~new_new_n45009__;
  assign new_new_n45011__ = ~ys__n28243 & new_new_n45010__;
  assign new_new_n45012__ = ys__n21510 & ~ys__n28243;
  assign new_new_n45013__ = ys__n21830 & ys__n28243;
  assign new_new_n45014__ = ~new_new_n45012__ & ~new_new_n45013__;
  assign new_new_n45015__ = ~ys__n28243 & ~new_new_n45014__;
  assign new_new_n45016__ = ys__n21990 & ~ys__n28243;
  assign new_new_n45017__ = ys__n22310 & ys__n28243;
  assign new_new_n45018__ = ~new_new_n45016__ & ~new_new_n45017__;
  assign new_new_n45019__ = ys__n28243 & ~new_new_n45018__;
  assign new_new_n45020__ = ~new_new_n45015__ & ~new_new_n45019__;
  assign new_new_n45021__ = ys__n28243 & ~new_new_n45020__;
  assign new_new_n45022__ = ~new_new_n45011__ & ~new_new_n45021__;
  assign new_new_n45023__ = new_new_n44813__ & ~new_new_n45022__;
  assign new_new_n45024__ = ys__n47796 & new_new_n44817__;
  assign new_new_n45025__ = ~new_new_n45023__ & ~new_new_n45024__;
  assign new_new_n45026__ = ~new_new_n45006__ & new_new_n45025__;
  assign new_new_n45027__ = ~new_new_n45005__ & new_new_n45026__;
  assign new_new_n45028__ = ~new_new_n45004__ & new_new_n45027__;
  assign ys__n32129 = ~new_new_n44845__ & ~new_new_n45028__;
  assign new_new_n45030__ = ~new_new_n22623__ & ~new_new_n37501__;
  assign new_new_n45031__ = ~new_new_n23232__ & ~new_new_n45030__;
  assign new_new_n45032__ = ~new_new_n44779__ & ~new_new_n45031__;
  assign new_new_n45033__ = ys__n27762 & new_new_n44779__;
  assign new_new_n45034__ = ~new_new_n45032__ & ~new_new_n45033__;
  assign new_new_n45035__ = new_new_n44788__ & ~new_new_n45034__;
  assign new_new_n45036__ = ys__n19896 & new_new_n44792__;
  assign new_new_n45037__ = ys__n47765 & new_new_n44823__;
  assign new_new_n45038__ = ys__n20968 & ~ys__n28243;
  assign new_new_n45039__ = ys__n21288 & ys__n28243;
  assign new_new_n45040__ = ~new_new_n45038__ & ~new_new_n45039__;
  assign new_new_n45041__ = ys__n28243 & ~new_new_n45040__;
  assign new_new_n45042__ = ~ys__n28243 & new_new_n45041__;
  assign new_new_n45043__ = ys__n21512 & ~ys__n28243;
  assign new_new_n45044__ = ys__n21832 & ys__n28243;
  assign new_new_n45045__ = ~new_new_n45043__ & ~new_new_n45044__;
  assign new_new_n45046__ = ~ys__n28243 & ~new_new_n45045__;
  assign new_new_n45047__ = ys__n21992 & ~ys__n28243;
  assign new_new_n45048__ = ys__n22312 & ys__n28243;
  assign new_new_n45049__ = ~new_new_n45047__ & ~new_new_n45048__;
  assign new_new_n45050__ = ys__n28243 & ~new_new_n45049__;
  assign new_new_n45051__ = ~new_new_n45046__ & ~new_new_n45050__;
  assign new_new_n45052__ = ys__n28243 & ~new_new_n45051__;
  assign new_new_n45053__ = ~new_new_n45042__ & ~new_new_n45052__;
  assign new_new_n45054__ = new_new_n44813__ & ~new_new_n45053__;
  assign new_new_n45055__ = ys__n47797 & new_new_n44817__;
  assign new_new_n45056__ = ~new_new_n45054__ & ~new_new_n45055__;
  assign new_new_n45057__ = ~new_new_n45037__ & new_new_n45056__;
  assign new_new_n45058__ = ~new_new_n45036__ & new_new_n45057__;
  assign new_new_n45059__ = ~new_new_n45035__ & new_new_n45058__;
  assign ys__n32130 = ~new_new_n44845__ & ~new_new_n45059__;
  assign new_new_n45061__ = ~new_new_n22623__ & ~new_new_n37509__;
  assign new_new_n45062__ = ~new_new_n23251__ & ~new_new_n45061__;
  assign new_new_n45063__ = ~new_new_n44779__ & ~new_new_n45062__;
  assign new_new_n45064__ = ys__n27765 & new_new_n44779__;
  assign new_new_n45065__ = ~new_new_n45063__ & ~new_new_n45064__;
  assign new_new_n45066__ = new_new_n44788__ & ~new_new_n45065__;
  assign new_new_n45067__ = ys__n19899 & new_new_n44792__;
  assign new_new_n45068__ = ys__n47766 & new_new_n44823__;
  assign new_new_n45069__ = ys__n20970 & ~ys__n28243;
  assign new_new_n45070__ = ys__n21290 & ys__n28243;
  assign new_new_n45071__ = ~new_new_n45069__ & ~new_new_n45070__;
  assign new_new_n45072__ = ys__n28243 & ~new_new_n45071__;
  assign new_new_n45073__ = ~ys__n28243 & new_new_n45072__;
  assign new_new_n45074__ = ys__n21514 & ~ys__n28243;
  assign new_new_n45075__ = ys__n21834 & ys__n28243;
  assign new_new_n45076__ = ~new_new_n45074__ & ~new_new_n45075__;
  assign new_new_n45077__ = ~ys__n28243 & ~new_new_n45076__;
  assign new_new_n45078__ = ys__n21994 & ~ys__n28243;
  assign new_new_n45079__ = ys__n22314 & ys__n28243;
  assign new_new_n45080__ = ~new_new_n45078__ & ~new_new_n45079__;
  assign new_new_n45081__ = ys__n28243 & ~new_new_n45080__;
  assign new_new_n45082__ = ~new_new_n45077__ & ~new_new_n45081__;
  assign new_new_n45083__ = ys__n28243 & ~new_new_n45082__;
  assign new_new_n45084__ = ~new_new_n45073__ & ~new_new_n45083__;
  assign new_new_n45085__ = new_new_n44813__ & ~new_new_n45084__;
  assign new_new_n45086__ = ys__n47798 & new_new_n44817__;
  assign new_new_n45087__ = ~new_new_n45085__ & ~new_new_n45086__;
  assign new_new_n45088__ = ~new_new_n45068__ & new_new_n45087__;
  assign new_new_n45089__ = ~new_new_n45067__ & new_new_n45088__;
  assign new_new_n45090__ = ~new_new_n45066__ & new_new_n45089__;
  assign ys__n32131 = ~new_new_n44845__ & ~new_new_n45090__;
  assign new_new_n45092__ = ~new_new_n22623__ & ~new_new_n37517__;
  assign new_new_n45093__ = ~new_new_n22932__ & ~new_new_n45092__;
  assign new_new_n45094__ = ~new_new_n44779__ & ~new_new_n45093__;
  assign new_new_n45095__ = ys__n27768 & new_new_n44779__;
  assign new_new_n45096__ = ~new_new_n45094__ & ~new_new_n45095__;
  assign new_new_n45097__ = new_new_n44788__ & ~new_new_n45096__;
  assign new_new_n45098__ = ys__n19902 & new_new_n44792__;
  assign new_new_n45099__ = ys__n47767 & new_new_n44823__;
  assign new_new_n45100__ = ys__n20972 & ~ys__n28243;
  assign new_new_n45101__ = ys__n21292 & ys__n28243;
  assign new_new_n45102__ = ~new_new_n45100__ & ~new_new_n45101__;
  assign new_new_n45103__ = ys__n28243 & ~new_new_n45102__;
  assign new_new_n45104__ = ~ys__n28243 & new_new_n45103__;
  assign new_new_n45105__ = ys__n21516 & ~ys__n28243;
  assign new_new_n45106__ = ys__n21836 & ys__n28243;
  assign new_new_n45107__ = ~new_new_n45105__ & ~new_new_n45106__;
  assign new_new_n45108__ = ~ys__n28243 & ~new_new_n45107__;
  assign new_new_n45109__ = ys__n21996 & ~ys__n28243;
  assign new_new_n45110__ = ys__n22316 & ys__n28243;
  assign new_new_n45111__ = ~new_new_n45109__ & ~new_new_n45110__;
  assign new_new_n45112__ = ys__n28243 & ~new_new_n45111__;
  assign new_new_n45113__ = ~new_new_n45108__ & ~new_new_n45112__;
  assign new_new_n45114__ = ys__n28243 & ~new_new_n45113__;
  assign new_new_n45115__ = ~new_new_n45104__ & ~new_new_n45114__;
  assign new_new_n45116__ = new_new_n44813__ & ~new_new_n45115__;
  assign new_new_n45117__ = ys__n47799 & new_new_n44817__;
  assign new_new_n45118__ = ~new_new_n45116__ & ~new_new_n45117__;
  assign new_new_n45119__ = ~new_new_n45099__ & new_new_n45118__;
  assign new_new_n45120__ = ~new_new_n45098__ & new_new_n45119__;
  assign new_new_n45121__ = ~new_new_n45097__ & new_new_n45120__;
  assign ys__n32132 = ~new_new_n44845__ & ~new_new_n45121__;
  assign new_new_n45123__ = ~new_new_n22623__ & ~new_new_n37525__;
  assign new_new_n45124__ = ~new_new_n22950__ & ~new_new_n45123__;
  assign new_new_n45125__ = ~new_new_n44779__ & ~new_new_n45124__;
  assign new_new_n45126__ = ys__n27771 & new_new_n44779__;
  assign new_new_n45127__ = ~new_new_n45125__ & ~new_new_n45126__;
  assign new_new_n45128__ = new_new_n44788__ & ~new_new_n45127__;
  assign new_new_n45129__ = ys__n19905 & new_new_n44792__;
  assign new_new_n45130__ = ys__n47768 & new_new_n44823__;
  assign new_new_n45131__ = ys__n20974 & ~ys__n28243;
  assign new_new_n45132__ = ys__n21294 & ys__n28243;
  assign new_new_n45133__ = ~new_new_n45131__ & ~new_new_n45132__;
  assign new_new_n45134__ = ys__n28243 & ~new_new_n45133__;
  assign new_new_n45135__ = ~ys__n28243 & new_new_n45134__;
  assign new_new_n45136__ = ys__n21518 & ~ys__n28243;
  assign new_new_n45137__ = ys__n21838 & ys__n28243;
  assign new_new_n45138__ = ~new_new_n45136__ & ~new_new_n45137__;
  assign new_new_n45139__ = ~ys__n28243 & ~new_new_n45138__;
  assign new_new_n45140__ = ys__n21998 & ~ys__n28243;
  assign new_new_n45141__ = ys__n22318 & ys__n28243;
  assign new_new_n45142__ = ~new_new_n45140__ & ~new_new_n45141__;
  assign new_new_n45143__ = ys__n28243 & ~new_new_n45142__;
  assign new_new_n45144__ = ~new_new_n45139__ & ~new_new_n45143__;
  assign new_new_n45145__ = ys__n28243 & ~new_new_n45144__;
  assign new_new_n45146__ = ~new_new_n45135__ & ~new_new_n45145__;
  assign new_new_n45147__ = new_new_n44813__ & ~new_new_n45146__;
  assign new_new_n45148__ = ys__n47800 & new_new_n44817__;
  assign new_new_n45149__ = ~new_new_n45147__ & ~new_new_n45148__;
  assign new_new_n45150__ = ~new_new_n45130__ & new_new_n45149__;
  assign new_new_n45151__ = ~new_new_n45129__ & new_new_n45150__;
  assign new_new_n45152__ = ~new_new_n45128__ & new_new_n45151__;
  assign ys__n32133 = ~new_new_n44845__ & ~new_new_n45152__;
  assign new_new_n45154__ = ~new_new_n22623__ & ~new_new_n37533__;
  assign new_new_n45155__ = ~new_new_n22968__ & ~new_new_n45154__;
  assign new_new_n45156__ = ~new_new_n44779__ & ~new_new_n45155__;
  assign new_new_n45157__ = ys__n27774 & new_new_n44779__;
  assign new_new_n45158__ = ~new_new_n45156__ & ~new_new_n45157__;
  assign new_new_n45159__ = new_new_n44788__ & ~new_new_n45158__;
  assign new_new_n45160__ = ys__n19908 & new_new_n44792__;
  assign new_new_n45161__ = ys__n47769 & new_new_n44823__;
  assign new_new_n45162__ = ys__n20976 & ~ys__n28243;
  assign new_new_n45163__ = ys__n21296 & ys__n28243;
  assign new_new_n45164__ = ~new_new_n45162__ & ~new_new_n45163__;
  assign new_new_n45165__ = ys__n28243 & ~new_new_n45164__;
  assign new_new_n45166__ = ~ys__n28243 & new_new_n45165__;
  assign new_new_n45167__ = ys__n21520 & ~ys__n28243;
  assign new_new_n45168__ = ys__n21840 & ys__n28243;
  assign new_new_n45169__ = ~new_new_n45167__ & ~new_new_n45168__;
  assign new_new_n45170__ = ~ys__n28243 & ~new_new_n45169__;
  assign new_new_n45171__ = ys__n22000 & ~ys__n28243;
  assign new_new_n45172__ = ys__n22320 & ys__n28243;
  assign new_new_n45173__ = ~new_new_n45171__ & ~new_new_n45172__;
  assign new_new_n45174__ = ys__n28243 & ~new_new_n45173__;
  assign new_new_n45175__ = ~new_new_n45170__ & ~new_new_n45174__;
  assign new_new_n45176__ = ys__n28243 & ~new_new_n45175__;
  assign new_new_n45177__ = ~new_new_n45166__ & ~new_new_n45176__;
  assign new_new_n45178__ = new_new_n44813__ & ~new_new_n45177__;
  assign new_new_n45179__ = ys__n47801 & new_new_n44817__;
  assign new_new_n45180__ = ~new_new_n45178__ & ~new_new_n45179__;
  assign new_new_n45181__ = ~new_new_n45161__ & new_new_n45180__;
  assign new_new_n45182__ = ~new_new_n45160__ & new_new_n45181__;
  assign new_new_n45183__ = ~new_new_n45159__ & new_new_n45182__;
  assign ys__n32134 = ~new_new_n44845__ & ~new_new_n45183__;
  assign new_new_n45185__ = ~new_new_n22623__ & ~new_new_n37541__;
  assign new_new_n45186__ = ~new_new_n22986__ & ~new_new_n45185__;
  assign new_new_n45187__ = ~new_new_n44779__ & ~new_new_n45186__;
  assign new_new_n45188__ = ys__n27777 & new_new_n44779__;
  assign new_new_n45189__ = ~new_new_n45187__ & ~new_new_n45188__;
  assign new_new_n45190__ = new_new_n44788__ & ~new_new_n45189__;
  assign new_new_n45191__ = ys__n19911 & new_new_n44792__;
  assign new_new_n45192__ = ys__n47770 & new_new_n44823__;
  assign new_new_n45193__ = ys__n20978 & ~ys__n28243;
  assign new_new_n45194__ = ys__n21298 & ys__n28243;
  assign new_new_n45195__ = ~new_new_n45193__ & ~new_new_n45194__;
  assign new_new_n45196__ = ys__n28243 & ~new_new_n45195__;
  assign new_new_n45197__ = ~ys__n28243 & new_new_n45196__;
  assign new_new_n45198__ = ys__n21522 & ~ys__n28243;
  assign new_new_n45199__ = ys__n21842 & ys__n28243;
  assign new_new_n45200__ = ~new_new_n45198__ & ~new_new_n45199__;
  assign new_new_n45201__ = ~ys__n28243 & ~new_new_n45200__;
  assign new_new_n45202__ = ys__n22002 & ~ys__n28243;
  assign new_new_n45203__ = ys__n22322 & ys__n28243;
  assign new_new_n45204__ = ~new_new_n45202__ & ~new_new_n45203__;
  assign new_new_n45205__ = ys__n28243 & ~new_new_n45204__;
  assign new_new_n45206__ = ~new_new_n45201__ & ~new_new_n45205__;
  assign new_new_n45207__ = ys__n28243 & ~new_new_n45206__;
  assign new_new_n45208__ = ~new_new_n45197__ & ~new_new_n45207__;
  assign new_new_n45209__ = new_new_n44813__ & ~new_new_n45208__;
  assign new_new_n45210__ = ys__n47802 & new_new_n44817__;
  assign new_new_n45211__ = ~new_new_n45209__ & ~new_new_n45210__;
  assign new_new_n45212__ = ~new_new_n45192__ & new_new_n45211__;
  assign new_new_n45213__ = ~new_new_n45191__ & new_new_n45212__;
  assign new_new_n45214__ = ~new_new_n45190__ & new_new_n45213__;
  assign ys__n32135 = ~new_new_n44845__ & ~new_new_n45214__;
  assign new_new_n45216__ = ~new_new_n22623__ & ~new_new_n37549__;
  assign new_new_n45217__ = ~new_new_n23004__ & ~new_new_n45216__;
  assign new_new_n45218__ = ~new_new_n44779__ & ~new_new_n45217__;
  assign new_new_n45219__ = ys__n27780 & new_new_n44779__;
  assign new_new_n45220__ = ~new_new_n45218__ & ~new_new_n45219__;
  assign new_new_n45221__ = new_new_n44788__ & ~new_new_n45220__;
  assign new_new_n45222__ = ys__n19914 & new_new_n44792__;
  assign new_new_n45223__ = ys__n47771 & new_new_n44823__;
  assign new_new_n45224__ = ys__n20980 & ~ys__n28243;
  assign new_new_n45225__ = ys__n21300 & ys__n28243;
  assign new_new_n45226__ = ~new_new_n45224__ & ~new_new_n45225__;
  assign new_new_n45227__ = ys__n28243 & ~new_new_n45226__;
  assign new_new_n45228__ = ~ys__n28243 & new_new_n45227__;
  assign new_new_n45229__ = ys__n21524 & ~ys__n28243;
  assign new_new_n45230__ = ys__n21844 & ys__n28243;
  assign new_new_n45231__ = ~new_new_n45229__ & ~new_new_n45230__;
  assign new_new_n45232__ = ~ys__n28243 & ~new_new_n45231__;
  assign new_new_n45233__ = ys__n22004 & ~ys__n28243;
  assign new_new_n45234__ = ys__n22324 & ys__n28243;
  assign new_new_n45235__ = ~new_new_n45233__ & ~new_new_n45234__;
  assign new_new_n45236__ = ys__n28243 & ~new_new_n45235__;
  assign new_new_n45237__ = ~new_new_n45232__ & ~new_new_n45236__;
  assign new_new_n45238__ = ys__n28243 & ~new_new_n45237__;
  assign new_new_n45239__ = ~new_new_n45228__ & ~new_new_n45238__;
  assign new_new_n45240__ = new_new_n44813__ & ~new_new_n45239__;
  assign new_new_n45241__ = ys__n47803 & new_new_n44817__;
  assign new_new_n45242__ = ~new_new_n45240__ & ~new_new_n45241__;
  assign new_new_n45243__ = ~new_new_n45223__ & new_new_n45242__;
  assign new_new_n45244__ = ~new_new_n45222__ & new_new_n45243__;
  assign new_new_n45245__ = ~new_new_n45221__ & new_new_n45244__;
  assign ys__n32136 = ~new_new_n44845__ & ~new_new_n45245__;
  assign new_new_n45247__ = ~new_new_n22623__ & ~new_new_n37557__;
  assign new_new_n45248__ = ~new_new_n23022__ & ~new_new_n45247__;
  assign new_new_n45249__ = ~new_new_n44779__ & ~new_new_n45248__;
  assign new_new_n45250__ = ys__n27783 & new_new_n44779__;
  assign new_new_n45251__ = ~new_new_n45249__ & ~new_new_n45250__;
  assign new_new_n45252__ = new_new_n44788__ & ~new_new_n45251__;
  assign new_new_n45253__ = ys__n19917 & new_new_n44792__;
  assign new_new_n45254__ = ys__n47772 & new_new_n44823__;
  assign new_new_n45255__ = ys__n20982 & ~ys__n28243;
  assign new_new_n45256__ = ys__n21302 & ys__n28243;
  assign new_new_n45257__ = ~new_new_n45255__ & ~new_new_n45256__;
  assign new_new_n45258__ = ys__n28243 & ~new_new_n45257__;
  assign new_new_n45259__ = ~ys__n28243 & new_new_n45258__;
  assign new_new_n45260__ = ys__n21526 & ~ys__n28243;
  assign new_new_n45261__ = ys__n21846 & ys__n28243;
  assign new_new_n45262__ = ~new_new_n45260__ & ~new_new_n45261__;
  assign new_new_n45263__ = ~ys__n28243 & ~new_new_n45262__;
  assign new_new_n45264__ = ys__n22006 & ~ys__n28243;
  assign new_new_n45265__ = ys__n22326 & ys__n28243;
  assign new_new_n45266__ = ~new_new_n45264__ & ~new_new_n45265__;
  assign new_new_n45267__ = ys__n28243 & ~new_new_n45266__;
  assign new_new_n45268__ = ~new_new_n45263__ & ~new_new_n45267__;
  assign new_new_n45269__ = ys__n28243 & ~new_new_n45268__;
  assign new_new_n45270__ = ~new_new_n45259__ & ~new_new_n45269__;
  assign new_new_n45271__ = new_new_n44813__ & ~new_new_n45270__;
  assign new_new_n45272__ = ys__n47804 & new_new_n44817__;
  assign new_new_n45273__ = ~new_new_n45271__ & ~new_new_n45272__;
  assign new_new_n45274__ = ~new_new_n45254__ & new_new_n45273__;
  assign new_new_n45275__ = ~new_new_n45253__ & new_new_n45274__;
  assign new_new_n45276__ = ~new_new_n45252__ & new_new_n45275__;
  assign ys__n32137 = ~new_new_n44845__ & ~new_new_n45276__;
  assign new_new_n45278__ = ~new_new_n22623__ & ~new_new_n37565__;
  assign new_new_n45279__ = ~new_new_n23040__ & ~new_new_n45278__;
  assign new_new_n45280__ = ~new_new_n44779__ & ~new_new_n45279__;
  assign new_new_n45281__ = ys__n27786 & new_new_n44779__;
  assign new_new_n45282__ = ~new_new_n45280__ & ~new_new_n45281__;
  assign new_new_n45283__ = new_new_n44788__ & ~new_new_n45282__;
  assign new_new_n45284__ = ys__n19920 & new_new_n44792__;
  assign new_new_n45285__ = ys__n47773 & new_new_n44823__;
  assign new_new_n45286__ = ys__n20984 & ~ys__n28243;
  assign new_new_n45287__ = ys__n21304 & ys__n28243;
  assign new_new_n45288__ = ~new_new_n45286__ & ~new_new_n45287__;
  assign new_new_n45289__ = ys__n28243 & ~new_new_n45288__;
  assign new_new_n45290__ = ~ys__n28243 & new_new_n45289__;
  assign new_new_n45291__ = ys__n21528 & ~ys__n28243;
  assign new_new_n45292__ = ys__n21848 & ys__n28243;
  assign new_new_n45293__ = ~new_new_n45291__ & ~new_new_n45292__;
  assign new_new_n45294__ = ~ys__n28243 & ~new_new_n45293__;
  assign new_new_n45295__ = ys__n22008 & ~ys__n28243;
  assign new_new_n45296__ = ys__n22328 & ys__n28243;
  assign new_new_n45297__ = ~new_new_n45295__ & ~new_new_n45296__;
  assign new_new_n45298__ = ys__n28243 & ~new_new_n45297__;
  assign new_new_n45299__ = ~new_new_n45294__ & ~new_new_n45298__;
  assign new_new_n45300__ = ys__n28243 & ~new_new_n45299__;
  assign new_new_n45301__ = ~new_new_n45290__ & ~new_new_n45300__;
  assign new_new_n45302__ = new_new_n44813__ & ~new_new_n45301__;
  assign new_new_n45303__ = ys__n47805 & new_new_n44817__;
  assign new_new_n45304__ = ~new_new_n45302__ & ~new_new_n45303__;
  assign new_new_n45305__ = ~new_new_n45285__ & new_new_n45304__;
  assign new_new_n45306__ = ~new_new_n45284__ & new_new_n45305__;
  assign new_new_n45307__ = ~new_new_n45283__ & new_new_n45306__;
  assign ys__n32138 = ~new_new_n44845__ & ~new_new_n45307__;
  assign new_new_n45309__ = ~new_new_n22623__ & ~new_new_n37573__;
  assign new_new_n45310__ = ~new_new_n23058__ & ~new_new_n45309__;
  assign new_new_n45311__ = ~new_new_n44779__ & ~new_new_n45310__;
  assign new_new_n45312__ = ys__n27789 & new_new_n44779__;
  assign new_new_n45313__ = ~new_new_n45311__ & ~new_new_n45312__;
  assign new_new_n45314__ = new_new_n44788__ & ~new_new_n45313__;
  assign new_new_n45315__ = ys__n19923 & new_new_n44792__;
  assign new_new_n45316__ = ys__n47774 & new_new_n44823__;
  assign new_new_n45317__ = ys__n20986 & ~ys__n28243;
  assign new_new_n45318__ = ys__n21306 & ys__n28243;
  assign new_new_n45319__ = ~new_new_n45317__ & ~new_new_n45318__;
  assign new_new_n45320__ = ys__n28243 & ~new_new_n45319__;
  assign new_new_n45321__ = ~ys__n28243 & new_new_n45320__;
  assign new_new_n45322__ = ys__n21530 & ~ys__n28243;
  assign new_new_n45323__ = ys__n21850 & ys__n28243;
  assign new_new_n45324__ = ~new_new_n45322__ & ~new_new_n45323__;
  assign new_new_n45325__ = ~ys__n28243 & ~new_new_n45324__;
  assign new_new_n45326__ = ys__n22010 & ~ys__n28243;
  assign new_new_n45327__ = ys__n22330 & ys__n28243;
  assign new_new_n45328__ = ~new_new_n45326__ & ~new_new_n45327__;
  assign new_new_n45329__ = ys__n28243 & ~new_new_n45328__;
  assign new_new_n45330__ = ~new_new_n45325__ & ~new_new_n45329__;
  assign new_new_n45331__ = ys__n28243 & ~new_new_n45330__;
  assign new_new_n45332__ = ~new_new_n45321__ & ~new_new_n45331__;
  assign new_new_n45333__ = new_new_n44813__ & ~new_new_n45332__;
  assign new_new_n45334__ = ys__n47806 & new_new_n44817__;
  assign new_new_n45335__ = ~new_new_n45333__ & ~new_new_n45334__;
  assign new_new_n45336__ = ~new_new_n45316__ & new_new_n45335__;
  assign new_new_n45337__ = ~new_new_n45315__ & new_new_n45336__;
  assign new_new_n45338__ = ~new_new_n45314__ & new_new_n45337__;
  assign ys__n32139 = ~new_new_n44845__ & ~new_new_n45338__;
  assign new_new_n45340__ = ~new_new_n22623__ & ~new_new_n37581__;
  assign new_new_n45341__ = ~new_new_n22772__ & ~new_new_n45340__;
  assign new_new_n45342__ = ~new_new_n44779__ & ~new_new_n45341__;
  assign new_new_n45343__ = ys__n27792 & new_new_n44779__;
  assign new_new_n45344__ = ~new_new_n45342__ & ~new_new_n45343__;
  assign new_new_n45345__ = new_new_n44788__ & ~new_new_n45344__;
  assign new_new_n45346__ = ys__n19926 & new_new_n44792__;
  assign new_new_n45347__ = ys__n47775 & new_new_n44823__;
  assign new_new_n45348__ = ys__n20988 & ~ys__n28243;
  assign new_new_n45349__ = ys__n21308 & ys__n28243;
  assign new_new_n45350__ = ~new_new_n45348__ & ~new_new_n45349__;
  assign new_new_n45351__ = ys__n28243 & ~new_new_n45350__;
  assign new_new_n45352__ = ~ys__n28243 & new_new_n45351__;
  assign new_new_n45353__ = ys__n21532 & ~ys__n28243;
  assign new_new_n45354__ = ys__n21852 & ys__n28243;
  assign new_new_n45355__ = ~new_new_n45353__ & ~new_new_n45354__;
  assign new_new_n45356__ = ~ys__n28243 & ~new_new_n45355__;
  assign new_new_n45357__ = ys__n22012 & ~ys__n28243;
  assign new_new_n45358__ = ys__n22332 & ys__n28243;
  assign new_new_n45359__ = ~new_new_n45357__ & ~new_new_n45358__;
  assign new_new_n45360__ = ys__n28243 & ~new_new_n45359__;
  assign new_new_n45361__ = ~new_new_n45356__ & ~new_new_n45360__;
  assign new_new_n45362__ = ys__n28243 & ~new_new_n45361__;
  assign new_new_n45363__ = ~new_new_n45352__ & ~new_new_n45362__;
  assign new_new_n45364__ = new_new_n44813__ & ~new_new_n45363__;
  assign new_new_n45365__ = ys__n47807 & new_new_n44817__;
  assign new_new_n45366__ = ~new_new_n45364__ & ~new_new_n45365__;
  assign new_new_n45367__ = ~new_new_n45347__ & new_new_n45366__;
  assign new_new_n45368__ = ~new_new_n45346__ & new_new_n45367__;
  assign new_new_n45369__ = ~new_new_n45345__ & new_new_n45368__;
  assign ys__n32140 = ~new_new_n44845__ & ~new_new_n45369__;
  assign new_new_n45371__ = ~new_new_n22623__ & ~new_new_n37589__;
  assign new_new_n45372__ = ~new_new_n22787__ & ~new_new_n45371__;
  assign new_new_n45373__ = ~new_new_n44779__ & ~new_new_n45372__;
  assign new_new_n45374__ = ys__n27795 & new_new_n44779__;
  assign new_new_n45375__ = ~new_new_n45373__ & ~new_new_n45374__;
  assign new_new_n45376__ = new_new_n44788__ & ~new_new_n45375__;
  assign new_new_n45377__ = ys__n19929 & new_new_n44792__;
  assign new_new_n45378__ = ys__n47776 & new_new_n44823__;
  assign new_new_n45379__ = ys__n20990 & ~ys__n28243;
  assign new_new_n45380__ = ys__n21310 & ys__n28243;
  assign new_new_n45381__ = ~new_new_n45379__ & ~new_new_n45380__;
  assign new_new_n45382__ = ys__n28243 & ~new_new_n45381__;
  assign new_new_n45383__ = ~ys__n28243 & new_new_n45382__;
  assign new_new_n45384__ = ys__n21534 & ~ys__n28243;
  assign new_new_n45385__ = ys__n21854 & ys__n28243;
  assign new_new_n45386__ = ~new_new_n45384__ & ~new_new_n45385__;
  assign new_new_n45387__ = ~ys__n28243 & ~new_new_n45386__;
  assign new_new_n45388__ = ys__n22014 & ~ys__n28243;
  assign new_new_n45389__ = ys__n22334 & ys__n28243;
  assign new_new_n45390__ = ~new_new_n45388__ & ~new_new_n45389__;
  assign new_new_n45391__ = ys__n28243 & ~new_new_n45390__;
  assign new_new_n45392__ = ~new_new_n45387__ & ~new_new_n45391__;
  assign new_new_n45393__ = ys__n28243 & ~new_new_n45392__;
  assign new_new_n45394__ = ~new_new_n45383__ & ~new_new_n45393__;
  assign new_new_n45395__ = new_new_n44813__ & ~new_new_n45394__;
  assign new_new_n45396__ = ys__n47808 & new_new_n44817__;
  assign new_new_n45397__ = ~new_new_n45395__ & ~new_new_n45396__;
  assign new_new_n45398__ = ~new_new_n45378__ & new_new_n45397__;
  assign new_new_n45399__ = ~new_new_n45377__ & new_new_n45398__;
  assign new_new_n45400__ = ~new_new_n45376__ & new_new_n45399__;
  assign ys__n32141 = ~new_new_n44845__ & ~new_new_n45400__;
  assign new_new_n45402__ = ~new_new_n22623__ & ~new_new_n37597__;
  assign new_new_n45403__ = ~new_new_n22802__ & ~new_new_n45402__;
  assign new_new_n45404__ = ~new_new_n44779__ & ~new_new_n45403__;
  assign new_new_n45405__ = ys__n27798 & new_new_n44779__;
  assign new_new_n45406__ = ~new_new_n45404__ & ~new_new_n45405__;
  assign new_new_n45407__ = new_new_n44788__ & ~new_new_n45406__;
  assign new_new_n45408__ = ys__n19932 & new_new_n44792__;
  assign new_new_n45409__ = ys__n47777 & new_new_n44823__;
  assign new_new_n45410__ = ys__n20992 & ~ys__n28243;
  assign new_new_n45411__ = ys__n21312 & ys__n28243;
  assign new_new_n45412__ = ~new_new_n45410__ & ~new_new_n45411__;
  assign new_new_n45413__ = ys__n28243 & ~new_new_n45412__;
  assign new_new_n45414__ = ~ys__n28243 & new_new_n45413__;
  assign new_new_n45415__ = ys__n21536 & ~ys__n28243;
  assign new_new_n45416__ = ys__n21856 & ys__n28243;
  assign new_new_n45417__ = ~new_new_n45415__ & ~new_new_n45416__;
  assign new_new_n45418__ = ~ys__n28243 & ~new_new_n45417__;
  assign new_new_n45419__ = ys__n22016 & ~ys__n28243;
  assign new_new_n45420__ = ys__n22336 & ys__n28243;
  assign new_new_n45421__ = ~new_new_n45419__ & ~new_new_n45420__;
  assign new_new_n45422__ = ys__n28243 & ~new_new_n45421__;
  assign new_new_n45423__ = ~new_new_n45418__ & ~new_new_n45422__;
  assign new_new_n45424__ = ys__n28243 & ~new_new_n45423__;
  assign new_new_n45425__ = ~new_new_n45414__ & ~new_new_n45424__;
  assign new_new_n45426__ = new_new_n44813__ & ~new_new_n45425__;
  assign new_new_n45427__ = ys__n47809 & new_new_n44817__;
  assign new_new_n45428__ = ~new_new_n45426__ & ~new_new_n45427__;
  assign new_new_n45429__ = ~new_new_n45409__ & new_new_n45428__;
  assign new_new_n45430__ = ~new_new_n45408__ & new_new_n45429__;
  assign new_new_n45431__ = ~new_new_n45407__ & new_new_n45430__;
  assign ys__n32142 = ~new_new_n44845__ & ~new_new_n45431__;
  assign new_new_n45433__ = ~new_new_n22623__ & ~new_new_n37605__;
  assign new_new_n45434__ = ~new_new_n22817__ & ~new_new_n45433__;
  assign new_new_n45435__ = ~new_new_n44779__ & ~new_new_n45434__;
  assign new_new_n45436__ = ys__n27801 & new_new_n44779__;
  assign new_new_n45437__ = ~new_new_n45435__ & ~new_new_n45436__;
  assign new_new_n45438__ = new_new_n44788__ & ~new_new_n45437__;
  assign new_new_n45439__ = ys__n19935 & new_new_n44792__;
  assign new_new_n45440__ = ys__n47778 & new_new_n44823__;
  assign new_new_n45441__ = ys__n20994 & ~ys__n28243;
  assign new_new_n45442__ = ys__n21314 & ys__n28243;
  assign new_new_n45443__ = ~new_new_n45441__ & ~new_new_n45442__;
  assign new_new_n45444__ = ys__n28243 & ~new_new_n45443__;
  assign new_new_n45445__ = ~ys__n28243 & new_new_n45444__;
  assign new_new_n45446__ = ys__n21538 & ~ys__n28243;
  assign new_new_n45447__ = ys__n21858 & ys__n28243;
  assign new_new_n45448__ = ~new_new_n45446__ & ~new_new_n45447__;
  assign new_new_n45449__ = ~ys__n28243 & ~new_new_n45448__;
  assign new_new_n45450__ = ys__n22018 & ~ys__n28243;
  assign new_new_n45451__ = ys__n22338 & ys__n28243;
  assign new_new_n45452__ = ~new_new_n45450__ & ~new_new_n45451__;
  assign new_new_n45453__ = ys__n28243 & ~new_new_n45452__;
  assign new_new_n45454__ = ~new_new_n45449__ & ~new_new_n45453__;
  assign new_new_n45455__ = ys__n28243 & ~new_new_n45454__;
  assign new_new_n45456__ = ~new_new_n45445__ & ~new_new_n45455__;
  assign new_new_n45457__ = new_new_n44813__ & ~new_new_n45456__;
  assign new_new_n45458__ = ys__n47810 & new_new_n44817__;
  assign new_new_n45459__ = ~new_new_n45457__ & ~new_new_n45458__;
  assign new_new_n45460__ = ~new_new_n45440__ & new_new_n45459__;
  assign new_new_n45461__ = ~new_new_n45439__ & new_new_n45460__;
  assign new_new_n45462__ = ~new_new_n45438__ & new_new_n45461__;
  assign ys__n32143 = ~new_new_n44845__ & ~new_new_n45462__;
  assign new_new_n45464__ = ~new_new_n22623__ & ~new_new_n37613__;
  assign new_new_n45465__ = ~new_new_n22832__ & ~new_new_n45464__;
  assign new_new_n45466__ = ~new_new_n44779__ & ~new_new_n45465__;
  assign new_new_n45467__ = ys__n27804 & new_new_n44779__;
  assign new_new_n45468__ = ~new_new_n45466__ & ~new_new_n45467__;
  assign new_new_n45469__ = new_new_n44788__ & ~new_new_n45468__;
  assign new_new_n45470__ = ys__n19938 & new_new_n44792__;
  assign new_new_n45471__ = ys__n47779 & new_new_n44823__;
  assign new_new_n45472__ = ys__n20996 & ~ys__n28243;
  assign new_new_n45473__ = ys__n21316 & ys__n28243;
  assign new_new_n45474__ = ~new_new_n45472__ & ~new_new_n45473__;
  assign new_new_n45475__ = ys__n28243 & ~new_new_n45474__;
  assign new_new_n45476__ = ~ys__n28243 & new_new_n45475__;
  assign new_new_n45477__ = ys__n21540 & ~ys__n28243;
  assign new_new_n45478__ = ys__n21860 & ys__n28243;
  assign new_new_n45479__ = ~new_new_n45477__ & ~new_new_n45478__;
  assign new_new_n45480__ = ~ys__n28243 & ~new_new_n45479__;
  assign new_new_n45481__ = ys__n22020 & ~ys__n28243;
  assign new_new_n45482__ = ys__n22340 & ys__n28243;
  assign new_new_n45483__ = ~new_new_n45481__ & ~new_new_n45482__;
  assign new_new_n45484__ = ys__n28243 & ~new_new_n45483__;
  assign new_new_n45485__ = ~new_new_n45480__ & ~new_new_n45484__;
  assign new_new_n45486__ = ys__n28243 & ~new_new_n45485__;
  assign new_new_n45487__ = ~new_new_n45476__ & ~new_new_n45486__;
  assign new_new_n45488__ = new_new_n44813__ & ~new_new_n45487__;
  assign new_new_n45489__ = ys__n47811 & new_new_n44817__;
  assign new_new_n45490__ = ~new_new_n45488__ & ~new_new_n45489__;
  assign new_new_n45491__ = ~new_new_n45471__ & new_new_n45490__;
  assign new_new_n45492__ = ~new_new_n45470__ & new_new_n45491__;
  assign new_new_n45493__ = ~new_new_n45469__ & new_new_n45492__;
  assign ys__n32144 = ~new_new_n44845__ & ~new_new_n45493__;
  assign new_new_n45495__ = ~new_new_n22623__ & ~new_new_n37621__;
  assign new_new_n45496__ = ~new_new_n22847__ & ~new_new_n45495__;
  assign new_new_n45497__ = ~new_new_n44779__ & ~new_new_n45496__;
  assign new_new_n45498__ = ys__n27807 & new_new_n44779__;
  assign new_new_n45499__ = ~new_new_n45497__ & ~new_new_n45498__;
  assign new_new_n45500__ = new_new_n44788__ & ~new_new_n45499__;
  assign new_new_n45501__ = ys__n19941 & new_new_n44792__;
  assign new_new_n45502__ = ys__n47780 & new_new_n44823__;
  assign new_new_n45503__ = ys__n20998 & ~ys__n28243;
  assign new_new_n45504__ = ys__n21318 & ys__n28243;
  assign new_new_n45505__ = ~new_new_n45503__ & ~new_new_n45504__;
  assign new_new_n45506__ = ys__n28243 & ~new_new_n45505__;
  assign new_new_n45507__ = ~ys__n28243 & new_new_n45506__;
  assign new_new_n45508__ = ys__n21542 & ~ys__n28243;
  assign new_new_n45509__ = ys__n21862 & ys__n28243;
  assign new_new_n45510__ = ~new_new_n45508__ & ~new_new_n45509__;
  assign new_new_n45511__ = ~ys__n28243 & ~new_new_n45510__;
  assign new_new_n45512__ = ys__n22022 & ~ys__n28243;
  assign new_new_n45513__ = ys__n22342 & ys__n28243;
  assign new_new_n45514__ = ~new_new_n45512__ & ~new_new_n45513__;
  assign new_new_n45515__ = ys__n28243 & ~new_new_n45514__;
  assign new_new_n45516__ = ~new_new_n45511__ & ~new_new_n45515__;
  assign new_new_n45517__ = ys__n28243 & ~new_new_n45516__;
  assign new_new_n45518__ = ~new_new_n45507__ & ~new_new_n45517__;
  assign new_new_n45519__ = new_new_n44813__ & ~new_new_n45518__;
  assign new_new_n45520__ = ys__n47812 & new_new_n44817__;
  assign new_new_n45521__ = ~new_new_n45519__ & ~new_new_n45520__;
  assign new_new_n45522__ = ~new_new_n45502__ & new_new_n45521__;
  assign new_new_n45523__ = ~new_new_n45501__ & new_new_n45522__;
  assign new_new_n45524__ = ~new_new_n45500__ & new_new_n45523__;
  assign ys__n32145 = ~new_new_n44845__ & ~new_new_n45524__;
  assign new_new_n45526__ = ~new_new_n22623__ & ~new_new_n37629__;
  assign new_new_n45527__ = ~new_new_n22862__ & ~new_new_n45526__;
  assign new_new_n45528__ = ~new_new_n44779__ & ~new_new_n45527__;
  assign new_new_n45529__ = ys__n27810 & new_new_n44779__;
  assign new_new_n45530__ = ~new_new_n45528__ & ~new_new_n45529__;
  assign new_new_n45531__ = new_new_n44788__ & ~new_new_n45530__;
  assign new_new_n45532__ = ys__n19944 & new_new_n44792__;
  assign new_new_n45533__ = ys__n47781 & new_new_n44823__;
  assign new_new_n45534__ = ys__n21000 & ~ys__n28243;
  assign new_new_n45535__ = ys__n21320 & ys__n28243;
  assign new_new_n45536__ = ~new_new_n45534__ & ~new_new_n45535__;
  assign new_new_n45537__ = ys__n28243 & ~new_new_n45536__;
  assign new_new_n45538__ = ~ys__n28243 & new_new_n45537__;
  assign new_new_n45539__ = ys__n21544 & ~ys__n28243;
  assign new_new_n45540__ = ys__n21864 & ys__n28243;
  assign new_new_n45541__ = ~new_new_n45539__ & ~new_new_n45540__;
  assign new_new_n45542__ = ~ys__n28243 & ~new_new_n45541__;
  assign new_new_n45543__ = ys__n22024 & ~ys__n28243;
  assign new_new_n45544__ = ys__n22344 & ys__n28243;
  assign new_new_n45545__ = ~new_new_n45543__ & ~new_new_n45544__;
  assign new_new_n45546__ = ys__n28243 & ~new_new_n45545__;
  assign new_new_n45547__ = ~new_new_n45542__ & ~new_new_n45546__;
  assign new_new_n45548__ = ys__n28243 & ~new_new_n45547__;
  assign new_new_n45549__ = ~new_new_n45538__ & ~new_new_n45548__;
  assign new_new_n45550__ = new_new_n44813__ & ~new_new_n45549__;
  assign new_new_n45551__ = ys__n47813 & new_new_n44817__;
  assign new_new_n45552__ = ~new_new_n45550__ & ~new_new_n45551__;
  assign new_new_n45553__ = ~new_new_n45533__ & new_new_n45552__;
  assign new_new_n45554__ = ~new_new_n45532__ & new_new_n45553__;
  assign new_new_n45555__ = ~new_new_n45531__ & new_new_n45554__;
  assign ys__n32146 = ~new_new_n44845__ & ~new_new_n45555__;
  assign new_new_n45557__ = ys__n19947 & new_new_n44792__;
  assign new_new_n45558__ = ~new_new_n22623__ & ~new_new_n37637__;
  assign new_new_n45559__ = ~new_new_n22877__ & ~new_new_n45558__;
  assign new_new_n45560__ = ~new_new_n44779__ & ~new_new_n45559__;
  assign new_new_n45561__ = ys__n27813 & new_new_n44779__;
  assign new_new_n45562__ = ~new_new_n45560__ & ~new_new_n45561__;
  assign new_new_n45563__ = new_new_n44788__ & ~new_new_n45562__;
  assign new_new_n45564__ = ys__n47782 & new_new_n44823__;
  assign new_new_n45565__ = ys__n21002 & ~ys__n28243;
  assign new_new_n45566__ = ys__n21322 & ys__n28243;
  assign new_new_n45567__ = ~new_new_n45565__ & ~new_new_n45566__;
  assign new_new_n45568__ = ys__n28243 & ~new_new_n45567__;
  assign new_new_n45569__ = ~ys__n28243 & new_new_n45568__;
  assign new_new_n45570__ = ys__n21546 & ~ys__n28243;
  assign new_new_n45571__ = ys__n21866 & ys__n28243;
  assign new_new_n45572__ = ~new_new_n45570__ & ~new_new_n45571__;
  assign new_new_n45573__ = ~ys__n28243 & ~new_new_n45572__;
  assign new_new_n45574__ = ys__n22026 & ~ys__n28243;
  assign new_new_n45575__ = ys__n22346 & ys__n28243;
  assign new_new_n45576__ = ~new_new_n45574__ & ~new_new_n45575__;
  assign new_new_n45577__ = ys__n28243 & ~new_new_n45576__;
  assign new_new_n45578__ = ~new_new_n45573__ & ~new_new_n45577__;
  assign new_new_n45579__ = ys__n28243 & ~new_new_n45578__;
  assign new_new_n45580__ = ~new_new_n45569__ & ~new_new_n45579__;
  assign new_new_n45581__ = new_new_n44813__ & ~new_new_n45580__;
  assign new_new_n45582__ = ys__n47814 & new_new_n44817__;
  assign new_new_n45583__ = ~new_new_n45581__ & ~new_new_n45582__;
  assign new_new_n45584__ = ~new_new_n45564__ & new_new_n45583__;
  assign new_new_n45585__ = ~new_new_n45563__ & new_new_n45584__;
  assign new_new_n45586__ = ~new_new_n45557__ & new_new_n45585__;
  assign ys__n32147 = ~new_new_n44845__ & ~new_new_n45586__;
  assign new_new_n45588__ = ~new_new_n22623__ & ~new_new_n37645__;
  assign new_new_n45589__ = ~new_new_n22624__ & ~new_new_n45588__;
  assign new_new_n45590__ = ~new_new_n44779__ & ~new_new_n45589__;
  assign new_new_n45591__ = ys__n27816 & new_new_n44779__;
  assign new_new_n45592__ = ~new_new_n45590__ & ~new_new_n45591__;
  assign new_new_n45593__ = new_new_n44788__ & ~new_new_n45592__;
  assign new_new_n45594__ = ys__n19950 & new_new_n44792__;
  assign new_new_n45595__ = ys__n47783 & new_new_n44823__;
  assign new_new_n45596__ = ys__n21004 & ~ys__n28243;
  assign new_new_n45597__ = ys__n21324 & ys__n28243;
  assign new_new_n45598__ = ~new_new_n45596__ & ~new_new_n45597__;
  assign new_new_n45599__ = ys__n28243 & ~new_new_n45598__;
  assign new_new_n45600__ = ~ys__n28243 & new_new_n45599__;
  assign new_new_n45601__ = ys__n21548 & ~ys__n28243;
  assign new_new_n45602__ = ys__n21868 & ys__n28243;
  assign new_new_n45603__ = ~new_new_n45601__ & ~new_new_n45602__;
  assign new_new_n45604__ = ~ys__n28243 & ~new_new_n45603__;
  assign new_new_n45605__ = ys__n22028 & ~ys__n28243;
  assign new_new_n45606__ = ys__n22348 & ys__n28243;
  assign new_new_n45607__ = ~new_new_n45605__ & ~new_new_n45606__;
  assign new_new_n45608__ = ys__n28243 & ~new_new_n45607__;
  assign new_new_n45609__ = ~new_new_n45604__ & ~new_new_n45608__;
  assign new_new_n45610__ = ys__n28243 & ~new_new_n45609__;
  assign new_new_n45611__ = ~new_new_n45600__ & ~new_new_n45610__;
  assign new_new_n45612__ = new_new_n44813__ & ~new_new_n45611__;
  assign new_new_n45613__ = ys__n47815 & new_new_n44817__;
  assign new_new_n45614__ = ~new_new_n45612__ & ~new_new_n45613__;
  assign new_new_n45615__ = ~new_new_n45595__ & new_new_n45614__;
  assign new_new_n45616__ = ~new_new_n45594__ & new_new_n45615__;
  assign new_new_n45617__ = ~new_new_n45593__ & new_new_n45616__;
  assign ys__n32148 = ~new_new_n44845__ & ~new_new_n45617__;
  assign new_new_n45619__ = ~new_new_n22623__ & ~new_new_n37653__;
  assign new_new_n45620__ = ~new_new_n22639__ & ~new_new_n45619__;
  assign new_new_n45621__ = ~new_new_n44779__ & ~new_new_n45620__;
  assign new_new_n45622__ = ys__n27819 & new_new_n44779__;
  assign new_new_n45623__ = ~new_new_n45621__ & ~new_new_n45622__;
  assign new_new_n45624__ = new_new_n44788__ & ~new_new_n45623__;
  assign new_new_n45625__ = ys__n19953 & new_new_n44792__;
  assign new_new_n45626__ = ys__n47784 & new_new_n44823__;
  assign new_new_n45627__ = ys__n21006 & ~ys__n28243;
  assign new_new_n45628__ = ys__n21326 & ys__n28243;
  assign new_new_n45629__ = ~new_new_n45627__ & ~new_new_n45628__;
  assign new_new_n45630__ = ys__n28243 & ~new_new_n45629__;
  assign new_new_n45631__ = ~ys__n28243 & new_new_n45630__;
  assign new_new_n45632__ = ys__n21550 & ~ys__n28243;
  assign new_new_n45633__ = ys__n21870 & ys__n28243;
  assign new_new_n45634__ = ~new_new_n45632__ & ~new_new_n45633__;
  assign new_new_n45635__ = ~ys__n28243 & ~new_new_n45634__;
  assign new_new_n45636__ = ys__n22030 & ~ys__n28243;
  assign new_new_n45637__ = ys__n22350 & ys__n28243;
  assign new_new_n45638__ = ~new_new_n45636__ & ~new_new_n45637__;
  assign new_new_n45639__ = ys__n28243 & ~new_new_n45638__;
  assign new_new_n45640__ = ~new_new_n45635__ & ~new_new_n45639__;
  assign new_new_n45641__ = ys__n28243 & ~new_new_n45640__;
  assign new_new_n45642__ = ~new_new_n45631__ & ~new_new_n45641__;
  assign new_new_n45643__ = new_new_n44813__ & ~new_new_n45642__;
  assign new_new_n45644__ = ys__n47816 & new_new_n44817__;
  assign new_new_n45645__ = ~new_new_n45643__ & ~new_new_n45644__;
  assign new_new_n45646__ = ~new_new_n45626__ & new_new_n45645__;
  assign new_new_n45647__ = ~new_new_n45625__ & new_new_n45646__;
  assign new_new_n45648__ = ~new_new_n45624__ & new_new_n45647__;
  assign ys__n32149 = ~new_new_n44845__ & ~new_new_n45648__;
  assign new_new_n45650__ = ~new_new_n22623__ & ~new_new_n37661__;
  assign new_new_n45651__ = ~new_new_n22654__ & ~new_new_n45650__;
  assign new_new_n45652__ = ~new_new_n44779__ & ~new_new_n45651__;
  assign new_new_n45653__ = ys__n27822 & new_new_n44779__;
  assign new_new_n45654__ = ~new_new_n45652__ & ~new_new_n45653__;
  assign new_new_n45655__ = new_new_n44788__ & ~new_new_n45654__;
  assign new_new_n45656__ = ys__n19956 & new_new_n44792__;
  assign new_new_n45657__ = ys__n47785 & new_new_n44823__;
  assign new_new_n45658__ = ys__n21008 & ~ys__n28243;
  assign new_new_n45659__ = ys__n21328 & ys__n28243;
  assign new_new_n45660__ = ~new_new_n45658__ & ~new_new_n45659__;
  assign new_new_n45661__ = ys__n28243 & ~new_new_n45660__;
  assign new_new_n45662__ = ~ys__n28243 & new_new_n45661__;
  assign new_new_n45663__ = ys__n21552 & ~ys__n28243;
  assign new_new_n45664__ = ys__n21872 & ys__n28243;
  assign new_new_n45665__ = ~new_new_n45663__ & ~new_new_n45664__;
  assign new_new_n45666__ = ~ys__n28243 & ~new_new_n45665__;
  assign new_new_n45667__ = ys__n22032 & ~ys__n28243;
  assign new_new_n45668__ = ys__n22352 & ys__n28243;
  assign new_new_n45669__ = ~new_new_n45667__ & ~new_new_n45668__;
  assign new_new_n45670__ = ys__n28243 & ~new_new_n45669__;
  assign new_new_n45671__ = ~new_new_n45666__ & ~new_new_n45670__;
  assign new_new_n45672__ = ys__n28243 & ~new_new_n45671__;
  assign new_new_n45673__ = ~new_new_n45662__ & ~new_new_n45672__;
  assign new_new_n45674__ = new_new_n44813__ & ~new_new_n45673__;
  assign new_new_n45675__ = ys__n47817 & new_new_n44817__;
  assign new_new_n45676__ = ~new_new_n45674__ & ~new_new_n45675__;
  assign new_new_n45677__ = ~new_new_n45657__ & new_new_n45676__;
  assign new_new_n45678__ = ~new_new_n45656__ & new_new_n45677__;
  assign new_new_n45679__ = ~new_new_n45655__ & new_new_n45678__;
  assign ys__n32150 = ~new_new_n44845__ & ~new_new_n45679__;
  assign new_new_n45681__ = ys__n19959 & new_new_n44792__;
  assign new_new_n45682__ = ~new_new_n22623__ & ~new_new_n37669__;
  assign new_new_n45683__ = ~new_new_n22669__ & ~new_new_n45682__;
  assign new_new_n45684__ = ~new_new_n44779__ & ~new_new_n45683__;
  assign new_new_n45685__ = ys__n27825 & new_new_n44779__;
  assign new_new_n45686__ = ~new_new_n45684__ & ~new_new_n45685__;
  assign new_new_n45687__ = new_new_n44788__ & ~new_new_n45686__;
  assign new_new_n45688__ = ys__n47786 & new_new_n44823__;
  assign new_new_n45689__ = ys__n21010 & ~ys__n28243;
  assign new_new_n45690__ = ys__n21330 & ys__n28243;
  assign new_new_n45691__ = ~new_new_n45689__ & ~new_new_n45690__;
  assign new_new_n45692__ = ys__n28243 & ~new_new_n45691__;
  assign new_new_n45693__ = ~ys__n28243 & new_new_n45692__;
  assign new_new_n45694__ = ys__n21554 & ~ys__n28243;
  assign new_new_n45695__ = ys__n21874 & ys__n28243;
  assign new_new_n45696__ = ~new_new_n45694__ & ~new_new_n45695__;
  assign new_new_n45697__ = ~ys__n28243 & ~new_new_n45696__;
  assign new_new_n45698__ = ys__n22034 & ~ys__n28243;
  assign new_new_n45699__ = ys__n22354 & ys__n28243;
  assign new_new_n45700__ = ~new_new_n45698__ & ~new_new_n45699__;
  assign new_new_n45701__ = ys__n28243 & ~new_new_n45700__;
  assign new_new_n45702__ = ~new_new_n45697__ & ~new_new_n45701__;
  assign new_new_n45703__ = ys__n28243 & ~new_new_n45702__;
  assign new_new_n45704__ = ~new_new_n45693__ & ~new_new_n45703__;
  assign new_new_n45705__ = new_new_n44813__ & ~new_new_n45704__;
  assign new_new_n45706__ = ys__n47818 & new_new_n44817__;
  assign new_new_n45707__ = ~new_new_n45705__ & ~new_new_n45706__;
  assign new_new_n45708__ = ~new_new_n45688__ & new_new_n45707__;
  assign new_new_n45709__ = ~new_new_n45687__ & new_new_n45708__;
  assign new_new_n45710__ = ~new_new_n45681__ & new_new_n45709__;
  assign ys__n32151 = ~new_new_n44845__ & ~new_new_n45710__;
  assign new_new_n45712__ = ~new_new_n22623__ & ~new_new_n37677__;
  assign new_new_n45713__ = ~new_new_n22684__ & ~new_new_n45712__;
  assign new_new_n45714__ = ~new_new_n44779__ & ~new_new_n45713__;
  assign new_new_n45715__ = ys__n27828 & new_new_n44779__;
  assign new_new_n45716__ = ~new_new_n45714__ & ~new_new_n45715__;
  assign new_new_n45717__ = new_new_n44788__ & ~new_new_n45716__;
  assign new_new_n45718__ = ys__n19962 & new_new_n44792__;
  assign new_new_n45719__ = ys__n47787 & new_new_n44823__;
  assign new_new_n45720__ = ys__n21012 & ~ys__n28243;
  assign new_new_n45721__ = ys__n21332 & ys__n28243;
  assign new_new_n45722__ = ~new_new_n45720__ & ~new_new_n45721__;
  assign new_new_n45723__ = ys__n28243 & ~new_new_n45722__;
  assign new_new_n45724__ = ~ys__n28243 & new_new_n45723__;
  assign new_new_n45725__ = ys__n21556 & ~ys__n28243;
  assign new_new_n45726__ = ys__n21876 & ys__n28243;
  assign new_new_n45727__ = ~new_new_n45725__ & ~new_new_n45726__;
  assign new_new_n45728__ = ~ys__n28243 & ~new_new_n45727__;
  assign new_new_n45729__ = ys__n22036 & ~ys__n28243;
  assign new_new_n45730__ = ys__n22356 & ys__n28243;
  assign new_new_n45731__ = ~new_new_n45729__ & ~new_new_n45730__;
  assign new_new_n45732__ = ys__n28243 & ~new_new_n45731__;
  assign new_new_n45733__ = ~new_new_n45728__ & ~new_new_n45732__;
  assign new_new_n45734__ = ys__n28243 & ~new_new_n45733__;
  assign new_new_n45735__ = ~new_new_n45724__ & ~new_new_n45734__;
  assign new_new_n45736__ = new_new_n44813__ & ~new_new_n45735__;
  assign new_new_n45737__ = ys__n47819 & new_new_n44817__;
  assign new_new_n45738__ = ~new_new_n45736__ & ~new_new_n45737__;
  assign new_new_n45739__ = ~new_new_n45719__ & new_new_n45738__;
  assign new_new_n45740__ = ~new_new_n45718__ & new_new_n45739__;
  assign new_new_n45741__ = ~new_new_n45717__ & new_new_n45740__;
  assign ys__n32152 = ~new_new_n44845__ & ~new_new_n45741__;
  assign new_new_n45743__ = ys__n19965 & new_new_n44792__;
  assign new_new_n45744__ = ~new_new_n22623__ & ~new_new_n37685__;
  assign new_new_n45745__ = ~new_new_n22699__ & ~new_new_n45744__;
  assign new_new_n45746__ = ~new_new_n44779__ & ~new_new_n45745__;
  assign new_new_n45747__ = ys__n27831 & new_new_n44779__;
  assign new_new_n45748__ = ~new_new_n45746__ & ~new_new_n45747__;
  assign new_new_n45749__ = new_new_n44788__ & ~new_new_n45748__;
  assign new_new_n45750__ = ys__n47788 & new_new_n44823__;
  assign new_new_n45751__ = ys__n21014 & ~ys__n28243;
  assign new_new_n45752__ = ys__n21334 & ys__n28243;
  assign new_new_n45753__ = ~new_new_n45751__ & ~new_new_n45752__;
  assign new_new_n45754__ = ys__n28243 & ~new_new_n45753__;
  assign new_new_n45755__ = ~ys__n28243 & new_new_n45754__;
  assign new_new_n45756__ = ys__n21558 & ~ys__n28243;
  assign new_new_n45757__ = ys__n21878 & ys__n28243;
  assign new_new_n45758__ = ~new_new_n45756__ & ~new_new_n45757__;
  assign new_new_n45759__ = ~ys__n28243 & ~new_new_n45758__;
  assign new_new_n45760__ = ys__n22038 & ~ys__n28243;
  assign new_new_n45761__ = ys__n22358 & ys__n28243;
  assign new_new_n45762__ = ~new_new_n45760__ & ~new_new_n45761__;
  assign new_new_n45763__ = ys__n28243 & ~new_new_n45762__;
  assign new_new_n45764__ = ~new_new_n45759__ & ~new_new_n45763__;
  assign new_new_n45765__ = ys__n28243 & ~new_new_n45764__;
  assign new_new_n45766__ = ~new_new_n45755__ & ~new_new_n45765__;
  assign new_new_n45767__ = new_new_n44813__ & ~new_new_n45766__;
  assign new_new_n45768__ = ys__n47820 & new_new_n44817__;
  assign new_new_n45769__ = ~new_new_n45767__ & ~new_new_n45768__;
  assign new_new_n45770__ = ~new_new_n45750__ & new_new_n45769__;
  assign new_new_n45771__ = ~new_new_n45749__ & new_new_n45770__;
  assign new_new_n45772__ = ~new_new_n45743__ & new_new_n45771__;
  assign ys__n32153 = ~new_new_n44845__ & ~new_new_n45772__;
  assign new_new_n45774__ = ys__n19968 & new_new_n44792__;
  assign new_new_n45775__ = ~new_new_n22623__ & ~new_new_n37693__;
  assign new_new_n45776__ = ~new_new_n22714__ & ~new_new_n45775__;
  assign new_new_n45777__ = ~new_new_n44779__ & ~new_new_n45776__;
  assign new_new_n45778__ = ys__n27834 & new_new_n44779__;
  assign new_new_n45779__ = ~new_new_n45777__ & ~new_new_n45778__;
  assign new_new_n45780__ = new_new_n44788__ & ~new_new_n45779__;
  assign new_new_n45781__ = ys__n47789 & new_new_n44823__;
  assign new_new_n45782__ = ys__n21016 & ~ys__n28243;
  assign new_new_n45783__ = ys__n21336 & ys__n28243;
  assign new_new_n45784__ = ~new_new_n45782__ & ~new_new_n45783__;
  assign new_new_n45785__ = ys__n28243 & ~new_new_n45784__;
  assign new_new_n45786__ = ~ys__n28243 & new_new_n45785__;
  assign new_new_n45787__ = ys__n21560 & ~ys__n28243;
  assign new_new_n45788__ = ys__n21880 & ys__n28243;
  assign new_new_n45789__ = ~new_new_n45787__ & ~new_new_n45788__;
  assign new_new_n45790__ = ~ys__n28243 & ~new_new_n45789__;
  assign new_new_n45791__ = ys__n22040 & ~ys__n28243;
  assign new_new_n45792__ = ys__n22360 & ys__n28243;
  assign new_new_n45793__ = ~new_new_n45791__ & ~new_new_n45792__;
  assign new_new_n45794__ = ys__n28243 & ~new_new_n45793__;
  assign new_new_n45795__ = ~new_new_n45790__ & ~new_new_n45794__;
  assign new_new_n45796__ = ys__n28243 & ~new_new_n45795__;
  assign new_new_n45797__ = ~new_new_n45786__ & ~new_new_n45796__;
  assign new_new_n45798__ = new_new_n44813__ & ~new_new_n45797__;
  assign new_new_n45799__ = ys__n47821 & new_new_n44817__;
  assign new_new_n45800__ = ~new_new_n45798__ & ~new_new_n45799__;
  assign new_new_n45801__ = ~new_new_n45781__ & new_new_n45800__;
  assign new_new_n45802__ = ~new_new_n45780__ & new_new_n45801__;
  assign new_new_n45803__ = ~new_new_n45774__ & new_new_n45802__;
  assign ys__n32154 = ~new_new_n44845__ & ~new_new_n45803__;
  assign new_new_n45805__ = ys__n19971 & new_new_n44792__;
  assign new_new_n45806__ = ~new_new_n22623__ & ~new_new_n37701__;
  assign new_new_n45807__ = ~new_new_n22729__ & ~new_new_n45806__;
  assign new_new_n45808__ = ~new_new_n44779__ & ~new_new_n45807__;
  assign new_new_n45809__ = ys__n27837 & new_new_n44779__;
  assign new_new_n45810__ = ~new_new_n45808__ & ~new_new_n45809__;
  assign new_new_n45811__ = new_new_n44788__ & ~new_new_n45810__;
  assign new_new_n45812__ = ys__n47790 & new_new_n44823__;
  assign new_new_n45813__ = ys__n21018 & ~ys__n28243;
  assign new_new_n45814__ = ys__n21338 & ys__n28243;
  assign new_new_n45815__ = ~new_new_n45813__ & ~new_new_n45814__;
  assign new_new_n45816__ = ys__n28243 & ~new_new_n45815__;
  assign new_new_n45817__ = ~ys__n28243 & new_new_n45816__;
  assign new_new_n45818__ = ys__n21562 & ~ys__n28243;
  assign new_new_n45819__ = ys__n21882 & ys__n28243;
  assign new_new_n45820__ = ~new_new_n45818__ & ~new_new_n45819__;
  assign new_new_n45821__ = ~ys__n28243 & ~new_new_n45820__;
  assign new_new_n45822__ = ys__n22042 & ~ys__n28243;
  assign new_new_n45823__ = ys__n22362 & ys__n28243;
  assign new_new_n45824__ = ~new_new_n45822__ & ~new_new_n45823__;
  assign new_new_n45825__ = ys__n28243 & ~new_new_n45824__;
  assign new_new_n45826__ = ~new_new_n45821__ & ~new_new_n45825__;
  assign new_new_n45827__ = ys__n28243 & ~new_new_n45826__;
  assign new_new_n45828__ = ~new_new_n45817__ & ~new_new_n45827__;
  assign new_new_n45829__ = new_new_n44813__ & ~new_new_n45828__;
  assign new_new_n45830__ = ys__n47822 & new_new_n44817__;
  assign new_new_n45831__ = ~new_new_n45829__ & ~new_new_n45830__;
  assign new_new_n45832__ = ~new_new_n45812__ & new_new_n45831__;
  assign new_new_n45833__ = ~new_new_n45811__ & new_new_n45832__;
  assign new_new_n45834__ = ~new_new_n45805__ & new_new_n45833__;
  assign ys__n32155 = ~new_new_n44845__ & ~new_new_n45834__;
  assign new_new_n45836__ = ~ys__n310 & new_new_n11708__;
  assign new_new_n45837__ = new_new_n11078__ & new_new_n45836__;
  assign ys__n32158 = ~new_new_n13966__ & new_new_n45837__;
  assign new_new_n45839__ = ys__n308 & ys__n310;
  assign new_new_n45840__ = ~new_new_n11774__ & ~new_new_n45839__;
  assign new_new_n45841__ = new_new_n11078__ & new_new_n11708__;
  assign new_new_n45842__ = ~new_new_n45840__ & new_new_n45841__;
  assign new_new_n45843__ = ~new_new_n11071__ & ~new_new_n45842__;
  assign ys__n32159 = ~new_new_n13966__ & ~new_new_n45843__;
  assign new_new_n45845__ = ys__n1301 & ~new_new_n11726__;
  assign new_new_n45846__ = ys__n47823 & new_new_n45845__;
  assign new_new_n45847__ = ~ys__n816 & new_new_n11726__;
  assign new_new_n45848__ = ~ys__n1301 & ~new_new_n11726__;
  assign new_new_n45849__ = ~new_new_n45847__ & ~new_new_n45848__;
  assign new_new_n45850__ = ys__n47857 & ~new_new_n45849__;
  assign new_new_n45851__ = ~new_new_n45846__ & ~new_new_n45850__;
  assign new_new_n45852__ = ~new_new_n45845__ & new_new_n45849__;
  assign ys__n32160 = ~new_new_n45851__ & ~new_new_n45852__;
  assign new_new_n45854__ = ys__n47824 & new_new_n45845__;
  assign new_new_n45855__ = ys__n47858 & ~new_new_n45849__;
  assign new_new_n45856__ = ~new_new_n45854__ & ~new_new_n45855__;
  assign ys__n32161 = ~new_new_n45852__ & ~new_new_n45856__;
  assign new_new_n45858__ = ys__n47825 & new_new_n45845__;
  assign new_new_n45859__ = ys__n47859 & ~new_new_n45849__;
  assign new_new_n45860__ = ~new_new_n45858__ & ~new_new_n45859__;
  assign ys__n32162 = ~new_new_n45852__ & ~new_new_n45860__;
  assign new_new_n45862__ = ys__n47826 & new_new_n45845__;
  assign new_new_n45863__ = ys__n47860 & ~new_new_n45849__;
  assign new_new_n45864__ = ~new_new_n45862__ & ~new_new_n45863__;
  assign ys__n32163 = ~new_new_n45852__ & ~new_new_n45864__;
  assign new_new_n45866__ = ys__n47827 & new_new_n45845__;
  assign new_new_n45867__ = ys__n47861 & ~new_new_n45849__;
  assign new_new_n45868__ = ~new_new_n45866__ & ~new_new_n45867__;
  assign ys__n32164 = ~new_new_n45852__ & ~new_new_n45868__;
  assign new_new_n45870__ = ys__n47828 & new_new_n45845__;
  assign new_new_n45871__ = ys__n47862 & ~new_new_n45849__;
  assign new_new_n45872__ = ~new_new_n45870__ & ~new_new_n45871__;
  assign ys__n32165 = ~new_new_n45852__ & ~new_new_n45872__;
  assign new_new_n45874__ = ys__n47829 & new_new_n45845__;
  assign new_new_n45875__ = ys__n47863 & ~new_new_n45849__;
  assign new_new_n45876__ = ~new_new_n45874__ & ~new_new_n45875__;
  assign ys__n32166 = ~new_new_n45852__ & ~new_new_n45876__;
  assign new_new_n45878__ = ys__n47830 & new_new_n45845__;
  assign new_new_n45879__ = ys__n47864 & ~new_new_n45849__;
  assign new_new_n45880__ = ~new_new_n45878__ & ~new_new_n45879__;
  assign ys__n32167 = ~new_new_n45852__ & ~new_new_n45880__;
  assign new_new_n45882__ = ys__n47831 & new_new_n45845__;
  assign new_new_n45883__ = ys__n47865 & ~new_new_n45849__;
  assign new_new_n45884__ = ~new_new_n45882__ & ~new_new_n45883__;
  assign ys__n32168 = ~new_new_n45852__ & ~new_new_n45884__;
  assign new_new_n45886__ = ys__n47832 & new_new_n45845__;
  assign new_new_n45887__ = ys__n47866 & ~new_new_n45849__;
  assign new_new_n45888__ = ~new_new_n45886__ & ~new_new_n45887__;
  assign ys__n32169 = ~new_new_n45852__ & ~new_new_n45888__;
  assign new_new_n45890__ = ys__n47833 & new_new_n45845__;
  assign new_new_n45891__ = ys__n47867 & ~new_new_n45849__;
  assign new_new_n45892__ = ~new_new_n45890__ & ~new_new_n45891__;
  assign ys__n32170 = ~new_new_n45852__ & ~new_new_n45892__;
  assign new_new_n45894__ = ys__n47834 & new_new_n45845__;
  assign new_new_n45895__ = ys__n47868 & ~new_new_n45849__;
  assign new_new_n45896__ = ~new_new_n45894__ & ~new_new_n45895__;
  assign ys__n32171 = ~new_new_n45852__ & ~new_new_n45896__;
  assign new_new_n45898__ = ys__n47835 & new_new_n45845__;
  assign new_new_n45899__ = ys__n47869 & ~new_new_n45849__;
  assign new_new_n45900__ = ~new_new_n45898__ & ~new_new_n45899__;
  assign ys__n32172 = ~new_new_n45852__ & ~new_new_n45900__;
  assign new_new_n45902__ = ys__n47836 & new_new_n45845__;
  assign new_new_n45903__ = ys__n47870 & ~new_new_n45849__;
  assign new_new_n45904__ = ~new_new_n45902__ & ~new_new_n45903__;
  assign ys__n32173 = ~new_new_n45852__ & ~new_new_n45904__;
  assign new_new_n45906__ = ys__n47837 & new_new_n45845__;
  assign new_new_n45907__ = ys__n47871 & ~new_new_n45849__;
  assign new_new_n45908__ = ~new_new_n45906__ & ~new_new_n45907__;
  assign ys__n32174 = ~new_new_n45852__ & ~new_new_n45908__;
  assign new_new_n45910__ = ys__n47838 & new_new_n45845__;
  assign new_new_n45911__ = ys__n47872 & ~new_new_n45849__;
  assign new_new_n45912__ = ~new_new_n45910__ & ~new_new_n45911__;
  assign ys__n32175 = ~new_new_n45852__ & ~new_new_n45912__;
  assign new_new_n45914__ = ys__n47839 & new_new_n45845__;
  assign new_new_n45915__ = ys__n47873 & ~new_new_n45849__;
  assign new_new_n45916__ = ~new_new_n45914__ & ~new_new_n45915__;
  assign ys__n32176 = ~new_new_n45852__ & ~new_new_n45916__;
  assign new_new_n45918__ = ys__n47840 & new_new_n45845__;
  assign new_new_n45919__ = ys__n47874 & ~new_new_n45849__;
  assign new_new_n45920__ = ~new_new_n45918__ & ~new_new_n45919__;
  assign ys__n32177 = ~new_new_n45852__ & ~new_new_n45920__;
  assign new_new_n45922__ = ys__n47841 & new_new_n45845__;
  assign new_new_n45923__ = ys__n47875 & ~new_new_n45849__;
  assign new_new_n45924__ = ~new_new_n45922__ & ~new_new_n45923__;
  assign ys__n32178 = ~new_new_n45852__ & ~new_new_n45924__;
  assign new_new_n45926__ = ys__n47842 & new_new_n45845__;
  assign new_new_n45927__ = ys__n47876 & ~new_new_n45849__;
  assign new_new_n45928__ = ~new_new_n45926__ & ~new_new_n45927__;
  assign ys__n32179 = ~new_new_n45852__ & ~new_new_n45928__;
  assign new_new_n45930__ = ys__n47843 & new_new_n45845__;
  assign new_new_n45931__ = ys__n47877 & ~new_new_n45849__;
  assign new_new_n45932__ = ~new_new_n45930__ & ~new_new_n45931__;
  assign ys__n32180 = ~new_new_n45852__ & ~new_new_n45932__;
  assign new_new_n45934__ = ys__n47844 & new_new_n45845__;
  assign new_new_n45935__ = ys__n47878 & ~new_new_n45849__;
  assign new_new_n45936__ = ~new_new_n45934__ & ~new_new_n45935__;
  assign ys__n32181 = ~new_new_n45852__ & ~new_new_n45936__;
  assign new_new_n45938__ = ys__n47845 & new_new_n45845__;
  assign new_new_n45939__ = ys__n47879 & ~new_new_n45849__;
  assign new_new_n45940__ = ~new_new_n45938__ & ~new_new_n45939__;
  assign ys__n32182 = ~new_new_n45852__ & ~new_new_n45940__;
  assign new_new_n45942__ = ys__n47846 & new_new_n45845__;
  assign new_new_n45943__ = ys__n47880 & ~new_new_n45849__;
  assign new_new_n45944__ = ~new_new_n45942__ & ~new_new_n45943__;
  assign ys__n32183 = ~new_new_n45852__ & ~new_new_n45944__;
  assign new_new_n45946__ = ys__n47847 & new_new_n45845__;
  assign new_new_n45947__ = ys__n47881 & ~new_new_n45849__;
  assign new_new_n45948__ = ~new_new_n45946__ & ~new_new_n45947__;
  assign ys__n32184 = ~new_new_n45852__ & ~new_new_n45948__;
  assign new_new_n45950__ = ys__n47848 & new_new_n45845__;
  assign new_new_n45951__ = ys__n47882 & ~new_new_n45849__;
  assign new_new_n45952__ = ~new_new_n45950__ & ~new_new_n45951__;
  assign ys__n32185 = ~new_new_n45852__ & ~new_new_n45952__;
  assign new_new_n45954__ = ys__n47849 & new_new_n45845__;
  assign new_new_n45955__ = ys__n47883 & ~new_new_n45849__;
  assign new_new_n45956__ = ~new_new_n45954__ & ~new_new_n45955__;
  assign ys__n32186 = ~new_new_n45852__ & ~new_new_n45956__;
  assign new_new_n45958__ = ys__n47850 & new_new_n45845__;
  assign new_new_n45959__ = ys__n47884 & ~new_new_n45849__;
  assign new_new_n45960__ = ~new_new_n45958__ & ~new_new_n45959__;
  assign ys__n32187 = ~new_new_n45852__ & ~new_new_n45960__;
  assign new_new_n45962__ = ys__n47851 & new_new_n45845__;
  assign new_new_n45963__ = ys__n47885 & ~new_new_n45849__;
  assign new_new_n45964__ = ~new_new_n45962__ & ~new_new_n45963__;
  assign ys__n32188 = ~new_new_n45852__ & ~new_new_n45964__;
  assign new_new_n45966__ = ys__n47852 & new_new_n45845__;
  assign new_new_n45967__ = ys__n47886 & ~new_new_n45849__;
  assign new_new_n45968__ = ~new_new_n45966__ & ~new_new_n45967__;
  assign ys__n32189 = ~new_new_n45852__ & ~new_new_n45968__;
  assign new_new_n45970__ = ys__n47853 & new_new_n45845__;
  assign new_new_n45971__ = ys__n47887 & ~new_new_n45849__;
  assign new_new_n45972__ = ~new_new_n45970__ & ~new_new_n45971__;
  assign ys__n32190 = ~new_new_n45852__ & ~new_new_n45972__;
  assign new_new_n45974__ = ys__n47854 & new_new_n45845__;
  assign new_new_n45975__ = ys__n47888 & ~new_new_n45849__;
  assign new_new_n45976__ = ~new_new_n45974__ & ~new_new_n45975__;
  assign ys__n32191 = ~new_new_n45852__ & ~new_new_n45976__;
  assign new_new_n45978__ = ys__n47855 & new_new_n45845__;
  assign new_new_n45979__ = ys__n19215 & ~new_new_n45849__;
  assign new_new_n45980__ = ~new_new_n45978__ & ~new_new_n45979__;
  assign ys__n32192 = ~new_new_n45852__ & ~new_new_n45980__;
  assign new_new_n45982__ = ys__n47856 & new_new_n45845__;
  assign new_new_n45983__ = ys__n47889 & ~new_new_n45849__;
  assign new_new_n45984__ = ~new_new_n45982__ & ~new_new_n45983__;
  assign ys__n32193 = ~new_new_n45852__ & ~new_new_n45984__;
  assign new_new_n45986__ = ys__n816 & ~new_new_n11726__;
  assign new_new_n45987__ = ys__n47890 & new_new_n45986__;
  assign new_new_n45988__ = ~ys__n818 & new_new_n11726__;
  assign new_new_n45989__ = ~ys__n816 & ~new_new_n11726__;
  assign new_new_n45990__ = ~new_new_n45988__ & ~new_new_n45989__;
  assign new_new_n45991__ = ys__n47857 & ~new_new_n45990__;
  assign new_new_n45992__ = ~new_new_n45987__ & ~new_new_n45991__;
  assign new_new_n45993__ = ~new_new_n45986__ & new_new_n45990__;
  assign ys__n32194 = ~new_new_n45992__ & ~new_new_n45993__;
  assign new_new_n45995__ = ys__n47891 & new_new_n45986__;
  assign new_new_n45996__ = ys__n47858 & ~new_new_n45990__;
  assign new_new_n45997__ = ~new_new_n45995__ & ~new_new_n45996__;
  assign ys__n32195 = ~new_new_n45993__ & ~new_new_n45997__;
  assign new_new_n45999__ = ys__n47892 & new_new_n45986__;
  assign new_new_n46000__ = ys__n47859 & ~new_new_n45990__;
  assign new_new_n46001__ = ~new_new_n45999__ & ~new_new_n46000__;
  assign ys__n32196 = ~new_new_n45993__ & ~new_new_n46001__;
  assign new_new_n46003__ = ys__n47893 & new_new_n45986__;
  assign new_new_n46004__ = ys__n47860 & ~new_new_n45990__;
  assign new_new_n46005__ = ~new_new_n46003__ & ~new_new_n46004__;
  assign ys__n32197 = ~new_new_n45993__ & ~new_new_n46005__;
  assign new_new_n46007__ = ys__n47894 & new_new_n45986__;
  assign new_new_n46008__ = ys__n47861 & ~new_new_n45990__;
  assign new_new_n46009__ = ~new_new_n46007__ & ~new_new_n46008__;
  assign ys__n32198 = ~new_new_n45993__ & ~new_new_n46009__;
  assign new_new_n46011__ = ys__n47895 & new_new_n45986__;
  assign new_new_n46012__ = ys__n47862 & ~new_new_n45990__;
  assign new_new_n46013__ = ~new_new_n46011__ & ~new_new_n46012__;
  assign ys__n32199 = ~new_new_n45993__ & ~new_new_n46013__;
  assign new_new_n46015__ = ys__n47896 & new_new_n45986__;
  assign new_new_n46016__ = ys__n47863 & ~new_new_n45990__;
  assign new_new_n46017__ = ~new_new_n46015__ & ~new_new_n46016__;
  assign ys__n32200 = ~new_new_n45993__ & ~new_new_n46017__;
  assign new_new_n46019__ = ys__n47897 & new_new_n45986__;
  assign new_new_n46020__ = ys__n47864 & ~new_new_n45990__;
  assign new_new_n46021__ = ~new_new_n46019__ & ~new_new_n46020__;
  assign ys__n32201 = ~new_new_n45993__ & ~new_new_n46021__;
  assign new_new_n46023__ = ys__n47898 & new_new_n45986__;
  assign new_new_n46024__ = ys__n47865 & ~new_new_n45990__;
  assign new_new_n46025__ = ~new_new_n46023__ & ~new_new_n46024__;
  assign ys__n32202 = ~new_new_n45993__ & ~new_new_n46025__;
  assign new_new_n46027__ = ys__n47899 & new_new_n45986__;
  assign new_new_n46028__ = ys__n47866 & ~new_new_n45990__;
  assign new_new_n46029__ = ~new_new_n46027__ & ~new_new_n46028__;
  assign ys__n32203 = ~new_new_n45993__ & ~new_new_n46029__;
  assign new_new_n46031__ = ys__n47900 & new_new_n45986__;
  assign new_new_n46032__ = ys__n47867 & ~new_new_n45990__;
  assign new_new_n46033__ = ~new_new_n46031__ & ~new_new_n46032__;
  assign ys__n32204 = ~new_new_n45993__ & ~new_new_n46033__;
  assign new_new_n46035__ = ys__n47901 & new_new_n45986__;
  assign new_new_n46036__ = ys__n47868 & ~new_new_n45990__;
  assign new_new_n46037__ = ~new_new_n46035__ & ~new_new_n46036__;
  assign ys__n32205 = ~new_new_n45993__ & ~new_new_n46037__;
  assign new_new_n46039__ = ys__n47902 & new_new_n45986__;
  assign new_new_n46040__ = ys__n47869 & ~new_new_n45990__;
  assign new_new_n46041__ = ~new_new_n46039__ & ~new_new_n46040__;
  assign ys__n32206 = ~new_new_n45993__ & ~new_new_n46041__;
  assign new_new_n46043__ = ys__n47903 & new_new_n45986__;
  assign new_new_n46044__ = ys__n47870 & ~new_new_n45990__;
  assign new_new_n46045__ = ~new_new_n46043__ & ~new_new_n46044__;
  assign ys__n32207 = ~new_new_n45993__ & ~new_new_n46045__;
  assign new_new_n46047__ = ys__n47904 & new_new_n45986__;
  assign new_new_n46048__ = ys__n47871 & ~new_new_n45990__;
  assign new_new_n46049__ = ~new_new_n46047__ & ~new_new_n46048__;
  assign ys__n32208 = ~new_new_n45993__ & ~new_new_n46049__;
  assign new_new_n46051__ = ys__n47905 & new_new_n45986__;
  assign new_new_n46052__ = ys__n47872 & ~new_new_n45990__;
  assign new_new_n46053__ = ~new_new_n46051__ & ~new_new_n46052__;
  assign ys__n32209 = ~new_new_n45993__ & ~new_new_n46053__;
  assign new_new_n46055__ = ys__n47906 & new_new_n45986__;
  assign new_new_n46056__ = ys__n47873 & ~new_new_n45990__;
  assign new_new_n46057__ = ~new_new_n46055__ & ~new_new_n46056__;
  assign ys__n32210 = ~new_new_n45993__ & ~new_new_n46057__;
  assign new_new_n46059__ = ys__n47907 & new_new_n45986__;
  assign new_new_n46060__ = ys__n47874 & ~new_new_n45990__;
  assign new_new_n46061__ = ~new_new_n46059__ & ~new_new_n46060__;
  assign ys__n32211 = ~new_new_n45993__ & ~new_new_n46061__;
  assign new_new_n46063__ = ys__n47908 & new_new_n45986__;
  assign new_new_n46064__ = ys__n47875 & ~new_new_n45990__;
  assign new_new_n46065__ = ~new_new_n46063__ & ~new_new_n46064__;
  assign ys__n32212 = ~new_new_n45993__ & ~new_new_n46065__;
  assign new_new_n46067__ = ys__n47909 & new_new_n45986__;
  assign new_new_n46068__ = ys__n47876 & ~new_new_n45990__;
  assign new_new_n46069__ = ~new_new_n46067__ & ~new_new_n46068__;
  assign ys__n32213 = ~new_new_n45993__ & ~new_new_n46069__;
  assign new_new_n46071__ = ys__n47910 & new_new_n45986__;
  assign new_new_n46072__ = ys__n47877 & ~new_new_n45990__;
  assign new_new_n46073__ = ~new_new_n46071__ & ~new_new_n46072__;
  assign ys__n32214 = ~new_new_n45993__ & ~new_new_n46073__;
  assign new_new_n46075__ = ys__n47911 & new_new_n45986__;
  assign new_new_n46076__ = ys__n47878 & ~new_new_n45990__;
  assign new_new_n46077__ = ~new_new_n46075__ & ~new_new_n46076__;
  assign ys__n32215 = ~new_new_n45993__ & ~new_new_n46077__;
  assign new_new_n46079__ = ys__n47912 & new_new_n45986__;
  assign new_new_n46080__ = ys__n47879 & ~new_new_n45990__;
  assign new_new_n46081__ = ~new_new_n46079__ & ~new_new_n46080__;
  assign ys__n32216 = ~new_new_n45993__ & ~new_new_n46081__;
  assign new_new_n46083__ = ys__n47913 & new_new_n45986__;
  assign new_new_n46084__ = ys__n47880 & ~new_new_n45990__;
  assign new_new_n46085__ = ~new_new_n46083__ & ~new_new_n46084__;
  assign ys__n32217 = ~new_new_n45993__ & ~new_new_n46085__;
  assign new_new_n46087__ = ys__n47914 & new_new_n45986__;
  assign new_new_n46088__ = ys__n47881 & ~new_new_n45990__;
  assign new_new_n46089__ = ~new_new_n46087__ & ~new_new_n46088__;
  assign ys__n32218 = ~new_new_n45993__ & ~new_new_n46089__;
  assign new_new_n46091__ = ys__n47915 & new_new_n45986__;
  assign new_new_n46092__ = ys__n47882 & ~new_new_n45990__;
  assign new_new_n46093__ = ~new_new_n46091__ & ~new_new_n46092__;
  assign ys__n32219 = ~new_new_n45993__ & ~new_new_n46093__;
  assign new_new_n46095__ = ys__n47916 & new_new_n45986__;
  assign new_new_n46096__ = ys__n47883 & ~new_new_n45990__;
  assign new_new_n46097__ = ~new_new_n46095__ & ~new_new_n46096__;
  assign ys__n32220 = ~new_new_n45993__ & ~new_new_n46097__;
  assign new_new_n46099__ = ys__n47917 & new_new_n45986__;
  assign new_new_n46100__ = ys__n47884 & ~new_new_n45990__;
  assign new_new_n46101__ = ~new_new_n46099__ & ~new_new_n46100__;
  assign ys__n32221 = ~new_new_n45993__ & ~new_new_n46101__;
  assign new_new_n46103__ = ys__n47918 & new_new_n45986__;
  assign new_new_n46104__ = ys__n47885 & ~new_new_n45990__;
  assign new_new_n46105__ = ~new_new_n46103__ & ~new_new_n46104__;
  assign ys__n32222 = ~new_new_n45993__ & ~new_new_n46105__;
  assign new_new_n46107__ = ys__n47919 & new_new_n45986__;
  assign new_new_n46108__ = ys__n47886 & ~new_new_n45990__;
  assign new_new_n46109__ = ~new_new_n46107__ & ~new_new_n46108__;
  assign ys__n32223 = ~new_new_n45993__ & ~new_new_n46109__;
  assign new_new_n46111__ = ys__n47920 & new_new_n45986__;
  assign new_new_n46112__ = ys__n47887 & ~new_new_n45990__;
  assign new_new_n46113__ = ~new_new_n46111__ & ~new_new_n46112__;
  assign ys__n32224 = ~new_new_n45993__ & ~new_new_n46113__;
  assign new_new_n46115__ = ys__n47921 & new_new_n45986__;
  assign new_new_n46116__ = ys__n47888 & ~new_new_n45990__;
  assign new_new_n46117__ = ~new_new_n46115__ & ~new_new_n46116__;
  assign ys__n32225 = ~new_new_n45993__ & ~new_new_n46117__;
  assign new_new_n46119__ = ys__n47922 & new_new_n45986__;
  assign new_new_n46120__ = ys__n19215 & ~new_new_n45990__;
  assign new_new_n46121__ = ~new_new_n46119__ & ~new_new_n46120__;
  assign ys__n32226 = ~new_new_n45993__ & ~new_new_n46121__;
  assign new_new_n46123__ = ys__n47923 & new_new_n45986__;
  assign new_new_n46124__ = ys__n47889 & ~new_new_n45990__;
  assign new_new_n46125__ = ~new_new_n46123__ & ~new_new_n46124__;
  assign ys__n32227 = ~new_new_n45993__ & ~new_new_n46125__;
  assign new_new_n46127__ = ys__n818 & ~new_new_n11726__;
  assign new_new_n46128__ = ys__n47924 & new_new_n46127__;
  assign new_new_n46129__ = ~ys__n820 & new_new_n11726__;
  assign new_new_n46130__ = ~ys__n818 & ~new_new_n11726__;
  assign new_new_n46131__ = ~new_new_n46129__ & ~new_new_n46130__;
  assign new_new_n46132__ = ys__n47857 & ~new_new_n46131__;
  assign new_new_n46133__ = ~new_new_n46128__ & ~new_new_n46132__;
  assign new_new_n46134__ = ~new_new_n46127__ & new_new_n46131__;
  assign ys__n32228 = ~new_new_n46133__ & ~new_new_n46134__;
  assign new_new_n46136__ = ys__n47925 & new_new_n46127__;
  assign new_new_n46137__ = ys__n47858 & ~new_new_n46131__;
  assign new_new_n46138__ = ~new_new_n46136__ & ~new_new_n46137__;
  assign ys__n32229 = ~new_new_n46134__ & ~new_new_n46138__;
  assign new_new_n46140__ = ys__n47926 & new_new_n46127__;
  assign new_new_n46141__ = ys__n47859 & ~new_new_n46131__;
  assign new_new_n46142__ = ~new_new_n46140__ & ~new_new_n46141__;
  assign ys__n32230 = ~new_new_n46134__ & ~new_new_n46142__;
  assign new_new_n46144__ = ys__n47927 & new_new_n46127__;
  assign new_new_n46145__ = ys__n47860 & ~new_new_n46131__;
  assign new_new_n46146__ = ~new_new_n46144__ & ~new_new_n46145__;
  assign ys__n32231 = ~new_new_n46134__ & ~new_new_n46146__;
  assign new_new_n46148__ = ys__n47928 & new_new_n46127__;
  assign new_new_n46149__ = ys__n47861 & ~new_new_n46131__;
  assign new_new_n46150__ = ~new_new_n46148__ & ~new_new_n46149__;
  assign ys__n32232 = ~new_new_n46134__ & ~new_new_n46150__;
  assign new_new_n46152__ = ys__n47929 & new_new_n46127__;
  assign new_new_n46153__ = ys__n47862 & ~new_new_n46131__;
  assign new_new_n46154__ = ~new_new_n46152__ & ~new_new_n46153__;
  assign ys__n32233 = ~new_new_n46134__ & ~new_new_n46154__;
  assign new_new_n46156__ = ys__n47930 & new_new_n46127__;
  assign new_new_n46157__ = ys__n47863 & ~new_new_n46131__;
  assign new_new_n46158__ = ~new_new_n46156__ & ~new_new_n46157__;
  assign ys__n32234 = ~new_new_n46134__ & ~new_new_n46158__;
  assign new_new_n46160__ = ys__n47931 & new_new_n46127__;
  assign new_new_n46161__ = ys__n47864 & ~new_new_n46131__;
  assign new_new_n46162__ = ~new_new_n46160__ & ~new_new_n46161__;
  assign ys__n32235 = ~new_new_n46134__ & ~new_new_n46162__;
  assign new_new_n46164__ = ys__n47932 & new_new_n46127__;
  assign new_new_n46165__ = ys__n47865 & ~new_new_n46131__;
  assign new_new_n46166__ = ~new_new_n46164__ & ~new_new_n46165__;
  assign ys__n32236 = ~new_new_n46134__ & ~new_new_n46166__;
  assign new_new_n46168__ = ys__n47933 & new_new_n46127__;
  assign new_new_n46169__ = ys__n47866 & ~new_new_n46131__;
  assign new_new_n46170__ = ~new_new_n46168__ & ~new_new_n46169__;
  assign ys__n32237 = ~new_new_n46134__ & ~new_new_n46170__;
  assign new_new_n46172__ = ys__n47934 & new_new_n46127__;
  assign new_new_n46173__ = ys__n47867 & ~new_new_n46131__;
  assign new_new_n46174__ = ~new_new_n46172__ & ~new_new_n46173__;
  assign ys__n32238 = ~new_new_n46134__ & ~new_new_n46174__;
  assign new_new_n46176__ = ys__n47935 & new_new_n46127__;
  assign new_new_n46177__ = ys__n47868 & ~new_new_n46131__;
  assign new_new_n46178__ = ~new_new_n46176__ & ~new_new_n46177__;
  assign ys__n32239 = ~new_new_n46134__ & ~new_new_n46178__;
  assign new_new_n46180__ = ys__n47936 & new_new_n46127__;
  assign new_new_n46181__ = ys__n47869 & ~new_new_n46131__;
  assign new_new_n46182__ = ~new_new_n46180__ & ~new_new_n46181__;
  assign ys__n32240 = ~new_new_n46134__ & ~new_new_n46182__;
  assign new_new_n46184__ = ys__n47937 & new_new_n46127__;
  assign new_new_n46185__ = ys__n47870 & ~new_new_n46131__;
  assign new_new_n46186__ = ~new_new_n46184__ & ~new_new_n46185__;
  assign ys__n32241 = ~new_new_n46134__ & ~new_new_n46186__;
  assign new_new_n46188__ = ys__n47938 & new_new_n46127__;
  assign new_new_n46189__ = ys__n47871 & ~new_new_n46131__;
  assign new_new_n46190__ = ~new_new_n46188__ & ~new_new_n46189__;
  assign ys__n32242 = ~new_new_n46134__ & ~new_new_n46190__;
  assign new_new_n46192__ = ys__n47939 & new_new_n46127__;
  assign new_new_n46193__ = ys__n47872 & ~new_new_n46131__;
  assign new_new_n46194__ = ~new_new_n46192__ & ~new_new_n46193__;
  assign ys__n32243 = ~new_new_n46134__ & ~new_new_n46194__;
  assign new_new_n46196__ = ys__n47940 & new_new_n46127__;
  assign new_new_n46197__ = ys__n47873 & ~new_new_n46131__;
  assign new_new_n46198__ = ~new_new_n46196__ & ~new_new_n46197__;
  assign ys__n32244 = ~new_new_n46134__ & ~new_new_n46198__;
  assign new_new_n46200__ = ys__n47941 & new_new_n46127__;
  assign new_new_n46201__ = ys__n47874 & ~new_new_n46131__;
  assign new_new_n46202__ = ~new_new_n46200__ & ~new_new_n46201__;
  assign ys__n32245 = ~new_new_n46134__ & ~new_new_n46202__;
  assign new_new_n46204__ = ys__n47942 & new_new_n46127__;
  assign new_new_n46205__ = ys__n47875 & ~new_new_n46131__;
  assign new_new_n46206__ = ~new_new_n46204__ & ~new_new_n46205__;
  assign ys__n32246 = ~new_new_n46134__ & ~new_new_n46206__;
  assign new_new_n46208__ = ys__n47943 & new_new_n46127__;
  assign new_new_n46209__ = ys__n47876 & ~new_new_n46131__;
  assign new_new_n46210__ = ~new_new_n46208__ & ~new_new_n46209__;
  assign ys__n32247 = ~new_new_n46134__ & ~new_new_n46210__;
  assign new_new_n46212__ = ys__n47944 & new_new_n46127__;
  assign new_new_n46213__ = ys__n47877 & ~new_new_n46131__;
  assign new_new_n46214__ = ~new_new_n46212__ & ~new_new_n46213__;
  assign ys__n32248 = ~new_new_n46134__ & ~new_new_n46214__;
  assign new_new_n46216__ = ys__n47945 & new_new_n46127__;
  assign new_new_n46217__ = ys__n47878 & ~new_new_n46131__;
  assign new_new_n46218__ = ~new_new_n46216__ & ~new_new_n46217__;
  assign ys__n32249 = ~new_new_n46134__ & ~new_new_n46218__;
  assign new_new_n46220__ = ys__n47946 & new_new_n46127__;
  assign new_new_n46221__ = ys__n47879 & ~new_new_n46131__;
  assign new_new_n46222__ = ~new_new_n46220__ & ~new_new_n46221__;
  assign ys__n32250 = ~new_new_n46134__ & ~new_new_n46222__;
  assign new_new_n46224__ = ys__n47947 & new_new_n46127__;
  assign new_new_n46225__ = ys__n47880 & ~new_new_n46131__;
  assign new_new_n46226__ = ~new_new_n46224__ & ~new_new_n46225__;
  assign ys__n32251 = ~new_new_n46134__ & ~new_new_n46226__;
  assign new_new_n46228__ = ys__n47948 & new_new_n46127__;
  assign new_new_n46229__ = ys__n47881 & ~new_new_n46131__;
  assign new_new_n46230__ = ~new_new_n46228__ & ~new_new_n46229__;
  assign ys__n32252 = ~new_new_n46134__ & ~new_new_n46230__;
  assign new_new_n46232__ = ys__n47949 & new_new_n46127__;
  assign new_new_n46233__ = ys__n47882 & ~new_new_n46131__;
  assign new_new_n46234__ = ~new_new_n46232__ & ~new_new_n46233__;
  assign ys__n32253 = ~new_new_n46134__ & ~new_new_n46234__;
  assign new_new_n46236__ = ys__n47950 & new_new_n46127__;
  assign new_new_n46237__ = ys__n47883 & ~new_new_n46131__;
  assign new_new_n46238__ = ~new_new_n46236__ & ~new_new_n46237__;
  assign ys__n32254 = ~new_new_n46134__ & ~new_new_n46238__;
  assign new_new_n46240__ = ys__n47951 & new_new_n46127__;
  assign new_new_n46241__ = ys__n47884 & ~new_new_n46131__;
  assign new_new_n46242__ = ~new_new_n46240__ & ~new_new_n46241__;
  assign ys__n32255 = ~new_new_n46134__ & ~new_new_n46242__;
  assign new_new_n46244__ = ys__n47952 & new_new_n46127__;
  assign new_new_n46245__ = ys__n47885 & ~new_new_n46131__;
  assign new_new_n46246__ = ~new_new_n46244__ & ~new_new_n46245__;
  assign ys__n32256 = ~new_new_n46134__ & ~new_new_n46246__;
  assign new_new_n46248__ = ys__n47953 & new_new_n46127__;
  assign new_new_n46249__ = ys__n47886 & ~new_new_n46131__;
  assign new_new_n46250__ = ~new_new_n46248__ & ~new_new_n46249__;
  assign ys__n32257 = ~new_new_n46134__ & ~new_new_n46250__;
  assign new_new_n46252__ = ys__n47954 & new_new_n46127__;
  assign new_new_n46253__ = ys__n47887 & ~new_new_n46131__;
  assign new_new_n46254__ = ~new_new_n46252__ & ~new_new_n46253__;
  assign ys__n32258 = ~new_new_n46134__ & ~new_new_n46254__;
  assign new_new_n46256__ = ys__n47955 & new_new_n46127__;
  assign new_new_n46257__ = ys__n47888 & ~new_new_n46131__;
  assign new_new_n46258__ = ~new_new_n46256__ & ~new_new_n46257__;
  assign ys__n32259 = ~new_new_n46134__ & ~new_new_n46258__;
  assign new_new_n46260__ = ys__n47956 & new_new_n46127__;
  assign new_new_n46261__ = ys__n19215 & ~new_new_n46131__;
  assign new_new_n46262__ = ~new_new_n46260__ & ~new_new_n46261__;
  assign ys__n32260 = ~new_new_n46134__ & ~new_new_n46262__;
  assign new_new_n46264__ = ys__n47957 & new_new_n46127__;
  assign new_new_n46265__ = ys__n47889 & ~new_new_n46131__;
  assign new_new_n46266__ = ~new_new_n46264__ & ~new_new_n46265__;
  assign ys__n32261 = ~new_new_n46134__ & ~new_new_n46266__;
  assign new_new_n46268__ = ys__n820 & ~new_new_n11726__;
  assign new_new_n46269__ = ys__n47958 & new_new_n46268__;
  assign new_new_n46270__ = ~ys__n822 & new_new_n11726__;
  assign new_new_n46271__ = ~ys__n820 & ~new_new_n11726__;
  assign new_new_n46272__ = ~new_new_n46270__ & ~new_new_n46271__;
  assign new_new_n46273__ = ys__n47857 & ~new_new_n46272__;
  assign new_new_n46274__ = ~new_new_n46269__ & ~new_new_n46273__;
  assign new_new_n46275__ = ~new_new_n46268__ & new_new_n46272__;
  assign ys__n32262 = ~new_new_n46274__ & ~new_new_n46275__;
  assign new_new_n46277__ = ys__n47959 & new_new_n46268__;
  assign new_new_n46278__ = ys__n47858 & ~new_new_n46272__;
  assign new_new_n46279__ = ~new_new_n46277__ & ~new_new_n46278__;
  assign ys__n32263 = ~new_new_n46275__ & ~new_new_n46279__;
  assign new_new_n46281__ = ys__n47960 & new_new_n46268__;
  assign new_new_n46282__ = ys__n47859 & ~new_new_n46272__;
  assign new_new_n46283__ = ~new_new_n46281__ & ~new_new_n46282__;
  assign ys__n32264 = ~new_new_n46275__ & ~new_new_n46283__;
  assign new_new_n46285__ = ys__n47961 & new_new_n46268__;
  assign new_new_n46286__ = ys__n47860 & ~new_new_n46272__;
  assign new_new_n46287__ = ~new_new_n46285__ & ~new_new_n46286__;
  assign ys__n32265 = ~new_new_n46275__ & ~new_new_n46287__;
  assign new_new_n46289__ = ys__n47962 & new_new_n46268__;
  assign new_new_n46290__ = ys__n47861 & ~new_new_n46272__;
  assign new_new_n46291__ = ~new_new_n46289__ & ~new_new_n46290__;
  assign ys__n32266 = ~new_new_n46275__ & ~new_new_n46291__;
  assign new_new_n46293__ = ys__n47963 & new_new_n46268__;
  assign new_new_n46294__ = ys__n47862 & ~new_new_n46272__;
  assign new_new_n46295__ = ~new_new_n46293__ & ~new_new_n46294__;
  assign ys__n32267 = ~new_new_n46275__ & ~new_new_n46295__;
  assign new_new_n46297__ = ys__n47964 & new_new_n46268__;
  assign new_new_n46298__ = ys__n47863 & ~new_new_n46272__;
  assign new_new_n46299__ = ~new_new_n46297__ & ~new_new_n46298__;
  assign ys__n32268 = ~new_new_n46275__ & ~new_new_n46299__;
  assign new_new_n46301__ = ys__n47965 & new_new_n46268__;
  assign new_new_n46302__ = ys__n47864 & ~new_new_n46272__;
  assign new_new_n46303__ = ~new_new_n46301__ & ~new_new_n46302__;
  assign ys__n32269 = ~new_new_n46275__ & ~new_new_n46303__;
  assign new_new_n46305__ = ys__n47966 & new_new_n46268__;
  assign new_new_n46306__ = ys__n47865 & ~new_new_n46272__;
  assign new_new_n46307__ = ~new_new_n46305__ & ~new_new_n46306__;
  assign ys__n32270 = ~new_new_n46275__ & ~new_new_n46307__;
  assign new_new_n46309__ = ys__n47967 & new_new_n46268__;
  assign new_new_n46310__ = ys__n47866 & ~new_new_n46272__;
  assign new_new_n46311__ = ~new_new_n46309__ & ~new_new_n46310__;
  assign ys__n32271 = ~new_new_n46275__ & ~new_new_n46311__;
  assign new_new_n46313__ = ys__n47968 & new_new_n46268__;
  assign new_new_n46314__ = ys__n47867 & ~new_new_n46272__;
  assign new_new_n46315__ = ~new_new_n46313__ & ~new_new_n46314__;
  assign ys__n32272 = ~new_new_n46275__ & ~new_new_n46315__;
  assign new_new_n46317__ = ys__n47969 & new_new_n46268__;
  assign new_new_n46318__ = ys__n47868 & ~new_new_n46272__;
  assign new_new_n46319__ = ~new_new_n46317__ & ~new_new_n46318__;
  assign ys__n32273 = ~new_new_n46275__ & ~new_new_n46319__;
  assign new_new_n46321__ = ys__n47970 & new_new_n46268__;
  assign new_new_n46322__ = ys__n47869 & ~new_new_n46272__;
  assign new_new_n46323__ = ~new_new_n46321__ & ~new_new_n46322__;
  assign ys__n32274 = ~new_new_n46275__ & ~new_new_n46323__;
  assign new_new_n46325__ = ys__n47971 & new_new_n46268__;
  assign new_new_n46326__ = ys__n47870 & ~new_new_n46272__;
  assign new_new_n46327__ = ~new_new_n46325__ & ~new_new_n46326__;
  assign ys__n32275 = ~new_new_n46275__ & ~new_new_n46327__;
  assign new_new_n46329__ = ys__n47972 & new_new_n46268__;
  assign new_new_n46330__ = ys__n47871 & ~new_new_n46272__;
  assign new_new_n46331__ = ~new_new_n46329__ & ~new_new_n46330__;
  assign ys__n32276 = ~new_new_n46275__ & ~new_new_n46331__;
  assign new_new_n46333__ = ys__n47973 & new_new_n46268__;
  assign new_new_n46334__ = ys__n47872 & ~new_new_n46272__;
  assign new_new_n46335__ = ~new_new_n46333__ & ~new_new_n46334__;
  assign ys__n32277 = ~new_new_n46275__ & ~new_new_n46335__;
  assign new_new_n46337__ = ys__n47974 & new_new_n46268__;
  assign new_new_n46338__ = ys__n47873 & ~new_new_n46272__;
  assign new_new_n46339__ = ~new_new_n46337__ & ~new_new_n46338__;
  assign ys__n32278 = ~new_new_n46275__ & ~new_new_n46339__;
  assign new_new_n46341__ = ys__n47975 & new_new_n46268__;
  assign new_new_n46342__ = ys__n47874 & ~new_new_n46272__;
  assign new_new_n46343__ = ~new_new_n46341__ & ~new_new_n46342__;
  assign ys__n32279 = ~new_new_n46275__ & ~new_new_n46343__;
  assign new_new_n46345__ = ys__n47976 & new_new_n46268__;
  assign new_new_n46346__ = ys__n47875 & ~new_new_n46272__;
  assign new_new_n46347__ = ~new_new_n46345__ & ~new_new_n46346__;
  assign ys__n32280 = ~new_new_n46275__ & ~new_new_n46347__;
  assign new_new_n46349__ = ys__n47977 & new_new_n46268__;
  assign new_new_n46350__ = ys__n47876 & ~new_new_n46272__;
  assign new_new_n46351__ = ~new_new_n46349__ & ~new_new_n46350__;
  assign ys__n32281 = ~new_new_n46275__ & ~new_new_n46351__;
  assign new_new_n46353__ = ys__n47978 & new_new_n46268__;
  assign new_new_n46354__ = ys__n47877 & ~new_new_n46272__;
  assign new_new_n46355__ = ~new_new_n46353__ & ~new_new_n46354__;
  assign ys__n32282 = ~new_new_n46275__ & ~new_new_n46355__;
  assign new_new_n46357__ = ys__n47979 & new_new_n46268__;
  assign new_new_n46358__ = ys__n47878 & ~new_new_n46272__;
  assign new_new_n46359__ = ~new_new_n46357__ & ~new_new_n46358__;
  assign ys__n32283 = ~new_new_n46275__ & ~new_new_n46359__;
  assign new_new_n46361__ = ys__n47980 & new_new_n46268__;
  assign new_new_n46362__ = ys__n47879 & ~new_new_n46272__;
  assign new_new_n46363__ = ~new_new_n46361__ & ~new_new_n46362__;
  assign ys__n32284 = ~new_new_n46275__ & ~new_new_n46363__;
  assign new_new_n46365__ = ys__n47981 & new_new_n46268__;
  assign new_new_n46366__ = ys__n47880 & ~new_new_n46272__;
  assign new_new_n46367__ = ~new_new_n46365__ & ~new_new_n46366__;
  assign ys__n32285 = ~new_new_n46275__ & ~new_new_n46367__;
  assign new_new_n46369__ = ys__n47982 & new_new_n46268__;
  assign new_new_n46370__ = ys__n47881 & ~new_new_n46272__;
  assign new_new_n46371__ = ~new_new_n46369__ & ~new_new_n46370__;
  assign ys__n32286 = ~new_new_n46275__ & ~new_new_n46371__;
  assign new_new_n46373__ = ys__n47983 & new_new_n46268__;
  assign new_new_n46374__ = ys__n47882 & ~new_new_n46272__;
  assign new_new_n46375__ = ~new_new_n46373__ & ~new_new_n46374__;
  assign ys__n32287 = ~new_new_n46275__ & ~new_new_n46375__;
  assign new_new_n46377__ = ys__n47984 & new_new_n46268__;
  assign new_new_n46378__ = ys__n47883 & ~new_new_n46272__;
  assign new_new_n46379__ = ~new_new_n46377__ & ~new_new_n46378__;
  assign ys__n32288 = ~new_new_n46275__ & ~new_new_n46379__;
  assign new_new_n46381__ = ys__n47985 & new_new_n46268__;
  assign new_new_n46382__ = ys__n47884 & ~new_new_n46272__;
  assign new_new_n46383__ = ~new_new_n46381__ & ~new_new_n46382__;
  assign ys__n32289 = ~new_new_n46275__ & ~new_new_n46383__;
  assign new_new_n46385__ = ys__n47986 & new_new_n46268__;
  assign new_new_n46386__ = ys__n47885 & ~new_new_n46272__;
  assign new_new_n46387__ = ~new_new_n46385__ & ~new_new_n46386__;
  assign ys__n32290 = ~new_new_n46275__ & ~new_new_n46387__;
  assign new_new_n46389__ = ys__n47987 & new_new_n46268__;
  assign new_new_n46390__ = ys__n47886 & ~new_new_n46272__;
  assign new_new_n46391__ = ~new_new_n46389__ & ~new_new_n46390__;
  assign ys__n32291 = ~new_new_n46275__ & ~new_new_n46391__;
  assign new_new_n46393__ = ys__n47988 & new_new_n46268__;
  assign new_new_n46394__ = ys__n47887 & ~new_new_n46272__;
  assign new_new_n46395__ = ~new_new_n46393__ & ~new_new_n46394__;
  assign ys__n32292 = ~new_new_n46275__ & ~new_new_n46395__;
  assign new_new_n46397__ = ys__n47989 & new_new_n46268__;
  assign new_new_n46398__ = ys__n47888 & ~new_new_n46272__;
  assign new_new_n46399__ = ~new_new_n46397__ & ~new_new_n46398__;
  assign ys__n32293 = ~new_new_n46275__ & ~new_new_n46399__;
  assign new_new_n46401__ = ys__n47990 & new_new_n46268__;
  assign new_new_n46402__ = ys__n19215 & ~new_new_n46272__;
  assign new_new_n46403__ = ~new_new_n46401__ & ~new_new_n46402__;
  assign ys__n32294 = ~new_new_n46275__ & ~new_new_n46403__;
  assign new_new_n46405__ = ys__n47991 & new_new_n46268__;
  assign new_new_n46406__ = ys__n47889 & ~new_new_n46272__;
  assign new_new_n46407__ = ~new_new_n46405__ & ~new_new_n46406__;
  assign ys__n32295 = ~new_new_n46275__ & ~new_new_n46407__;
  assign new_new_n46409__ = ys__n822 & ~new_new_n11726__;
  assign new_new_n46410__ = ys__n47992 & new_new_n46409__;
  assign new_new_n46411__ = ~ys__n824 & new_new_n11726__;
  assign new_new_n46412__ = ~ys__n822 & ~new_new_n11726__;
  assign new_new_n46413__ = ~new_new_n46411__ & ~new_new_n46412__;
  assign new_new_n46414__ = ys__n47857 & ~new_new_n46413__;
  assign new_new_n46415__ = ~new_new_n46410__ & ~new_new_n46414__;
  assign new_new_n46416__ = ~new_new_n46409__ & new_new_n46413__;
  assign ys__n32296 = ~new_new_n46415__ & ~new_new_n46416__;
  assign new_new_n46418__ = ys__n47993 & new_new_n46409__;
  assign new_new_n46419__ = ys__n47858 & ~new_new_n46413__;
  assign new_new_n46420__ = ~new_new_n46418__ & ~new_new_n46419__;
  assign ys__n32297 = ~new_new_n46416__ & ~new_new_n46420__;
  assign new_new_n46422__ = ys__n47994 & new_new_n46409__;
  assign new_new_n46423__ = ys__n47859 & ~new_new_n46413__;
  assign new_new_n46424__ = ~new_new_n46422__ & ~new_new_n46423__;
  assign ys__n32298 = ~new_new_n46416__ & ~new_new_n46424__;
  assign new_new_n46426__ = ys__n47995 & new_new_n46409__;
  assign new_new_n46427__ = ys__n47860 & ~new_new_n46413__;
  assign new_new_n46428__ = ~new_new_n46426__ & ~new_new_n46427__;
  assign ys__n32299 = ~new_new_n46416__ & ~new_new_n46428__;
  assign new_new_n46430__ = ys__n47996 & new_new_n46409__;
  assign new_new_n46431__ = ys__n47861 & ~new_new_n46413__;
  assign new_new_n46432__ = ~new_new_n46430__ & ~new_new_n46431__;
  assign ys__n32300 = ~new_new_n46416__ & ~new_new_n46432__;
  assign new_new_n46434__ = ys__n47997 & new_new_n46409__;
  assign new_new_n46435__ = ys__n47862 & ~new_new_n46413__;
  assign new_new_n46436__ = ~new_new_n46434__ & ~new_new_n46435__;
  assign ys__n32301 = ~new_new_n46416__ & ~new_new_n46436__;
  assign new_new_n46438__ = ys__n47998 & new_new_n46409__;
  assign new_new_n46439__ = ys__n47863 & ~new_new_n46413__;
  assign new_new_n46440__ = ~new_new_n46438__ & ~new_new_n46439__;
  assign ys__n32302 = ~new_new_n46416__ & ~new_new_n46440__;
  assign new_new_n46442__ = ys__n47999 & new_new_n46409__;
  assign new_new_n46443__ = ys__n47864 & ~new_new_n46413__;
  assign new_new_n46444__ = ~new_new_n46442__ & ~new_new_n46443__;
  assign ys__n32303 = ~new_new_n46416__ & ~new_new_n46444__;
  assign new_new_n46446__ = ys__n48000 & new_new_n46409__;
  assign new_new_n46447__ = ys__n47865 & ~new_new_n46413__;
  assign new_new_n46448__ = ~new_new_n46446__ & ~new_new_n46447__;
  assign ys__n32304 = ~new_new_n46416__ & ~new_new_n46448__;
  assign new_new_n46450__ = ys__n48001 & new_new_n46409__;
  assign new_new_n46451__ = ys__n47866 & ~new_new_n46413__;
  assign new_new_n46452__ = ~new_new_n46450__ & ~new_new_n46451__;
  assign ys__n32305 = ~new_new_n46416__ & ~new_new_n46452__;
  assign new_new_n46454__ = ys__n48002 & new_new_n46409__;
  assign new_new_n46455__ = ys__n47867 & ~new_new_n46413__;
  assign new_new_n46456__ = ~new_new_n46454__ & ~new_new_n46455__;
  assign ys__n32306 = ~new_new_n46416__ & ~new_new_n46456__;
  assign new_new_n46458__ = ys__n48003 & new_new_n46409__;
  assign new_new_n46459__ = ys__n47868 & ~new_new_n46413__;
  assign new_new_n46460__ = ~new_new_n46458__ & ~new_new_n46459__;
  assign ys__n32307 = ~new_new_n46416__ & ~new_new_n46460__;
  assign new_new_n46462__ = ys__n48004 & new_new_n46409__;
  assign new_new_n46463__ = ys__n47869 & ~new_new_n46413__;
  assign new_new_n46464__ = ~new_new_n46462__ & ~new_new_n46463__;
  assign ys__n32308 = ~new_new_n46416__ & ~new_new_n46464__;
  assign new_new_n46466__ = ys__n48005 & new_new_n46409__;
  assign new_new_n46467__ = ys__n47870 & ~new_new_n46413__;
  assign new_new_n46468__ = ~new_new_n46466__ & ~new_new_n46467__;
  assign ys__n32309 = ~new_new_n46416__ & ~new_new_n46468__;
  assign new_new_n46470__ = ys__n48006 & new_new_n46409__;
  assign new_new_n46471__ = ys__n47871 & ~new_new_n46413__;
  assign new_new_n46472__ = ~new_new_n46470__ & ~new_new_n46471__;
  assign ys__n32310 = ~new_new_n46416__ & ~new_new_n46472__;
  assign new_new_n46474__ = ys__n48007 & new_new_n46409__;
  assign new_new_n46475__ = ys__n47872 & ~new_new_n46413__;
  assign new_new_n46476__ = ~new_new_n46474__ & ~new_new_n46475__;
  assign ys__n32311 = ~new_new_n46416__ & ~new_new_n46476__;
  assign new_new_n46478__ = ys__n48008 & new_new_n46409__;
  assign new_new_n46479__ = ys__n47873 & ~new_new_n46413__;
  assign new_new_n46480__ = ~new_new_n46478__ & ~new_new_n46479__;
  assign ys__n32312 = ~new_new_n46416__ & ~new_new_n46480__;
  assign new_new_n46482__ = ys__n48009 & new_new_n46409__;
  assign new_new_n46483__ = ys__n47874 & ~new_new_n46413__;
  assign new_new_n46484__ = ~new_new_n46482__ & ~new_new_n46483__;
  assign ys__n32313 = ~new_new_n46416__ & ~new_new_n46484__;
  assign new_new_n46486__ = ys__n48010 & new_new_n46409__;
  assign new_new_n46487__ = ys__n47875 & ~new_new_n46413__;
  assign new_new_n46488__ = ~new_new_n46486__ & ~new_new_n46487__;
  assign ys__n32314 = ~new_new_n46416__ & ~new_new_n46488__;
  assign new_new_n46490__ = ys__n48011 & new_new_n46409__;
  assign new_new_n46491__ = ys__n47876 & ~new_new_n46413__;
  assign new_new_n46492__ = ~new_new_n46490__ & ~new_new_n46491__;
  assign ys__n32315 = ~new_new_n46416__ & ~new_new_n46492__;
  assign new_new_n46494__ = ys__n48012 & new_new_n46409__;
  assign new_new_n46495__ = ys__n47877 & ~new_new_n46413__;
  assign new_new_n46496__ = ~new_new_n46494__ & ~new_new_n46495__;
  assign ys__n32316 = ~new_new_n46416__ & ~new_new_n46496__;
  assign new_new_n46498__ = ys__n48013 & new_new_n46409__;
  assign new_new_n46499__ = ys__n47878 & ~new_new_n46413__;
  assign new_new_n46500__ = ~new_new_n46498__ & ~new_new_n46499__;
  assign ys__n32317 = ~new_new_n46416__ & ~new_new_n46500__;
  assign new_new_n46502__ = ys__n48014 & new_new_n46409__;
  assign new_new_n46503__ = ys__n47879 & ~new_new_n46413__;
  assign new_new_n46504__ = ~new_new_n46502__ & ~new_new_n46503__;
  assign ys__n32318 = ~new_new_n46416__ & ~new_new_n46504__;
  assign new_new_n46506__ = ys__n48015 & new_new_n46409__;
  assign new_new_n46507__ = ys__n47880 & ~new_new_n46413__;
  assign new_new_n46508__ = ~new_new_n46506__ & ~new_new_n46507__;
  assign ys__n32319 = ~new_new_n46416__ & ~new_new_n46508__;
  assign new_new_n46510__ = ys__n48016 & new_new_n46409__;
  assign new_new_n46511__ = ys__n47881 & ~new_new_n46413__;
  assign new_new_n46512__ = ~new_new_n46510__ & ~new_new_n46511__;
  assign ys__n32320 = ~new_new_n46416__ & ~new_new_n46512__;
  assign new_new_n46514__ = ys__n48017 & new_new_n46409__;
  assign new_new_n46515__ = ys__n47882 & ~new_new_n46413__;
  assign new_new_n46516__ = ~new_new_n46514__ & ~new_new_n46515__;
  assign ys__n32321 = ~new_new_n46416__ & ~new_new_n46516__;
  assign new_new_n46518__ = ys__n48018 & new_new_n46409__;
  assign new_new_n46519__ = ys__n47883 & ~new_new_n46413__;
  assign new_new_n46520__ = ~new_new_n46518__ & ~new_new_n46519__;
  assign ys__n32322 = ~new_new_n46416__ & ~new_new_n46520__;
  assign new_new_n46522__ = ys__n48019 & new_new_n46409__;
  assign new_new_n46523__ = ys__n47884 & ~new_new_n46413__;
  assign new_new_n46524__ = ~new_new_n46522__ & ~new_new_n46523__;
  assign ys__n32323 = ~new_new_n46416__ & ~new_new_n46524__;
  assign new_new_n46526__ = ys__n48020 & new_new_n46409__;
  assign new_new_n46527__ = ys__n47885 & ~new_new_n46413__;
  assign new_new_n46528__ = ~new_new_n46526__ & ~new_new_n46527__;
  assign ys__n32324 = ~new_new_n46416__ & ~new_new_n46528__;
  assign new_new_n46530__ = ys__n48021 & new_new_n46409__;
  assign new_new_n46531__ = ys__n47886 & ~new_new_n46413__;
  assign new_new_n46532__ = ~new_new_n46530__ & ~new_new_n46531__;
  assign ys__n32325 = ~new_new_n46416__ & ~new_new_n46532__;
  assign new_new_n46534__ = ys__n48022 & new_new_n46409__;
  assign new_new_n46535__ = ys__n47887 & ~new_new_n46413__;
  assign new_new_n46536__ = ~new_new_n46534__ & ~new_new_n46535__;
  assign ys__n32326 = ~new_new_n46416__ & ~new_new_n46536__;
  assign new_new_n46538__ = ys__n48023 & new_new_n46409__;
  assign new_new_n46539__ = ys__n47888 & ~new_new_n46413__;
  assign new_new_n46540__ = ~new_new_n46538__ & ~new_new_n46539__;
  assign ys__n32327 = ~new_new_n46416__ & ~new_new_n46540__;
  assign new_new_n46542__ = ys__n48024 & new_new_n46409__;
  assign new_new_n46543__ = ys__n19215 & ~new_new_n46413__;
  assign new_new_n46544__ = ~new_new_n46542__ & ~new_new_n46543__;
  assign ys__n32328 = ~new_new_n46416__ & ~new_new_n46544__;
  assign new_new_n46546__ = ys__n48025 & new_new_n46409__;
  assign new_new_n46547__ = ys__n47889 & ~new_new_n46413__;
  assign new_new_n46548__ = ~new_new_n46546__ & ~new_new_n46547__;
  assign ys__n32329 = ~new_new_n46416__ & ~new_new_n46548__;
  assign new_new_n46550__ = ys__n824 & ~new_new_n11726__;
  assign new_new_n46551__ = ys__n48026 & new_new_n46550__;
  assign new_new_n46552__ = ~ys__n826 & new_new_n11726__;
  assign new_new_n46553__ = ~ys__n824 & ~new_new_n11726__;
  assign new_new_n46554__ = ~new_new_n46552__ & ~new_new_n46553__;
  assign new_new_n46555__ = ys__n47857 & ~new_new_n46554__;
  assign new_new_n46556__ = ~new_new_n46551__ & ~new_new_n46555__;
  assign new_new_n46557__ = ~new_new_n46550__ & new_new_n46554__;
  assign ys__n32330 = ~new_new_n46556__ & ~new_new_n46557__;
  assign new_new_n46559__ = ys__n48027 & new_new_n46550__;
  assign new_new_n46560__ = ys__n47858 & ~new_new_n46554__;
  assign new_new_n46561__ = ~new_new_n46559__ & ~new_new_n46560__;
  assign ys__n32331 = ~new_new_n46557__ & ~new_new_n46561__;
  assign new_new_n46563__ = ys__n48028 & new_new_n46550__;
  assign new_new_n46564__ = ys__n47859 & ~new_new_n46554__;
  assign new_new_n46565__ = ~new_new_n46563__ & ~new_new_n46564__;
  assign ys__n32332 = ~new_new_n46557__ & ~new_new_n46565__;
  assign new_new_n46567__ = ys__n48029 & new_new_n46550__;
  assign new_new_n46568__ = ys__n47860 & ~new_new_n46554__;
  assign new_new_n46569__ = ~new_new_n46567__ & ~new_new_n46568__;
  assign ys__n32333 = ~new_new_n46557__ & ~new_new_n46569__;
  assign new_new_n46571__ = ys__n48030 & new_new_n46550__;
  assign new_new_n46572__ = ys__n47861 & ~new_new_n46554__;
  assign new_new_n46573__ = ~new_new_n46571__ & ~new_new_n46572__;
  assign ys__n32334 = ~new_new_n46557__ & ~new_new_n46573__;
  assign new_new_n46575__ = ys__n48031 & new_new_n46550__;
  assign new_new_n46576__ = ys__n47862 & ~new_new_n46554__;
  assign new_new_n46577__ = ~new_new_n46575__ & ~new_new_n46576__;
  assign ys__n32335 = ~new_new_n46557__ & ~new_new_n46577__;
  assign new_new_n46579__ = ys__n48032 & new_new_n46550__;
  assign new_new_n46580__ = ys__n47863 & ~new_new_n46554__;
  assign new_new_n46581__ = ~new_new_n46579__ & ~new_new_n46580__;
  assign ys__n32336 = ~new_new_n46557__ & ~new_new_n46581__;
  assign new_new_n46583__ = ys__n48033 & new_new_n46550__;
  assign new_new_n46584__ = ys__n47864 & ~new_new_n46554__;
  assign new_new_n46585__ = ~new_new_n46583__ & ~new_new_n46584__;
  assign ys__n32337 = ~new_new_n46557__ & ~new_new_n46585__;
  assign new_new_n46587__ = ys__n48034 & new_new_n46550__;
  assign new_new_n46588__ = ys__n47865 & ~new_new_n46554__;
  assign new_new_n46589__ = ~new_new_n46587__ & ~new_new_n46588__;
  assign ys__n32338 = ~new_new_n46557__ & ~new_new_n46589__;
  assign new_new_n46591__ = ys__n48035 & new_new_n46550__;
  assign new_new_n46592__ = ys__n47866 & ~new_new_n46554__;
  assign new_new_n46593__ = ~new_new_n46591__ & ~new_new_n46592__;
  assign ys__n32339 = ~new_new_n46557__ & ~new_new_n46593__;
  assign new_new_n46595__ = ys__n48036 & new_new_n46550__;
  assign new_new_n46596__ = ys__n47867 & ~new_new_n46554__;
  assign new_new_n46597__ = ~new_new_n46595__ & ~new_new_n46596__;
  assign ys__n32340 = ~new_new_n46557__ & ~new_new_n46597__;
  assign new_new_n46599__ = ys__n48037 & new_new_n46550__;
  assign new_new_n46600__ = ys__n47868 & ~new_new_n46554__;
  assign new_new_n46601__ = ~new_new_n46599__ & ~new_new_n46600__;
  assign ys__n32341 = ~new_new_n46557__ & ~new_new_n46601__;
  assign new_new_n46603__ = ys__n48038 & new_new_n46550__;
  assign new_new_n46604__ = ys__n47869 & ~new_new_n46554__;
  assign new_new_n46605__ = ~new_new_n46603__ & ~new_new_n46604__;
  assign ys__n32342 = ~new_new_n46557__ & ~new_new_n46605__;
  assign new_new_n46607__ = ys__n48039 & new_new_n46550__;
  assign new_new_n46608__ = ys__n47870 & ~new_new_n46554__;
  assign new_new_n46609__ = ~new_new_n46607__ & ~new_new_n46608__;
  assign ys__n32343 = ~new_new_n46557__ & ~new_new_n46609__;
  assign new_new_n46611__ = ys__n48040 & new_new_n46550__;
  assign new_new_n46612__ = ys__n47871 & ~new_new_n46554__;
  assign new_new_n46613__ = ~new_new_n46611__ & ~new_new_n46612__;
  assign ys__n32344 = ~new_new_n46557__ & ~new_new_n46613__;
  assign new_new_n46615__ = ys__n48041 & new_new_n46550__;
  assign new_new_n46616__ = ys__n47872 & ~new_new_n46554__;
  assign new_new_n46617__ = ~new_new_n46615__ & ~new_new_n46616__;
  assign ys__n32345 = ~new_new_n46557__ & ~new_new_n46617__;
  assign new_new_n46619__ = ys__n48042 & new_new_n46550__;
  assign new_new_n46620__ = ys__n47873 & ~new_new_n46554__;
  assign new_new_n46621__ = ~new_new_n46619__ & ~new_new_n46620__;
  assign ys__n32346 = ~new_new_n46557__ & ~new_new_n46621__;
  assign new_new_n46623__ = ys__n48043 & new_new_n46550__;
  assign new_new_n46624__ = ys__n47874 & ~new_new_n46554__;
  assign new_new_n46625__ = ~new_new_n46623__ & ~new_new_n46624__;
  assign ys__n32347 = ~new_new_n46557__ & ~new_new_n46625__;
  assign new_new_n46627__ = ys__n48044 & new_new_n46550__;
  assign new_new_n46628__ = ys__n47875 & ~new_new_n46554__;
  assign new_new_n46629__ = ~new_new_n46627__ & ~new_new_n46628__;
  assign ys__n32348 = ~new_new_n46557__ & ~new_new_n46629__;
  assign new_new_n46631__ = ys__n48045 & new_new_n46550__;
  assign new_new_n46632__ = ys__n47876 & ~new_new_n46554__;
  assign new_new_n46633__ = ~new_new_n46631__ & ~new_new_n46632__;
  assign ys__n32349 = ~new_new_n46557__ & ~new_new_n46633__;
  assign new_new_n46635__ = ys__n48046 & new_new_n46550__;
  assign new_new_n46636__ = ys__n47877 & ~new_new_n46554__;
  assign new_new_n46637__ = ~new_new_n46635__ & ~new_new_n46636__;
  assign ys__n32350 = ~new_new_n46557__ & ~new_new_n46637__;
  assign new_new_n46639__ = ys__n48047 & new_new_n46550__;
  assign new_new_n46640__ = ys__n47878 & ~new_new_n46554__;
  assign new_new_n46641__ = ~new_new_n46639__ & ~new_new_n46640__;
  assign ys__n32351 = ~new_new_n46557__ & ~new_new_n46641__;
  assign new_new_n46643__ = ys__n48048 & new_new_n46550__;
  assign new_new_n46644__ = ys__n47879 & ~new_new_n46554__;
  assign new_new_n46645__ = ~new_new_n46643__ & ~new_new_n46644__;
  assign ys__n32352 = ~new_new_n46557__ & ~new_new_n46645__;
  assign new_new_n46647__ = ys__n48049 & new_new_n46550__;
  assign new_new_n46648__ = ys__n47880 & ~new_new_n46554__;
  assign new_new_n46649__ = ~new_new_n46647__ & ~new_new_n46648__;
  assign ys__n32353 = ~new_new_n46557__ & ~new_new_n46649__;
  assign new_new_n46651__ = ys__n48050 & new_new_n46550__;
  assign new_new_n46652__ = ys__n47881 & ~new_new_n46554__;
  assign new_new_n46653__ = ~new_new_n46651__ & ~new_new_n46652__;
  assign ys__n32354 = ~new_new_n46557__ & ~new_new_n46653__;
  assign new_new_n46655__ = ys__n48051 & new_new_n46550__;
  assign new_new_n46656__ = ys__n47882 & ~new_new_n46554__;
  assign new_new_n46657__ = ~new_new_n46655__ & ~new_new_n46656__;
  assign ys__n32355 = ~new_new_n46557__ & ~new_new_n46657__;
  assign new_new_n46659__ = ys__n48052 & new_new_n46550__;
  assign new_new_n46660__ = ys__n47883 & ~new_new_n46554__;
  assign new_new_n46661__ = ~new_new_n46659__ & ~new_new_n46660__;
  assign ys__n32356 = ~new_new_n46557__ & ~new_new_n46661__;
  assign new_new_n46663__ = ys__n48053 & new_new_n46550__;
  assign new_new_n46664__ = ys__n47884 & ~new_new_n46554__;
  assign new_new_n46665__ = ~new_new_n46663__ & ~new_new_n46664__;
  assign ys__n32357 = ~new_new_n46557__ & ~new_new_n46665__;
  assign new_new_n46667__ = ys__n48054 & new_new_n46550__;
  assign new_new_n46668__ = ys__n47885 & ~new_new_n46554__;
  assign new_new_n46669__ = ~new_new_n46667__ & ~new_new_n46668__;
  assign ys__n32358 = ~new_new_n46557__ & ~new_new_n46669__;
  assign new_new_n46671__ = ys__n48055 & new_new_n46550__;
  assign new_new_n46672__ = ys__n47886 & ~new_new_n46554__;
  assign new_new_n46673__ = ~new_new_n46671__ & ~new_new_n46672__;
  assign ys__n32359 = ~new_new_n46557__ & ~new_new_n46673__;
  assign new_new_n46675__ = ys__n48056 & new_new_n46550__;
  assign new_new_n46676__ = ys__n47887 & ~new_new_n46554__;
  assign new_new_n46677__ = ~new_new_n46675__ & ~new_new_n46676__;
  assign ys__n32360 = ~new_new_n46557__ & ~new_new_n46677__;
  assign new_new_n46679__ = ys__n48057 & new_new_n46550__;
  assign new_new_n46680__ = ys__n47888 & ~new_new_n46554__;
  assign new_new_n46681__ = ~new_new_n46679__ & ~new_new_n46680__;
  assign ys__n32361 = ~new_new_n46557__ & ~new_new_n46681__;
  assign new_new_n46683__ = ys__n48058 & new_new_n46550__;
  assign new_new_n46684__ = ys__n19215 & ~new_new_n46554__;
  assign new_new_n46685__ = ~new_new_n46683__ & ~new_new_n46684__;
  assign ys__n32362 = ~new_new_n46557__ & ~new_new_n46685__;
  assign new_new_n46687__ = ys__n48059 & new_new_n46550__;
  assign new_new_n46688__ = ys__n47889 & ~new_new_n46554__;
  assign new_new_n46689__ = ~new_new_n46687__ & ~new_new_n46688__;
  assign ys__n32363 = ~new_new_n46557__ & ~new_new_n46689__;
  assign new_new_n46691__ = ys__n826 & ~new_new_n11726__;
  assign new_new_n46692__ = ys__n48060 & new_new_n46691__;
  assign new_new_n46693__ = ~ys__n828 & new_new_n11726__;
  assign new_new_n46694__ = ~ys__n826 & ~new_new_n11726__;
  assign new_new_n46695__ = ~new_new_n46693__ & ~new_new_n46694__;
  assign new_new_n46696__ = ys__n47857 & ~new_new_n46695__;
  assign new_new_n46697__ = ~new_new_n46692__ & ~new_new_n46696__;
  assign new_new_n46698__ = ~new_new_n46691__ & new_new_n46695__;
  assign ys__n32364 = ~new_new_n46697__ & ~new_new_n46698__;
  assign new_new_n46700__ = ys__n48061 & new_new_n46691__;
  assign new_new_n46701__ = ys__n47858 & ~new_new_n46695__;
  assign new_new_n46702__ = ~new_new_n46700__ & ~new_new_n46701__;
  assign ys__n32365 = ~new_new_n46698__ & ~new_new_n46702__;
  assign new_new_n46704__ = ys__n48062 & new_new_n46691__;
  assign new_new_n46705__ = ys__n47859 & ~new_new_n46695__;
  assign new_new_n46706__ = ~new_new_n46704__ & ~new_new_n46705__;
  assign ys__n32366 = ~new_new_n46698__ & ~new_new_n46706__;
  assign new_new_n46708__ = ys__n48063 & new_new_n46691__;
  assign new_new_n46709__ = ys__n47860 & ~new_new_n46695__;
  assign new_new_n46710__ = ~new_new_n46708__ & ~new_new_n46709__;
  assign ys__n32367 = ~new_new_n46698__ & ~new_new_n46710__;
  assign new_new_n46712__ = ys__n48064 & new_new_n46691__;
  assign new_new_n46713__ = ys__n47861 & ~new_new_n46695__;
  assign new_new_n46714__ = ~new_new_n46712__ & ~new_new_n46713__;
  assign ys__n32368 = ~new_new_n46698__ & ~new_new_n46714__;
  assign new_new_n46716__ = ys__n48065 & new_new_n46691__;
  assign new_new_n46717__ = ys__n47862 & ~new_new_n46695__;
  assign new_new_n46718__ = ~new_new_n46716__ & ~new_new_n46717__;
  assign ys__n32369 = ~new_new_n46698__ & ~new_new_n46718__;
  assign new_new_n46720__ = ys__n48066 & new_new_n46691__;
  assign new_new_n46721__ = ys__n47863 & ~new_new_n46695__;
  assign new_new_n46722__ = ~new_new_n46720__ & ~new_new_n46721__;
  assign ys__n32370 = ~new_new_n46698__ & ~new_new_n46722__;
  assign new_new_n46724__ = ys__n48067 & new_new_n46691__;
  assign new_new_n46725__ = ys__n47864 & ~new_new_n46695__;
  assign new_new_n46726__ = ~new_new_n46724__ & ~new_new_n46725__;
  assign ys__n32371 = ~new_new_n46698__ & ~new_new_n46726__;
  assign new_new_n46728__ = ys__n48068 & new_new_n46691__;
  assign new_new_n46729__ = ys__n47865 & ~new_new_n46695__;
  assign new_new_n46730__ = ~new_new_n46728__ & ~new_new_n46729__;
  assign ys__n32372 = ~new_new_n46698__ & ~new_new_n46730__;
  assign new_new_n46732__ = ys__n48069 & new_new_n46691__;
  assign new_new_n46733__ = ys__n47866 & ~new_new_n46695__;
  assign new_new_n46734__ = ~new_new_n46732__ & ~new_new_n46733__;
  assign ys__n32373 = ~new_new_n46698__ & ~new_new_n46734__;
  assign new_new_n46736__ = ys__n48070 & new_new_n46691__;
  assign new_new_n46737__ = ys__n47867 & ~new_new_n46695__;
  assign new_new_n46738__ = ~new_new_n46736__ & ~new_new_n46737__;
  assign ys__n32374 = ~new_new_n46698__ & ~new_new_n46738__;
  assign new_new_n46740__ = ys__n48071 & new_new_n46691__;
  assign new_new_n46741__ = ys__n47868 & ~new_new_n46695__;
  assign new_new_n46742__ = ~new_new_n46740__ & ~new_new_n46741__;
  assign ys__n32375 = ~new_new_n46698__ & ~new_new_n46742__;
  assign new_new_n46744__ = ys__n48072 & new_new_n46691__;
  assign new_new_n46745__ = ys__n47869 & ~new_new_n46695__;
  assign new_new_n46746__ = ~new_new_n46744__ & ~new_new_n46745__;
  assign ys__n32376 = ~new_new_n46698__ & ~new_new_n46746__;
  assign new_new_n46748__ = ys__n48073 & new_new_n46691__;
  assign new_new_n46749__ = ys__n47870 & ~new_new_n46695__;
  assign new_new_n46750__ = ~new_new_n46748__ & ~new_new_n46749__;
  assign ys__n32377 = ~new_new_n46698__ & ~new_new_n46750__;
  assign new_new_n46752__ = ys__n48074 & new_new_n46691__;
  assign new_new_n46753__ = ys__n47871 & ~new_new_n46695__;
  assign new_new_n46754__ = ~new_new_n46752__ & ~new_new_n46753__;
  assign ys__n32378 = ~new_new_n46698__ & ~new_new_n46754__;
  assign new_new_n46756__ = ys__n48075 & new_new_n46691__;
  assign new_new_n46757__ = ys__n47872 & ~new_new_n46695__;
  assign new_new_n46758__ = ~new_new_n46756__ & ~new_new_n46757__;
  assign ys__n32379 = ~new_new_n46698__ & ~new_new_n46758__;
  assign new_new_n46760__ = ys__n48076 & new_new_n46691__;
  assign new_new_n46761__ = ys__n47873 & ~new_new_n46695__;
  assign new_new_n46762__ = ~new_new_n46760__ & ~new_new_n46761__;
  assign ys__n32380 = ~new_new_n46698__ & ~new_new_n46762__;
  assign new_new_n46764__ = ys__n48077 & new_new_n46691__;
  assign new_new_n46765__ = ys__n47874 & ~new_new_n46695__;
  assign new_new_n46766__ = ~new_new_n46764__ & ~new_new_n46765__;
  assign ys__n32381 = ~new_new_n46698__ & ~new_new_n46766__;
  assign new_new_n46768__ = ys__n48078 & new_new_n46691__;
  assign new_new_n46769__ = ys__n47875 & ~new_new_n46695__;
  assign new_new_n46770__ = ~new_new_n46768__ & ~new_new_n46769__;
  assign ys__n32382 = ~new_new_n46698__ & ~new_new_n46770__;
  assign new_new_n46772__ = ys__n48079 & new_new_n46691__;
  assign new_new_n46773__ = ys__n47876 & ~new_new_n46695__;
  assign new_new_n46774__ = ~new_new_n46772__ & ~new_new_n46773__;
  assign ys__n32383 = ~new_new_n46698__ & ~new_new_n46774__;
  assign new_new_n46776__ = ys__n48080 & new_new_n46691__;
  assign new_new_n46777__ = ys__n47877 & ~new_new_n46695__;
  assign new_new_n46778__ = ~new_new_n46776__ & ~new_new_n46777__;
  assign ys__n32384 = ~new_new_n46698__ & ~new_new_n46778__;
  assign new_new_n46780__ = ys__n48081 & new_new_n46691__;
  assign new_new_n46781__ = ys__n47878 & ~new_new_n46695__;
  assign new_new_n46782__ = ~new_new_n46780__ & ~new_new_n46781__;
  assign ys__n32385 = ~new_new_n46698__ & ~new_new_n46782__;
  assign new_new_n46784__ = ys__n48082 & new_new_n46691__;
  assign new_new_n46785__ = ys__n47879 & ~new_new_n46695__;
  assign new_new_n46786__ = ~new_new_n46784__ & ~new_new_n46785__;
  assign ys__n32386 = ~new_new_n46698__ & ~new_new_n46786__;
  assign new_new_n46788__ = ys__n48083 & new_new_n46691__;
  assign new_new_n46789__ = ys__n47880 & ~new_new_n46695__;
  assign new_new_n46790__ = ~new_new_n46788__ & ~new_new_n46789__;
  assign ys__n32387 = ~new_new_n46698__ & ~new_new_n46790__;
  assign new_new_n46792__ = ys__n48084 & new_new_n46691__;
  assign new_new_n46793__ = ys__n47881 & ~new_new_n46695__;
  assign new_new_n46794__ = ~new_new_n46792__ & ~new_new_n46793__;
  assign ys__n32388 = ~new_new_n46698__ & ~new_new_n46794__;
  assign new_new_n46796__ = ys__n48085 & new_new_n46691__;
  assign new_new_n46797__ = ys__n47882 & ~new_new_n46695__;
  assign new_new_n46798__ = ~new_new_n46796__ & ~new_new_n46797__;
  assign ys__n32389 = ~new_new_n46698__ & ~new_new_n46798__;
  assign new_new_n46800__ = ys__n48086 & new_new_n46691__;
  assign new_new_n46801__ = ys__n47883 & ~new_new_n46695__;
  assign new_new_n46802__ = ~new_new_n46800__ & ~new_new_n46801__;
  assign ys__n32390 = ~new_new_n46698__ & ~new_new_n46802__;
  assign new_new_n46804__ = ys__n48087 & new_new_n46691__;
  assign new_new_n46805__ = ys__n47884 & ~new_new_n46695__;
  assign new_new_n46806__ = ~new_new_n46804__ & ~new_new_n46805__;
  assign ys__n32391 = ~new_new_n46698__ & ~new_new_n46806__;
  assign new_new_n46808__ = ys__n48088 & new_new_n46691__;
  assign new_new_n46809__ = ys__n47885 & ~new_new_n46695__;
  assign new_new_n46810__ = ~new_new_n46808__ & ~new_new_n46809__;
  assign ys__n32392 = ~new_new_n46698__ & ~new_new_n46810__;
  assign new_new_n46812__ = ys__n48089 & new_new_n46691__;
  assign new_new_n46813__ = ys__n47886 & ~new_new_n46695__;
  assign new_new_n46814__ = ~new_new_n46812__ & ~new_new_n46813__;
  assign ys__n32393 = ~new_new_n46698__ & ~new_new_n46814__;
  assign new_new_n46816__ = ys__n48090 & new_new_n46691__;
  assign new_new_n46817__ = ys__n47887 & ~new_new_n46695__;
  assign new_new_n46818__ = ~new_new_n46816__ & ~new_new_n46817__;
  assign ys__n32394 = ~new_new_n46698__ & ~new_new_n46818__;
  assign new_new_n46820__ = ys__n48091 & new_new_n46691__;
  assign new_new_n46821__ = ys__n47888 & ~new_new_n46695__;
  assign new_new_n46822__ = ~new_new_n46820__ & ~new_new_n46821__;
  assign ys__n32395 = ~new_new_n46698__ & ~new_new_n46822__;
  assign new_new_n46824__ = ys__n48092 & new_new_n46691__;
  assign new_new_n46825__ = ys__n19215 & ~new_new_n46695__;
  assign new_new_n46826__ = ~new_new_n46824__ & ~new_new_n46825__;
  assign ys__n32396 = ~new_new_n46698__ & ~new_new_n46826__;
  assign new_new_n46828__ = ys__n48093 & new_new_n46691__;
  assign new_new_n46829__ = ys__n47889 & ~new_new_n46695__;
  assign new_new_n46830__ = ~new_new_n46828__ & ~new_new_n46829__;
  assign ys__n32397 = ~new_new_n46698__ & ~new_new_n46830__;
  assign new_new_n46832__ = ys__n116 & new_new_n12106__;
  assign new_new_n46833__ = ys__n48094 & new_new_n46832__;
  assign new_new_n46834__ = ~ys__n846 & ~new_new_n12106__;
  assign new_new_n46835__ = ~ys__n116 & new_new_n12106__;
  assign new_new_n46836__ = ~new_new_n46834__ & ~new_new_n46835__;
  assign new_new_n46837__ = ys__n18654 & ~new_new_n46836__;
  assign new_new_n46838__ = ~new_new_n46833__ & ~new_new_n46837__;
  assign new_new_n46839__ = ~new_new_n46832__ & new_new_n46836__;
  assign ys__n32398 = ~new_new_n46838__ & ~new_new_n46839__;
  assign new_new_n46841__ = ys__n48095 & new_new_n46832__;
  assign new_new_n46842__ = ys__n18657 & ~new_new_n46836__;
  assign new_new_n46843__ = ~new_new_n46841__ & ~new_new_n46842__;
  assign ys__n32399 = ~new_new_n46839__ & ~new_new_n46843__;
  assign new_new_n46845__ = ys__n48096 & new_new_n46832__;
  assign new_new_n46846__ = ys__n18660 & ~new_new_n46836__;
  assign new_new_n46847__ = ~new_new_n46845__ & ~new_new_n46846__;
  assign ys__n32400 = ~new_new_n46839__ & ~new_new_n46847__;
  assign new_new_n46849__ = ys__n48097 & new_new_n46832__;
  assign new_new_n46850__ = ys__n18663 & ~new_new_n46836__;
  assign new_new_n46851__ = ~new_new_n46849__ & ~new_new_n46850__;
  assign ys__n32401 = ~new_new_n46839__ & ~new_new_n46851__;
  assign new_new_n46853__ = ys__n37758 & new_new_n46832__;
  assign new_new_n46854__ = ys__n18666 & ~new_new_n46836__;
  assign new_new_n46855__ = ~new_new_n46853__ & ~new_new_n46854__;
  assign ys__n32402 = ~new_new_n46839__ & ~new_new_n46855__;
  assign new_new_n46857__ = ys__n37759 & new_new_n46832__;
  assign new_new_n46858__ = ys__n18669 & ~new_new_n46836__;
  assign new_new_n46859__ = ~new_new_n46857__ & ~new_new_n46858__;
  assign ys__n32403 = ~new_new_n46839__ & ~new_new_n46859__;
  assign new_new_n46861__ = ys__n37760 & new_new_n46832__;
  assign new_new_n46862__ = ys__n18672 & ~new_new_n46836__;
  assign new_new_n46863__ = ~new_new_n46861__ & ~new_new_n46862__;
  assign ys__n32404 = ~new_new_n46839__ & ~new_new_n46863__;
  assign new_new_n46865__ = ys__n37761 & new_new_n46832__;
  assign new_new_n46866__ = ys__n18675 & ~new_new_n46836__;
  assign new_new_n46867__ = ~new_new_n46865__ & ~new_new_n46866__;
  assign ys__n32405 = ~new_new_n46839__ & ~new_new_n46867__;
  assign new_new_n46869__ = ys__n37762 & new_new_n46832__;
  assign new_new_n46870__ = ys__n18678 & ~new_new_n46836__;
  assign new_new_n46871__ = ~new_new_n46869__ & ~new_new_n46870__;
  assign ys__n32406 = ~new_new_n46839__ & ~new_new_n46871__;
  assign new_new_n46873__ = ys__n37763 & new_new_n46832__;
  assign new_new_n46874__ = ys__n18681 & ~new_new_n46836__;
  assign new_new_n46875__ = ~new_new_n46873__ & ~new_new_n46874__;
  assign ys__n32407 = ~new_new_n46839__ & ~new_new_n46875__;
  assign new_new_n46877__ = ys__n37764 & new_new_n46832__;
  assign new_new_n46878__ = ys__n18684 & ~new_new_n46836__;
  assign new_new_n46879__ = ~new_new_n46877__ & ~new_new_n46878__;
  assign ys__n32408 = ~new_new_n46839__ & ~new_new_n46879__;
  assign new_new_n46881__ = ys__n37765 & new_new_n46832__;
  assign new_new_n46882__ = ys__n18687 & ~new_new_n46836__;
  assign new_new_n46883__ = ~new_new_n46881__ & ~new_new_n46882__;
  assign ys__n32409 = ~new_new_n46839__ & ~new_new_n46883__;
  assign new_new_n46885__ = ys__n37766 & new_new_n46832__;
  assign new_new_n46886__ = ys__n18690 & ~new_new_n46836__;
  assign new_new_n46887__ = ~new_new_n46885__ & ~new_new_n46886__;
  assign ys__n32410 = ~new_new_n46839__ & ~new_new_n46887__;
  assign new_new_n46889__ = ys__n37767 & new_new_n46832__;
  assign new_new_n46890__ = ys__n18693 & ~new_new_n46836__;
  assign new_new_n46891__ = ~new_new_n46889__ & ~new_new_n46890__;
  assign ys__n32411 = ~new_new_n46839__ & ~new_new_n46891__;
  assign new_new_n46893__ = ys__n37768 & new_new_n46832__;
  assign new_new_n46894__ = ys__n18696 & ~new_new_n46836__;
  assign new_new_n46895__ = ~new_new_n46893__ & ~new_new_n46894__;
  assign ys__n32412 = ~new_new_n46839__ & ~new_new_n46895__;
  assign new_new_n46897__ = ys__n37769 & new_new_n46832__;
  assign new_new_n46898__ = ys__n18699 & ~new_new_n46836__;
  assign new_new_n46899__ = ~new_new_n46897__ & ~new_new_n46898__;
  assign ys__n32413 = ~new_new_n46839__ & ~new_new_n46899__;
  assign new_new_n46901__ = ys__n37770 & new_new_n46832__;
  assign new_new_n46902__ = ys__n18702 & ~new_new_n46836__;
  assign new_new_n46903__ = ~new_new_n46901__ & ~new_new_n46902__;
  assign ys__n32414 = ~new_new_n46839__ & ~new_new_n46903__;
  assign new_new_n46905__ = ys__n37771 & new_new_n46832__;
  assign new_new_n46906__ = ys__n18705 & ~new_new_n46836__;
  assign new_new_n46907__ = ~new_new_n46905__ & ~new_new_n46906__;
  assign ys__n32415 = ~new_new_n46839__ & ~new_new_n46907__;
  assign new_new_n46909__ = ys__n37772 & new_new_n46832__;
  assign new_new_n46910__ = ys__n18708 & ~new_new_n46836__;
  assign new_new_n46911__ = ~new_new_n46909__ & ~new_new_n46910__;
  assign ys__n32416 = ~new_new_n46839__ & ~new_new_n46911__;
  assign new_new_n46913__ = ys__n37773 & new_new_n46832__;
  assign new_new_n46914__ = ys__n18711 & ~new_new_n46836__;
  assign new_new_n46915__ = ~new_new_n46913__ & ~new_new_n46914__;
  assign ys__n32417 = ~new_new_n46839__ & ~new_new_n46915__;
  assign new_new_n46917__ = ys__n37774 & new_new_n46832__;
  assign new_new_n46918__ = ys__n18714 & ~new_new_n46836__;
  assign new_new_n46919__ = ~new_new_n46917__ & ~new_new_n46918__;
  assign ys__n32418 = ~new_new_n46839__ & ~new_new_n46919__;
  assign new_new_n46921__ = ys__n37775 & new_new_n46832__;
  assign new_new_n46922__ = ys__n18717 & ~new_new_n46836__;
  assign new_new_n46923__ = ~new_new_n46921__ & ~new_new_n46922__;
  assign ys__n32419 = ~new_new_n46839__ & ~new_new_n46923__;
  assign new_new_n46925__ = ys__n37776 & new_new_n46832__;
  assign new_new_n46926__ = ys__n18720 & ~new_new_n46836__;
  assign new_new_n46927__ = ~new_new_n46925__ & ~new_new_n46926__;
  assign ys__n32420 = ~new_new_n46839__ & ~new_new_n46927__;
  assign new_new_n46929__ = ys__n37777 & new_new_n46832__;
  assign new_new_n46930__ = ys__n18723 & ~new_new_n46836__;
  assign new_new_n46931__ = ~new_new_n46929__ & ~new_new_n46930__;
  assign ys__n32421 = ~new_new_n46839__ & ~new_new_n46931__;
  assign new_new_n46933__ = ys__n37778 & new_new_n46832__;
  assign new_new_n46934__ = ys__n18726 & ~new_new_n46836__;
  assign new_new_n46935__ = ~new_new_n46933__ & ~new_new_n46934__;
  assign ys__n32422 = ~new_new_n46839__ & ~new_new_n46935__;
  assign new_new_n46937__ = ys__n37779 & new_new_n46832__;
  assign new_new_n46938__ = ys__n18729 & ~new_new_n46836__;
  assign new_new_n46939__ = ~new_new_n46937__ & ~new_new_n46938__;
  assign ys__n32423 = ~new_new_n46839__ & ~new_new_n46939__;
  assign new_new_n46941__ = ys__n37780 & new_new_n46832__;
  assign new_new_n46942__ = ys__n18732 & ~new_new_n46836__;
  assign new_new_n46943__ = ~new_new_n46941__ & ~new_new_n46942__;
  assign ys__n32424 = ~new_new_n46839__ & ~new_new_n46943__;
  assign new_new_n46945__ = ys__n37781 & new_new_n46832__;
  assign new_new_n46946__ = ys__n18735 & ~new_new_n46836__;
  assign new_new_n46947__ = ~new_new_n46945__ & ~new_new_n46946__;
  assign ys__n32425 = ~new_new_n46839__ & ~new_new_n46947__;
  assign new_new_n46949__ = ys__n37782 & new_new_n46832__;
  assign new_new_n46950__ = ys__n18738 & ~new_new_n46836__;
  assign new_new_n46951__ = ~new_new_n46949__ & ~new_new_n46950__;
  assign ys__n32426 = ~new_new_n46839__ & ~new_new_n46951__;
  assign new_new_n46953__ = ys__n37783 & new_new_n46832__;
  assign new_new_n46954__ = ys__n18741 & ~new_new_n46836__;
  assign new_new_n46955__ = ~new_new_n46953__ & ~new_new_n46954__;
  assign ys__n32427 = ~new_new_n46839__ & ~new_new_n46955__;
  assign new_new_n46957__ = ys__n37784 & new_new_n46832__;
  assign new_new_n46958__ = ys__n18744 & ~new_new_n46836__;
  assign new_new_n46959__ = ~new_new_n46957__ & ~new_new_n46958__;
  assign ys__n32428 = ~new_new_n46839__ & ~new_new_n46959__;
  assign new_new_n46961__ = ys__n37785 & new_new_n46832__;
  assign new_new_n46962__ = ys__n18747 & ~new_new_n46836__;
  assign new_new_n46963__ = ~new_new_n46961__ & ~new_new_n46962__;
  assign ys__n32429 = ~new_new_n46839__ & ~new_new_n46963__;
  assign new_new_n46965__ = ys__n846 & new_new_n12106__;
  assign new_new_n46966__ = ys__n48098 & new_new_n46965__;
  assign new_new_n46967__ = ~ys__n848 & ~new_new_n12106__;
  assign new_new_n46968__ = ~ys__n846 & new_new_n12106__;
  assign new_new_n46969__ = ~new_new_n46967__ & ~new_new_n46968__;
  assign new_new_n46970__ = ys__n18654 & ~new_new_n46969__;
  assign new_new_n46971__ = ~new_new_n46966__ & ~new_new_n46970__;
  assign new_new_n46972__ = ~new_new_n46965__ & new_new_n46969__;
  assign ys__n32430 = ~new_new_n46971__ & ~new_new_n46972__;
  assign new_new_n46974__ = ys__n48099 & new_new_n46965__;
  assign new_new_n46975__ = ys__n18657 & ~new_new_n46969__;
  assign new_new_n46976__ = ~new_new_n46974__ & ~new_new_n46975__;
  assign ys__n32431 = ~new_new_n46972__ & ~new_new_n46976__;
  assign new_new_n46978__ = ys__n48100 & new_new_n46965__;
  assign new_new_n46979__ = ys__n18660 & ~new_new_n46969__;
  assign new_new_n46980__ = ~new_new_n46978__ & ~new_new_n46979__;
  assign ys__n32432 = ~new_new_n46972__ & ~new_new_n46980__;
  assign new_new_n46982__ = ys__n48101 & new_new_n46965__;
  assign new_new_n46983__ = ys__n18663 & ~new_new_n46969__;
  assign new_new_n46984__ = ~new_new_n46982__ & ~new_new_n46983__;
  assign ys__n32433 = ~new_new_n46972__ & ~new_new_n46984__;
  assign new_new_n46986__ = ys__n37786 & new_new_n46965__;
  assign new_new_n46987__ = ys__n18666 & ~new_new_n46969__;
  assign new_new_n46988__ = ~new_new_n46986__ & ~new_new_n46987__;
  assign ys__n32434 = ~new_new_n46972__ & ~new_new_n46988__;
  assign new_new_n46990__ = ys__n37787 & new_new_n46965__;
  assign new_new_n46991__ = ys__n18669 & ~new_new_n46969__;
  assign new_new_n46992__ = ~new_new_n46990__ & ~new_new_n46991__;
  assign ys__n32435 = ~new_new_n46972__ & ~new_new_n46992__;
  assign new_new_n46994__ = ys__n37788 & new_new_n46965__;
  assign new_new_n46995__ = ys__n18672 & ~new_new_n46969__;
  assign new_new_n46996__ = ~new_new_n46994__ & ~new_new_n46995__;
  assign ys__n32436 = ~new_new_n46972__ & ~new_new_n46996__;
  assign new_new_n46998__ = ys__n37789 & new_new_n46965__;
  assign new_new_n46999__ = ys__n18675 & ~new_new_n46969__;
  assign new_new_n47000__ = ~new_new_n46998__ & ~new_new_n46999__;
  assign ys__n32437 = ~new_new_n46972__ & ~new_new_n47000__;
  assign new_new_n47002__ = ys__n37790 & new_new_n46965__;
  assign new_new_n47003__ = ys__n18678 & ~new_new_n46969__;
  assign new_new_n47004__ = ~new_new_n47002__ & ~new_new_n47003__;
  assign ys__n32438 = ~new_new_n46972__ & ~new_new_n47004__;
  assign new_new_n47006__ = ys__n37791 & new_new_n46965__;
  assign new_new_n47007__ = ys__n18681 & ~new_new_n46969__;
  assign new_new_n47008__ = ~new_new_n47006__ & ~new_new_n47007__;
  assign ys__n32439 = ~new_new_n46972__ & ~new_new_n47008__;
  assign new_new_n47010__ = ys__n37792 & new_new_n46965__;
  assign new_new_n47011__ = ys__n18684 & ~new_new_n46969__;
  assign new_new_n47012__ = ~new_new_n47010__ & ~new_new_n47011__;
  assign ys__n32440 = ~new_new_n46972__ & ~new_new_n47012__;
  assign new_new_n47014__ = ys__n37793 & new_new_n46965__;
  assign new_new_n47015__ = ys__n18687 & ~new_new_n46969__;
  assign new_new_n47016__ = ~new_new_n47014__ & ~new_new_n47015__;
  assign ys__n32441 = ~new_new_n46972__ & ~new_new_n47016__;
  assign new_new_n47018__ = ys__n37794 & new_new_n46965__;
  assign new_new_n47019__ = ys__n18690 & ~new_new_n46969__;
  assign new_new_n47020__ = ~new_new_n47018__ & ~new_new_n47019__;
  assign ys__n32442 = ~new_new_n46972__ & ~new_new_n47020__;
  assign new_new_n47022__ = ys__n37795 & new_new_n46965__;
  assign new_new_n47023__ = ys__n18693 & ~new_new_n46969__;
  assign new_new_n47024__ = ~new_new_n47022__ & ~new_new_n47023__;
  assign ys__n32443 = ~new_new_n46972__ & ~new_new_n47024__;
  assign new_new_n47026__ = ys__n37796 & new_new_n46965__;
  assign new_new_n47027__ = ys__n18696 & ~new_new_n46969__;
  assign new_new_n47028__ = ~new_new_n47026__ & ~new_new_n47027__;
  assign ys__n32444 = ~new_new_n46972__ & ~new_new_n47028__;
  assign new_new_n47030__ = ys__n37797 & new_new_n46965__;
  assign new_new_n47031__ = ys__n18699 & ~new_new_n46969__;
  assign new_new_n47032__ = ~new_new_n47030__ & ~new_new_n47031__;
  assign ys__n32445 = ~new_new_n46972__ & ~new_new_n47032__;
  assign new_new_n47034__ = ys__n37798 & new_new_n46965__;
  assign new_new_n47035__ = ys__n18702 & ~new_new_n46969__;
  assign new_new_n47036__ = ~new_new_n47034__ & ~new_new_n47035__;
  assign ys__n32446 = ~new_new_n46972__ & ~new_new_n47036__;
  assign new_new_n47038__ = ys__n37799 & new_new_n46965__;
  assign new_new_n47039__ = ys__n18705 & ~new_new_n46969__;
  assign new_new_n47040__ = ~new_new_n47038__ & ~new_new_n47039__;
  assign ys__n32447 = ~new_new_n46972__ & ~new_new_n47040__;
  assign new_new_n47042__ = ys__n37800 & new_new_n46965__;
  assign new_new_n47043__ = ys__n18708 & ~new_new_n46969__;
  assign new_new_n47044__ = ~new_new_n47042__ & ~new_new_n47043__;
  assign ys__n32448 = ~new_new_n46972__ & ~new_new_n47044__;
  assign new_new_n47046__ = ys__n37801 & new_new_n46965__;
  assign new_new_n47047__ = ys__n18711 & ~new_new_n46969__;
  assign new_new_n47048__ = ~new_new_n47046__ & ~new_new_n47047__;
  assign ys__n32449 = ~new_new_n46972__ & ~new_new_n47048__;
  assign new_new_n47050__ = ys__n37802 & new_new_n46965__;
  assign new_new_n47051__ = ys__n18714 & ~new_new_n46969__;
  assign new_new_n47052__ = ~new_new_n47050__ & ~new_new_n47051__;
  assign ys__n32450 = ~new_new_n46972__ & ~new_new_n47052__;
  assign new_new_n47054__ = ys__n37803 & new_new_n46965__;
  assign new_new_n47055__ = ys__n18717 & ~new_new_n46969__;
  assign new_new_n47056__ = ~new_new_n47054__ & ~new_new_n47055__;
  assign ys__n32451 = ~new_new_n46972__ & ~new_new_n47056__;
  assign new_new_n47058__ = ys__n37804 & new_new_n46965__;
  assign new_new_n47059__ = ys__n18720 & ~new_new_n46969__;
  assign new_new_n47060__ = ~new_new_n47058__ & ~new_new_n47059__;
  assign ys__n32452 = ~new_new_n46972__ & ~new_new_n47060__;
  assign new_new_n47062__ = ys__n37805 & new_new_n46965__;
  assign new_new_n47063__ = ys__n18723 & ~new_new_n46969__;
  assign new_new_n47064__ = ~new_new_n47062__ & ~new_new_n47063__;
  assign ys__n32453 = ~new_new_n46972__ & ~new_new_n47064__;
  assign new_new_n47066__ = ys__n37806 & new_new_n46965__;
  assign new_new_n47067__ = ys__n18726 & ~new_new_n46969__;
  assign new_new_n47068__ = ~new_new_n47066__ & ~new_new_n47067__;
  assign ys__n32454 = ~new_new_n46972__ & ~new_new_n47068__;
  assign new_new_n47070__ = ys__n37807 & new_new_n46965__;
  assign new_new_n47071__ = ys__n18729 & ~new_new_n46969__;
  assign new_new_n47072__ = ~new_new_n47070__ & ~new_new_n47071__;
  assign ys__n32455 = ~new_new_n46972__ & ~new_new_n47072__;
  assign new_new_n47074__ = ys__n37808 & new_new_n46965__;
  assign new_new_n47075__ = ys__n18732 & ~new_new_n46969__;
  assign new_new_n47076__ = ~new_new_n47074__ & ~new_new_n47075__;
  assign ys__n32456 = ~new_new_n46972__ & ~new_new_n47076__;
  assign new_new_n47078__ = ys__n37809 & new_new_n46965__;
  assign new_new_n47079__ = ys__n18735 & ~new_new_n46969__;
  assign new_new_n47080__ = ~new_new_n47078__ & ~new_new_n47079__;
  assign ys__n32457 = ~new_new_n46972__ & ~new_new_n47080__;
  assign new_new_n47082__ = ys__n37810 & new_new_n46965__;
  assign new_new_n47083__ = ys__n18738 & ~new_new_n46969__;
  assign new_new_n47084__ = ~new_new_n47082__ & ~new_new_n47083__;
  assign ys__n32458 = ~new_new_n46972__ & ~new_new_n47084__;
  assign new_new_n47086__ = ys__n37811 & new_new_n46965__;
  assign new_new_n47087__ = ys__n18741 & ~new_new_n46969__;
  assign new_new_n47088__ = ~new_new_n47086__ & ~new_new_n47087__;
  assign ys__n32459 = ~new_new_n46972__ & ~new_new_n47088__;
  assign new_new_n47090__ = ys__n37812 & new_new_n46965__;
  assign new_new_n47091__ = ys__n18744 & ~new_new_n46969__;
  assign new_new_n47092__ = ~new_new_n47090__ & ~new_new_n47091__;
  assign ys__n32460 = ~new_new_n46972__ & ~new_new_n47092__;
  assign new_new_n47094__ = ys__n37813 & new_new_n46965__;
  assign new_new_n47095__ = ys__n18747 & ~new_new_n46969__;
  assign new_new_n47096__ = ~new_new_n47094__ & ~new_new_n47095__;
  assign ys__n32461 = ~new_new_n46972__ & ~new_new_n47096__;
  assign new_new_n47098__ = ys__n848 & new_new_n12106__;
  assign new_new_n47099__ = ys__n48102 & new_new_n47098__;
  assign new_new_n47100__ = ~ys__n850 & ~new_new_n12106__;
  assign new_new_n47101__ = ~ys__n848 & new_new_n12106__;
  assign new_new_n47102__ = ~new_new_n47100__ & ~new_new_n47101__;
  assign new_new_n47103__ = ys__n18654 & ~new_new_n47102__;
  assign new_new_n47104__ = ~new_new_n47099__ & ~new_new_n47103__;
  assign new_new_n47105__ = ~new_new_n47098__ & new_new_n47102__;
  assign ys__n32462 = ~new_new_n47104__ & ~new_new_n47105__;
  assign new_new_n47107__ = ys__n48103 & new_new_n47098__;
  assign new_new_n47108__ = ys__n18657 & ~new_new_n47102__;
  assign new_new_n47109__ = ~new_new_n47107__ & ~new_new_n47108__;
  assign ys__n32463 = ~new_new_n47105__ & ~new_new_n47109__;
  assign new_new_n47111__ = ys__n48104 & new_new_n47098__;
  assign new_new_n47112__ = ys__n18660 & ~new_new_n47102__;
  assign new_new_n47113__ = ~new_new_n47111__ & ~new_new_n47112__;
  assign ys__n32464 = ~new_new_n47105__ & ~new_new_n47113__;
  assign new_new_n47115__ = ys__n48105 & new_new_n47098__;
  assign new_new_n47116__ = ys__n18663 & ~new_new_n47102__;
  assign new_new_n47117__ = ~new_new_n47115__ & ~new_new_n47116__;
  assign ys__n32465 = ~new_new_n47105__ & ~new_new_n47117__;
  assign new_new_n47119__ = ys__n37814 & new_new_n47098__;
  assign new_new_n47120__ = ys__n18666 & ~new_new_n47102__;
  assign new_new_n47121__ = ~new_new_n47119__ & ~new_new_n47120__;
  assign ys__n32466 = ~new_new_n47105__ & ~new_new_n47121__;
  assign new_new_n47123__ = ys__n37815 & new_new_n47098__;
  assign new_new_n47124__ = ys__n18669 & ~new_new_n47102__;
  assign new_new_n47125__ = ~new_new_n47123__ & ~new_new_n47124__;
  assign ys__n32467 = ~new_new_n47105__ & ~new_new_n47125__;
  assign new_new_n47127__ = ys__n37816 & new_new_n47098__;
  assign new_new_n47128__ = ys__n18672 & ~new_new_n47102__;
  assign new_new_n47129__ = ~new_new_n47127__ & ~new_new_n47128__;
  assign ys__n32468 = ~new_new_n47105__ & ~new_new_n47129__;
  assign new_new_n47131__ = ys__n37817 & new_new_n47098__;
  assign new_new_n47132__ = ys__n18675 & ~new_new_n47102__;
  assign new_new_n47133__ = ~new_new_n47131__ & ~new_new_n47132__;
  assign ys__n32469 = ~new_new_n47105__ & ~new_new_n47133__;
  assign new_new_n47135__ = ys__n37818 & new_new_n47098__;
  assign new_new_n47136__ = ys__n18678 & ~new_new_n47102__;
  assign new_new_n47137__ = ~new_new_n47135__ & ~new_new_n47136__;
  assign ys__n32470 = ~new_new_n47105__ & ~new_new_n47137__;
  assign new_new_n47139__ = ys__n37819 & new_new_n47098__;
  assign new_new_n47140__ = ys__n18681 & ~new_new_n47102__;
  assign new_new_n47141__ = ~new_new_n47139__ & ~new_new_n47140__;
  assign ys__n32471 = ~new_new_n47105__ & ~new_new_n47141__;
  assign new_new_n47143__ = ys__n37820 & new_new_n47098__;
  assign new_new_n47144__ = ys__n18684 & ~new_new_n47102__;
  assign new_new_n47145__ = ~new_new_n47143__ & ~new_new_n47144__;
  assign ys__n32472 = ~new_new_n47105__ & ~new_new_n47145__;
  assign new_new_n47147__ = ys__n37821 & new_new_n47098__;
  assign new_new_n47148__ = ys__n18687 & ~new_new_n47102__;
  assign new_new_n47149__ = ~new_new_n47147__ & ~new_new_n47148__;
  assign ys__n32473 = ~new_new_n47105__ & ~new_new_n47149__;
  assign new_new_n47151__ = ys__n37822 & new_new_n47098__;
  assign new_new_n47152__ = ys__n18690 & ~new_new_n47102__;
  assign new_new_n47153__ = ~new_new_n47151__ & ~new_new_n47152__;
  assign ys__n32474 = ~new_new_n47105__ & ~new_new_n47153__;
  assign new_new_n47155__ = ys__n37823 & new_new_n47098__;
  assign new_new_n47156__ = ys__n18693 & ~new_new_n47102__;
  assign new_new_n47157__ = ~new_new_n47155__ & ~new_new_n47156__;
  assign ys__n32475 = ~new_new_n47105__ & ~new_new_n47157__;
  assign new_new_n47159__ = ys__n37824 & new_new_n47098__;
  assign new_new_n47160__ = ys__n18696 & ~new_new_n47102__;
  assign new_new_n47161__ = ~new_new_n47159__ & ~new_new_n47160__;
  assign ys__n32476 = ~new_new_n47105__ & ~new_new_n47161__;
  assign new_new_n47163__ = ys__n37825 & new_new_n47098__;
  assign new_new_n47164__ = ys__n18699 & ~new_new_n47102__;
  assign new_new_n47165__ = ~new_new_n47163__ & ~new_new_n47164__;
  assign ys__n32477 = ~new_new_n47105__ & ~new_new_n47165__;
  assign new_new_n47167__ = ys__n37826 & new_new_n47098__;
  assign new_new_n47168__ = ys__n18702 & ~new_new_n47102__;
  assign new_new_n47169__ = ~new_new_n47167__ & ~new_new_n47168__;
  assign ys__n32478 = ~new_new_n47105__ & ~new_new_n47169__;
  assign new_new_n47171__ = ys__n37827 & new_new_n47098__;
  assign new_new_n47172__ = ys__n18705 & ~new_new_n47102__;
  assign new_new_n47173__ = ~new_new_n47171__ & ~new_new_n47172__;
  assign ys__n32479 = ~new_new_n47105__ & ~new_new_n47173__;
  assign new_new_n47175__ = ys__n37828 & new_new_n47098__;
  assign new_new_n47176__ = ys__n18708 & ~new_new_n47102__;
  assign new_new_n47177__ = ~new_new_n47175__ & ~new_new_n47176__;
  assign ys__n32480 = ~new_new_n47105__ & ~new_new_n47177__;
  assign new_new_n47179__ = ys__n37829 & new_new_n47098__;
  assign new_new_n47180__ = ys__n18711 & ~new_new_n47102__;
  assign new_new_n47181__ = ~new_new_n47179__ & ~new_new_n47180__;
  assign ys__n32481 = ~new_new_n47105__ & ~new_new_n47181__;
  assign new_new_n47183__ = ys__n37830 & new_new_n47098__;
  assign new_new_n47184__ = ys__n18714 & ~new_new_n47102__;
  assign new_new_n47185__ = ~new_new_n47183__ & ~new_new_n47184__;
  assign ys__n32482 = ~new_new_n47105__ & ~new_new_n47185__;
  assign new_new_n47187__ = ys__n37831 & new_new_n47098__;
  assign new_new_n47188__ = ys__n18717 & ~new_new_n47102__;
  assign new_new_n47189__ = ~new_new_n47187__ & ~new_new_n47188__;
  assign ys__n32483 = ~new_new_n47105__ & ~new_new_n47189__;
  assign new_new_n47191__ = ys__n37832 & new_new_n47098__;
  assign new_new_n47192__ = ys__n18720 & ~new_new_n47102__;
  assign new_new_n47193__ = ~new_new_n47191__ & ~new_new_n47192__;
  assign ys__n32484 = ~new_new_n47105__ & ~new_new_n47193__;
  assign new_new_n47195__ = ys__n37833 & new_new_n47098__;
  assign new_new_n47196__ = ys__n18723 & ~new_new_n47102__;
  assign new_new_n47197__ = ~new_new_n47195__ & ~new_new_n47196__;
  assign ys__n32485 = ~new_new_n47105__ & ~new_new_n47197__;
  assign new_new_n47199__ = ys__n37834 & new_new_n47098__;
  assign new_new_n47200__ = ys__n18726 & ~new_new_n47102__;
  assign new_new_n47201__ = ~new_new_n47199__ & ~new_new_n47200__;
  assign ys__n32486 = ~new_new_n47105__ & ~new_new_n47201__;
  assign new_new_n47203__ = ys__n37835 & new_new_n47098__;
  assign new_new_n47204__ = ys__n18729 & ~new_new_n47102__;
  assign new_new_n47205__ = ~new_new_n47203__ & ~new_new_n47204__;
  assign ys__n32487 = ~new_new_n47105__ & ~new_new_n47205__;
  assign new_new_n47207__ = ys__n37836 & new_new_n47098__;
  assign new_new_n47208__ = ys__n18732 & ~new_new_n47102__;
  assign new_new_n47209__ = ~new_new_n47207__ & ~new_new_n47208__;
  assign ys__n32488 = ~new_new_n47105__ & ~new_new_n47209__;
  assign new_new_n47211__ = ys__n37837 & new_new_n47098__;
  assign new_new_n47212__ = ys__n18735 & ~new_new_n47102__;
  assign new_new_n47213__ = ~new_new_n47211__ & ~new_new_n47212__;
  assign ys__n32489 = ~new_new_n47105__ & ~new_new_n47213__;
  assign new_new_n47215__ = ys__n37838 & new_new_n47098__;
  assign new_new_n47216__ = ys__n18738 & ~new_new_n47102__;
  assign new_new_n47217__ = ~new_new_n47215__ & ~new_new_n47216__;
  assign ys__n32490 = ~new_new_n47105__ & ~new_new_n47217__;
  assign new_new_n47219__ = ys__n37839 & new_new_n47098__;
  assign new_new_n47220__ = ys__n18741 & ~new_new_n47102__;
  assign new_new_n47221__ = ~new_new_n47219__ & ~new_new_n47220__;
  assign ys__n32491 = ~new_new_n47105__ & ~new_new_n47221__;
  assign new_new_n47223__ = ys__n37840 & new_new_n47098__;
  assign new_new_n47224__ = ys__n18744 & ~new_new_n47102__;
  assign new_new_n47225__ = ~new_new_n47223__ & ~new_new_n47224__;
  assign ys__n32492 = ~new_new_n47105__ & ~new_new_n47225__;
  assign new_new_n47227__ = ys__n37841 & new_new_n47098__;
  assign new_new_n47228__ = ys__n18747 & ~new_new_n47102__;
  assign new_new_n47229__ = ~new_new_n47227__ & ~new_new_n47228__;
  assign ys__n32493 = ~new_new_n47105__ & ~new_new_n47229__;
  assign new_new_n47231__ = ys__n48106 & new_new_n43944__;
  assign new_new_n47232__ = ys__n18654 & ~new_new_n43948__;
  assign new_new_n47233__ = ~new_new_n47231__ & ~new_new_n47232__;
  assign ys__n32494 = ~new_new_n43951__ & ~new_new_n47233__;
  assign new_new_n47235__ = ys__n48107 & new_new_n43944__;
  assign new_new_n47236__ = ys__n18657 & ~new_new_n43948__;
  assign new_new_n47237__ = ~new_new_n47235__ & ~new_new_n47236__;
  assign ys__n32495 = ~new_new_n43951__ & ~new_new_n47237__;
  assign new_new_n47239__ = ys__n48108 & new_new_n43944__;
  assign new_new_n47240__ = ys__n18660 & ~new_new_n43948__;
  assign new_new_n47241__ = ~new_new_n47239__ & ~new_new_n47240__;
  assign ys__n32496 = ~new_new_n43951__ & ~new_new_n47241__;
  assign new_new_n47243__ = ys__n48109 & new_new_n43944__;
  assign new_new_n47244__ = ys__n18663 & ~new_new_n43948__;
  assign new_new_n47245__ = ~new_new_n47243__ & ~new_new_n47244__;
  assign ys__n32497 = ~new_new_n43951__ & ~new_new_n47245__;
  assign new_new_n47247__ = ys__n37842 & new_new_n43944__;
  assign new_new_n47248__ = ys__n18666 & ~new_new_n43948__;
  assign new_new_n47249__ = ~new_new_n47247__ & ~new_new_n47248__;
  assign ys__n32498 = ~new_new_n43951__ & ~new_new_n47249__;
  assign new_new_n47251__ = ys__n37843 & new_new_n43944__;
  assign new_new_n47252__ = ys__n18669 & ~new_new_n43948__;
  assign new_new_n47253__ = ~new_new_n47251__ & ~new_new_n47252__;
  assign ys__n32499 = ~new_new_n43951__ & ~new_new_n47253__;
  assign new_new_n47255__ = ys__n37844 & new_new_n43944__;
  assign new_new_n47256__ = ys__n18672 & ~new_new_n43948__;
  assign new_new_n47257__ = ~new_new_n47255__ & ~new_new_n47256__;
  assign ys__n32500 = ~new_new_n43951__ & ~new_new_n47257__;
  assign new_new_n47259__ = ys__n37845 & new_new_n43944__;
  assign new_new_n47260__ = ys__n18675 & ~new_new_n43948__;
  assign new_new_n47261__ = ~new_new_n47259__ & ~new_new_n47260__;
  assign ys__n32501 = ~new_new_n43951__ & ~new_new_n47261__;
  assign new_new_n47263__ = ys__n37846 & new_new_n43944__;
  assign new_new_n47264__ = ys__n18678 & ~new_new_n43948__;
  assign new_new_n47265__ = ~new_new_n47263__ & ~new_new_n47264__;
  assign ys__n32502 = ~new_new_n43951__ & ~new_new_n47265__;
  assign new_new_n47267__ = ys__n37847 & new_new_n43944__;
  assign new_new_n47268__ = ys__n18681 & ~new_new_n43948__;
  assign new_new_n47269__ = ~new_new_n47267__ & ~new_new_n47268__;
  assign ys__n32503 = ~new_new_n43951__ & ~new_new_n47269__;
  assign new_new_n47271__ = ys__n37848 & new_new_n43944__;
  assign new_new_n47272__ = ys__n18684 & ~new_new_n43948__;
  assign new_new_n47273__ = ~new_new_n47271__ & ~new_new_n47272__;
  assign ys__n32504 = ~new_new_n43951__ & ~new_new_n47273__;
  assign new_new_n47275__ = ys__n37849 & new_new_n43944__;
  assign new_new_n47276__ = ys__n18687 & ~new_new_n43948__;
  assign new_new_n47277__ = ~new_new_n47275__ & ~new_new_n47276__;
  assign ys__n32505 = ~new_new_n43951__ & ~new_new_n47277__;
  assign new_new_n47279__ = ys__n37850 & new_new_n43944__;
  assign new_new_n47280__ = ys__n18690 & ~new_new_n43948__;
  assign new_new_n47281__ = ~new_new_n47279__ & ~new_new_n47280__;
  assign ys__n32506 = ~new_new_n43951__ & ~new_new_n47281__;
  assign new_new_n47283__ = ys__n37851 & new_new_n43944__;
  assign new_new_n47284__ = ys__n18693 & ~new_new_n43948__;
  assign new_new_n47285__ = ~new_new_n47283__ & ~new_new_n47284__;
  assign ys__n32507 = ~new_new_n43951__ & ~new_new_n47285__;
  assign new_new_n47287__ = ys__n37852 & new_new_n43944__;
  assign new_new_n47288__ = ys__n18696 & ~new_new_n43948__;
  assign new_new_n47289__ = ~new_new_n47287__ & ~new_new_n47288__;
  assign ys__n32508 = ~new_new_n43951__ & ~new_new_n47289__;
  assign new_new_n47291__ = ys__n37853 & new_new_n43944__;
  assign new_new_n47292__ = ys__n18699 & ~new_new_n43948__;
  assign new_new_n47293__ = ~new_new_n47291__ & ~new_new_n47292__;
  assign ys__n32509 = ~new_new_n43951__ & ~new_new_n47293__;
  assign new_new_n47295__ = ys__n37854 & new_new_n43944__;
  assign new_new_n47296__ = ys__n18702 & ~new_new_n43948__;
  assign new_new_n47297__ = ~new_new_n47295__ & ~new_new_n47296__;
  assign ys__n32510 = ~new_new_n43951__ & ~new_new_n47297__;
  assign new_new_n47299__ = ys__n37855 & new_new_n43944__;
  assign new_new_n47300__ = ys__n18705 & ~new_new_n43948__;
  assign new_new_n47301__ = ~new_new_n47299__ & ~new_new_n47300__;
  assign ys__n32511 = ~new_new_n43951__ & ~new_new_n47301__;
  assign new_new_n47303__ = ys__n37856 & new_new_n43944__;
  assign new_new_n47304__ = ys__n18708 & ~new_new_n43948__;
  assign new_new_n47305__ = ~new_new_n47303__ & ~new_new_n47304__;
  assign ys__n32512 = ~new_new_n43951__ & ~new_new_n47305__;
  assign new_new_n47307__ = ys__n37857 & new_new_n43944__;
  assign new_new_n47308__ = ys__n18711 & ~new_new_n43948__;
  assign new_new_n47309__ = ~new_new_n47307__ & ~new_new_n47308__;
  assign ys__n32513 = ~new_new_n43951__ & ~new_new_n47309__;
  assign new_new_n47311__ = ys__n37858 & new_new_n43944__;
  assign new_new_n47312__ = ys__n18714 & ~new_new_n43948__;
  assign new_new_n47313__ = ~new_new_n47311__ & ~new_new_n47312__;
  assign ys__n32514 = ~new_new_n43951__ & ~new_new_n47313__;
  assign new_new_n47315__ = ys__n37859 & new_new_n43944__;
  assign new_new_n47316__ = ys__n18717 & ~new_new_n43948__;
  assign new_new_n47317__ = ~new_new_n47315__ & ~new_new_n47316__;
  assign ys__n32515 = ~new_new_n43951__ & ~new_new_n47317__;
  assign new_new_n47319__ = ys__n37860 & new_new_n43944__;
  assign new_new_n47320__ = ys__n18720 & ~new_new_n43948__;
  assign new_new_n47321__ = ~new_new_n47319__ & ~new_new_n47320__;
  assign ys__n32516 = ~new_new_n43951__ & ~new_new_n47321__;
  assign new_new_n47323__ = ys__n37861 & new_new_n43944__;
  assign new_new_n47324__ = ys__n18723 & ~new_new_n43948__;
  assign new_new_n47325__ = ~new_new_n47323__ & ~new_new_n47324__;
  assign ys__n32517 = ~new_new_n43951__ & ~new_new_n47325__;
  assign new_new_n47327__ = ys__n37862 & new_new_n43944__;
  assign new_new_n47328__ = ys__n18726 & ~new_new_n43948__;
  assign new_new_n47329__ = ~new_new_n47327__ & ~new_new_n47328__;
  assign ys__n32518 = ~new_new_n43951__ & ~new_new_n47329__;
  assign new_new_n47331__ = ys__n37863 & new_new_n43944__;
  assign new_new_n47332__ = ys__n18729 & ~new_new_n43948__;
  assign new_new_n47333__ = ~new_new_n47331__ & ~new_new_n47332__;
  assign ys__n32519 = ~new_new_n43951__ & ~new_new_n47333__;
  assign new_new_n47335__ = ys__n37864 & new_new_n43944__;
  assign new_new_n47336__ = ys__n18732 & ~new_new_n43948__;
  assign new_new_n47337__ = ~new_new_n47335__ & ~new_new_n47336__;
  assign ys__n32520 = ~new_new_n43951__ & ~new_new_n47337__;
  assign new_new_n47339__ = ys__n37865 & new_new_n43944__;
  assign new_new_n47340__ = ys__n18735 & ~new_new_n43948__;
  assign new_new_n47341__ = ~new_new_n47339__ & ~new_new_n47340__;
  assign ys__n32521 = ~new_new_n43951__ & ~new_new_n47341__;
  assign new_new_n47343__ = ys__n37866 & new_new_n43944__;
  assign new_new_n47344__ = ys__n18738 & ~new_new_n43948__;
  assign new_new_n47345__ = ~new_new_n47343__ & ~new_new_n47344__;
  assign ys__n32522 = ~new_new_n43951__ & ~new_new_n47345__;
  assign new_new_n47347__ = ys__n37867 & new_new_n43944__;
  assign new_new_n47348__ = ys__n18741 & ~new_new_n43948__;
  assign new_new_n47349__ = ~new_new_n47347__ & ~new_new_n47348__;
  assign ys__n32523 = ~new_new_n43951__ & ~new_new_n47349__;
  assign new_new_n47351__ = ys__n37868 & new_new_n43944__;
  assign new_new_n47352__ = ys__n18744 & ~new_new_n43948__;
  assign new_new_n47353__ = ~new_new_n47351__ & ~new_new_n47352__;
  assign ys__n32524 = ~new_new_n43951__ & ~new_new_n47353__;
  assign new_new_n47355__ = ys__n37869 & new_new_n43944__;
  assign new_new_n47356__ = ys__n18747 & ~new_new_n43948__;
  assign new_new_n47357__ = ~new_new_n47355__ & ~new_new_n47356__;
  assign ys__n32525 = ~new_new_n43951__ & ~new_new_n47357__;
  assign new_new_n47359__ = ys__n48110 & new_new_n43799__;
  assign new_new_n47360__ = ys__n18654 & ~new_new_n43803__;
  assign new_new_n47361__ = ~new_new_n47359__ & ~new_new_n47360__;
  assign ys__n32526 = ~new_new_n43806__ & ~new_new_n47361__;
  assign new_new_n47363__ = ys__n48111 & new_new_n43799__;
  assign new_new_n47364__ = ys__n18657 & ~new_new_n43803__;
  assign new_new_n47365__ = ~new_new_n47363__ & ~new_new_n47364__;
  assign ys__n32527 = ~new_new_n43806__ & ~new_new_n47365__;
  assign new_new_n47367__ = ys__n48112 & new_new_n43799__;
  assign new_new_n47368__ = ys__n18660 & ~new_new_n43803__;
  assign new_new_n47369__ = ~new_new_n47367__ & ~new_new_n47368__;
  assign ys__n32528 = ~new_new_n43806__ & ~new_new_n47369__;
  assign new_new_n47371__ = ys__n48113 & new_new_n43799__;
  assign new_new_n47372__ = ys__n18663 & ~new_new_n43803__;
  assign new_new_n47373__ = ~new_new_n47371__ & ~new_new_n47372__;
  assign ys__n32529 = ~new_new_n43806__ & ~new_new_n47373__;
  assign new_new_n47375__ = ys__n37870 & new_new_n43799__;
  assign new_new_n47376__ = ys__n18666 & ~new_new_n43803__;
  assign new_new_n47377__ = ~new_new_n47375__ & ~new_new_n47376__;
  assign ys__n32530 = ~new_new_n43806__ & ~new_new_n47377__;
  assign new_new_n47379__ = ys__n37871 & new_new_n43799__;
  assign new_new_n47380__ = ys__n18669 & ~new_new_n43803__;
  assign new_new_n47381__ = ~new_new_n47379__ & ~new_new_n47380__;
  assign ys__n32531 = ~new_new_n43806__ & ~new_new_n47381__;
  assign new_new_n47383__ = ys__n37872 & new_new_n43799__;
  assign new_new_n47384__ = ys__n18672 & ~new_new_n43803__;
  assign new_new_n47385__ = ~new_new_n47383__ & ~new_new_n47384__;
  assign ys__n32532 = ~new_new_n43806__ & ~new_new_n47385__;
  assign new_new_n47387__ = ys__n37873 & new_new_n43799__;
  assign new_new_n47388__ = ys__n18675 & ~new_new_n43803__;
  assign new_new_n47389__ = ~new_new_n47387__ & ~new_new_n47388__;
  assign ys__n32533 = ~new_new_n43806__ & ~new_new_n47389__;
  assign new_new_n47391__ = ys__n37874 & new_new_n43799__;
  assign new_new_n47392__ = ys__n18678 & ~new_new_n43803__;
  assign new_new_n47393__ = ~new_new_n47391__ & ~new_new_n47392__;
  assign ys__n32534 = ~new_new_n43806__ & ~new_new_n47393__;
  assign new_new_n47395__ = ys__n37875 & new_new_n43799__;
  assign new_new_n47396__ = ys__n18681 & ~new_new_n43803__;
  assign new_new_n47397__ = ~new_new_n47395__ & ~new_new_n47396__;
  assign ys__n32535 = ~new_new_n43806__ & ~new_new_n47397__;
  assign new_new_n47399__ = ys__n37876 & new_new_n43799__;
  assign new_new_n47400__ = ys__n18684 & ~new_new_n43803__;
  assign new_new_n47401__ = ~new_new_n47399__ & ~new_new_n47400__;
  assign ys__n32536 = ~new_new_n43806__ & ~new_new_n47401__;
  assign new_new_n47403__ = ys__n37877 & new_new_n43799__;
  assign new_new_n47404__ = ys__n18687 & ~new_new_n43803__;
  assign new_new_n47405__ = ~new_new_n47403__ & ~new_new_n47404__;
  assign ys__n32537 = ~new_new_n43806__ & ~new_new_n47405__;
  assign new_new_n47407__ = ys__n37878 & new_new_n43799__;
  assign new_new_n47408__ = ys__n18690 & ~new_new_n43803__;
  assign new_new_n47409__ = ~new_new_n47407__ & ~new_new_n47408__;
  assign ys__n32538 = ~new_new_n43806__ & ~new_new_n47409__;
  assign new_new_n47411__ = ys__n37879 & new_new_n43799__;
  assign new_new_n47412__ = ys__n18693 & ~new_new_n43803__;
  assign new_new_n47413__ = ~new_new_n47411__ & ~new_new_n47412__;
  assign ys__n32539 = ~new_new_n43806__ & ~new_new_n47413__;
  assign new_new_n47415__ = ys__n37880 & new_new_n43799__;
  assign new_new_n47416__ = ys__n18696 & ~new_new_n43803__;
  assign new_new_n47417__ = ~new_new_n47415__ & ~new_new_n47416__;
  assign ys__n32540 = ~new_new_n43806__ & ~new_new_n47417__;
  assign new_new_n47419__ = ys__n37881 & new_new_n43799__;
  assign new_new_n47420__ = ys__n18699 & ~new_new_n43803__;
  assign new_new_n47421__ = ~new_new_n47419__ & ~new_new_n47420__;
  assign ys__n32541 = ~new_new_n43806__ & ~new_new_n47421__;
  assign new_new_n47423__ = ys__n37882 & new_new_n43799__;
  assign new_new_n47424__ = ys__n18702 & ~new_new_n43803__;
  assign new_new_n47425__ = ~new_new_n47423__ & ~new_new_n47424__;
  assign ys__n32542 = ~new_new_n43806__ & ~new_new_n47425__;
  assign new_new_n47427__ = ys__n37883 & new_new_n43799__;
  assign new_new_n47428__ = ys__n18705 & ~new_new_n43803__;
  assign new_new_n47429__ = ~new_new_n47427__ & ~new_new_n47428__;
  assign ys__n32543 = ~new_new_n43806__ & ~new_new_n47429__;
  assign new_new_n47431__ = ys__n37884 & new_new_n43799__;
  assign new_new_n47432__ = ys__n18708 & ~new_new_n43803__;
  assign new_new_n47433__ = ~new_new_n47431__ & ~new_new_n47432__;
  assign ys__n32544 = ~new_new_n43806__ & ~new_new_n47433__;
  assign new_new_n47435__ = ys__n37885 & new_new_n43799__;
  assign new_new_n47436__ = ys__n18711 & ~new_new_n43803__;
  assign new_new_n47437__ = ~new_new_n47435__ & ~new_new_n47436__;
  assign ys__n32545 = ~new_new_n43806__ & ~new_new_n47437__;
  assign new_new_n47439__ = ys__n37886 & new_new_n43799__;
  assign new_new_n47440__ = ys__n18714 & ~new_new_n43803__;
  assign new_new_n47441__ = ~new_new_n47439__ & ~new_new_n47440__;
  assign ys__n32546 = ~new_new_n43806__ & ~new_new_n47441__;
  assign new_new_n47443__ = ys__n37887 & new_new_n43799__;
  assign new_new_n47444__ = ys__n18717 & ~new_new_n43803__;
  assign new_new_n47445__ = ~new_new_n47443__ & ~new_new_n47444__;
  assign ys__n32547 = ~new_new_n43806__ & ~new_new_n47445__;
  assign new_new_n47447__ = ys__n37888 & new_new_n43799__;
  assign new_new_n47448__ = ys__n18720 & ~new_new_n43803__;
  assign new_new_n47449__ = ~new_new_n47447__ & ~new_new_n47448__;
  assign ys__n32548 = ~new_new_n43806__ & ~new_new_n47449__;
  assign new_new_n47451__ = ys__n37889 & new_new_n43799__;
  assign new_new_n47452__ = ys__n18723 & ~new_new_n43803__;
  assign new_new_n47453__ = ~new_new_n47451__ & ~new_new_n47452__;
  assign ys__n32549 = ~new_new_n43806__ & ~new_new_n47453__;
  assign new_new_n47455__ = ys__n37890 & new_new_n43799__;
  assign new_new_n47456__ = ys__n18726 & ~new_new_n43803__;
  assign new_new_n47457__ = ~new_new_n47455__ & ~new_new_n47456__;
  assign ys__n32550 = ~new_new_n43806__ & ~new_new_n47457__;
  assign new_new_n47459__ = ys__n37891 & new_new_n43799__;
  assign new_new_n47460__ = ys__n18729 & ~new_new_n43803__;
  assign new_new_n47461__ = ~new_new_n47459__ & ~new_new_n47460__;
  assign ys__n32551 = ~new_new_n43806__ & ~new_new_n47461__;
  assign new_new_n47463__ = ys__n37892 & new_new_n43799__;
  assign new_new_n47464__ = ys__n18732 & ~new_new_n43803__;
  assign new_new_n47465__ = ~new_new_n47463__ & ~new_new_n47464__;
  assign ys__n32552 = ~new_new_n43806__ & ~new_new_n47465__;
  assign new_new_n47467__ = ys__n37893 & new_new_n43799__;
  assign new_new_n47468__ = ys__n18735 & ~new_new_n43803__;
  assign new_new_n47469__ = ~new_new_n47467__ & ~new_new_n47468__;
  assign ys__n32553 = ~new_new_n43806__ & ~new_new_n47469__;
  assign new_new_n47471__ = ys__n37894 & new_new_n43799__;
  assign new_new_n47472__ = ys__n18738 & ~new_new_n43803__;
  assign new_new_n47473__ = ~new_new_n47471__ & ~new_new_n47472__;
  assign ys__n32554 = ~new_new_n43806__ & ~new_new_n47473__;
  assign new_new_n47475__ = ys__n37895 & new_new_n43799__;
  assign new_new_n47476__ = ys__n18741 & ~new_new_n43803__;
  assign new_new_n47477__ = ~new_new_n47475__ & ~new_new_n47476__;
  assign ys__n32555 = ~new_new_n43806__ & ~new_new_n47477__;
  assign new_new_n47479__ = ys__n37896 & new_new_n43799__;
  assign new_new_n47480__ = ys__n18744 & ~new_new_n43803__;
  assign new_new_n47481__ = ~new_new_n47479__ & ~new_new_n47480__;
  assign ys__n32556 = ~new_new_n43806__ & ~new_new_n47481__;
  assign new_new_n47483__ = ys__n37897 & new_new_n43799__;
  assign new_new_n47484__ = ys__n18747 & ~new_new_n43803__;
  assign new_new_n47485__ = ~new_new_n47483__ & ~new_new_n47484__;
  assign ys__n32557 = ~new_new_n43806__ & ~new_new_n47485__;
  assign new_new_n47487__ = ys__n48114 & new_new_n43654__;
  assign new_new_n47488__ = ys__n18654 & ~new_new_n43658__;
  assign new_new_n47489__ = ~new_new_n47487__ & ~new_new_n47488__;
  assign ys__n32558 = ~new_new_n43661__ & ~new_new_n47489__;
  assign new_new_n47491__ = ys__n48115 & new_new_n43654__;
  assign new_new_n47492__ = ys__n18657 & ~new_new_n43658__;
  assign new_new_n47493__ = ~new_new_n47491__ & ~new_new_n47492__;
  assign ys__n32559 = ~new_new_n43661__ & ~new_new_n47493__;
  assign new_new_n47495__ = ys__n48116 & new_new_n43654__;
  assign new_new_n47496__ = ys__n18660 & ~new_new_n43658__;
  assign new_new_n47497__ = ~new_new_n47495__ & ~new_new_n47496__;
  assign ys__n32560 = ~new_new_n43661__ & ~new_new_n47497__;
  assign new_new_n47499__ = ys__n48117 & new_new_n43654__;
  assign new_new_n47500__ = ys__n18663 & ~new_new_n43658__;
  assign new_new_n47501__ = ~new_new_n47499__ & ~new_new_n47500__;
  assign ys__n32561 = ~new_new_n43661__ & ~new_new_n47501__;
  assign new_new_n47503__ = ys__n37898 & new_new_n43654__;
  assign new_new_n47504__ = ys__n18666 & ~new_new_n43658__;
  assign new_new_n47505__ = ~new_new_n47503__ & ~new_new_n47504__;
  assign ys__n32562 = ~new_new_n43661__ & ~new_new_n47505__;
  assign new_new_n47507__ = ys__n37899 & new_new_n43654__;
  assign new_new_n47508__ = ys__n18669 & ~new_new_n43658__;
  assign new_new_n47509__ = ~new_new_n47507__ & ~new_new_n47508__;
  assign ys__n32563 = ~new_new_n43661__ & ~new_new_n47509__;
  assign new_new_n47511__ = ys__n37900 & new_new_n43654__;
  assign new_new_n47512__ = ys__n18672 & ~new_new_n43658__;
  assign new_new_n47513__ = ~new_new_n47511__ & ~new_new_n47512__;
  assign ys__n32564 = ~new_new_n43661__ & ~new_new_n47513__;
  assign new_new_n47515__ = ys__n37901 & new_new_n43654__;
  assign new_new_n47516__ = ys__n18675 & ~new_new_n43658__;
  assign new_new_n47517__ = ~new_new_n47515__ & ~new_new_n47516__;
  assign ys__n32565 = ~new_new_n43661__ & ~new_new_n47517__;
  assign new_new_n47519__ = ys__n37902 & new_new_n43654__;
  assign new_new_n47520__ = ys__n18678 & ~new_new_n43658__;
  assign new_new_n47521__ = ~new_new_n47519__ & ~new_new_n47520__;
  assign ys__n32566 = ~new_new_n43661__ & ~new_new_n47521__;
  assign new_new_n47523__ = ys__n37903 & new_new_n43654__;
  assign new_new_n47524__ = ys__n18681 & ~new_new_n43658__;
  assign new_new_n47525__ = ~new_new_n47523__ & ~new_new_n47524__;
  assign ys__n32567 = ~new_new_n43661__ & ~new_new_n47525__;
  assign new_new_n47527__ = ys__n37904 & new_new_n43654__;
  assign new_new_n47528__ = ys__n18684 & ~new_new_n43658__;
  assign new_new_n47529__ = ~new_new_n47527__ & ~new_new_n47528__;
  assign ys__n32568 = ~new_new_n43661__ & ~new_new_n47529__;
  assign new_new_n47531__ = ys__n37905 & new_new_n43654__;
  assign new_new_n47532__ = ys__n18687 & ~new_new_n43658__;
  assign new_new_n47533__ = ~new_new_n47531__ & ~new_new_n47532__;
  assign ys__n32569 = ~new_new_n43661__ & ~new_new_n47533__;
  assign new_new_n47535__ = ys__n37906 & new_new_n43654__;
  assign new_new_n47536__ = ys__n18690 & ~new_new_n43658__;
  assign new_new_n47537__ = ~new_new_n47535__ & ~new_new_n47536__;
  assign ys__n32570 = ~new_new_n43661__ & ~new_new_n47537__;
  assign new_new_n47539__ = ys__n37907 & new_new_n43654__;
  assign new_new_n47540__ = ys__n18693 & ~new_new_n43658__;
  assign new_new_n47541__ = ~new_new_n47539__ & ~new_new_n47540__;
  assign ys__n32571 = ~new_new_n43661__ & ~new_new_n47541__;
  assign new_new_n47543__ = ys__n37908 & new_new_n43654__;
  assign new_new_n47544__ = ys__n18696 & ~new_new_n43658__;
  assign new_new_n47545__ = ~new_new_n47543__ & ~new_new_n47544__;
  assign ys__n32572 = ~new_new_n43661__ & ~new_new_n47545__;
  assign new_new_n47547__ = ys__n37909 & new_new_n43654__;
  assign new_new_n47548__ = ys__n18699 & ~new_new_n43658__;
  assign new_new_n47549__ = ~new_new_n47547__ & ~new_new_n47548__;
  assign ys__n32573 = ~new_new_n43661__ & ~new_new_n47549__;
  assign new_new_n47551__ = ys__n37910 & new_new_n43654__;
  assign new_new_n47552__ = ys__n18702 & ~new_new_n43658__;
  assign new_new_n47553__ = ~new_new_n47551__ & ~new_new_n47552__;
  assign ys__n32574 = ~new_new_n43661__ & ~new_new_n47553__;
  assign new_new_n47555__ = ys__n37911 & new_new_n43654__;
  assign new_new_n47556__ = ys__n18705 & ~new_new_n43658__;
  assign new_new_n47557__ = ~new_new_n47555__ & ~new_new_n47556__;
  assign ys__n32575 = ~new_new_n43661__ & ~new_new_n47557__;
  assign new_new_n47559__ = ys__n37912 & new_new_n43654__;
  assign new_new_n47560__ = ys__n18708 & ~new_new_n43658__;
  assign new_new_n47561__ = ~new_new_n47559__ & ~new_new_n47560__;
  assign ys__n32576 = ~new_new_n43661__ & ~new_new_n47561__;
  assign new_new_n47563__ = ys__n37913 & new_new_n43654__;
  assign new_new_n47564__ = ys__n18711 & ~new_new_n43658__;
  assign new_new_n47565__ = ~new_new_n47563__ & ~new_new_n47564__;
  assign ys__n32577 = ~new_new_n43661__ & ~new_new_n47565__;
  assign new_new_n47567__ = ys__n37914 & new_new_n43654__;
  assign new_new_n47568__ = ys__n18714 & ~new_new_n43658__;
  assign new_new_n47569__ = ~new_new_n47567__ & ~new_new_n47568__;
  assign ys__n32578 = ~new_new_n43661__ & ~new_new_n47569__;
  assign new_new_n47571__ = ys__n37915 & new_new_n43654__;
  assign new_new_n47572__ = ys__n18717 & ~new_new_n43658__;
  assign new_new_n47573__ = ~new_new_n47571__ & ~new_new_n47572__;
  assign ys__n32579 = ~new_new_n43661__ & ~new_new_n47573__;
  assign new_new_n47575__ = ys__n37916 & new_new_n43654__;
  assign new_new_n47576__ = ys__n18720 & ~new_new_n43658__;
  assign new_new_n47577__ = ~new_new_n47575__ & ~new_new_n47576__;
  assign ys__n32580 = ~new_new_n43661__ & ~new_new_n47577__;
  assign new_new_n47579__ = ys__n37917 & new_new_n43654__;
  assign new_new_n47580__ = ys__n18723 & ~new_new_n43658__;
  assign new_new_n47581__ = ~new_new_n47579__ & ~new_new_n47580__;
  assign ys__n32581 = ~new_new_n43661__ & ~new_new_n47581__;
  assign new_new_n47583__ = ys__n37918 & new_new_n43654__;
  assign new_new_n47584__ = ys__n18726 & ~new_new_n43658__;
  assign new_new_n47585__ = ~new_new_n47583__ & ~new_new_n47584__;
  assign ys__n32582 = ~new_new_n43661__ & ~new_new_n47585__;
  assign new_new_n47587__ = ys__n37919 & new_new_n43654__;
  assign new_new_n47588__ = ys__n18729 & ~new_new_n43658__;
  assign new_new_n47589__ = ~new_new_n47587__ & ~new_new_n47588__;
  assign ys__n32583 = ~new_new_n43661__ & ~new_new_n47589__;
  assign new_new_n47591__ = ys__n37920 & new_new_n43654__;
  assign new_new_n47592__ = ys__n18732 & ~new_new_n43658__;
  assign new_new_n47593__ = ~new_new_n47591__ & ~new_new_n47592__;
  assign ys__n32584 = ~new_new_n43661__ & ~new_new_n47593__;
  assign new_new_n47595__ = ys__n37921 & new_new_n43654__;
  assign new_new_n47596__ = ys__n18735 & ~new_new_n43658__;
  assign new_new_n47597__ = ~new_new_n47595__ & ~new_new_n47596__;
  assign ys__n32585 = ~new_new_n43661__ & ~new_new_n47597__;
  assign new_new_n47599__ = ys__n37922 & new_new_n43654__;
  assign new_new_n47600__ = ys__n18738 & ~new_new_n43658__;
  assign new_new_n47601__ = ~new_new_n47599__ & ~new_new_n47600__;
  assign ys__n32586 = ~new_new_n43661__ & ~new_new_n47601__;
  assign new_new_n47603__ = ys__n37923 & new_new_n43654__;
  assign new_new_n47604__ = ys__n18741 & ~new_new_n43658__;
  assign new_new_n47605__ = ~new_new_n47603__ & ~new_new_n47604__;
  assign ys__n32587 = ~new_new_n43661__ & ~new_new_n47605__;
  assign new_new_n47607__ = ys__n37924 & new_new_n43654__;
  assign new_new_n47608__ = ys__n18744 & ~new_new_n43658__;
  assign new_new_n47609__ = ~new_new_n47607__ & ~new_new_n47608__;
  assign ys__n32588 = ~new_new_n43661__ & ~new_new_n47609__;
  assign new_new_n47611__ = ys__n37925 & new_new_n43654__;
  assign new_new_n47612__ = ys__n18747 & ~new_new_n43658__;
  assign new_new_n47613__ = ~new_new_n47611__ & ~new_new_n47612__;
  assign ys__n32589 = ~new_new_n43661__ & ~new_new_n47613__;
  assign new_new_n47615__ = ys__n48118 & new_new_n43509__;
  assign new_new_n47616__ = ys__n18654 & ~new_new_n43513__;
  assign new_new_n47617__ = ~new_new_n47615__ & ~new_new_n47616__;
  assign ys__n32590 = ~new_new_n43516__ & ~new_new_n47617__;
  assign new_new_n47619__ = ys__n48119 & new_new_n43509__;
  assign new_new_n47620__ = ys__n18657 & ~new_new_n43513__;
  assign new_new_n47621__ = ~new_new_n47619__ & ~new_new_n47620__;
  assign ys__n32591 = ~new_new_n43516__ & ~new_new_n47621__;
  assign new_new_n47623__ = ys__n48120 & new_new_n43509__;
  assign new_new_n47624__ = ys__n18660 & ~new_new_n43513__;
  assign new_new_n47625__ = ~new_new_n47623__ & ~new_new_n47624__;
  assign ys__n32592 = ~new_new_n43516__ & ~new_new_n47625__;
  assign new_new_n47627__ = ys__n48121 & new_new_n43509__;
  assign new_new_n47628__ = ys__n18663 & ~new_new_n43513__;
  assign new_new_n47629__ = ~new_new_n47627__ & ~new_new_n47628__;
  assign ys__n32593 = ~new_new_n43516__ & ~new_new_n47629__;
  assign new_new_n47631__ = ys__n37926 & new_new_n43509__;
  assign new_new_n47632__ = ys__n18666 & ~new_new_n43513__;
  assign new_new_n47633__ = ~new_new_n47631__ & ~new_new_n47632__;
  assign ys__n32594 = ~new_new_n43516__ & ~new_new_n47633__;
  assign new_new_n47635__ = ys__n37927 & new_new_n43509__;
  assign new_new_n47636__ = ys__n18669 & ~new_new_n43513__;
  assign new_new_n47637__ = ~new_new_n47635__ & ~new_new_n47636__;
  assign ys__n32595 = ~new_new_n43516__ & ~new_new_n47637__;
  assign new_new_n47639__ = ys__n37928 & new_new_n43509__;
  assign new_new_n47640__ = ys__n18672 & ~new_new_n43513__;
  assign new_new_n47641__ = ~new_new_n47639__ & ~new_new_n47640__;
  assign ys__n32596 = ~new_new_n43516__ & ~new_new_n47641__;
  assign new_new_n47643__ = ys__n37929 & new_new_n43509__;
  assign new_new_n47644__ = ys__n18675 & ~new_new_n43513__;
  assign new_new_n47645__ = ~new_new_n47643__ & ~new_new_n47644__;
  assign ys__n32597 = ~new_new_n43516__ & ~new_new_n47645__;
  assign new_new_n47647__ = ys__n37930 & new_new_n43509__;
  assign new_new_n47648__ = ys__n18678 & ~new_new_n43513__;
  assign new_new_n47649__ = ~new_new_n47647__ & ~new_new_n47648__;
  assign ys__n32598 = ~new_new_n43516__ & ~new_new_n47649__;
  assign new_new_n47651__ = ys__n37931 & new_new_n43509__;
  assign new_new_n47652__ = ys__n18681 & ~new_new_n43513__;
  assign new_new_n47653__ = ~new_new_n47651__ & ~new_new_n47652__;
  assign ys__n32599 = ~new_new_n43516__ & ~new_new_n47653__;
  assign new_new_n47655__ = ys__n37932 & new_new_n43509__;
  assign new_new_n47656__ = ys__n18684 & ~new_new_n43513__;
  assign new_new_n47657__ = ~new_new_n47655__ & ~new_new_n47656__;
  assign ys__n32600 = ~new_new_n43516__ & ~new_new_n47657__;
  assign new_new_n47659__ = ys__n37933 & new_new_n43509__;
  assign new_new_n47660__ = ys__n18687 & ~new_new_n43513__;
  assign new_new_n47661__ = ~new_new_n47659__ & ~new_new_n47660__;
  assign ys__n32601 = ~new_new_n43516__ & ~new_new_n47661__;
  assign new_new_n47663__ = ys__n37934 & new_new_n43509__;
  assign new_new_n47664__ = ys__n18690 & ~new_new_n43513__;
  assign new_new_n47665__ = ~new_new_n47663__ & ~new_new_n47664__;
  assign ys__n32602 = ~new_new_n43516__ & ~new_new_n47665__;
  assign new_new_n47667__ = ys__n37935 & new_new_n43509__;
  assign new_new_n47668__ = ys__n18693 & ~new_new_n43513__;
  assign new_new_n47669__ = ~new_new_n47667__ & ~new_new_n47668__;
  assign ys__n32603 = ~new_new_n43516__ & ~new_new_n47669__;
  assign new_new_n47671__ = ys__n37936 & new_new_n43509__;
  assign new_new_n47672__ = ys__n18696 & ~new_new_n43513__;
  assign new_new_n47673__ = ~new_new_n47671__ & ~new_new_n47672__;
  assign ys__n32604 = ~new_new_n43516__ & ~new_new_n47673__;
  assign new_new_n47675__ = ys__n37937 & new_new_n43509__;
  assign new_new_n47676__ = ys__n18699 & ~new_new_n43513__;
  assign new_new_n47677__ = ~new_new_n47675__ & ~new_new_n47676__;
  assign ys__n32605 = ~new_new_n43516__ & ~new_new_n47677__;
  assign new_new_n47679__ = ys__n37938 & new_new_n43509__;
  assign new_new_n47680__ = ys__n18702 & ~new_new_n43513__;
  assign new_new_n47681__ = ~new_new_n47679__ & ~new_new_n47680__;
  assign ys__n32606 = ~new_new_n43516__ & ~new_new_n47681__;
  assign new_new_n47683__ = ys__n37939 & new_new_n43509__;
  assign new_new_n47684__ = ys__n18705 & ~new_new_n43513__;
  assign new_new_n47685__ = ~new_new_n47683__ & ~new_new_n47684__;
  assign ys__n32607 = ~new_new_n43516__ & ~new_new_n47685__;
  assign new_new_n47687__ = ys__n37940 & new_new_n43509__;
  assign new_new_n47688__ = ys__n18708 & ~new_new_n43513__;
  assign new_new_n47689__ = ~new_new_n47687__ & ~new_new_n47688__;
  assign ys__n32608 = ~new_new_n43516__ & ~new_new_n47689__;
  assign new_new_n47691__ = ys__n37941 & new_new_n43509__;
  assign new_new_n47692__ = ys__n18711 & ~new_new_n43513__;
  assign new_new_n47693__ = ~new_new_n47691__ & ~new_new_n47692__;
  assign ys__n32609 = ~new_new_n43516__ & ~new_new_n47693__;
  assign new_new_n47695__ = ys__n37942 & new_new_n43509__;
  assign new_new_n47696__ = ys__n18714 & ~new_new_n43513__;
  assign new_new_n47697__ = ~new_new_n47695__ & ~new_new_n47696__;
  assign ys__n32610 = ~new_new_n43516__ & ~new_new_n47697__;
  assign new_new_n47699__ = ys__n37943 & new_new_n43509__;
  assign new_new_n47700__ = ys__n18717 & ~new_new_n43513__;
  assign new_new_n47701__ = ~new_new_n47699__ & ~new_new_n47700__;
  assign ys__n32611 = ~new_new_n43516__ & ~new_new_n47701__;
  assign new_new_n47703__ = ys__n37944 & new_new_n43509__;
  assign new_new_n47704__ = ys__n18720 & ~new_new_n43513__;
  assign new_new_n47705__ = ~new_new_n47703__ & ~new_new_n47704__;
  assign ys__n32612 = ~new_new_n43516__ & ~new_new_n47705__;
  assign new_new_n47707__ = ys__n37945 & new_new_n43509__;
  assign new_new_n47708__ = ys__n18723 & ~new_new_n43513__;
  assign new_new_n47709__ = ~new_new_n47707__ & ~new_new_n47708__;
  assign ys__n32613 = ~new_new_n43516__ & ~new_new_n47709__;
  assign new_new_n47711__ = ys__n37946 & new_new_n43509__;
  assign new_new_n47712__ = ys__n18726 & ~new_new_n43513__;
  assign new_new_n47713__ = ~new_new_n47711__ & ~new_new_n47712__;
  assign ys__n32614 = ~new_new_n43516__ & ~new_new_n47713__;
  assign new_new_n47715__ = ys__n37947 & new_new_n43509__;
  assign new_new_n47716__ = ys__n18729 & ~new_new_n43513__;
  assign new_new_n47717__ = ~new_new_n47715__ & ~new_new_n47716__;
  assign ys__n32615 = ~new_new_n43516__ & ~new_new_n47717__;
  assign new_new_n47719__ = ys__n37948 & new_new_n43509__;
  assign new_new_n47720__ = ys__n18732 & ~new_new_n43513__;
  assign new_new_n47721__ = ~new_new_n47719__ & ~new_new_n47720__;
  assign ys__n32616 = ~new_new_n43516__ & ~new_new_n47721__;
  assign new_new_n47723__ = ys__n37949 & new_new_n43509__;
  assign new_new_n47724__ = ys__n18735 & ~new_new_n43513__;
  assign new_new_n47725__ = ~new_new_n47723__ & ~new_new_n47724__;
  assign ys__n32617 = ~new_new_n43516__ & ~new_new_n47725__;
  assign new_new_n47727__ = ys__n37950 & new_new_n43509__;
  assign new_new_n47728__ = ys__n18738 & ~new_new_n43513__;
  assign new_new_n47729__ = ~new_new_n47727__ & ~new_new_n47728__;
  assign ys__n32618 = ~new_new_n43516__ & ~new_new_n47729__;
  assign new_new_n47731__ = ys__n37951 & new_new_n43509__;
  assign new_new_n47732__ = ys__n18741 & ~new_new_n43513__;
  assign new_new_n47733__ = ~new_new_n47731__ & ~new_new_n47732__;
  assign ys__n32619 = ~new_new_n43516__ & ~new_new_n47733__;
  assign new_new_n47735__ = ys__n37952 & new_new_n43509__;
  assign new_new_n47736__ = ys__n18744 & ~new_new_n43513__;
  assign new_new_n47737__ = ~new_new_n47735__ & ~new_new_n47736__;
  assign ys__n32620 = ~new_new_n43516__ & ~new_new_n47737__;
  assign new_new_n47739__ = ys__n37953 & new_new_n43509__;
  assign new_new_n47740__ = ys__n18747 & ~new_new_n43513__;
  assign new_new_n47741__ = ~new_new_n47739__ & ~new_new_n47740__;
  assign ys__n32621 = ~new_new_n43516__ & ~new_new_n47741__;
  assign new_new_n47743__ = ys__n48122 & new_new_n43364__;
  assign new_new_n47744__ = ys__n18654 & ~new_new_n43368__;
  assign new_new_n47745__ = ~new_new_n47743__ & ~new_new_n47744__;
  assign ys__n32622 = ~new_new_n43371__ & ~new_new_n47745__;
  assign new_new_n47747__ = ys__n48123 & new_new_n43364__;
  assign new_new_n47748__ = ys__n18657 & ~new_new_n43368__;
  assign new_new_n47749__ = ~new_new_n47747__ & ~new_new_n47748__;
  assign ys__n32623 = ~new_new_n43371__ & ~new_new_n47749__;
  assign new_new_n47751__ = ys__n48124 & new_new_n43364__;
  assign new_new_n47752__ = ys__n18660 & ~new_new_n43368__;
  assign new_new_n47753__ = ~new_new_n47751__ & ~new_new_n47752__;
  assign ys__n32624 = ~new_new_n43371__ & ~new_new_n47753__;
  assign new_new_n47755__ = ys__n48125 & new_new_n43364__;
  assign new_new_n47756__ = ys__n18663 & ~new_new_n43368__;
  assign new_new_n47757__ = ~new_new_n47755__ & ~new_new_n47756__;
  assign ys__n32625 = ~new_new_n43371__ & ~new_new_n47757__;
  assign new_new_n47759__ = ys__n37954 & new_new_n43364__;
  assign new_new_n47760__ = ys__n18666 & ~new_new_n43368__;
  assign new_new_n47761__ = ~new_new_n47759__ & ~new_new_n47760__;
  assign ys__n32626 = ~new_new_n43371__ & ~new_new_n47761__;
  assign new_new_n47763__ = ys__n37955 & new_new_n43364__;
  assign new_new_n47764__ = ys__n18669 & ~new_new_n43368__;
  assign new_new_n47765__ = ~new_new_n47763__ & ~new_new_n47764__;
  assign ys__n32627 = ~new_new_n43371__ & ~new_new_n47765__;
  assign new_new_n47767__ = ys__n37956 & new_new_n43364__;
  assign new_new_n47768__ = ys__n18672 & ~new_new_n43368__;
  assign new_new_n47769__ = ~new_new_n47767__ & ~new_new_n47768__;
  assign ys__n32628 = ~new_new_n43371__ & ~new_new_n47769__;
  assign new_new_n47771__ = ys__n37957 & new_new_n43364__;
  assign new_new_n47772__ = ys__n18675 & ~new_new_n43368__;
  assign new_new_n47773__ = ~new_new_n47771__ & ~new_new_n47772__;
  assign ys__n32629 = ~new_new_n43371__ & ~new_new_n47773__;
  assign new_new_n47775__ = ys__n37958 & new_new_n43364__;
  assign new_new_n47776__ = ys__n18678 & ~new_new_n43368__;
  assign new_new_n47777__ = ~new_new_n47775__ & ~new_new_n47776__;
  assign ys__n32630 = ~new_new_n43371__ & ~new_new_n47777__;
  assign new_new_n47779__ = ys__n37959 & new_new_n43364__;
  assign new_new_n47780__ = ys__n18681 & ~new_new_n43368__;
  assign new_new_n47781__ = ~new_new_n47779__ & ~new_new_n47780__;
  assign ys__n32631 = ~new_new_n43371__ & ~new_new_n47781__;
  assign new_new_n47783__ = ys__n37960 & new_new_n43364__;
  assign new_new_n47784__ = ys__n18684 & ~new_new_n43368__;
  assign new_new_n47785__ = ~new_new_n47783__ & ~new_new_n47784__;
  assign ys__n32632 = ~new_new_n43371__ & ~new_new_n47785__;
  assign new_new_n47787__ = ys__n37961 & new_new_n43364__;
  assign new_new_n47788__ = ys__n18687 & ~new_new_n43368__;
  assign new_new_n47789__ = ~new_new_n47787__ & ~new_new_n47788__;
  assign ys__n32633 = ~new_new_n43371__ & ~new_new_n47789__;
  assign new_new_n47791__ = ys__n37962 & new_new_n43364__;
  assign new_new_n47792__ = ys__n18690 & ~new_new_n43368__;
  assign new_new_n47793__ = ~new_new_n47791__ & ~new_new_n47792__;
  assign ys__n32634 = ~new_new_n43371__ & ~new_new_n47793__;
  assign new_new_n47795__ = ys__n37963 & new_new_n43364__;
  assign new_new_n47796__ = ys__n18693 & ~new_new_n43368__;
  assign new_new_n47797__ = ~new_new_n47795__ & ~new_new_n47796__;
  assign ys__n32635 = ~new_new_n43371__ & ~new_new_n47797__;
  assign new_new_n47799__ = ys__n37964 & new_new_n43364__;
  assign new_new_n47800__ = ys__n18696 & ~new_new_n43368__;
  assign new_new_n47801__ = ~new_new_n47799__ & ~new_new_n47800__;
  assign ys__n32636 = ~new_new_n43371__ & ~new_new_n47801__;
  assign new_new_n47803__ = ys__n37965 & new_new_n43364__;
  assign new_new_n47804__ = ys__n18699 & ~new_new_n43368__;
  assign new_new_n47805__ = ~new_new_n47803__ & ~new_new_n47804__;
  assign ys__n32637 = ~new_new_n43371__ & ~new_new_n47805__;
  assign new_new_n47807__ = ys__n37966 & new_new_n43364__;
  assign new_new_n47808__ = ys__n18702 & ~new_new_n43368__;
  assign new_new_n47809__ = ~new_new_n47807__ & ~new_new_n47808__;
  assign ys__n32638 = ~new_new_n43371__ & ~new_new_n47809__;
  assign new_new_n47811__ = ys__n37967 & new_new_n43364__;
  assign new_new_n47812__ = ys__n18705 & ~new_new_n43368__;
  assign new_new_n47813__ = ~new_new_n47811__ & ~new_new_n47812__;
  assign ys__n32639 = ~new_new_n43371__ & ~new_new_n47813__;
  assign new_new_n47815__ = ys__n37968 & new_new_n43364__;
  assign new_new_n47816__ = ys__n18708 & ~new_new_n43368__;
  assign new_new_n47817__ = ~new_new_n47815__ & ~new_new_n47816__;
  assign ys__n32640 = ~new_new_n43371__ & ~new_new_n47817__;
  assign new_new_n47819__ = ys__n37969 & new_new_n43364__;
  assign new_new_n47820__ = ys__n18711 & ~new_new_n43368__;
  assign new_new_n47821__ = ~new_new_n47819__ & ~new_new_n47820__;
  assign ys__n32641 = ~new_new_n43371__ & ~new_new_n47821__;
  assign new_new_n47823__ = ys__n37970 & new_new_n43364__;
  assign new_new_n47824__ = ys__n18714 & ~new_new_n43368__;
  assign new_new_n47825__ = ~new_new_n47823__ & ~new_new_n47824__;
  assign ys__n32642 = ~new_new_n43371__ & ~new_new_n47825__;
  assign new_new_n47827__ = ys__n37971 & new_new_n43364__;
  assign new_new_n47828__ = ys__n18717 & ~new_new_n43368__;
  assign new_new_n47829__ = ~new_new_n47827__ & ~new_new_n47828__;
  assign ys__n32643 = ~new_new_n43371__ & ~new_new_n47829__;
  assign new_new_n47831__ = ys__n37972 & new_new_n43364__;
  assign new_new_n47832__ = ys__n18720 & ~new_new_n43368__;
  assign new_new_n47833__ = ~new_new_n47831__ & ~new_new_n47832__;
  assign ys__n32644 = ~new_new_n43371__ & ~new_new_n47833__;
  assign new_new_n47835__ = ys__n37973 & new_new_n43364__;
  assign new_new_n47836__ = ys__n18723 & ~new_new_n43368__;
  assign new_new_n47837__ = ~new_new_n47835__ & ~new_new_n47836__;
  assign ys__n32645 = ~new_new_n43371__ & ~new_new_n47837__;
  assign new_new_n47839__ = ys__n37974 & new_new_n43364__;
  assign new_new_n47840__ = ys__n18726 & ~new_new_n43368__;
  assign new_new_n47841__ = ~new_new_n47839__ & ~new_new_n47840__;
  assign ys__n32646 = ~new_new_n43371__ & ~new_new_n47841__;
  assign new_new_n47843__ = ys__n37975 & new_new_n43364__;
  assign new_new_n47844__ = ys__n18729 & ~new_new_n43368__;
  assign new_new_n47845__ = ~new_new_n47843__ & ~new_new_n47844__;
  assign ys__n32647 = ~new_new_n43371__ & ~new_new_n47845__;
  assign new_new_n47847__ = ys__n37976 & new_new_n43364__;
  assign new_new_n47848__ = ys__n18732 & ~new_new_n43368__;
  assign new_new_n47849__ = ~new_new_n47847__ & ~new_new_n47848__;
  assign ys__n32648 = ~new_new_n43371__ & ~new_new_n47849__;
  assign new_new_n47851__ = ys__n37977 & new_new_n43364__;
  assign new_new_n47852__ = ys__n18735 & ~new_new_n43368__;
  assign new_new_n47853__ = ~new_new_n47851__ & ~new_new_n47852__;
  assign ys__n32649 = ~new_new_n43371__ & ~new_new_n47853__;
  assign new_new_n47855__ = ys__n37978 & new_new_n43364__;
  assign new_new_n47856__ = ys__n18738 & ~new_new_n43368__;
  assign new_new_n47857__ = ~new_new_n47855__ & ~new_new_n47856__;
  assign ys__n32650 = ~new_new_n43371__ & ~new_new_n47857__;
  assign new_new_n47859__ = ys__n37979 & new_new_n43364__;
  assign new_new_n47860__ = ys__n18741 & ~new_new_n43368__;
  assign new_new_n47861__ = ~new_new_n47859__ & ~new_new_n47860__;
  assign ys__n32651 = ~new_new_n43371__ & ~new_new_n47861__;
  assign new_new_n47863__ = ys__n37980 & new_new_n43364__;
  assign new_new_n47864__ = ys__n18744 & ~new_new_n43368__;
  assign new_new_n47865__ = ~new_new_n47863__ & ~new_new_n47864__;
  assign ys__n32652 = ~new_new_n43371__ & ~new_new_n47865__;
  assign new_new_n47867__ = ys__n37981 & new_new_n43364__;
  assign new_new_n47868__ = ys__n18747 & ~new_new_n43368__;
  assign new_new_n47869__ = ~new_new_n47867__ & ~new_new_n47868__;
  assign ys__n32653 = ~new_new_n43371__ & ~new_new_n47869__;
  assign new_new_n47871__ = ys__n48126 & new_new_n43219__;
  assign new_new_n47872__ = ys__n18654 & ~new_new_n43223__;
  assign new_new_n47873__ = ~new_new_n47871__ & ~new_new_n47872__;
  assign ys__n32654 = ~new_new_n43226__ & ~new_new_n47873__;
  assign new_new_n47875__ = ys__n48127 & new_new_n43219__;
  assign new_new_n47876__ = ys__n18657 & ~new_new_n43223__;
  assign new_new_n47877__ = ~new_new_n47875__ & ~new_new_n47876__;
  assign ys__n32655 = ~new_new_n43226__ & ~new_new_n47877__;
  assign new_new_n47879__ = ys__n48128 & new_new_n43219__;
  assign new_new_n47880__ = ys__n18660 & ~new_new_n43223__;
  assign new_new_n47881__ = ~new_new_n47879__ & ~new_new_n47880__;
  assign ys__n32656 = ~new_new_n43226__ & ~new_new_n47881__;
  assign new_new_n47883__ = ys__n48129 & new_new_n43219__;
  assign new_new_n47884__ = ys__n18663 & ~new_new_n43223__;
  assign new_new_n47885__ = ~new_new_n47883__ & ~new_new_n47884__;
  assign ys__n32657 = ~new_new_n43226__ & ~new_new_n47885__;
  assign new_new_n47887__ = ys__n37982 & new_new_n43219__;
  assign new_new_n47888__ = ys__n18666 & ~new_new_n43223__;
  assign new_new_n47889__ = ~new_new_n47887__ & ~new_new_n47888__;
  assign ys__n32658 = ~new_new_n43226__ & ~new_new_n47889__;
  assign new_new_n47891__ = ys__n37983 & new_new_n43219__;
  assign new_new_n47892__ = ys__n18669 & ~new_new_n43223__;
  assign new_new_n47893__ = ~new_new_n47891__ & ~new_new_n47892__;
  assign ys__n32659 = ~new_new_n43226__ & ~new_new_n47893__;
  assign new_new_n47895__ = ys__n37984 & new_new_n43219__;
  assign new_new_n47896__ = ys__n18672 & ~new_new_n43223__;
  assign new_new_n47897__ = ~new_new_n47895__ & ~new_new_n47896__;
  assign ys__n32660 = ~new_new_n43226__ & ~new_new_n47897__;
  assign new_new_n47899__ = ys__n37985 & new_new_n43219__;
  assign new_new_n47900__ = ys__n18675 & ~new_new_n43223__;
  assign new_new_n47901__ = ~new_new_n47899__ & ~new_new_n47900__;
  assign ys__n32661 = ~new_new_n43226__ & ~new_new_n47901__;
  assign new_new_n47903__ = ys__n37986 & new_new_n43219__;
  assign new_new_n47904__ = ys__n18678 & ~new_new_n43223__;
  assign new_new_n47905__ = ~new_new_n47903__ & ~new_new_n47904__;
  assign ys__n32662 = ~new_new_n43226__ & ~new_new_n47905__;
  assign new_new_n47907__ = ys__n37987 & new_new_n43219__;
  assign new_new_n47908__ = ys__n18681 & ~new_new_n43223__;
  assign new_new_n47909__ = ~new_new_n47907__ & ~new_new_n47908__;
  assign ys__n32663 = ~new_new_n43226__ & ~new_new_n47909__;
  assign new_new_n47911__ = ys__n37988 & new_new_n43219__;
  assign new_new_n47912__ = ys__n18684 & ~new_new_n43223__;
  assign new_new_n47913__ = ~new_new_n47911__ & ~new_new_n47912__;
  assign ys__n32664 = ~new_new_n43226__ & ~new_new_n47913__;
  assign new_new_n47915__ = ys__n37989 & new_new_n43219__;
  assign new_new_n47916__ = ys__n18687 & ~new_new_n43223__;
  assign new_new_n47917__ = ~new_new_n47915__ & ~new_new_n47916__;
  assign ys__n32665 = ~new_new_n43226__ & ~new_new_n47917__;
  assign new_new_n47919__ = ys__n37990 & new_new_n43219__;
  assign new_new_n47920__ = ys__n18690 & ~new_new_n43223__;
  assign new_new_n47921__ = ~new_new_n47919__ & ~new_new_n47920__;
  assign ys__n32666 = ~new_new_n43226__ & ~new_new_n47921__;
  assign new_new_n47923__ = ys__n37991 & new_new_n43219__;
  assign new_new_n47924__ = ys__n18693 & ~new_new_n43223__;
  assign new_new_n47925__ = ~new_new_n47923__ & ~new_new_n47924__;
  assign ys__n32667 = ~new_new_n43226__ & ~new_new_n47925__;
  assign new_new_n47927__ = ys__n37992 & new_new_n43219__;
  assign new_new_n47928__ = ys__n18696 & ~new_new_n43223__;
  assign new_new_n47929__ = ~new_new_n47927__ & ~new_new_n47928__;
  assign ys__n32668 = ~new_new_n43226__ & ~new_new_n47929__;
  assign new_new_n47931__ = ys__n37993 & new_new_n43219__;
  assign new_new_n47932__ = ys__n18699 & ~new_new_n43223__;
  assign new_new_n47933__ = ~new_new_n47931__ & ~new_new_n47932__;
  assign ys__n32669 = ~new_new_n43226__ & ~new_new_n47933__;
  assign new_new_n47935__ = ys__n37994 & new_new_n43219__;
  assign new_new_n47936__ = ys__n18702 & ~new_new_n43223__;
  assign new_new_n47937__ = ~new_new_n47935__ & ~new_new_n47936__;
  assign ys__n32670 = ~new_new_n43226__ & ~new_new_n47937__;
  assign new_new_n47939__ = ys__n37995 & new_new_n43219__;
  assign new_new_n47940__ = ys__n18705 & ~new_new_n43223__;
  assign new_new_n47941__ = ~new_new_n47939__ & ~new_new_n47940__;
  assign ys__n32671 = ~new_new_n43226__ & ~new_new_n47941__;
  assign new_new_n47943__ = ys__n37996 & new_new_n43219__;
  assign new_new_n47944__ = ys__n18708 & ~new_new_n43223__;
  assign new_new_n47945__ = ~new_new_n47943__ & ~new_new_n47944__;
  assign ys__n32672 = ~new_new_n43226__ & ~new_new_n47945__;
  assign new_new_n47947__ = ys__n37997 & new_new_n43219__;
  assign new_new_n47948__ = ys__n18711 & ~new_new_n43223__;
  assign new_new_n47949__ = ~new_new_n47947__ & ~new_new_n47948__;
  assign ys__n32673 = ~new_new_n43226__ & ~new_new_n47949__;
  assign new_new_n47951__ = ys__n37998 & new_new_n43219__;
  assign new_new_n47952__ = ys__n18714 & ~new_new_n43223__;
  assign new_new_n47953__ = ~new_new_n47951__ & ~new_new_n47952__;
  assign ys__n32674 = ~new_new_n43226__ & ~new_new_n47953__;
  assign new_new_n47955__ = ys__n37999 & new_new_n43219__;
  assign new_new_n47956__ = ys__n18717 & ~new_new_n43223__;
  assign new_new_n47957__ = ~new_new_n47955__ & ~new_new_n47956__;
  assign ys__n32675 = ~new_new_n43226__ & ~new_new_n47957__;
  assign new_new_n47959__ = ys__n38000 & new_new_n43219__;
  assign new_new_n47960__ = ys__n18720 & ~new_new_n43223__;
  assign new_new_n47961__ = ~new_new_n47959__ & ~new_new_n47960__;
  assign ys__n32676 = ~new_new_n43226__ & ~new_new_n47961__;
  assign new_new_n47963__ = ys__n38001 & new_new_n43219__;
  assign new_new_n47964__ = ys__n18723 & ~new_new_n43223__;
  assign new_new_n47965__ = ~new_new_n47963__ & ~new_new_n47964__;
  assign ys__n32677 = ~new_new_n43226__ & ~new_new_n47965__;
  assign new_new_n47967__ = ys__n38002 & new_new_n43219__;
  assign new_new_n47968__ = ys__n18726 & ~new_new_n43223__;
  assign new_new_n47969__ = ~new_new_n47967__ & ~new_new_n47968__;
  assign ys__n32678 = ~new_new_n43226__ & ~new_new_n47969__;
  assign new_new_n47971__ = ys__n38003 & new_new_n43219__;
  assign new_new_n47972__ = ys__n18729 & ~new_new_n43223__;
  assign new_new_n47973__ = ~new_new_n47971__ & ~new_new_n47972__;
  assign ys__n32679 = ~new_new_n43226__ & ~new_new_n47973__;
  assign new_new_n47975__ = ys__n38004 & new_new_n43219__;
  assign new_new_n47976__ = ys__n18732 & ~new_new_n43223__;
  assign new_new_n47977__ = ~new_new_n47975__ & ~new_new_n47976__;
  assign ys__n32680 = ~new_new_n43226__ & ~new_new_n47977__;
  assign new_new_n47979__ = ys__n38005 & new_new_n43219__;
  assign new_new_n47980__ = ys__n18735 & ~new_new_n43223__;
  assign new_new_n47981__ = ~new_new_n47979__ & ~new_new_n47980__;
  assign ys__n32681 = ~new_new_n43226__ & ~new_new_n47981__;
  assign new_new_n47983__ = ys__n38006 & new_new_n43219__;
  assign new_new_n47984__ = ys__n18738 & ~new_new_n43223__;
  assign new_new_n47985__ = ~new_new_n47983__ & ~new_new_n47984__;
  assign ys__n32682 = ~new_new_n43226__ & ~new_new_n47985__;
  assign new_new_n47987__ = ys__n38007 & new_new_n43219__;
  assign new_new_n47988__ = ys__n18741 & ~new_new_n43223__;
  assign new_new_n47989__ = ~new_new_n47987__ & ~new_new_n47988__;
  assign ys__n32683 = ~new_new_n43226__ & ~new_new_n47989__;
  assign new_new_n47991__ = ys__n38008 & new_new_n43219__;
  assign new_new_n47992__ = ys__n18744 & ~new_new_n43223__;
  assign new_new_n47993__ = ~new_new_n47991__ & ~new_new_n47992__;
  assign ys__n32684 = ~new_new_n43226__ & ~new_new_n47993__;
  assign new_new_n47995__ = ys__n38009 & new_new_n43219__;
  assign new_new_n47996__ = ys__n18747 & ~new_new_n43223__;
  assign new_new_n47997__ = ~new_new_n47995__ & ~new_new_n47996__;
  assign ys__n32685 = ~new_new_n43226__ & ~new_new_n47997__;
  assign new_new_n47999__ = ys__n48130 & new_new_n42895__;
  assign new_new_n48000__ = ys__n18654 & ~new_new_n42899__;
  assign new_new_n48001__ = ~new_new_n47999__ & ~new_new_n48000__;
  assign ys__n32686 = ~new_new_n42902__ & ~new_new_n48001__;
  assign new_new_n48003__ = ys__n48131 & new_new_n42895__;
  assign new_new_n48004__ = ys__n18657 & ~new_new_n42899__;
  assign new_new_n48005__ = ~new_new_n48003__ & ~new_new_n48004__;
  assign ys__n32687 = ~new_new_n42902__ & ~new_new_n48005__;
  assign new_new_n48007__ = ys__n48132 & new_new_n42895__;
  assign new_new_n48008__ = ys__n18660 & ~new_new_n42899__;
  assign new_new_n48009__ = ~new_new_n48007__ & ~new_new_n48008__;
  assign ys__n32688 = ~new_new_n42902__ & ~new_new_n48009__;
  assign new_new_n48011__ = ys__n48133 & new_new_n42895__;
  assign new_new_n48012__ = ys__n18663 & ~new_new_n42899__;
  assign new_new_n48013__ = ~new_new_n48011__ & ~new_new_n48012__;
  assign ys__n32689 = ~new_new_n42902__ & ~new_new_n48013__;
  assign new_new_n48015__ = ys__n38010 & new_new_n42895__;
  assign new_new_n48016__ = ys__n18666 & ~new_new_n42899__;
  assign new_new_n48017__ = ~new_new_n48015__ & ~new_new_n48016__;
  assign ys__n32690 = ~new_new_n42902__ & ~new_new_n48017__;
  assign new_new_n48019__ = ys__n38011 & new_new_n42895__;
  assign new_new_n48020__ = ys__n18669 & ~new_new_n42899__;
  assign new_new_n48021__ = ~new_new_n48019__ & ~new_new_n48020__;
  assign ys__n32691 = ~new_new_n42902__ & ~new_new_n48021__;
  assign new_new_n48023__ = ys__n38012 & new_new_n42895__;
  assign new_new_n48024__ = ys__n18672 & ~new_new_n42899__;
  assign new_new_n48025__ = ~new_new_n48023__ & ~new_new_n48024__;
  assign ys__n32692 = ~new_new_n42902__ & ~new_new_n48025__;
  assign new_new_n48027__ = ys__n38013 & new_new_n42895__;
  assign new_new_n48028__ = ys__n18675 & ~new_new_n42899__;
  assign new_new_n48029__ = ~new_new_n48027__ & ~new_new_n48028__;
  assign ys__n32693 = ~new_new_n42902__ & ~new_new_n48029__;
  assign new_new_n48031__ = ys__n38014 & new_new_n42895__;
  assign new_new_n48032__ = ys__n18678 & ~new_new_n42899__;
  assign new_new_n48033__ = ~new_new_n48031__ & ~new_new_n48032__;
  assign ys__n32694 = ~new_new_n42902__ & ~new_new_n48033__;
  assign new_new_n48035__ = ys__n38015 & new_new_n42895__;
  assign new_new_n48036__ = ys__n18681 & ~new_new_n42899__;
  assign new_new_n48037__ = ~new_new_n48035__ & ~new_new_n48036__;
  assign ys__n32695 = ~new_new_n42902__ & ~new_new_n48037__;
  assign new_new_n48039__ = ys__n38016 & new_new_n42895__;
  assign new_new_n48040__ = ys__n18684 & ~new_new_n42899__;
  assign new_new_n48041__ = ~new_new_n48039__ & ~new_new_n48040__;
  assign ys__n32696 = ~new_new_n42902__ & ~new_new_n48041__;
  assign new_new_n48043__ = ys__n38017 & new_new_n42895__;
  assign new_new_n48044__ = ys__n18687 & ~new_new_n42899__;
  assign new_new_n48045__ = ~new_new_n48043__ & ~new_new_n48044__;
  assign ys__n32697 = ~new_new_n42902__ & ~new_new_n48045__;
  assign new_new_n48047__ = ys__n38018 & new_new_n42895__;
  assign new_new_n48048__ = ys__n18690 & ~new_new_n42899__;
  assign new_new_n48049__ = ~new_new_n48047__ & ~new_new_n48048__;
  assign ys__n32698 = ~new_new_n42902__ & ~new_new_n48049__;
  assign new_new_n48051__ = ys__n38019 & new_new_n42895__;
  assign new_new_n48052__ = ys__n18693 & ~new_new_n42899__;
  assign new_new_n48053__ = ~new_new_n48051__ & ~new_new_n48052__;
  assign ys__n32699 = ~new_new_n42902__ & ~new_new_n48053__;
  assign new_new_n48055__ = ys__n38020 & new_new_n42895__;
  assign new_new_n48056__ = ys__n18696 & ~new_new_n42899__;
  assign new_new_n48057__ = ~new_new_n48055__ & ~new_new_n48056__;
  assign ys__n32700 = ~new_new_n42902__ & ~new_new_n48057__;
  assign new_new_n48059__ = ys__n38021 & new_new_n42895__;
  assign new_new_n48060__ = ys__n18699 & ~new_new_n42899__;
  assign new_new_n48061__ = ~new_new_n48059__ & ~new_new_n48060__;
  assign ys__n32701 = ~new_new_n42902__ & ~new_new_n48061__;
  assign new_new_n48063__ = ys__n38022 & new_new_n42895__;
  assign new_new_n48064__ = ys__n18702 & ~new_new_n42899__;
  assign new_new_n48065__ = ~new_new_n48063__ & ~new_new_n48064__;
  assign ys__n32702 = ~new_new_n42902__ & ~new_new_n48065__;
  assign new_new_n48067__ = ys__n38023 & new_new_n42895__;
  assign new_new_n48068__ = ys__n18705 & ~new_new_n42899__;
  assign new_new_n48069__ = ~new_new_n48067__ & ~new_new_n48068__;
  assign ys__n32703 = ~new_new_n42902__ & ~new_new_n48069__;
  assign new_new_n48071__ = ys__n38024 & new_new_n42895__;
  assign new_new_n48072__ = ys__n18708 & ~new_new_n42899__;
  assign new_new_n48073__ = ~new_new_n48071__ & ~new_new_n48072__;
  assign ys__n32704 = ~new_new_n42902__ & ~new_new_n48073__;
  assign new_new_n48075__ = ys__n38025 & new_new_n42895__;
  assign new_new_n48076__ = ys__n18711 & ~new_new_n42899__;
  assign new_new_n48077__ = ~new_new_n48075__ & ~new_new_n48076__;
  assign ys__n32705 = ~new_new_n42902__ & ~new_new_n48077__;
  assign new_new_n48079__ = ys__n38026 & new_new_n42895__;
  assign new_new_n48080__ = ys__n18714 & ~new_new_n42899__;
  assign new_new_n48081__ = ~new_new_n48079__ & ~new_new_n48080__;
  assign ys__n32706 = ~new_new_n42902__ & ~new_new_n48081__;
  assign new_new_n48083__ = ys__n38027 & new_new_n42895__;
  assign new_new_n48084__ = ys__n18717 & ~new_new_n42899__;
  assign new_new_n48085__ = ~new_new_n48083__ & ~new_new_n48084__;
  assign ys__n32707 = ~new_new_n42902__ & ~new_new_n48085__;
  assign new_new_n48087__ = ys__n38028 & new_new_n42895__;
  assign new_new_n48088__ = ys__n18720 & ~new_new_n42899__;
  assign new_new_n48089__ = ~new_new_n48087__ & ~new_new_n48088__;
  assign ys__n32708 = ~new_new_n42902__ & ~new_new_n48089__;
  assign new_new_n48091__ = ys__n38029 & new_new_n42895__;
  assign new_new_n48092__ = ys__n18723 & ~new_new_n42899__;
  assign new_new_n48093__ = ~new_new_n48091__ & ~new_new_n48092__;
  assign ys__n32709 = ~new_new_n42902__ & ~new_new_n48093__;
  assign new_new_n48095__ = ys__n38030 & new_new_n42895__;
  assign new_new_n48096__ = ys__n18726 & ~new_new_n42899__;
  assign new_new_n48097__ = ~new_new_n48095__ & ~new_new_n48096__;
  assign ys__n32710 = ~new_new_n42902__ & ~new_new_n48097__;
  assign new_new_n48099__ = ys__n38031 & new_new_n42895__;
  assign new_new_n48100__ = ys__n18729 & ~new_new_n42899__;
  assign new_new_n48101__ = ~new_new_n48099__ & ~new_new_n48100__;
  assign ys__n32711 = ~new_new_n42902__ & ~new_new_n48101__;
  assign new_new_n48103__ = ys__n38032 & new_new_n42895__;
  assign new_new_n48104__ = ys__n18732 & ~new_new_n42899__;
  assign new_new_n48105__ = ~new_new_n48103__ & ~new_new_n48104__;
  assign ys__n32712 = ~new_new_n42902__ & ~new_new_n48105__;
  assign new_new_n48107__ = ys__n38033 & new_new_n42895__;
  assign new_new_n48108__ = ys__n18735 & ~new_new_n42899__;
  assign new_new_n48109__ = ~new_new_n48107__ & ~new_new_n48108__;
  assign ys__n32713 = ~new_new_n42902__ & ~new_new_n48109__;
  assign new_new_n48111__ = ys__n38034 & new_new_n42895__;
  assign new_new_n48112__ = ys__n18738 & ~new_new_n42899__;
  assign new_new_n48113__ = ~new_new_n48111__ & ~new_new_n48112__;
  assign ys__n32714 = ~new_new_n42902__ & ~new_new_n48113__;
  assign new_new_n48115__ = ys__n38035 & new_new_n42895__;
  assign new_new_n48116__ = ys__n18741 & ~new_new_n42899__;
  assign new_new_n48117__ = ~new_new_n48115__ & ~new_new_n48116__;
  assign ys__n32715 = ~new_new_n42902__ & ~new_new_n48117__;
  assign new_new_n48119__ = ys__n38036 & new_new_n42895__;
  assign new_new_n48120__ = ys__n18744 & ~new_new_n42899__;
  assign new_new_n48121__ = ~new_new_n48119__ & ~new_new_n48120__;
  assign ys__n32716 = ~new_new_n42902__ & ~new_new_n48121__;
  assign new_new_n48123__ = ys__n38037 & new_new_n42895__;
  assign new_new_n48124__ = ys__n18747 & ~new_new_n42899__;
  assign new_new_n48125__ = ~new_new_n48123__ & ~new_new_n48124__;
  assign ys__n32717 = ~new_new_n42902__ & ~new_new_n48125__;
  assign new_new_n48127__ = ys__n48134 & new_new_n43040__;
  assign new_new_n48128__ = ys__n18654 & ~new_new_n43044__;
  assign new_new_n48129__ = ~new_new_n48127__ & ~new_new_n48128__;
  assign ys__n32718 = ~new_new_n43047__ & ~new_new_n48129__;
  assign new_new_n48131__ = ys__n48135 & new_new_n43040__;
  assign new_new_n48132__ = ys__n18657 & ~new_new_n43044__;
  assign new_new_n48133__ = ~new_new_n48131__ & ~new_new_n48132__;
  assign ys__n32719 = ~new_new_n43047__ & ~new_new_n48133__;
  assign new_new_n48135__ = ys__n48136 & new_new_n43040__;
  assign new_new_n48136__ = ys__n18660 & ~new_new_n43044__;
  assign new_new_n48137__ = ~new_new_n48135__ & ~new_new_n48136__;
  assign ys__n32720 = ~new_new_n43047__ & ~new_new_n48137__;
  assign new_new_n48139__ = ys__n48137 & new_new_n43040__;
  assign new_new_n48140__ = ys__n18663 & ~new_new_n43044__;
  assign new_new_n48141__ = ~new_new_n48139__ & ~new_new_n48140__;
  assign ys__n32721 = ~new_new_n43047__ & ~new_new_n48141__;
  assign new_new_n48143__ = ys__n38038 & new_new_n43040__;
  assign new_new_n48144__ = ys__n18666 & ~new_new_n43044__;
  assign new_new_n48145__ = ~new_new_n48143__ & ~new_new_n48144__;
  assign ys__n32722 = ~new_new_n43047__ & ~new_new_n48145__;
  assign new_new_n48147__ = ys__n38039 & new_new_n43040__;
  assign new_new_n48148__ = ys__n18669 & ~new_new_n43044__;
  assign new_new_n48149__ = ~new_new_n48147__ & ~new_new_n48148__;
  assign ys__n32723 = ~new_new_n43047__ & ~new_new_n48149__;
  assign new_new_n48151__ = ys__n38040 & new_new_n43040__;
  assign new_new_n48152__ = ys__n18672 & ~new_new_n43044__;
  assign new_new_n48153__ = ~new_new_n48151__ & ~new_new_n48152__;
  assign ys__n32724 = ~new_new_n43047__ & ~new_new_n48153__;
  assign new_new_n48155__ = ys__n38041 & new_new_n43040__;
  assign new_new_n48156__ = ys__n18675 & ~new_new_n43044__;
  assign new_new_n48157__ = ~new_new_n48155__ & ~new_new_n48156__;
  assign ys__n32725 = ~new_new_n43047__ & ~new_new_n48157__;
  assign new_new_n48159__ = ys__n38042 & new_new_n43040__;
  assign new_new_n48160__ = ys__n18678 & ~new_new_n43044__;
  assign new_new_n48161__ = ~new_new_n48159__ & ~new_new_n48160__;
  assign ys__n32726 = ~new_new_n43047__ & ~new_new_n48161__;
  assign new_new_n48163__ = ys__n38043 & new_new_n43040__;
  assign new_new_n48164__ = ys__n18681 & ~new_new_n43044__;
  assign new_new_n48165__ = ~new_new_n48163__ & ~new_new_n48164__;
  assign ys__n32727 = ~new_new_n43047__ & ~new_new_n48165__;
  assign new_new_n48167__ = ys__n38044 & new_new_n43040__;
  assign new_new_n48168__ = ys__n18684 & ~new_new_n43044__;
  assign new_new_n48169__ = ~new_new_n48167__ & ~new_new_n48168__;
  assign ys__n32728 = ~new_new_n43047__ & ~new_new_n48169__;
  assign new_new_n48171__ = ys__n38045 & new_new_n43040__;
  assign new_new_n48172__ = ys__n18687 & ~new_new_n43044__;
  assign new_new_n48173__ = ~new_new_n48171__ & ~new_new_n48172__;
  assign ys__n32729 = ~new_new_n43047__ & ~new_new_n48173__;
  assign new_new_n48175__ = ys__n38046 & new_new_n43040__;
  assign new_new_n48176__ = ys__n18690 & ~new_new_n43044__;
  assign new_new_n48177__ = ~new_new_n48175__ & ~new_new_n48176__;
  assign ys__n32730 = ~new_new_n43047__ & ~new_new_n48177__;
  assign new_new_n48179__ = ys__n38047 & new_new_n43040__;
  assign new_new_n48180__ = ys__n18693 & ~new_new_n43044__;
  assign new_new_n48181__ = ~new_new_n48179__ & ~new_new_n48180__;
  assign ys__n32731 = ~new_new_n43047__ & ~new_new_n48181__;
  assign new_new_n48183__ = ys__n38048 & new_new_n43040__;
  assign new_new_n48184__ = ys__n18696 & ~new_new_n43044__;
  assign new_new_n48185__ = ~new_new_n48183__ & ~new_new_n48184__;
  assign ys__n32732 = ~new_new_n43047__ & ~new_new_n48185__;
  assign new_new_n48187__ = ys__n38049 & new_new_n43040__;
  assign new_new_n48188__ = ys__n18699 & ~new_new_n43044__;
  assign new_new_n48189__ = ~new_new_n48187__ & ~new_new_n48188__;
  assign ys__n32733 = ~new_new_n43047__ & ~new_new_n48189__;
  assign new_new_n48191__ = ys__n38050 & new_new_n43040__;
  assign new_new_n48192__ = ys__n18702 & ~new_new_n43044__;
  assign new_new_n48193__ = ~new_new_n48191__ & ~new_new_n48192__;
  assign ys__n32734 = ~new_new_n43047__ & ~new_new_n48193__;
  assign new_new_n48195__ = ys__n38051 & new_new_n43040__;
  assign new_new_n48196__ = ys__n18705 & ~new_new_n43044__;
  assign new_new_n48197__ = ~new_new_n48195__ & ~new_new_n48196__;
  assign ys__n32735 = ~new_new_n43047__ & ~new_new_n48197__;
  assign new_new_n48199__ = ys__n38052 & new_new_n43040__;
  assign new_new_n48200__ = ys__n18708 & ~new_new_n43044__;
  assign new_new_n48201__ = ~new_new_n48199__ & ~new_new_n48200__;
  assign ys__n32736 = ~new_new_n43047__ & ~new_new_n48201__;
  assign new_new_n48203__ = ys__n38053 & new_new_n43040__;
  assign new_new_n48204__ = ys__n18711 & ~new_new_n43044__;
  assign new_new_n48205__ = ~new_new_n48203__ & ~new_new_n48204__;
  assign ys__n32737 = ~new_new_n43047__ & ~new_new_n48205__;
  assign new_new_n48207__ = ys__n38054 & new_new_n43040__;
  assign new_new_n48208__ = ys__n18714 & ~new_new_n43044__;
  assign new_new_n48209__ = ~new_new_n48207__ & ~new_new_n48208__;
  assign ys__n32738 = ~new_new_n43047__ & ~new_new_n48209__;
  assign new_new_n48211__ = ys__n38055 & new_new_n43040__;
  assign new_new_n48212__ = ys__n18717 & ~new_new_n43044__;
  assign new_new_n48213__ = ~new_new_n48211__ & ~new_new_n48212__;
  assign ys__n32739 = ~new_new_n43047__ & ~new_new_n48213__;
  assign new_new_n48215__ = ys__n38056 & new_new_n43040__;
  assign new_new_n48216__ = ys__n18720 & ~new_new_n43044__;
  assign new_new_n48217__ = ~new_new_n48215__ & ~new_new_n48216__;
  assign ys__n32740 = ~new_new_n43047__ & ~new_new_n48217__;
  assign new_new_n48219__ = ys__n38057 & new_new_n43040__;
  assign new_new_n48220__ = ys__n18723 & ~new_new_n43044__;
  assign new_new_n48221__ = ~new_new_n48219__ & ~new_new_n48220__;
  assign ys__n32741 = ~new_new_n43047__ & ~new_new_n48221__;
  assign new_new_n48223__ = ys__n38058 & new_new_n43040__;
  assign new_new_n48224__ = ys__n18726 & ~new_new_n43044__;
  assign new_new_n48225__ = ~new_new_n48223__ & ~new_new_n48224__;
  assign ys__n32742 = ~new_new_n43047__ & ~new_new_n48225__;
  assign new_new_n48227__ = ys__n38059 & new_new_n43040__;
  assign new_new_n48228__ = ys__n18729 & ~new_new_n43044__;
  assign new_new_n48229__ = ~new_new_n48227__ & ~new_new_n48228__;
  assign ys__n32743 = ~new_new_n43047__ & ~new_new_n48229__;
  assign new_new_n48231__ = ys__n38060 & new_new_n43040__;
  assign new_new_n48232__ = ys__n18732 & ~new_new_n43044__;
  assign new_new_n48233__ = ~new_new_n48231__ & ~new_new_n48232__;
  assign ys__n32744 = ~new_new_n43047__ & ~new_new_n48233__;
  assign new_new_n48235__ = ys__n38061 & new_new_n43040__;
  assign new_new_n48236__ = ys__n18735 & ~new_new_n43044__;
  assign new_new_n48237__ = ~new_new_n48235__ & ~new_new_n48236__;
  assign ys__n32745 = ~new_new_n43047__ & ~new_new_n48237__;
  assign new_new_n48239__ = ys__n38062 & new_new_n43040__;
  assign new_new_n48240__ = ys__n18738 & ~new_new_n43044__;
  assign new_new_n48241__ = ~new_new_n48239__ & ~new_new_n48240__;
  assign ys__n32746 = ~new_new_n43047__ & ~new_new_n48241__;
  assign new_new_n48243__ = ys__n38063 & new_new_n43040__;
  assign new_new_n48244__ = ys__n18741 & ~new_new_n43044__;
  assign new_new_n48245__ = ~new_new_n48243__ & ~new_new_n48244__;
  assign ys__n32747 = ~new_new_n43047__ & ~new_new_n48245__;
  assign new_new_n48247__ = ys__n38064 & new_new_n43040__;
  assign new_new_n48248__ = ys__n18744 & ~new_new_n43044__;
  assign new_new_n48249__ = ~new_new_n48247__ & ~new_new_n48248__;
  assign ys__n32748 = ~new_new_n43047__ & ~new_new_n48249__;
  assign new_new_n48251__ = ys__n38065 & new_new_n43040__;
  assign new_new_n48252__ = ys__n18747 & ~new_new_n43044__;
  assign new_new_n48253__ = ~new_new_n48251__ & ~new_new_n48252__;
  assign ys__n32749 = ~new_new_n43047__ & ~new_new_n48253__;
  assign new_new_n48255__ = ys__n48138 & new_new_n42750__;
  assign new_new_n48256__ = ys__n18654 & ~new_new_n42754__;
  assign new_new_n48257__ = ~new_new_n48255__ & ~new_new_n48256__;
  assign ys__n32750 = ~new_new_n42757__ & ~new_new_n48257__;
  assign new_new_n48259__ = ys__n48139 & new_new_n42750__;
  assign new_new_n48260__ = ys__n18657 & ~new_new_n42754__;
  assign new_new_n48261__ = ~new_new_n48259__ & ~new_new_n48260__;
  assign ys__n32751 = ~new_new_n42757__ & ~new_new_n48261__;
  assign new_new_n48263__ = ys__n48140 & new_new_n42750__;
  assign new_new_n48264__ = ys__n18660 & ~new_new_n42754__;
  assign new_new_n48265__ = ~new_new_n48263__ & ~new_new_n48264__;
  assign ys__n32752 = ~new_new_n42757__ & ~new_new_n48265__;
  assign new_new_n48267__ = ys__n48141 & new_new_n42750__;
  assign new_new_n48268__ = ys__n18663 & ~new_new_n42754__;
  assign new_new_n48269__ = ~new_new_n48267__ & ~new_new_n48268__;
  assign ys__n32753 = ~new_new_n42757__ & ~new_new_n48269__;
  assign new_new_n48271__ = ys__n38066 & new_new_n42750__;
  assign new_new_n48272__ = ys__n18666 & ~new_new_n42754__;
  assign new_new_n48273__ = ~new_new_n48271__ & ~new_new_n48272__;
  assign ys__n32754 = ~new_new_n42757__ & ~new_new_n48273__;
  assign new_new_n48275__ = ys__n38067 & new_new_n42750__;
  assign new_new_n48276__ = ys__n18669 & ~new_new_n42754__;
  assign new_new_n48277__ = ~new_new_n48275__ & ~new_new_n48276__;
  assign ys__n32755 = ~new_new_n42757__ & ~new_new_n48277__;
  assign new_new_n48279__ = ys__n38068 & new_new_n42750__;
  assign new_new_n48280__ = ys__n18672 & ~new_new_n42754__;
  assign new_new_n48281__ = ~new_new_n48279__ & ~new_new_n48280__;
  assign ys__n32756 = ~new_new_n42757__ & ~new_new_n48281__;
  assign new_new_n48283__ = ys__n38069 & new_new_n42750__;
  assign new_new_n48284__ = ys__n18675 & ~new_new_n42754__;
  assign new_new_n48285__ = ~new_new_n48283__ & ~new_new_n48284__;
  assign ys__n32757 = ~new_new_n42757__ & ~new_new_n48285__;
  assign new_new_n48287__ = ys__n38070 & new_new_n42750__;
  assign new_new_n48288__ = ys__n18678 & ~new_new_n42754__;
  assign new_new_n48289__ = ~new_new_n48287__ & ~new_new_n48288__;
  assign ys__n32758 = ~new_new_n42757__ & ~new_new_n48289__;
  assign new_new_n48291__ = ys__n38071 & new_new_n42750__;
  assign new_new_n48292__ = ys__n18681 & ~new_new_n42754__;
  assign new_new_n48293__ = ~new_new_n48291__ & ~new_new_n48292__;
  assign ys__n32759 = ~new_new_n42757__ & ~new_new_n48293__;
  assign new_new_n48295__ = ys__n38072 & new_new_n42750__;
  assign new_new_n48296__ = ys__n18684 & ~new_new_n42754__;
  assign new_new_n48297__ = ~new_new_n48295__ & ~new_new_n48296__;
  assign ys__n32760 = ~new_new_n42757__ & ~new_new_n48297__;
  assign new_new_n48299__ = ys__n38073 & new_new_n42750__;
  assign new_new_n48300__ = ys__n18687 & ~new_new_n42754__;
  assign new_new_n48301__ = ~new_new_n48299__ & ~new_new_n48300__;
  assign ys__n32761 = ~new_new_n42757__ & ~new_new_n48301__;
  assign new_new_n48303__ = ys__n38074 & new_new_n42750__;
  assign new_new_n48304__ = ys__n18690 & ~new_new_n42754__;
  assign new_new_n48305__ = ~new_new_n48303__ & ~new_new_n48304__;
  assign ys__n32762 = ~new_new_n42757__ & ~new_new_n48305__;
  assign new_new_n48307__ = ys__n38075 & new_new_n42750__;
  assign new_new_n48308__ = ys__n18693 & ~new_new_n42754__;
  assign new_new_n48309__ = ~new_new_n48307__ & ~new_new_n48308__;
  assign ys__n32763 = ~new_new_n42757__ & ~new_new_n48309__;
  assign new_new_n48311__ = ys__n38076 & new_new_n42750__;
  assign new_new_n48312__ = ys__n18696 & ~new_new_n42754__;
  assign new_new_n48313__ = ~new_new_n48311__ & ~new_new_n48312__;
  assign ys__n32764 = ~new_new_n42757__ & ~new_new_n48313__;
  assign new_new_n48315__ = ys__n38077 & new_new_n42750__;
  assign new_new_n48316__ = ys__n18699 & ~new_new_n42754__;
  assign new_new_n48317__ = ~new_new_n48315__ & ~new_new_n48316__;
  assign ys__n32765 = ~new_new_n42757__ & ~new_new_n48317__;
  assign new_new_n48319__ = ys__n38078 & new_new_n42750__;
  assign new_new_n48320__ = ys__n18702 & ~new_new_n42754__;
  assign new_new_n48321__ = ~new_new_n48319__ & ~new_new_n48320__;
  assign ys__n32766 = ~new_new_n42757__ & ~new_new_n48321__;
  assign new_new_n48323__ = ys__n38079 & new_new_n42750__;
  assign new_new_n48324__ = ys__n18705 & ~new_new_n42754__;
  assign new_new_n48325__ = ~new_new_n48323__ & ~new_new_n48324__;
  assign ys__n32767 = ~new_new_n42757__ & ~new_new_n48325__;
  assign new_new_n48327__ = ys__n38080 & new_new_n42750__;
  assign new_new_n48328__ = ys__n18708 & ~new_new_n42754__;
  assign new_new_n48329__ = ~new_new_n48327__ & ~new_new_n48328__;
  assign ys__n32768 = ~new_new_n42757__ & ~new_new_n48329__;
  assign new_new_n48331__ = ys__n38081 & new_new_n42750__;
  assign new_new_n48332__ = ys__n18711 & ~new_new_n42754__;
  assign new_new_n48333__ = ~new_new_n48331__ & ~new_new_n48332__;
  assign ys__n32769 = ~new_new_n42757__ & ~new_new_n48333__;
  assign new_new_n48335__ = ys__n38082 & new_new_n42750__;
  assign new_new_n48336__ = ys__n18714 & ~new_new_n42754__;
  assign new_new_n48337__ = ~new_new_n48335__ & ~new_new_n48336__;
  assign ys__n32770 = ~new_new_n42757__ & ~new_new_n48337__;
  assign new_new_n48339__ = ys__n38083 & new_new_n42750__;
  assign new_new_n48340__ = ys__n18717 & ~new_new_n42754__;
  assign new_new_n48341__ = ~new_new_n48339__ & ~new_new_n48340__;
  assign ys__n32771 = ~new_new_n42757__ & ~new_new_n48341__;
  assign new_new_n48343__ = ys__n38084 & new_new_n42750__;
  assign new_new_n48344__ = ys__n18720 & ~new_new_n42754__;
  assign new_new_n48345__ = ~new_new_n48343__ & ~new_new_n48344__;
  assign ys__n32772 = ~new_new_n42757__ & ~new_new_n48345__;
  assign new_new_n48347__ = ys__n38085 & new_new_n42750__;
  assign new_new_n48348__ = ys__n18723 & ~new_new_n42754__;
  assign new_new_n48349__ = ~new_new_n48347__ & ~new_new_n48348__;
  assign ys__n32773 = ~new_new_n42757__ & ~new_new_n48349__;
  assign new_new_n48351__ = ys__n38086 & new_new_n42750__;
  assign new_new_n48352__ = ys__n18726 & ~new_new_n42754__;
  assign new_new_n48353__ = ~new_new_n48351__ & ~new_new_n48352__;
  assign ys__n32774 = ~new_new_n42757__ & ~new_new_n48353__;
  assign new_new_n48355__ = ys__n38087 & new_new_n42750__;
  assign new_new_n48356__ = ys__n18729 & ~new_new_n42754__;
  assign new_new_n48357__ = ~new_new_n48355__ & ~new_new_n48356__;
  assign ys__n32775 = ~new_new_n42757__ & ~new_new_n48357__;
  assign new_new_n48359__ = ys__n38088 & new_new_n42750__;
  assign new_new_n48360__ = ys__n18732 & ~new_new_n42754__;
  assign new_new_n48361__ = ~new_new_n48359__ & ~new_new_n48360__;
  assign ys__n32776 = ~new_new_n42757__ & ~new_new_n48361__;
  assign new_new_n48363__ = ys__n38089 & new_new_n42750__;
  assign new_new_n48364__ = ys__n18735 & ~new_new_n42754__;
  assign new_new_n48365__ = ~new_new_n48363__ & ~new_new_n48364__;
  assign ys__n32777 = ~new_new_n42757__ & ~new_new_n48365__;
  assign new_new_n48367__ = ys__n38090 & new_new_n42750__;
  assign new_new_n48368__ = ys__n18738 & ~new_new_n42754__;
  assign new_new_n48369__ = ~new_new_n48367__ & ~new_new_n48368__;
  assign ys__n32778 = ~new_new_n42757__ & ~new_new_n48369__;
  assign new_new_n48371__ = ys__n38091 & new_new_n42750__;
  assign new_new_n48372__ = ys__n18741 & ~new_new_n42754__;
  assign new_new_n48373__ = ~new_new_n48371__ & ~new_new_n48372__;
  assign ys__n32779 = ~new_new_n42757__ & ~new_new_n48373__;
  assign new_new_n48375__ = ys__n38092 & new_new_n42750__;
  assign new_new_n48376__ = ys__n18744 & ~new_new_n42754__;
  assign new_new_n48377__ = ~new_new_n48375__ & ~new_new_n48376__;
  assign ys__n32780 = ~new_new_n42757__ & ~new_new_n48377__;
  assign new_new_n48379__ = ys__n38093 & new_new_n42750__;
  assign new_new_n48380__ = ys__n18747 & ~new_new_n42754__;
  assign new_new_n48381__ = ~new_new_n48379__ & ~new_new_n48380__;
  assign ys__n32781 = ~new_new_n42757__ & ~new_new_n48381__;
  assign new_new_n48383__ = ys__n48142 & new_new_n42522__;
  assign new_new_n48384__ = ys__n18654 & ~new_new_n42526__;
  assign new_new_n48385__ = ~new_new_n48383__ & ~new_new_n48384__;
  assign ys__n32782 = ~new_new_n42529__ & ~new_new_n48385__;
  assign new_new_n48387__ = ys__n48143 & new_new_n42522__;
  assign new_new_n48388__ = ys__n18657 & ~new_new_n42526__;
  assign new_new_n48389__ = ~new_new_n48387__ & ~new_new_n48388__;
  assign ys__n32783 = ~new_new_n42529__ & ~new_new_n48389__;
  assign new_new_n48391__ = ys__n48144 & new_new_n42522__;
  assign new_new_n48392__ = ys__n18660 & ~new_new_n42526__;
  assign new_new_n48393__ = ~new_new_n48391__ & ~new_new_n48392__;
  assign ys__n32784 = ~new_new_n42529__ & ~new_new_n48393__;
  assign new_new_n48395__ = ys__n48145 & new_new_n42522__;
  assign new_new_n48396__ = ys__n18663 & ~new_new_n42526__;
  assign new_new_n48397__ = ~new_new_n48395__ & ~new_new_n48396__;
  assign ys__n32785 = ~new_new_n42529__ & ~new_new_n48397__;
  assign new_new_n48399__ = ys__n38094 & new_new_n42522__;
  assign new_new_n48400__ = ys__n18666 & ~new_new_n42526__;
  assign new_new_n48401__ = ~new_new_n48399__ & ~new_new_n48400__;
  assign ys__n32786 = ~new_new_n42529__ & ~new_new_n48401__;
  assign new_new_n48403__ = ys__n38095 & new_new_n42522__;
  assign new_new_n48404__ = ys__n18669 & ~new_new_n42526__;
  assign new_new_n48405__ = ~new_new_n48403__ & ~new_new_n48404__;
  assign ys__n32787 = ~new_new_n42529__ & ~new_new_n48405__;
  assign new_new_n48407__ = ys__n38096 & new_new_n42522__;
  assign new_new_n48408__ = ys__n18672 & ~new_new_n42526__;
  assign new_new_n48409__ = ~new_new_n48407__ & ~new_new_n48408__;
  assign ys__n32788 = ~new_new_n42529__ & ~new_new_n48409__;
  assign new_new_n48411__ = ys__n38097 & new_new_n42522__;
  assign new_new_n48412__ = ys__n18675 & ~new_new_n42526__;
  assign new_new_n48413__ = ~new_new_n48411__ & ~new_new_n48412__;
  assign ys__n32789 = ~new_new_n42529__ & ~new_new_n48413__;
  assign new_new_n48415__ = ys__n38098 & new_new_n42522__;
  assign new_new_n48416__ = ys__n18678 & ~new_new_n42526__;
  assign new_new_n48417__ = ~new_new_n48415__ & ~new_new_n48416__;
  assign ys__n32790 = ~new_new_n42529__ & ~new_new_n48417__;
  assign new_new_n48419__ = ys__n38099 & new_new_n42522__;
  assign new_new_n48420__ = ys__n18681 & ~new_new_n42526__;
  assign new_new_n48421__ = ~new_new_n48419__ & ~new_new_n48420__;
  assign ys__n32791 = ~new_new_n42529__ & ~new_new_n48421__;
  assign new_new_n48423__ = ys__n38100 & new_new_n42522__;
  assign new_new_n48424__ = ys__n18684 & ~new_new_n42526__;
  assign new_new_n48425__ = ~new_new_n48423__ & ~new_new_n48424__;
  assign ys__n32792 = ~new_new_n42529__ & ~new_new_n48425__;
  assign new_new_n48427__ = ys__n38101 & new_new_n42522__;
  assign new_new_n48428__ = ys__n18687 & ~new_new_n42526__;
  assign new_new_n48429__ = ~new_new_n48427__ & ~new_new_n48428__;
  assign ys__n32793 = ~new_new_n42529__ & ~new_new_n48429__;
  assign new_new_n48431__ = ys__n38102 & new_new_n42522__;
  assign new_new_n48432__ = ys__n18690 & ~new_new_n42526__;
  assign new_new_n48433__ = ~new_new_n48431__ & ~new_new_n48432__;
  assign ys__n32794 = ~new_new_n42529__ & ~new_new_n48433__;
  assign new_new_n48435__ = ys__n38103 & new_new_n42522__;
  assign new_new_n48436__ = ys__n18693 & ~new_new_n42526__;
  assign new_new_n48437__ = ~new_new_n48435__ & ~new_new_n48436__;
  assign ys__n32795 = ~new_new_n42529__ & ~new_new_n48437__;
  assign new_new_n48439__ = ys__n38104 & new_new_n42522__;
  assign new_new_n48440__ = ys__n18696 & ~new_new_n42526__;
  assign new_new_n48441__ = ~new_new_n48439__ & ~new_new_n48440__;
  assign ys__n32796 = ~new_new_n42529__ & ~new_new_n48441__;
  assign new_new_n48443__ = ys__n38105 & new_new_n42522__;
  assign new_new_n48444__ = ys__n18699 & ~new_new_n42526__;
  assign new_new_n48445__ = ~new_new_n48443__ & ~new_new_n48444__;
  assign ys__n32797 = ~new_new_n42529__ & ~new_new_n48445__;
  assign new_new_n48447__ = ys__n38106 & new_new_n42522__;
  assign new_new_n48448__ = ys__n18702 & ~new_new_n42526__;
  assign new_new_n48449__ = ~new_new_n48447__ & ~new_new_n48448__;
  assign ys__n32798 = ~new_new_n42529__ & ~new_new_n48449__;
  assign new_new_n48451__ = ys__n38107 & new_new_n42522__;
  assign new_new_n48452__ = ys__n18705 & ~new_new_n42526__;
  assign new_new_n48453__ = ~new_new_n48451__ & ~new_new_n48452__;
  assign ys__n32799 = ~new_new_n42529__ & ~new_new_n48453__;
  assign new_new_n48455__ = ys__n38108 & new_new_n42522__;
  assign new_new_n48456__ = ys__n18708 & ~new_new_n42526__;
  assign new_new_n48457__ = ~new_new_n48455__ & ~new_new_n48456__;
  assign ys__n32800 = ~new_new_n42529__ & ~new_new_n48457__;
  assign new_new_n48459__ = ys__n38109 & new_new_n42522__;
  assign new_new_n48460__ = ys__n18711 & ~new_new_n42526__;
  assign new_new_n48461__ = ~new_new_n48459__ & ~new_new_n48460__;
  assign ys__n32801 = ~new_new_n42529__ & ~new_new_n48461__;
  assign new_new_n48463__ = ys__n38110 & new_new_n42522__;
  assign new_new_n48464__ = ys__n18714 & ~new_new_n42526__;
  assign new_new_n48465__ = ~new_new_n48463__ & ~new_new_n48464__;
  assign ys__n32802 = ~new_new_n42529__ & ~new_new_n48465__;
  assign new_new_n48467__ = ys__n38111 & new_new_n42522__;
  assign new_new_n48468__ = ys__n18717 & ~new_new_n42526__;
  assign new_new_n48469__ = ~new_new_n48467__ & ~new_new_n48468__;
  assign ys__n32803 = ~new_new_n42529__ & ~new_new_n48469__;
  assign new_new_n48471__ = ys__n38112 & new_new_n42522__;
  assign new_new_n48472__ = ys__n18720 & ~new_new_n42526__;
  assign new_new_n48473__ = ~new_new_n48471__ & ~new_new_n48472__;
  assign ys__n32804 = ~new_new_n42529__ & ~new_new_n48473__;
  assign new_new_n48475__ = ys__n38113 & new_new_n42522__;
  assign new_new_n48476__ = ys__n18723 & ~new_new_n42526__;
  assign new_new_n48477__ = ~new_new_n48475__ & ~new_new_n48476__;
  assign ys__n32805 = ~new_new_n42529__ & ~new_new_n48477__;
  assign new_new_n48479__ = ys__n38114 & new_new_n42522__;
  assign new_new_n48480__ = ys__n18726 & ~new_new_n42526__;
  assign new_new_n48481__ = ~new_new_n48479__ & ~new_new_n48480__;
  assign ys__n32806 = ~new_new_n42529__ & ~new_new_n48481__;
  assign new_new_n48483__ = ys__n38115 & new_new_n42522__;
  assign new_new_n48484__ = ys__n18729 & ~new_new_n42526__;
  assign new_new_n48485__ = ~new_new_n48483__ & ~new_new_n48484__;
  assign ys__n32807 = ~new_new_n42529__ & ~new_new_n48485__;
  assign new_new_n48487__ = ys__n38116 & new_new_n42522__;
  assign new_new_n48488__ = ys__n18732 & ~new_new_n42526__;
  assign new_new_n48489__ = ~new_new_n48487__ & ~new_new_n48488__;
  assign ys__n32808 = ~new_new_n42529__ & ~new_new_n48489__;
  assign new_new_n48491__ = ys__n38117 & new_new_n42522__;
  assign new_new_n48492__ = ys__n18735 & ~new_new_n42526__;
  assign new_new_n48493__ = ~new_new_n48491__ & ~new_new_n48492__;
  assign ys__n32809 = ~new_new_n42529__ & ~new_new_n48493__;
  assign new_new_n48495__ = ys__n38118 & new_new_n42522__;
  assign new_new_n48496__ = ys__n18738 & ~new_new_n42526__;
  assign new_new_n48497__ = ~new_new_n48495__ & ~new_new_n48496__;
  assign ys__n32810 = ~new_new_n42529__ & ~new_new_n48497__;
  assign new_new_n48499__ = ys__n38119 & new_new_n42522__;
  assign new_new_n48500__ = ys__n18741 & ~new_new_n42526__;
  assign new_new_n48501__ = ~new_new_n48499__ & ~new_new_n48500__;
  assign ys__n32811 = ~new_new_n42529__ & ~new_new_n48501__;
  assign new_new_n48503__ = ys__n38120 & new_new_n42522__;
  assign new_new_n48504__ = ys__n18744 & ~new_new_n42526__;
  assign new_new_n48505__ = ~new_new_n48503__ & ~new_new_n48504__;
  assign ys__n32812 = ~new_new_n42529__ & ~new_new_n48505__;
  assign new_new_n48507__ = ys__n38121 & new_new_n42522__;
  assign new_new_n48508__ = ys__n18747 & ~new_new_n42526__;
  assign new_new_n48509__ = ~new_new_n48507__ & ~new_new_n48508__;
  assign ys__n32813 = ~new_new_n42529__ & ~new_new_n48509__;
  assign new_new_n48511__ = ys__n48146 & new_new_n42377__;
  assign new_new_n48512__ = ys__n18654 & ~new_new_n42381__;
  assign new_new_n48513__ = ~new_new_n48511__ & ~new_new_n48512__;
  assign ys__n32814 = ~new_new_n42384__ & ~new_new_n48513__;
  assign new_new_n48515__ = ys__n48147 & new_new_n42377__;
  assign new_new_n48516__ = ys__n18657 & ~new_new_n42381__;
  assign new_new_n48517__ = ~new_new_n48515__ & ~new_new_n48516__;
  assign ys__n32815 = ~new_new_n42384__ & ~new_new_n48517__;
  assign new_new_n48519__ = ys__n48148 & new_new_n42377__;
  assign new_new_n48520__ = ys__n18660 & ~new_new_n42381__;
  assign new_new_n48521__ = ~new_new_n48519__ & ~new_new_n48520__;
  assign ys__n32816 = ~new_new_n42384__ & ~new_new_n48521__;
  assign new_new_n48523__ = ys__n48149 & new_new_n42377__;
  assign new_new_n48524__ = ys__n18663 & ~new_new_n42381__;
  assign new_new_n48525__ = ~new_new_n48523__ & ~new_new_n48524__;
  assign ys__n32817 = ~new_new_n42384__ & ~new_new_n48525__;
  assign new_new_n48527__ = ys__n38122 & new_new_n42377__;
  assign new_new_n48528__ = ys__n18666 & ~new_new_n42381__;
  assign new_new_n48529__ = ~new_new_n48527__ & ~new_new_n48528__;
  assign ys__n32818 = ~new_new_n42384__ & ~new_new_n48529__;
  assign new_new_n48531__ = ys__n38123 & new_new_n42377__;
  assign new_new_n48532__ = ys__n18669 & ~new_new_n42381__;
  assign new_new_n48533__ = ~new_new_n48531__ & ~new_new_n48532__;
  assign ys__n32819 = ~new_new_n42384__ & ~new_new_n48533__;
  assign new_new_n48535__ = ys__n38124 & new_new_n42377__;
  assign new_new_n48536__ = ys__n18672 & ~new_new_n42381__;
  assign new_new_n48537__ = ~new_new_n48535__ & ~new_new_n48536__;
  assign ys__n32820 = ~new_new_n42384__ & ~new_new_n48537__;
  assign new_new_n48539__ = ys__n38125 & new_new_n42377__;
  assign new_new_n48540__ = ys__n18675 & ~new_new_n42381__;
  assign new_new_n48541__ = ~new_new_n48539__ & ~new_new_n48540__;
  assign ys__n32821 = ~new_new_n42384__ & ~new_new_n48541__;
  assign new_new_n48543__ = ys__n38126 & new_new_n42377__;
  assign new_new_n48544__ = ys__n18678 & ~new_new_n42381__;
  assign new_new_n48545__ = ~new_new_n48543__ & ~new_new_n48544__;
  assign ys__n32822 = ~new_new_n42384__ & ~new_new_n48545__;
  assign new_new_n48547__ = ys__n38127 & new_new_n42377__;
  assign new_new_n48548__ = ys__n18681 & ~new_new_n42381__;
  assign new_new_n48549__ = ~new_new_n48547__ & ~new_new_n48548__;
  assign ys__n32823 = ~new_new_n42384__ & ~new_new_n48549__;
  assign new_new_n48551__ = ys__n38128 & new_new_n42377__;
  assign new_new_n48552__ = ys__n18684 & ~new_new_n42381__;
  assign new_new_n48553__ = ~new_new_n48551__ & ~new_new_n48552__;
  assign ys__n32824 = ~new_new_n42384__ & ~new_new_n48553__;
  assign new_new_n48555__ = ys__n38129 & new_new_n42377__;
  assign new_new_n48556__ = ys__n18687 & ~new_new_n42381__;
  assign new_new_n48557__ = ~new_new_n48555__ & ~new_new_n48556__;
  assign ys__n32825 = ~new_new_n42384__ & ~new_new_n48557__;
  assign new_new_n48559__ = ys__n38130 & new_new_n42377__;
  assign new_new_n48560__ = ys__n18690 & ~new_new_n42381__;
  assign new_new_n48561__ = ~new_new_n48559__ & ~new_new_n48560__;
  assign ys__n32826 = ~new_new_n42384__ & ~new_new_n48561__;
  assign new_new_n48563__ = ys__n38131 & new_new_n42377__;
  assign new_new_n48564__ = ys__n18693 & ~new_new_n42381__;
  assign new_new_n48565__ = ~new_new_n48563__ & ~new_new_n48564__;
  assign ys__n32827 = ~new_new_n42384__ & ~new_new_n48565__;
  assign new_new_n48567__ = ys__n38132 & new_new_n42377__;
  assign new_new_n48568__ = ys__n18696 & ~new_new_n42381__;
  assign new_new_n48569__ = ~new_new_n48567__ & ~new_new_n48568__;
  assign ys__n32828 = ~new_new_n42384__ & ~new_new_n48569__;
  assign new_new_n48571__ = ys__n38133 & new_new_n42377__;
  assign new_new_n48572__ = ys__n18699 & ~new_new_n42381__;
  assign new_new_n48573__ = ~new_new_n48571__ & ~new_new_n48572__;
  assign ys__n32829 = ~new_new_n42384__ & ~new_new_n48573__;
  assign new_new_n48575__ = ys__n38134 & new_new_n42377__;
  assign new_new_n48576__ = ys__n18702 & ~new_new_n42381__;
  assign new_new_n48577__ = ~new_new_n48575__ & ~new_new_n48576__;
  assign ys__n32830 = ~new_new_n42384__ & ~new_new_n48577__;
  assign new_new_n48579__ = ys__n38135 & new_new_n42377__;
  assign new_new_n48580__ = ys__n18705 & ~new_new_n42381__;
  assign new_new_n48581__ = ~new_new_n48579__ & ~new_new_n48580__;
  assign ys__n32831 = ~new_new_n42384__ & ~new_new_n48581__;
  assign new_new_n48583__ = ys__n38136 & new_new_n42377__;
  assign new_new_n48584__ = ys__n18708 & ~new_new_n42381__;
  assign new_new_n48585__ = ~new_new_n48583__ & ~new_new_n48584__;
  assign ys__n32832 = ~new_new_n42384__ & ~new_new_n48585__;
  assign new_new_n48587__ = ys__n38137 & new_new_n42377__;
  assign new_new_n48588__ = ys__n18711 & ~new_new_n42381__;
  assign new_new_n48589__ = ~new_new_n48587__ & ~new_new_n48588__;
  assign ys__n32833 = ~new_new_n42384__ & ~new_new_n48589__;
  assign new_new_n48591__ = ys__n38138 & new_new_n42377__;
  assign new_new_n48592__ = ys__n18714 & ~new_new_n42381__;
  assign new_new_n48593__ = ~new_new_n48591__ & ~new_new_n48592__;
  assign ys__n32834 = ~new_new_n42384__ & ~new_new_n48593__;
  assign new_new_n48595__ = ys__n38139 & new_new_n42377__;
  assign new_new_n48596__ = ys__n18717 & ~new_new_n42381__;
  assign new_new_n48597__ = ~new_new_n48595__ & ~new_new_n48596__;
  assign ys__n32835 = ~new_new_n42384__ & ~new_new_n48597__;
  assign new_new_n48599__ = ys__n38140 & new_new_n42377__;
  assign new_new_n48600__ = ys__n18720 & ~new_new_n42381__;
  assign new_new_n48601__ = ~new_new_n48599__ & ~new_new_n48600__;
  assign ys__n32836 = ~new_new_n42384__ & ~new_new_n48601__;
  assign new_new_n48603__ = ys__n38141 & new_new_n42377__;
  assign new_new_n48604__ = ys__n18723 & ~new_new_n42381__;
  assign new_new_n48605__ = ~new_new_n48603__ & ~new_new_n48604__;
  assign ys__n32837 = ~new_new_n42384__ & ~new_new_n48605__;
  assign new_new_n48607__ = ys__n38142 & new_new_n42377__;
  assign new_new_n48608__ = ys__n18726 & ~new_new_n42381__;
  assign new_new_n48609__ = ~new_new_n48607__ & ~new_new_n48608__;
  assign ys__n32838 = ~new_new_n42384__ & ~new_new_n48609__;
  assign new_new_n48611__ = ys__n38143 & new_new_n42377__;
  assign new_new_n48612__ = ys__n18729 & ~new_new_n42381__;
  assign new_new_n48613__ = ~new_new_n48611__ & ~new_new_n48612__;
  assign ys__n32839 = ~new_new_n42384__ & ~new_new_n48613__;
  assign new_new_n48615__ = ys__n38144 & new_new_n42377__;
  assign new_new_n48616__ = ys__n18732 & ~new_new_n42381__;
  assign new_new_n48617__ = ~new_new_n48615__ & ~new_new_n48616__;
  assign ys__n32840 = ~new_new_n42384__ & ~new_new_n48617__;
  assign new_new_n48619__ = ys__n38145 & new_new_n42377__;
  assign new_new_n48620__ = ys__n18735 & ~new_new_n42381__;
  assign new_new_n48621__ = ~new_new_n48619__ & ~new_new_n48620__;
  assign ys__n32841 = ~new_new_n42384__ & ~new_new_n48621__;
  assign new_new_n48623__ = ys__n38146 & new_new_n42377__;
  assign new_new_n48624__ = ys__n18738 & ~new_new_n42381__;
  assign new_new_n48625__ = ~new_new_n48623__ & ~new_new_n48624__;
  assign ys__n32842 = ~new_new_n42384__ & ~new_new_n48625__;
  assign new_new_n48627__ = ys__n38147 & new_new_n42377__;
  assign new_new_n48628__ = ys__n18741 & ~new_new_n42381__;
  assign new_new_n48629__ = ~new_new_n48627__ & ~new_new_n48628__;
  assign ys__n32843 = ~new_new_n42384__ & ~new_new_n48629__;
  assign new_new_n48631__ = ys__n38148 & new_new_n42377__;
  assign new_new_n48632__ = ys__n18744 & ~new_new_n42381__;
  assign new_new_n48633__ = ~new_new_n48631__ & ~new_new_n48632__;
  assign ys__n32844 = ~new_new_n42384__ & ~new_new_n48633__;
  assign new_new_n48635__ = ys__n38149 & new_new_n42377__;
  assign new_new_n48636__ = ys__n18747 & ~new_new_n42381__;
  assign new_new_n48637__ = ~new_new_n48635__ & ~new_new_n48636__;
  assign ys__n32845 = ~new_new_n42384__ & ~new_new_n48637__;
  assign new_new_n48639__ = ys__n48150 & new_new_n42232__;
  assign new_new_n48640__ = ys__n18654 & ~new_new_n42236__;
  assign new_new_n48641__ = ~new_new_n48639__ & ~new_new_n48640__;
  assign ys__n32846 = ~new_new_n42239__ & ~new_new_n48641__;
  assign new_new_n48643__ = ys__n48151 & new_new_n42232__;
  assign new_new_n48644__ = ys__n18657 & ~new_new_n42236__;
  assign new_new_n48645__ = ~new_new_n48643__ & ~new_new_n48644__;
  assign ys__n32847 = ~new_new_n42239__ & ~new_new_n48645__;
  assign new_new_n48647__ = ys__n48152 & new_new_n42232__;
  assign new_new_n48648__ = ys__n18660 & ~new_new_n42236__;
  assign new_new_n48649__ = ~new_new_n48647__ & ~new_new_n48648__;
  assign ys__n32848 = ~new_new_n42239__ & ~new_new_n48649__;
  assign new_new_n48651__ = ys__n48153 & new_new_n42232__;
  assign new_new_n48652__ = ys__n18663 & ~new_new_n42236__;
  assign new_new_n48653__ = ~new_new_n48651__ & ~new_new_n48652__;
  assign ys__n32849 = ~new_new_n42239__ & ~new_new_n48653__;
  assign new_new_n48655__ = ys__n38150 & new_new_n42232__;
  assign new_new_n48656__ = ys__n18666 & ~new_new_n42236__;
  assign new_new_n48657__ = ~new_new_n48655__ & ~new_new_n48656__;
  assign ys__n32850 = ~new_new_n42239__ & ~new_new_n48657__;
  assign new_new_n48659__ = ys__n38151 & new_new_n42232__;
  assign new_new_n48660__ = ys__n18669 & ~new_new_n42236__;
  assign new_new_n48661__ = ~new_new_n48659__ & ~new_new_n48660__;
  assign ys__n32851 = ~new_new_n42239__ & ~new_new_n48661__;
  assign new_new_n48663__ = ys__n38152 & new_new_n42232__;
  assign new_new_n48664__ = ys__n18672 & ~new_new_n42236__;
  assign new_new_n48665__ = ~new_new_n48663__ & ~new_new_n48664__;
  assign ys__n32852 = ~new_new_n42239__ & ~new_new_n48665__;
  assign new_new_n48667__ = ys__n38153 & new_new_n42232__;
  assign new_new_n48668__ = ys__n18675 & ~new_new_n42236__;
  assign new_new_n48669__ = ~new_new_n48667__ & ~new_new_n48668__;
  assign ys__n32853 = ~new_new_n42239__ & ~new_new_n48669__;
  assign new_new_n48671__ = ys__n38154 & new_new_n42232__;
  assign new_new_n48672__ = ys__n18678 & ~new_new_n42236__;
  assign new_new_n48673__ = ~new_new_n48671__ & ~new_new_n48672__;
  assign ys__n32854 = ~new_new_n42239__ & ~new_new_n48673__;
  assign new_new_n48675__ = ys__n38155 & new_new_n42232__;
  assign new_new_n48676__ = ys__n18681 & ~new_new_n42236__;
  assign new_new_n48677__ = ~new_new_n48675__ & ~new_new_n48676__;
  assign ys__n32855 = ~new_new_n42239__ & ~new_new_n48677__;
  assign new_new_n48679__ = ys__n38156 & new_new_n42232__;
  assign new_new_n48680__ = ys__n18684 & ~new_new_n42236__;
  assign new_new_n48681__ = ~new_new_n48679__ & ~new_new_n48680__;
  assign ys__n32856 = ~new_new_n42239__ & ~new_new_n48681__;
  assign new_new_n48683__ = ys__n38157 & new_new_n42232__;
  assign new_new_n48684__ = ys__n18687 & ~new_new_n42236__;
  assign new_new_n48685__ = ~new_new_n48683__ & ~new_new_n48684__;
  assign ys__n32857 = ~new_new_n42239__ & ~new_new_n48685__;
  assign new_new_n48687__ = ys__n38158 & new_new_n42232__;
  assign new_new_n48688__ = ys__n18690 & ~new_new_n42236__;
  assign new_new_n48689__ = ~new_new_n48687__ & ~new_new_n48688__;
  assign ys__n32858 = ~new_new_n42239__ & ~new_new_n48689__;
  assign new_new_n48691__ = ys__n38159 & new_new_n42232__;
  assign new_new_n48692__ = ys__n18693 & ~new_new_n42236__;
  assign new_new_n48693__ = ~new_new_n48691__ & ~new_new_n48692__;
  assign ys__n32859 = ~new_new_n42239__ & ~new_new_n48693__;
  assign new_new_n48695__ = ys__n38160 & new_new_n42232__;
  assign new_new_n48696__ = ys__n18696 & ~new_new_n42236__;
  assign new_new_n48697__ = ~new_new_n48695__ & ~new_new_n48696__;
  assign ys__n32860 = ~new_new_n42239__ & ~new_new_n48697__;
  assign new_new_n48699__ = ys__n38161 & new_new_n42232__;
  assign new_new_n48700__ = ys__n18699 & ~new_new_n42236__;
  assign new_new_n48701__ = ~new_new_n48699__ & ~new_new_n48700__;
  assign ys__n32861 = ~new_new_n42239__ & ~new_new_n48701__;
  assign new_new_n48703__ = ys__n38162 & new_new_n42232__;
  assign new_new_n48704__ = ys__n18702 & ~new_new_n42236__;
  assign new_new_n48705__ = ~new_new_n48703__ & ~new_new_n48704__;
  assign ys__n32862 = ~new_new_n42239__ & ~new_new_n48705__;
  assign new_new_n48707__ = ys__n38163 & new_new_n42232__;
  assign new_new_n48708__ = ys__n18705 & ~new_new_n42236__;
  assign new_new_n48709__ = ~new_new_n48707__ & ~new_new_n48708__;
  assign ys__n32863 = ~new_new_n42239__ & ~new_new_n48709__;
  assign new_new_n48711__ = ys__n38164 & new_new_n42232__;
  assign new_new_n48712__ = ys__n18708 & ~new_new_n42236__;
  assign new_new_n48713__ = ~new_new_n48711__ & ~new_new_n48712__;
  assign ys__n32864 = ~new_new_n42239__ & ~new_new_n48713__;
  assign new_new_n48715__ = ys__n38165 & new_new_n42232__;
  assign new_new_n48716__ = ys__n18711 & ~new_new_n42236__;
  assign new_new_n48717__ = ~new_new_n48715__ & ~new_new_n48716__;
  assign ys__n32865 = ~new_new_n42239__ & ~new_new_n48717__;
  assign new_new_n48719__ = ys__n38166 & new_new_n42232__;
  assign new_new_n48720__ = ys__n18714 & ~new_new_n42236__;
  assign new_new_n48721__ = ~new_new_n48719__ & ~new_new_n48720__;
  assign ys__n32866 = ~new_new_n42239__ & ~new_new_n48721__;
  assign new_new_n48723__ = ys__n38167 & new_new_n42232__;
  assign new_new_n48724__ = ys__n18717 & ~new_new_n42236__;
  assign new_new_n48725__ = ~new_new_n48723__ & ~new_new_n48724__;
  assign ys__n32867 = ~new_new_n42239__ & ~new_new_n48725__;
  assign new_new_n48727__ = ys__n38168 & new_new_n42232__;
  assign new_new_n48728__ = ys__n18720 & ~new_new_n42236__;
  assign new_new_n48729__ = ~new_new_n48727__ & ~new_new_n48728__;
  assign ys__n32868 = ~new_new_n42239__ & ~new_new_n48729__;
  assign new_new_n48731__ = ys__n38169 & new_new_n42232__;
  assign new_new_n48732__ = ys__n18723 & ~new_new_n42236__;
  assign new_new_n48733__ = ~new_new_n48731__ & ~new_new_n48732__;
  assign ys__n32869 = ~new_new_n42239__ & ~new_new_n48733__;
  assign new_new_n48735__ = ys__n38170 & new_new_n42232__;
  assign new_new_n48736__ = ys__n18726 & ~new_new_n42236__;
  assign new_new_n48737__ = ~new_new_n48735__ & ~new_new_n48736__;
  assign ys__n32870 = ~new_new_n42239__ & ~new_new_n48737__;
  assign new_new_n48739__ = ys__n38171 & new_new_n42232__;
  assign new_new_n48740__ = ys__n18729 & ~new_new_n42236__;
  assign new_new_n48741__ = ~new_new_n48739__ & ~new_new_n48740__;
  assign ys__n32871 = ~new_new_n42239__ & ~new_new_n48741__;
  assign new_new_n48743__ = ys__n38172 & new_new_n42232__;
  assign new_new_n48744__ = ys__n18732 & ~new_new_n42236__;
  assign new_new_n48745__ = ~new_new_n48743__ & ~new_new_n48744__;
  assign ys__n32872 = ~new_new_n42239__ & ~new_new_n48745__;
  assign new_new_n48747__ = ys__n38173 & new_new_n42232__;
  assign new_new_n48748__ = ys__n18735 & ~new_new_n42236__;
  assign new_new_n48749__ = ~new_new_n48747__ & ~new_new_n48748__;
  assign ys__n32873 = ~new_new_n42239__ & ~new_new_n48749__;
  assign new_new_n48751__ = ys__n38174 & new_new_n42232__;
  assign new_new_n48752__ = ys__n18738 & ~new_new_n42236__;
  assign new_new_n48753__ = ~new_new_n48751__ & ~new_new_n48752__;
  assign ys__n32874 = ~new_new_n42239__ & ~new_new_n48753__;
  assign new_new_n48755__ = ys__n38175 & new_new_n42232__;
  assign new_new_n48756__ = ys__n18741 & ~new_new_n42236__;
  assign new_new_n48757__ = ~new_new_n48755__ & ~new_new_n48756__;
  assign ys__n32875 = ~new_new_n42239__ & ~new_new_n48757__;
  assign new_new_n48759__ = ys__n38176 & new_new_n42232__;
  assign new_new_n48760__ = ys__n18744 & ~new_new_n42236__;
  assign new_new_n48761__ = ~new_new_n48759__ & ~new_new_n48760__;
  assign ys__n32876 = ~new_new_n42239__ & ~new_new_n48761__;
  assign new_new_n48763__ = ys__n38177 & new_new_n42232__;
  assign new_new_n48764__ = ys__n18747 & ~new_new_n42236__;
  assign new_new_n48765__ = ~new_new_n48763__ & ~new_new_n48764__;
  assign ys__n32877 = ~new_new_n42239__ & ~new_new_n48765__;
  assign new_new_n48767__ = ys__n37757 & new_new_n46832__;
  assign new_new_n48768__ = ys__n18759 & ~new_new_n46836__;
  assign new_new_n48769__ = ~new_new_n48767__ & ~new_new_n48768__;
  assign ys__n32878 = ~new_new_n46839__ & ~new_new_n48769__;
  assign new_new_n48771__ = ys__n37756 & new_new_n46965__;
  assign new_new_n48772__ = ys__n18759 & ~new_new_n46969__;
  assign new_new_n48773__ = ~new_new_n48771__ & ~new_new_n48772__;
  assign ys__n32879 = ~new_new_n46972__ & ~new_new_n48773__;
  assign new_new_n48775__ = ys__n37755 & new_new_n47098__;
  assign new_new_n48776__ = ys__n18759 & ~new_new_n47102__;
  assign new_new_n48777__ = ~new_new_n48775__ & ~new_new_n48776__;
  assign ys__n32880 = ~new_new_n47105__ & ~new_new_n48777__;
  assign new_new_n48779__ = ys__n37754 & new_new_n43944__;
  assign new_new_n48780__ = ys__n18759 & ~new_new_n43948__;
  assign new_new_n48781__ = ~new_new_n48779__ & ~new_new_n48780__;
  assign ys__n32881 = ~new_new_n43951__ & ~new_new_n48781__;
  assign new_new_n48783__ = ys__n37753 & new_new_n43799__;
  assign new_new_n48784__ = ys__n18759 & ~new_new_n43803__;
  assign new_new_n48785__ = ~new_new_n48783__ & ~new_new_n48784__;
  assign ys__n32882 = ~new_new_n43806__ & ~new_new_n48785__;
  assign new_new_n48787__ = ys__n37752 & new_new_n43654__;
  assign new_new_n48788__ = ys__n18759 & ~new_new_n43658__;
  assign new_new_n48789__ = ~new_new_n48787__ & ~new_new_n48788__;
  assign ys__n32883 = ~new_new_n43661__ & ~new_new_n48789__;
  assign new_new_n48791__ = ys__n37751 & new_new_n43509__;
  assign new_new_n48792__ = ys__n18759 & ~new_new_n43513__;
  assign new_new_n48793__ = ~new_new_n48791__ & ~new_new_n48792__;
  assign ys__n32884 = ~new_new_n43516__ & ~new_new_n48793__;
  assign new_new_n48795__ = ys__n37750 & new_new_n43364__;
  assign new_new_n48796__ = ys__n18759 & ~new_new_n43368__;
  assign new_new_n48797__ = ~new_new_n48795__ & ~new_new_n48796__;
  assign ys__n32885 = ~new_new_n43371__ & ~new_new_n48797__;
  assign new_new_n48799__ = ys__n37749 & new_new_n43219__;
  assign new_new_n48800__ = ys__n18759 & ~new_new_n43223__;
  assign new_new_n48801__ = ~new_new_n48799__ & ~new_new_n48800__;
  assign ys__n32886 = ~new_new_n43226__ & ~new_new_n48801__;
  assign new_new_n48803__ = ys__n37748 & new_new_n42895__;
  assign new_new_n48804__ = ys__n18759 & ~new_new_n42899__;
  assign new_new_n48805__ = ~new_new_n48803__ & ~new_new_n48804__;
  assign ys__n32887 = ~new_new_n42902__ & ~new_new_n48805__;
  assign new_new_n48807__ = ys__n37747 & new_new_n43040__;
  assign new_new_n48808__ = ys__n18759 & ~new_new_n43044__;
  assign new_new_n48809__ = ~new_new_n48807__ & ~new_new_n48808__;
  assign ys__n32888 = ~new_new_n43047__ & ~new_new_n48809__;
  assign new_new_n48811__ = ys__n37746 & new_new_n42750__;
  assign new_new_n48812__ = ys__n18759 & ~new_new_n42754__;
  assign new_new_n48813__ = ~new_new_n48811__ & ~new_new_n48812__;
  assign ys__n32889 = ~new_new_n42757__ & ~new_new_n48813__;
  assign new_new_n48815__ = ys__n37745 & new_new_n42522__;
  assign new_new_n48816__ = ys__n18759 & ~new_new_n42526__;
  assign new_new_n48817__ = ~new_new_n48815__ & ~new_new_n48816__;
  assign ys__n32890 = ~new_new_n42529__ & ~new_new_n48817__;
  assign new_new_n48819__ = ys__n37744 & new_new_n42377__;
  assign new_new_n48820__ = ys__n18759 & ~new_new_n42381__;
  assign new_new_n48821__ = ~new_new_n48819__ & ~new_new_n48820__;
  assign ys__n32891 = ~new_new_n42384__ & ~new_new_n48821__;
  assign new_new_n48823__ = ys__n37743 & new_new_n42232__;
  assign new_new_n48824__ = ys__n18759 & ~new_new_n42236__;
  assign new_new_n48825__ = ~new_new_n48823__ & ~new_new_n48824__;
  assign ys__n32892 = ~new_new_n42239__ & ~new_new_n48825__;
  assign new_new_n48827__ = ys__n48154 & new_new_n46832__;
  assign new_new_n48828__ = ys__n47202 & ~new_new_n46836__;
  assign new_new_n48829__ = ~new_new_n48827__ & ~new_new_n48828__;
  assign ys__n32893 = ~new_new_n46839__ & ~new_new_n48829__;
  assign new_new_n48831__ = ys__n48155 & new_new_n46832__;
  assign new_new_n48832__ = ys__n47203 & ~new_new_n46836__;
  assign new_new_n48833__ = ~new_new_n48831__ & ~new_new_n48832__;
  assign ys__n32894 = ~new_new_n46839__ & ~new_new_n48833__;
  assign new_new_n48835__ = ys__n48156 & new_new_n46832__;
  assign new_new_n48836__ = ys__n47204 & ~new_new_n46836__;
  assign new_new_n48837__ = ~new_new_n48835__ & ~new_new_n48836__;
  assign ys__n32895 = ~new_new_n46839__ & ~new_new_n48837__;
  assign new_new_n48839__ = ys__n48157 & new_new_n46832__;
  assign new_new_n48840__ = ys__n47205 & ~new_new_n46836__;
  assign new_new_n48841__ = ~new_new_n48839__ & ~new_new_n48840__;
  assign ys__n32896 = ~new_new_n46839__ & ~new_new_n48841__;
  assign new_new_n48843__ = ys__n48158 & new_new_n46832__;
  assign new_new_n48844__ = ys__n47206 & ~new_new_n46836__;
  assign new_new_n48845__ = ~new_new_n48843__ & ~new_new_n48844__;
  assign ys__n32897 = ~new_new_n46839__ & ~new_new_n48845__;
  assign new_new_n48847__ = ys__n48159 & new_new_n46832__;
  assign new_new_n48848__ = ys__n47207 & ~new_new_n46836__;
  assign new_new_n48849__ = ~new_new_n48847__ & ~new_new_n48848__;
  assign ys__n32898 = ~new_new_n46839__ & ~new_new_n48849__;
  assign new_new_n48851__ = ys__n48160 & new_new_n46832__;
  assign new_new_n48852__ = ys__n47208 & ~new_new_n46836__;
  assign new_new_n48853__ = ~new_new_n48851__ & ~new_new_n48852__;
  assign ys__n32899 = ~new_new_n46839__ & ~new_new_n48853__;
  assign new_new_n48855__ = ys__n48161 & new_new_n46832__;
  assign new_new_n48856__ = ys__n47209 & ~new_new_n46836__;
  assign new_new_n48857__ = ~new_new_n48855__ & ~new_new_n48856__;
  assign ys__n32900 = ~new_new_n46839__ & ~new_new_n48857__;
  assign new_new_n48859__ = ys__n48162 & new_new_n46832__;
  assign new_new_n48860__ = ys__n47210 & ~new_new_n46836__;
  assign new_new_n48861__ = ~new_new_n48859__ & ~new_new_n48860__;
  assign ys__n32901 = ~new_new_n46839__ & ~new_new_n48861__;
  assign new_new_n48863__ = ys__n48163 & new_new_n46832__;
  assign new_new_n48864__ = ys__n47211 & ~new_new_n46836__;
  assign new_new_n48865__ = ~new_new_n48863__ & ~new_new_n48864__;
  assign ys__n32902 = ~new_new_n46839__ & ~new_new_n48865__;
  assign new_new_n48867__ = ys__n48164 & new_new_n46832__;
  assign new_new_n48868__ = ys__n47212 & ~new_new_n46836__;
  assign new_new_n48869__ = ~new_new_n48867__ & ~new_new_n48868__;
  assign ys__n32903 = ~new_new_n46839__ & ~new_new_n48869__;
  assign new_new_n48871__ = ys__n48165 & new_new_n46832__;
  assign new_new_n48872__ = ys__n47213 & ~new_new_n46836__;
  assign new_new_n48873__ = ~new_new_n48871__ & ~new_new_n48872__;
  assign ys__n32904 = ~new_new_n46839__ & ~new_new_n48873__;
  assign new_new_n48875__ = ys__n48166 & new_new_n46832__;
  assign new_new_n48876__ = ys__n47214 & ~new_new_n46836__;
  assign new_new_n48877__ = ~new_new_n48875__ & ~new_new_n48876__;
  assign ys__n32905 = ~new_new_n46839__ & ~new_new_n48877__;
  assign new_new_n48879__ = ys__n48167 & new_new_n46832__;
  assign new_new_n48880__ = ys__n47215 & ~new_new_n46836__;
  assign new_new_n48881__ = ~new_new_n48879__ & ~new_new_n48880__;
  assign ys__n32906 = ~new_new_n46839__ & ~new_new_n48881__;
  assign new_new_n48883__ = ys__n48168 & new_new_n46832__;
  assign new_new_n48884__ = ys__n47216 & ~new_new_n46836__;
  assign new_new_n48885__ = ~new_new_n48883__ & ~new_new_n48884__;
  assign ys__n32907 = ~new_new_n46839__ & ~new_new_n48885__;
  assign new_new_n48887__ = ys__n48169 & new_new_n46832__;
  assign new_new_n48888__ = ys__n47217 & ~new_new_n46836__;
  assign new_new_n48889__ = ~new_new_n48887__ & ~new_new_n48888__;
  assign ys__n32908 = ~new_new_n46839__ & ~new_new_n48889__;
  assign new_new_n48891__ = ys__n48170 & new_new_n46832__;
  assign new_new_n48892__ = ys__n47218 & ~new_new_n46836__;
  assign new_new_n48893__ = ~new_new_n48891__ & ~new_new_n48892__;
  assign ys__n32909 = ~new_new_n46839__ & ~new_new_n48893__;
  assign new_new_n48895__ = ys__n48171 & new_new_n46832__;
  assign new_new_n48896__ = ys__n47219 & ~new_new_n46836__;
  assign new_new_n48897__ = ~new_new_n48895__ & ~new_new_n48896__;
  assign ys__n32910 = ~new_new_n46839__ & ~new_new_n48897__;
  assign new_new_n48899__ = ys__n48172 & new_new_n46832__;
  assign new_new_n48900__ = ys__n47220 & ~new_new_n46836__;
  assign new_new_n48901__ = ~new_new_n48899__ & ~new_new_n48900__;
  assign ys__n32911 = ~new_new_n46839__ & ~new_new_n48901__;
  assign new_new_n48903__ = ys__n48173 & new_new_n46832__;
  assign new_new_n48904__ = ys__n47221 & ~new_new_n46836__;
  assign new_new_n48905__ = ~new_new_n48903__ & ~new_new_n48904__;
  assign ys__n32912 = ~new_new_n46839__ & ~new_new_n48905__;
  assign new_new_n48907__ = ys__n48174 & new_new_n46832__;
  assign new_new_n48908__ = ys__n47222 & ~new_new_n46836__;
  assign new_new_n48909__ = ~new_new_n48907__ & ~new_new_n48908__;
  assign ys__n32913 = ~new_new_n46839__ & ~new_new_n48909__;
  assign new_new_n48911__ = ys__n48175 & new_new_n46832__;
  assign new_new_n48912__ = ys__n47223 & ~new_new_n46836__;
  assign new_new_n48913__ = ~new_new_n48911__ & ~new_new_n48912__;
  assign ys__n32914 = ~new_new_n46839__ & ~new_new_n48913__;
  assign new_new_n48915__ = ys__n48176 & new_new_n46832__;
  assign new_new_n48916__ = ys__n47224 & ~new_new_n46836__;
  assign new_new_n48917__ = ~new_new_n48915__ & ~new_new_n48916__;
  assign ys__n32915 = ~new_new_n46839__ & ~new_new_n48917__;
  assign new_new_n48919__ = ys__n48177 & new_new_n46832__;
  assign new_new_n48920__ = ys__n47225 & ~new_new_n46836__;
  assign new_new_n48921__ = ~new_new_n48919__ & ~new_new_n48920__;
  assign ys__n32916 = ~new_new_n46839__ & ~new_new_n48921__;
  assign new_new_n48923__ = ys__n48178 & new_new_n46832__;
  assign new_new_n48924__ = ys__n47226 & ~new_new_n46836__;
  assign new_new_n48925__ = ~new_new_n48923__ & ~new_new_n48924__;
  assign ys__n32917 = ~new_new_n46839__ & ~new_new_n48925__;
  assign new_new_n48927__ = ys__n48179 & new_new_n46832__;
  assign new_new_n48928__ = ys__n47227 & ~new_new_n46836__;
  assign new_new_n48929__ = ~new_new_n48927__ & ~new_new_n48928__;
  assign ys__n32918 = ~new_new_n46839__ & ~new_new_n48929__;
  assign new_new_n48931__ = ys__n48180 & new_new_n46832__;
  assign new_new_n48932__ = ys__n47228 & ~new_new_n46836__;
  assign new_new_n48933__ = ~new_new_n48931__ & ~new_new_n48932__;
  assign ys__n32919 = ~new_new_n46839__ & ~new_new_n48933__;
  assign new_new_n48935__ = ys__n48181 & new_new_n46832__;
  assign new_new_n48936__ = ys__n47229 & ~new_new_n46836__;
  assign new_new_n48937__ = ~new_new_n48935__ & ~new_new_n48936__;
  assign ys__n32920 = ~new_new_n46839__ & ~new_new_n48937__;
  assign new_new_n48939__ = ys__n48182 & new_new_n46832__;
  assign new_new_n48940__ = ys__n47230 & ~new_new_n46836__;
  assign new_new_n48941__ = ~new_new_n48939__ & ~new_new_n48940__;
  assign ys__n32921 = ~new_new_n46839__ & ~new_new_n48941__;
  assign new_new_n48943__ = ys__n48183 & new_new_n46832__;
  assign new_new_n48944__ = ys__n47231 & ~new_new_n46836__;
  assign new_new_n48945__ = ~new_new_n48943__ & ~new_new_n48944__;
  assign ys__n32922 = ~new_new_n46839__ & ~new_new_n48945__;
  assign new_new_n48947__ = ys__n48184 & new_new_n46832__;
  assign new_new_n48948__ = ys__n47232 & ~new_new_n46836__;
  assign new_new_n48949__ = ~new_new_n48947__ & ~new_new_n48948__;
  assign ys__n32923 = ~new_new_n46839__ & ~new_new_n48949__;
  assign new_new_n48951__ = ys__n48185 & new_new_n46832__;
  assign new_new_n48952__ = ys__n47233 & ~new_new_n46836__;
  assign new_new_n48953__ = ~new_new_n48951__ & ~new_new_n48952__;
  assign ys__n32924 = ~new_new_n46839__ & ~new_new_n48953__;
  assign new_new_n48955__ = ys__n48186 & new_new_n46832__;
  assign new_new_n48956__ = ys__n18762 & ~new_new_n46836__;
  assign new_new_n48957__ = ~new_new_n48955__ & ~new_new_n48956__;
  assign ys__n32925 = ~new_new_n46839__ & ~new_new_n48957__;
  assign new_new_n48959__ = ys__n48187 & new_new_n46832__;
  assign new_new_n48960__ = ys__n18750 & ~new_new_n46836__;
  assign new_new_n48961__ = ~new_new_n48959__ & ~new_new_n48960__;
  assign ys__n32926 = ~new_new_n46839__ & ~new_new_n48961__;
  assign new_new_n48963__ = ys__n48188 & new_new_n46832__;
  assign new_new_n48964__ = ys__n18753 & ~new_new_n46836__;
  assign new_new_n48965__ = ~new_new_n48963__ & ~new_new_n48964__;
  assign ys__n32927 = ~new_new_n46839__ & ~new_new_n48965__;
  assign new_new_n48967__ = ys__n48189 & new_new_n46965__;
  assign new_new_n48968__ = ys__n47202 & ~new_new_n46969__;
  assign new_new_n48969__ = ~new_new_n48967__ & ~new_new_n48968__;
  assign ys__n32928 = ~new_new_n46972__ & ~new_new_n48969__;
  assign new_new_n48971__ = ys__n48190 & new_new_n46965__;
  assign new_new_n48972__ = ys__n47203 & ~new_new_n46969__;
  assign new_new_n48973__ = ~new_new_n48971__ & ~new_new_n48972__;
  assign ys__n32929 = ~new_new_n46972__ & ~new_new_n48973__;
  assign new_new_n48975__ = ys__n48191 & new_new_n46965__;
  assign new_new_n48976__ = ys__n47204 & ~new_new_n46969__;
  assign new_new_n48977__ = ~new_new_n48975__ & ~new_new_n48976__;
  assign ys__n32930 = ~new_new_n46972__ & ~new_new_n48977__;
  assign new_new_n48979__ = ys__n48192 & new_new_n46965__;
  assign new_new_n48980__ = ys__n47205 & ~new_new_n46969__;
  assign new_new_n48981__ = ~new_new_n48979__ & ~new_new_n48980__;
  assign ys__n32931 = ~new_new_n46972__ & ~new_new_n48981__;
  assign new_new_n48983__ = ys__n48193 & new_new_n46965__;
  assign new_new_n48984__ = ys__n47206 & ~new_new_n46969__;
  assign new_new_n48985__ = ~new_new_n48983__ & ~new_new_n48984__;
  assign ys__n32932 = ~new_new_n46972__ & ~new_new_n48985__;
  assign new_new_n48987__ = ys__n48194 & new_new_n46965__;
  assign new_new_n48988__ = ys__n47207 & ~new_new_n46969__;
  assign new_new_n48989__ = ~new_new_n48987__ & ~new_new_n48988__;
  assign ys__n32933 = ~new_new_n46972__ & ~new_new_n48989__;
  assign new_new_n48991__ = ys__n48195 & new_new_n46965__;
  assign new_new_n48992__ = ys__n47208 & ~new_new_n46969__;
  assign new_new_n48993__ = ~new_new_n48991__ & ~new_new_n48992__;
  assign ys__n32934 = ~new_new_n46972__ & ~new_new_n48993__;
  assign new_new_n48995__ = ys__n48196 & new_new_n46965__;
  assign new_new_n48996__ = ys__n47209 & ~new_new_n46969__;
  assign new_new_n48997__ = ~new_new_n48995__ & ~new_new_n48996__;
  assign ys__n32935 = ~new_new_n46972__ & ~new_new_n48997__;
  assign new_new_n48999__ = ys__n48197 & new_new_n46965__;
  assign new_new_n49000__ = ys__n47210 & ~new_new_n46969__;
  assign new_new_n49001__ = ~new_new_n48999__ & ~new_new_n49000__;
  assign ys__n32936 = ~new_new_n46972__ & ~new_new_n49001__;
  assign new_new_n49003__ = ys__n48198 & new_new_n46965__;
  assign new_new_n49004__ = ys__n47211 & ~new_new_n46969__;
  assign new_new_n49005__ = ~new_new_n49003__ & ~new_new_n49004__;
  assign ys__n32937 = ~new_new_n46972__ & ~new_new_n49005__;
  assign new_new_n49007__ = ys__n48199 & new_new_n46965__;
  assign new_new_n49008__ = ys__n47212 & ~new_new_n46969__;
  assign new_new_n49009__ = ~new_new_n49007__ & ~new_new_n49008__;
  assign ys__n32938 = ~new_new_n46972__ & ~new_new_n49009__;
  assign new_new_n49011__ = ys__n48200 & new_new_n46965__;
  assign new_new_n49012__ = ys__n47213 & ~new_new_n46969__;
  assign new_new_n49013__ = ~new_new_n49011__ & ~new_new_n49012__;
  assign ys__n32939 = ~new_new_n46972__ & ~new_new_n49013__;
  assign new_new_n49015__ = ys__n48201 & new_new_n46965__;
  assign new_new_n49016__ = ys__n47214 & ~new_new_n46969__;
  assign new_new_n49017__ = ~new_new_n49015__ & ~new_new_n49016__;
  assign ys__n32940 = ~new_new_n46972__ & ~new_new_n49017__;
  assign new_new_n49019__ = ys__n48202 & new_new_n46965__;
  assign new_new_n49020__ = ys__n47215 & ~new_new_n46969__;
  assign new_new_n49021__ = ~new_new_n49019__ & ~new_new_n49020__;
  assign ys__n32941 = ~new_new_n46972__ & ~new_new_n49021__;
  assign new_new_n49023__ = ys__n48203 & new_new_n46965__;
  assign new_new_n49024__ = ys__n47216 & ~new_new_n46969__;
  assign new_new_n49025__ = ~new_new_n49023__ & ~new_new_n49024__;
  assign ys__n32942 = ~new_new_n46972__ & ~new_new_n49025__;
  assign new_new_n49027__ = ys__n48204 & new_new_n46965__;
  assign new_new_n49028__ = ys__n47217 & ~new_new_n46969__;
  assign new_new_n49029__ = ~new_new_n49027__ & ~new_new_n49028__;
  assign ys__n32943 = ~new_new_n46972__ & ~new_new_n49029__;
  assign new_new_n49031__ = ys__n48205 & new_new_n46965__;
  assign new_new_n49032__ = ys__n47218 & ~new_new_n46969__;
  assign new_new_n49033__ = ~new_new_n49031__ & ~new_new_n49032__;
  assign ys__n32944 = ~new_new_n46972__ & ~new_new_n49033__;
  assign new_new_n49035__ = ys__n48206 & new_new_n46965__;
  assign new_new_n49036__ = ys__n47219 & ~new_new_n46969__;
  assign new_new_n49037__ = ~new_new_n49035__ & ~new_new_n49036__;
  assign ys__n32945 = ~new_new_n46972__ & ~new_new_n49037__;
  assign new_new_n49039__ = ys__n48207 & new_new_n46965__;
  assign new_new_n49040__ = ys__n47220 & ~new_new_n46969__;
  assign new_new_n49041__ = ~new_new_n49039__ & ~new_new_n49040__;
  assign ys__n32946 = ~new_new_n46972__ & ~new_new_n49041__;
  assign new_new_n49043__ = ys__n48208 & new_new_n46965__;
  assign new_new_n49044__ = ys__n47221 & ~new_new_n46969__;
  assign new_new_n49045__ = ~new_new_n49043__ & ~new_new_n49044__;
  assign ys__n32947 = ~new_new_n46972__ & ~new_new_n49045__;
  assign new_new_n49047__ = ys__n48209 & new_new_n46965__;
  assign new_new_n49048__ = ys__n47222 & ~new_new_n46969__;
  assign new_new_n49049__ = ~new_new_n49047__ & ~new_new_n49048__;
  assign ys__n32948 = ~new_new_n46972__ & ~new_new_n49049__;
  assign new_new_n49051__ = ys__n48210 & new_new_n46965__;
  assign new_new_n49052__ = ys__n47223 & ~new_new_n46969__;
  assign new_new_n49053__ = ~new_new_n49051__ & ~new_new_n49052__;
  assign ys__n32949 = ~new_new_n46972__ & ~new_new_n49053__;
  assign new_new_n49055__ = ys__n48211 & new_new_n46965__;
  assign new_new_n49056__ = ys__n47224 & ~new_new_n46969__;
  assign new_new_n49057__ = ~new_new_n49055__ & ~new_new_n49056__;
  assign ys__n32950 = ~new_new_n46972__ & ~new_new_n49057__;
  assign new_new_n49059__ = ys__n48212 & new_new_n46965__;
  assign new_new_n49060__ = ys__n47225 & ~new_new_n46969__;
  assign new_new_n49061__ = ~new_new_n49059__ & ~new_new_n49060__;
  assign ys__n32951 = ~new_new_n46972__ & ~new_new_n49061__;
  assign new_new_n49063__ = ys__n48213 & new_new_n46965__;
  assign new_new_n49064__ = ys__n47226 & ~new_new_n46969__;
  assign new_new_n49065__ = ~new_new_n49063__ & ~new_new_n49064__;
  assign ys__n32952 = ~new_new_n46972__ & ~new_new_n49065__;
  assign new_new_n49067__ = ys__n48214 & new_new_n46965__;
  assign new_new_n49068__ = ys__n47227 & ~new_new_n46969__;
  assign new_new_n49069__ = ~new_new_n49067__ & ~new_new_n49068__;
  assign ys__n32953 = ~new_new_n46972__ & ~new_new_n49069__;
  assign new_new_n49071__ = ys__n48215 & new_new_n46965__;
  assign new_new_n49072__ = ys__n47228 & ~new_new_n46969__;
  assign new_new_n49073__ = ~new_new_n49071__ & ~new_new_n49072__;
  assign ys__n32954 = ~new_new_n46972__ & ~new_new_n49073__;
  assign new_new_n49075__ = ys__n48216 & new_new_n46965__;
  assign new_new_n49076__ = ys__n47229 & ~new_new_n46969__;
  assign new_new_n49077__ = ~new_new_n49075__ & ~new_new_n49076__;
  assign ys__n32955 = ~new_new_n46972__ & ~new_new_n49077__;
  assign new_new_n49079__ = ys__n48217 & new_new_n46965__;
  assign new_new_n49080__ = ys__n47230 & ~new_new_n46969__;
  assign new_new_n49081__ = ~new_new_n49079__ & ~new_new_n49080__;
  assign ys__n32956 = ~new_new_n46972__ & ~new_new_n49081__;
  assign new_new_n49083__ = ys__n48218 & new_new_n46965__;
  assign new_new_n49084__ = ys__n47231 & ~new_new_n46969__;
  assign new_new_n49085__ = ~new_new_n49083__ & ~new_new_n49084__;
  assign ys__n32957 = ~new_new_n46972__ & ~new_new_n49085__;
  assign new_new_n49087__ = ys__n48219 & new_new_n46965__;
  assign new_new_n49088__ = ys__n47232 & ~new_new_n46969__;
  assign new_new_n49089__ = ~new_new_n49087__ & ~new_new_n49088__;
  assign ys__n32958 = ~new_new_n46972__ & ~new_new_n49089__;
  assign new_new_n49091__ = ys__n48220 & new_new_n46965__;
  assign new_new_n49092__ = ys__n47233 & ~new_new_n46969__;
  assign new_new_n49093__ = ~new_new_n49091__ & ~new_new_n49092__;
  assign ys__n32959 = ~new_new_n46972__ & ~new_new_n49093__;
  assign new_new_n49095__ = ys__n48221 & new_new_n46965__;
  assign new_new_n49096__ = ys__n18762 & ~new_new_n46969__;
  assign new_new_n49097__ = ~new_new_n49095__ & ~new_new_n49096__;
  assign ys__n32960 = ~new_new_n46972__ & ~new_new_n49097__;
  assign new_new_n49099__ = ys__n48222 & new_new_n46965__;
  assign new_new_n49100__ = ys__n18750 & ~new_new_n46969__;
  assign new_new_n49101__ = ~new_new_n49099__ & ~new_new_n49100__;
  assign ys__n32961 = ~new_new_n46972__ & ~new_new_n49101__;
  assign new_new_n49103__ = ys__n48223 & new_new_n46965__;
  assign new_new_n49104__ = ys__n18753 & ~new_new_n46969__;
  assign new_new_n49105__ = ~new_new_n49103__ & ~new_new_n49104__;
  assign ys__n32962 = ~new_new_n46972__ & ~new_new_n49105__;
  assign new_new_n49107__ = ys__n48224 & new_new_n47098__;
  assign new_new_n49108__ = ys__n47202 & ~new_new_n47102__;
  assign new_new_n49109__ = ~new_new_n49107__ & ~new_new_n49108__;
  assign ys__n32963 = ~new_new_n47105__ & ~new_new_n49109__;
  assign new_new_n49111__ = ys__n48225 & new_new_n47098__;
  assign new_new_n49112__ = ys__n47203 & ~new_new_n47102__;
  assign new_new_n49113__ = ~new_new_n49111__ & ~new_new_n49112__;
  assign ys__n32964 = ~new_new_n47105__ & ~new_new_n49113__;
  assign new_new_n49115__ = ys__n48226 & new_new_n47098__;
  assign new_new_n49116__ = ys__n47204 & ~new_new_n47102__;
  assign new_new_n49117__ = ~new_new_n49115__ & ~new_new_n49116__;
  assign ys__n32965 = ~new_new_n47105__ & ~new_new_n49117__;
  assign new_new_n49119__ = ys__n48227 & new_new_n47098__;
  assign new_new_n49120__ = ys__n47205 & ~new_new_n47102__;
  assign new_new_n49121__ = ~new_new_n49119__ & ~new_new_n49120__;
  assign ys__n32966 = ~new_new_n47105__ & ~new_new_n49121__;
  assign new_new_n49123__ = ys__n48228 & new_new_n47098__;
  assign new_new_n49124__ = ys__n47206 & ~new_new_n47102__;
  assign new_new_n49125__ = ~new_new_n49123__ & ~new_new_n49124__;
  assign ys__n32967 = ~new_new_n47105__ & ~new_new_n49125__;
  assign new_new_n49127__ = ys__n48229 & new_new_n47098__;
  assign new_new_n49128__ = ys__n47207 & ~new_new_n47102__;
  assign new_new_n49129__ = ~new_new_n49127__ & ~new_new_n49128__;
  assign ys__n32968 = ~new_new_n47105__ & ~new_new_n49129__;
  assign new_new_n49131__ = ys__n48230 & new_new_n47098__;
  assign new_new_n49132__ = ys__n47208 & ~new_new_n47102__;
  assign new_new_n49133__ = ~new_new_n49131__ & ~new_new_n49132__;
  assign ys__n32969 = ~new_new_n47105__ & ~new_new_n49133__;
  assign new_new_n49135__ = ys__n48231 & new_new_n47098__;
  assign new_new_n49136__ = ys__n47209 & ~new_new_n47102__;
  assign new_new_n49137__ = ~new_new_n49135__ & ~new_new_n49136__;
  assign ys__n32970 = ~new_new_n47105__ & ~new_new_n49137__;
  assign new_new_n49139__ = ys__n48232 & new_new_n47098__;
  assign new_new_n49140__ = ys__n47210 & ~new_new_n47102__;
  assign new_new_n49141__ = ~new_new_n49139__ & ~new_new_n49140__;
  assign ys__n32971 = ~new_new_n47105__ & ~new_new_n49141__;
  assign new_new_n49143__ = ys__n48233 & new_new_n47098__;
  assign new_new_n49144__ = ys__n47211 & ~new_new_n47102__;
  assign new_new_n49145__ = ~new_new_n49143__ & ~new_new_n49144__;
  assign ys__n32972 = ~new_new_n47105__ & ~new_new_n49145__;
  assign new_new_n49147__ = ys__n48234 & new_new_n47098__;
  assign new_new_n49148__ = ys__n47212 & ~new_new_n47102__;
  assign new_new_n49149__ = ~new_new_n49147__ & ~new_new_n49148__;
  assign ys__n32973 = ~new_new_n47105__ & ~new_new_n49149__;
  assign new_new_n49151__ = ys__n48235 & new_new_n47098__;
  assign new_new_n49152__ = ys__n47213 & ~new_new_n47102__;
  assign new_new_n49153__ = ~new_new_n49151__ & ~new_new_n49152__;
  assign ys__n32974 = ~new_new_n47105__ & ~new_new_n49153__;
  assign new_new_n49155__ = ys__n48236 & new_new_n47098__;
  assign new_new_n49156__ = ys__n47214 & ~new_new_n47102__;
  assign new_new_n49157__ = ~new_new_n49155__ & ~new_new_n49156__;
  assign ys__n32975 = ~new_new_n47105__ & ~new_new_n49157__;
  assign new_new_n49159__ = ys__n48237 & new_new_n47098__;
  assign new_new_n49160__ = ys__n47215 & ~new_new_n47102__;
  assign new_new_n49161__ = ~new_new_n49159__ & ~new_new_n49160__;
  assign ys__n32976 = ~new_new_n47105__ & ~new_new_n49161__;
  assign new_new_n49163__ = ys__n48238 & new_new_n47098__;
  assign new_new_n49164__ = ys__n47216 & ~new_new_n47102__;
  assign new_new_n49165__ = ~new_new_n49163__ & ~new_new_n49164__;
  assign ys__n32977 = ~new_new_n47105__ & ~new_new_n49165__;
  assign new_new_n49167__ = ys__n48239 & new_new_n47098__;
  assign new_new_n49168__ = ys__n47217 & ~new_new_n47102__;
  assign new_new_n49169__ = ~new_new_n49167__ & ~new_new_n49168__;
  assign ys__n32978 = ~new_new_n47105__ & ~new_new_n49169__;
  assign new_new_n49171__ = ys__n48240 & new_new_n47098__;
  assign new_new_n49172__ = ys__n47218 & ~new_new_n47102__;
  assign new_new_n49173__ = ~new_new_n49171__ & ~new_new_n49172__;
  assign ys__n32979 = ~new_new_n47105__ & ~new_new_n49173__;
  assign new_new_n49175__ = ys__n48241 & new_new_n47098__;
  assign new_new_n49176__ = ys__n47219 & ~new_new_n47102__;
  assign new_new_n49177__ = ~new_new_n49175__ & ~new_new_n49176__;
  assign ys__n32980 = ~new_new_n47105__ & ~new_new_n49177__;
  assign new_new_n49179__ = ys__n48242 & new_new_n47098__;
  assign new_new_n49180__ = ys__n47220 & ~new_new_n47102__;
  assign new_new_n49181__ = ~new_new_n49179__ & ~new_new_n49180__;
  assign ys__n32981 = ~new_new_n47105__ & ~new_new_n49181__;
  assign new_new_n49183__ = ys__n48243 & new_new_n47098__;
  assign new_new_n49184__ = ys__n47221 & ~new_new_n47102__;
  assign new_new_n49185__ = ~new_new_n49183__ & ~new_new_n49184__;
  assign ys__n32982 = ~new_new_n47105__ & ~new_new_n49185__;
  assign new_new_n49187__ = ys__n48244 & new_new_n47098__;
  assign new_new_n49188__ = ys__n47222 & ~new_new_n47102__;
  assign new_new_n49189__ = ~new_new_n49187__ & ~new_new_n49188__;
  assign ys__n32983 = ~new_new_n47105__ & ~new_new_n49189__;
  assign new_new_n49191__ = ys__n48245 & new_new_n47098__;
  assign new_new_n49192__ = ys__n47223 & ~new_new_n47102__;
  assign new_new_n49193__ = ~new_new_n49191__ & ~new_new_n49192__;
  assign ys__n32984 = ~new_new_n47105__ & ~new_new_n49193__;
  assign new_new_n49195__ = ys__n48246 & new_new_n47098__;
  assign new_new_n49196__ = ys__n47224 & ~new_new_n47102__;
  assign new_new_n49197__ = ~new_new_n49195__ & ~new_new_n49196__;
  assign ys__n32985 = ~new_new_n47105__ & ~new_new_n49197__;
  assign new_new_n49199__ = ys__n48247 & new_new_n47098__;
  assign new_new_n49200__ = ys__n47225 & ~new_new_n47102__;
  assign new_new_n49201__ = ~new_new_n49199__ & ~new_new_n49200__;
  assign ys__n32986 = ~new_new_n47105__ & ~new_new_n49201__;
  assign new_new_n49203__ = ys__n48248 & new_new_n47098__;
  assign new_new_n49204__ = ys__n47226 & ~new_new_n47102__;
  assign new_new_n49205__ = ~new_new_n49203__ & ~new_new_n49204__;
  assign ys__n32987 = ~new_new_n47105__ & ~new_new_n49205__;
  assign new_new_n49207__ = ys__n48249 & new_new_n47098__;
  assign new_new_n49208__ = ys__n47227 & ~new_new_n47102__;
  assign new_new_n49209__ = ~new_new_n49207__ & ~new_new_n49208__;
  assign ys__n32988 = ~new_new_n47105__ & ~new_new_n49209__;
  assign new_new_n49211__ = ys__n48250 & new_new_n47098__;
  assign new_new_n49212__ = ys__n47228 & ~new_new_n47102__;
  assign new_new_n49213__ = ~new_new_n49211__ & ~new_new_n49212__;
  assign ys__n32989 = ~new_new_n47105__ & ~new_new_n49213__;
  assign new_new_n49215__ = ys__n48251 & new_new_n47098__;
  assign new_new_n49216__ = ys__n47229 & ~new_new_n47102__;
  assign new_new_n49217__ = ~new_new_n49215__ & ~new_new_n49216__;
  assign ys__n32990 = ~new_new_n47105__ & ~new_new_n49217__;
  assign new_new_n49219__ = ys__n48252 & new_new_n47098__;
  assign new_new_n49220__ = ys__n47230 & ~new_new_n47102__;
  assign new_new_n49221__ = ~new_new_n49219__ & ~new_new_n49220__;
  assign ys__n32991 = ~new_new_n47105__ & ~new_new_n49221__;
  assign new_new_n49223__ = ys__n48253 & new_new_n47098__;
  assign new_new_n49224__ = ys__n47231 & ~new_new_n47102__;
  assign new_new_n49225__ = ~new_new_n49223__ & ~new_new_n49224__;
  assign ys__n32992 = ~new_new_n47105__ & ~new_new_n49225__;
  assign new_new_n49227__ = ys__n48254 & new_new_n47098__;
  assign new_new_n49228__ = ys__n47232 & ~new_new_n47102__;
  assign new_new_n49229__ = ~new_new_n49227__ & ~new_new_n49228__;
  assign ys__n32993 = ~new_new_n47105__ & ~new_new_n49229__;
  assign new_new_n49231__ = ys__n48255 & new_new_n47098__;
  assign new_new_n49232__ = ys__n47233 & ~new_new_n47102__;
  assign new_new_n49233__ = ~new_new_n49231__ & ~new_new_n49232__;
  assign ys__n32994 = ~new_new_n47105__ & ~new_new_n49233__;
  assign new_new_n49235__ = ys__n48256 & new_new_n47098__;
  assign new_new_n49236__ = ys__n18762 & ~new_new_n47102__;
  assign new_new_n49237__ = ~new_new_n49235__ & ~new_new_n49236__;
  assign ys__n32995 = ~new_new_n47105__ & ~new_new_n49237__;
  assign new_new_n49239__ = ys__n48257 & new_new_n47098__;
  assign new_new_n49240__ = ys__n18750 & ~new_new_n47102__;
  assign new_new_n49241__ = ~new_new_n49239__ & ~new_new_n49240__;
  assign ys__n32996 = ~new_new_n47105__ & ~new_new_n49241__;
  assign new_new_n49243__ = ys__n48258 & new_new_n47098__;
  assign new_new_n49244__ = ys__n18753 & ~new_new_n47102__;
  assign new_new_n49245__ = ~new_new_n49243__ & ~new_new_n49244__;
  assign ys__n32997 = ~new_new_n47105__ & ~new_new_n49245__;
  assign ys__n32998 = new_new_n12343__ & ~new_new_n12352__;
  assign new_new_n49248__ = ys__n140 & ~ys__n214;
  assign new_new_n49249__ = new_new_n12154__ & new_new_n49248__;
  assign new_new_n49250__ = ~new_new_n12156__ & ~new_new_n49249__;
  assign new_new_n49251__ = new_new_n12153__ & new_new_n49250__;
  assign new_new_n49252__ = new_new_n16904__ & new_new_n49251__;
  assign new_new_n49253__ = ~ys__n740 & new_new_n16904__;
  assign new_new_n49254__ = new_new_n12150__ & new_new_n49253__;
  assign new_new_n49255__ = ys__n30223 & new_new_n16904__;
  assign new_new_n49256__ = new_new_n12152__ & new_new_n49255__;
  assign new_new_n49257__ = ~new_new_n49254__ & ~new_new_n49256__;
  assign new_new_n49258__ = ~ys__n1020 & new_new_n12429__;
  assign new_new_n49259__ = new_new_n16904__ & new_new_n49258__;
  assign new_new_n49260__ = new_new_n12156__ & new_new_n49259__;
  assign new_new_n49261__ = new_new_n49249__ & new_new_n49253__;
  assign new_new_n49262__ = ~new_new_n49260__ & ~new_new_n49261__;
  assign new_new_n49263__ = new_new_n49257__ & new_new_n49262__;
  assign new_new_n49264__ = ~new_new_n49251__ & ~new_new_n49263__;
  assign ys__n33014 = new_new_n49252__ | new_new_n49264__;
  assign new_new_n49266__ = new_new_n12130__ & new_new_n49251__;
  assign new_new_n49267__ = ~ys__n740 & new_new_n12130__;
  assign new_new_n49268__ = new_new_n12150__ & new_new_n49267__;
  assign new_new_n49269__ = ys__n30223 & new_new_n12130__;
  assign new_new_n49270__ = new_new_n12152__ & new_new_n49269__;
  assign new_new_n49271__ = ~new_new_n49268__ & ~new_new_n49270__;
  assign new_new_n49272__ = new_new_n12130__ & new_new_n49258__;
  assign new_new_n49273__ = new_new_n12156__ & new_new_n49272__;
  assign new_new_n49274__ = new_new_n49249__ & new_new_n49267__;
  assign new_new_n49275__ = ~new_new_n49273__ & ~new_new_n49274__;
  assign new_new_n49276__ = new_new_n49271__ & new_new_n49275__;
  assign new_new_n49277__ = ~new_new_n49251__ & ~new_new_n49276__;
  assign ys__n33015 = new_new_n49266__ | new_new_n49277__;
  assign new_new_n49279__ = new_new_n12112__ & new_new_n49251__;
  assign new_new_n49280__ = ~ys__n740 & new_new_n12112__;
  assign new_new_n49281__ = new_new_n12150__ & new_new_n49280__;
  assign new_new_n49282__ = ys__n30223 & new_new_n12112__;
  assign new_new_n49283__ = new_new_n12152__ & new_new_n49282__;
  assign new_new_n49284__ = ~new_new_n49281__ & ~new_new_n49283__;
  assign new_new_n49285__ = new_new_n12112__ & new_new_n49258__;
  assign new_new_n49286__ = new_new_n12156__ & new_new_n49285__;
  assign new_new_n49287__ = new_new_n49249__ & new_new_n49280__;
  assign new_new_n49288__ = ~new_new_n49286__ & ~new_new_n49287__;
  assign new_new_n49289__ = new_new_n49284__ & new_new_n49288__;
  assign new_new_n49290__ = ~new_new_n49251__ & ~new_new_n49289__;
  assign ys__n33016 = new_new_n49279__ | new_new_n49290__;
  assign new_new_n49292__ = new_new_n12054__ & new_new_n49251__;
  assign new_new_n49293__ = ~ys__n740 & new_new_n12054__;
  assign new_new_n49294__ = new_new_n12150__ & new_new_n49293__;
  assign new_new_n49295__ = ys__n30223 & new_new_n12054__;
  assign new_new_n49296__ = new_new_n12152__ & new_new_n49295__;
  assign new_new_n49297__ = ~new_new_n49294__ & ~new_new_n49296__;
  assign new_new_n49298__ = new_new_n12054__ & new_new_n49258__;
  assign new_new_n49299__ = new_new_n12156__ & new_new_n49298__;
  assign new_new_n49300__ = new_new_n49249__ & new_new_n49293__;
  assign new_new_n49301__ = ~new_new_n49299__ & ~new_new_n49300__;
  assign new_new_n49302__ = new_new_n49297__ & new_new_n49301__;
  assign new_new_n49303__ = ~new_new_n49251__ & ~new_new_n49302__;
  assign ys__n33017 = new_new_n49292__ | new_new_n49303__;
  assign new_new_n49305__ = new_new_n10605__ & new_new_n49251__;
  assign new_new_n49306__ = new_new_n10605__ & ~ys__n740;
  assign new_new_n49307__ = new_new_n12150__ & new_new_n49306__;
  assign new_new_n49308__ = new_new_n10605__ & ys__n30223;
  assign new_new_n49309__ = new_new_n12152__ & new_new_n49308__;
  assign new_new_n49310__ = ~new_new_n49307__ & ~new_new_n49309__;
  assign new_new_n49311__ = new_new_n10605__ & new_new_n49258__;
  assign new_new_n49312__ = new_new_n12156__ & new_new_n49311__;
  assign new_new_n49313__ = new_new_n49249__ & new_new_n49306__;
  assign new_new_n49314__ = ~new_new_n49312__ & ~new_new_n49313__;
  assign new_new_n49315__ = new_new_n49310__ & new_new_n49314__;
  assign new_new_n49316__ = ~new_new_n49251__ & ~new_new_n49315__;
  assign ys__n33018 = new_new_n49305__ | new_new_n49316__;
  assign new_new_n49318__ = new_new_n44241__ & new_new_n49251__;
  assign new_new_n49319__ = ~ys__n740 & new_new_n44241__;
  assign new_new_n49320__ = new_new_n12150__ & new_new_n49319__;
  assign new_new_n49321__ = ys__n30223 & new_new_n44241__;
  assign new_new_n49322__ = new_new_n12152__ & new_new_n49321__;
  assign new_new_n49323__ = ~new_new_n49320__ & ~new_new_n49322__;
  assign new_new_n49324__ = new_new_n44241__ & new_new_n49258__;
  assign new_new_n49325__ = new_new_n12156__ & new_new_n49324__;
  assign new_new_n49326__ = new_new_n49249__ & new_new_n49319__;
  assign new_new_n49327__ = ~new_new_n49325__ & ~new_new_n49326__;
  assign new_new_n49328__ = new_new_n49323__ & new_new_n49327__;
  assign new_new_n49329__ = ~new_new_n49251__ & ~new_new_n49328__;
  assign ys__n33019 = new_new_n49318__ | new_new_n49329__;
  assign new_new_n49331__ = new_new_n26170__ & new_new_n49251__;
  assign new_new_n49332__ = ~ys__n740 & new_new_n26170__;
  assign new_new_n49333__ = new_new_n12150__ & new_new_n49332__;
  assign new_new_n49334__ = ys__n30223 & new_new_n26170__;
  assign new_new_n49335__ = new_new_n12152__ & new_new_n49334__;
  assign new_new_n49336__ = ~new_new_n49333__ & ~new_new_n49335__;
  assign new_new_n49337__ = new_new_n26170__ & new_new_n49258__;
  assign new_new_n49338__ = new_new_n12156__ & new_new_n49337__;
  assign new_new_n49339__ = new_new_n49249__ & new_new_n49332__;
  assign new_new_n49340__ = ~new_new_n49338__ & ~new_new_n49339__;
  assign new_new_n49341__ = new_new_n49336__ & new_new_n49340__;
  assign new_new_n49342__ = ~new_new_n49251__ & ~new_new_n49341__;
  assign ys__n33020 = new_new_n49331__ | new_new_n49342__;
  assign new_new_n49344__ = new_new_n26181__ & new_new_n49251__;
  assign new_new_n49345__ = ~ys__n740 & new_new_n26181__;
  assign new_new_n49346__ = new_new_n12150__ & new_new_n49345__;
  assign new_new_n49347__ = ys__n30223 & new_new_n26181__;
  assign new_new_n49348__ = new_new_n12152__ & new_new_n49347__;
  assign new_new_n49349__ = ~new_new_n49346__ & ~new_new_n49348__;
  assign new_new_n49350__ = new_new_n26181__ & new_new_n49258__;
  assign new_new_n49351__ = new_new_n12156__ & new_new_n49350__;
  assign new_new_n49352__ = new_new_n49249__ & new_new_n49345__;
  assign new_new_n49353__ = ~new_new_n49351__ & ~new_new_n49352__;
  assign new_new_n49354__ = new_new_n49349__ & new_new_n49353__;
  assign new_new_n49355__ = ~new_new_n49251__ & ~new_new_n49354__;
  assign ys__n33021 = new_new_n49344__ | new_new_n49355__;
  assign new_new_n49357__ = new_new_n26192__ & new_new_n49251__;
  assign new_new_n49358__ = ~ys__n740 & new_new_n26192__;
  assign new_new_n49359__ = new_new_n12150__ & new_new_n49358__;
  assign new_new_n49360__ = ys__n30223 & new_new_n26192__;
  assign new_new_n49361__ = new_new_n12152__ & new_new_n49360__;
  assign new_new_n49362__ = ~new_new_n49359__ & ~new_new_n49361__;
  assign new_new_n49363__ = new_new_n26192__ & new_new_n49258__;
  assign new_new_n49364__ = new_new_n12156__ & new_new_n49363__;
  assign new_new_n49365__ = new_new_n49249__ & new_new_n49358__;
  assign new_new_n49366__ = ~new_new_n49364__ & ~new_new_n49365__;
  assign new_new_n49367__ = new_new_n49362__ & new_new_n49366__;
  assign new_new_n49368__ = ~new_new_n49251__ & ~new_new_n49367__;
  assign ys__n33022 = new_new_n49357__ | new_new_n49368__;
  assign new_new_n49370__ = new_new_n16892__ & new_new_n49251__;
  assign new_new_n49371__ = ~ys__n740 & new_new_n16892__;
  assign new_new_n49372__ = new_new_n12150__ & new_new_n49371__;
  assign new_new_n49373__ = ys__n30223 & new_new_n16892__;
  assign new_new_n49374__ = new_new_n12152__ & new_new_n49373__;
  assign new_new_n49375__ = ~new_new_n49372__ & ~new_new_n49374__;
  assign new_new_n49376__ = new_new_n16892__ & new_new_n49258__;
  assign new_new_n49377__ = new_new_n12156__ & new_new_n49376__;
  assign new_new_n49378__ = new_new_n49249__ & new_new_n49371__;
  assign new_new_n49379__ = ~new_new_n49377__ & ~new_new_n49378__;
  assign new_new_n49380__ = new_new_n49375__ & new_new_n49379__;
  assign new_new_n49381__ = ~new_new_n49251__ & ~new_new_n49380__;
  assign ys__n33023 = new_new_n49370__ | new_new_n49381__;
  assign new_new_n49383__ = new_new_n44252__ & new_new_n49251__;
  assign new_new_n49384__ = ~ys__n740 & new_new_n44252__;
  assign new_new_n49385__ = new_new_n12150__ & new_new_n49384__;
  assign new_new_n49386__ = ys__n30223 & new_new_n44252__;
  assign new_new_n49387__ = new_new_n12152__ & new_new_n49386__;
  assign new_new_n49388__ = ~new_new_n49385__ & ~new_new_n49387__;
  assign new_new_n49389__ = new_new_n44252__ & new_new_n49258__;
  assign new_new_n49390__ = new_new_n12156__ & new_new_n49389__;
  assign new_new_n49391__ = new_new_n49249__ & new_new_n49384__;
  assign new_new_n49392__ = ~new_new_n49390__ & ~new_new_n49391__;
  assign new_new_n49393__ = new_new_n49388__ & new_new_n49392__;
  assign new_new_n49394__ = ~new_new_n49251__ & ~new_new_n49393__;
  assign ys__n33024 = new_new_n49383__ | new_new_n49394__;
  assign new_new_n49396__ = new_new_n44263__ & new_new_n49251__;
  assign new_new_n49397__ = ~ys__n740 & new_new_n44263__;
  assign new_new_n49398__ = new_new_n12150__ & new_new_n49397__;
  assign new_new_n49399__ = ys__n30223 & new_new_n44263__;
  assign new_new_n49400__ = new_new_n12152__ & new_new_n49399__;
  assign new_new_n49401__ = ~new_new_n49398__ & ~new_new_n49400__;
  assign new_new_n49402__ = new_new_n44263__ & new_new_n49258__;
  assign new_new_n49403__ = new_new_n12156__ & new_new_n49402__;
  assign new_new_n49404__ = new_new_n49249__ & new_new_n49397__;
  assign new_new_n49405__ = ~new_new_n49403__ & ~new_new_n49404__;
  assign new_new_n49406__ = new_new_n49401__ & new_new_n49405__;
  assign new_new_n49407__ = ~new_new_n49251__ & ~new_new_n49406__;
  assign ys__n33025 = new_new_n49396__ | new_new_n49407__;
  assign new_new_n49409__ = new_new_n44274__ & new_new_n49251__;
  assign new_new_n49410__ = ~ys__n740 & new_new_n44274__;
  assign new_new_n49411__ = new_new_n12150__ & new_new_n49410__;
  assign new_new_n49412__ = ys__n30223 & new_new_n44274__;
  assign new_new_n49413__ = new_new_n12152__ & new_new_n49412__;
  assign new_new_n49414__ = ~new_new_n49411__ & ~new_new_n49413__;
  assign new_new_n49415__ = new_new_n44274__ & new_new_n49258__;
  assign new_new_n49416__ = new_new_n12156__ & new_new_n49415__;
  assign new_new_n49417__ = new_new_n49249__ & new_new_n49410__;
  assign new_new_n49418__ = ~new_new_n49416__ & ~new_new_n49417__;
  assign new_new_n49419__ = new_new_n49414__ & new_new_n49418__;
  assign new_new_n49420__ = ~new_new_n49251__ & ~new_new_n49419__;
  assign ys__n33026 = new_new_n49409__ | new_new_n49420__;
  assign new_new_n49422__ = new_new_n44285__ & new_new_n49251__;
  assign new_new_n49423__ = ~ys__n740 & new_new_n44285__;
  assign new_new_n49424__ = new_new_n12150__ & new_new_n49423__;
  assign new_new_n49425__ = ys__n30223 & new_new_n44285__;
  assign new_new_n49426__ = new_new_n12152__ & new_new_n49425__;
  assign new_new_n49427__ = ~new_new_n49424__ & ~new_new_n49426__;
  assign new_new_n49428__ = new_new_n44285__ & new_new_n49258__;
  assign new_new_n49429__ = new_new_n12156__ & new_new_n49428__;
  assign new_new_n49430__ = new_new_n49249__ & new_new_n49423__;
  assign new_new_n49431__ = ~new_new_n49429__ & ~new_new_n49430__;
  assign new_new_n49432__ = new_new_n49427__ & new_new_n49431__;
  assign new_new_n49433__ = ~new_new_n49251__ & ~new_new_n49432__;
  assign ys__n33027 = new_new_n49422__ | new_new_n49433__;
  assign new_new_n49435__ = new_new_n44298__ & new_new_n49251__;
  assign new_new_n49436__ = ~ys__n740 & new_new_n44298__;
  assign new_new_n49437__ = new_new_n12150__ & new_new_n49436__;
  assign new_new_n49438__ = ys__n30223 & new_new_n44298__;
  assign new_new_n49439__ = new_new_n12152__ & new_new_n49438__;
  assign new_new_n49440__ = ~new_new_n49437__ & ~new_new_n49439__;
  assign new_new_n49441__ = new_new_n44298__ & new_new_n49258__;
  assign new_new_n49442__ = new_new_n12156__ & new_new_n49441__;
  assign new_new_n49443__ = new_new_n49249__ & new_new_n49436__;
  assign new_new_n49444__ = ~new_new_n49442__ & ~new_new_n49443__;
  assign new_new_n49445__ = new_new_n49440__ & new_new_n49444__;
  assign new_new_n49446__ = ~new_new_n49251__ & ~new_new_n49445__;
  assign ys__n33028 = new_new_n49435__ | new_new_n49446__;
  assign new_new_n49448__ = new_new_n44309__ & new_new_n49251__;
  assign new_new_n49449__ = ~ys__n740 & new_new_n44309__;
  assign new_new_n49450__ = new_new_n12150__ & new_new_n49449__;
  assign new_new_n49451__ = ys__n30223 & new_new_n44309__;
  assign new_new_n49452__ = new_new_n12152__ & new_new_n49451__;
  assign new_new_n49453__ = ~new_new_n49450__ & ~new_new_n49452__;
  assign new_new_n49454__ = new_new_n44309__ & new_new_n49258__;
  assign new_new_n49455__ = new_new_n12156__ & new_new_n49454__;
  assign new_new_n49456__ = new_new_n49249__ & new_new_n49449__;
  assign new_new_n49457__ = ~new_new_n49455__ & ~new_new_n49456__;
  assign new_new_n49458__ = new_new_n49453__ & new_new_n49457__;
  assign new_new_n49459__ = ~new_new_n49251__ & ~new_new_n49458__;
  assign ys__n33029 = new_new_n49448__ | new_new_n49459__;
  assign new_new_n49461__ = new_new_n16907__ & new_new_n49251__;
  assign new_new_n49462__ = ~ys__n740 & new_new_n16907__;
  assign new_new_n49463__ = new_new_n12150__ & new_new_n49462__;
  assign new_new_n49464__ = ys__n30223 & new_new_n16907__;
  assign new_new_n49465__ = new_new_n12152__ & new_new_n49464__;
  assign new_new_n49466__ = ~new_new_n49463__ & ~new_new_n49465__;
  assign new_new_n49467__ = new_new_n16907__ & new_new_n49258__;
  assign new_new_n49468__ = new_new_n12156__ & new_new_n49467__;
  assign new_new_n49469__ = new_new_n49249__ & new_new_n49462__;
  assign new_new_n49470__ = ~new_new_n49468__ & ~new_new_n49469__;
  assign new_new_n49471__ = new_new_n49466__ & new_new_n49470__;
  assign new_new_n49472__ = ~new_new_n49251__ & ~new_new_n49471__;
  assign ys__n33030 = new_new_n49461__ | new_new_n49472__;
  assign new_new_n49474__ = new_new_n12133__ & new_new_n49251__;
  assign new_new_n49475__ = ~ys__n740 & new_new_n12133__;
  assign new_new_n49476__ = new_new_n12150__ & new_new_n49475__;
  assign new_new_n49477__ = ys__n30223 & new_new_n12133__;
  assign new_new_n49478__ = new_new_n12152__ & new_new_n49477__;
  assign new_new_n49479__ = ~new_new_n49476__ & ~new_new_n49478__;
  assign new_new_n49480__ = new_new_n12133__ & new_new_n49258__;
  assign new_new_n49481__ = new_new_n12156__ & new_new_n49480__;
  assign new_new_n49482__ = new_new_n49249__ & new_new_n49475__;
  assign new_new_n49483__ = ~new_new_n49481__ & ~new_new_n49482__;
  assign new_new_n49484__ = new_new_n49479__ & new_new_n49483__;
  assign new_new_n49485__ = ~new_new_n49251__ & ~new_new_n49484__;
  assign ys__n33031 = new_new_n49474__ | new_new_n49485__;
  assign new_new_n49487__ = new_new_n12115__ & new_new_n49251__;
  assign new_new_n49488__ = ~ys__n740 & new_new_n12115__;
  assign new_new_n49489__ = new_new_n12150__ & new_new_n49488__;
  assign new_new_n49490__ = ys__n30223 & new_new_n12115__;
  assign new_new_n49491__ = new_new_n12152__ & new_new_n49490__;
  assign new_new_n49492__ = ~new_new_n49489__ & ~new_new_n49491__;
  assign new_new_n49493__ = new_new_n12115__ & new_new_n49258__;
  assign new_new_n49494__ = new_new_n12156__ & new_new_n49493__;
  assign new_new_n49495__ = new_new_n49249__ & new_new_n49488__;
  assign new_new_n49496__ = ~new_new_n49494__ & ~new_new_n49495__;
  assign new_new_n49497__ = new_new_n49492__ & new_new_n49496__;
  assign new_new_n49498__ = ~new_new_n49251__ & ~new_new_n49497__;
  assign ys__n33032 = new_new_n49487__ | new_new_n49498__;
  assign new_new_n49500__ = new_new_n12057__ & new_new_n49251__;
  assign new_new_n49501__ = ~ys__n740 & new_new_n12057__;
  assign new_new_n49502__ = new_new_n12150__ & new_new_n49501__;
  assign new_new_n49503__ = ys__n30223 & new_new_n12057__;
  assign new_new_n49504__ = new_new_n12152__ & new_new_n49503__;
  assign new_new_n49505__ = ~new_new_n49502__ & ~new_new_n49504__;
  assign new_new_n49506__ = new_new_n12057__ & new_new_n49258__;
  assign new_new_n49507__ = new_new_n12156__ & new_new_n49506__;
  assign new_new_n49508__ = new_new_n49249__ & new_new_n49501__;
  assign new_new_n49509__ = ~new_new_n49507__ & ~new_new_n49508__;
  assign new_new_n49510__ = new_new_n49505__ & new_new_n49509__;
  assign new_new_n49511__ = ~new_new_n49251__ & ~new_new_n49510__;
  assign ys__n33033 = new_new_n49500__ | new_new_n49511__;
  assign new_new_n49513__ = new_new_n10620__ & new_new_n49251__;
  assign new_new_n49514__ = new_new_n10620__ & ~ys__n740;
  assign new_new_n49515__ = new_new_n12150__ & new_new_n49514__;
  assign new_new_n49516__ = new_new_n10620__ & ys__n30223;
  assign new_new_n49517__ = new_new_n12152__ & new_new_n49516__;
  assign new_new_n49518__ = ~new_new_n49515__ & ~new_new_n49517__;
  assign new_new_n49519__ = new_new_n10620__ & new_new_n49258__;
  assign new_new_n49520__ = new_new_n12156__ & new_new_n49519__;
  assign new_new_n49521__ = new_new_n49249__ & new_new_n49514__;
  assign new_new_n49522__ = ~new_new_n49520__ & ~new_new_n49521__;
  assign new_new_n49523__ = new_new_n49518__ & new_new_n49522__;
  assign new_new_n49524__ = ~new_new_n49251__ & ~new_new_n49523__;
  assign ys__n33034 = new_new_n49513__ | new_new_n49524__;
  assign new_new_n49526__ = ~ys__n740 & new_new_n12186__;
  assign new_new_n49527__ = ~ys__n23850 & new_new_n12183__;
  assign new_new_n49528__ = ~new_new_n49526__ & ~new_new_n49527__;
  assign new_new_n49529__ = ~new_new_n12190__ & ~new_new_n49528__;
  assign ys__n33035 = new_new_n12190__ | new_new_n49529__;
  assign new_new_n49531__ = ys__n140 & ~ys__n210;
  assign new_new_n49532__ = new_new_n12165__ & new_new_n49531__;
  assign new_new_n49533__ = ~new_new_n12167__ & ~new_new_n49532__;
  assign new_new_n49534__ = new_new_n12164__ & new_new_n49533__;
  assign new_new_n49535__ = new_new_n16904__ & new_new_n49534__;
  assign new_new_n49536__ = new_new_n12161__ & new_new_n49253__;
  assign new_new_n49537__ = new_new_n12163__ & new_new_n49255__;
  assign new_new_n49538__ = ~new_new_n49536__ & ~new_new_n49537__;
  assign new_new_n49539__ = new_new_n12167__ & new_new_n49259__;
  assign new_new_n49540__ = new_new_n49253__ & new_new_n49532__;
  assign new_new_n49541__ = ~new_new_n49539__ & ~new_new_n49540__;
  assign new_new_n49542__ = new_new_n49538__ & new_new_n49541__;
  assign new_new_n49543__ = ~new_new_n49534__ & ~new_new_n49542__;
  assign ys__n33036 = new_new_n49535__ | new_new_n49543__;
  assign new_new_n49545__ = new_new_n12130__ & new_new_n49534__;
  assign new_new_n49546__ = new_new_n12161__ & new_new_n49267__;
  assign new_new_n49547__ = new_new_n12163__ & new_new_n49269__;
  assign new_new_n49548__ = ~new_new_n49546__ & ~new_new_n49547__;
  assign new_new_n49549__ = new_new_n12167__ & new_new_n49272__;
  assign new_new_n49550__ = new_new_n49267__ & new_new_n49532__;
  assign new_new_n49551__ = ~new_new_n49549__ & ~new_new_n49550__;
  assign new_new_n49552__ = new_new_n49548__ & new_new_n49551__;
  assign new_new_n49553__ = ~new_new_n49534__ & ~new_new_n49552__;
  assign ys__n33037 = new_new_n49545__ | new_new_n49553__;
  assign new_new_n49555__ = new_new_n12112__ & new_new_n49534__;
  assign new_new_n49556__ = new_new_n12161__ & new_new_n49280__;
  assign new_new_n49557__ = new_new_n12163__ & new_new_n49282__;
  assign new_new_n49558__ = ~new_new_n49556__ & ~new_new_n49557__;
  assign new_new_n49559__ = new_new_n12167__ & new_new_n49285__;
  assign new_new_n49560__ = new_new_n49280__ & new_new_n49532__;
  assign new_new_n49561__ = ~new_new_n49559__ & ~new_new_n49560__;
  assign new_new_n49562__ = new_new_n49558__ & new_new_n49561__;
  assign new_new_n49563__ = ~new_new_n49534__ & ~new_new_n49562__;
  assign ys__n33038 = new_new_n49555__ | new_new_n49563__;
  assign new_new_n49565__ = new_new_n12054__ & new_new_n49534__;
  assign new_new_n49566__ = new_new_n12161__ & new_new_n49293__;
  assign new_new_n49567__ = new_new_n12163__ & new_new_n49295__;
  assign new_new_n49568__ = ~new_new_n49566__ & ~new_new_n49567__;
  assign new_new_n49569__ = new_new_n12167__ & new_new_n49298__;
  assign new_new_n49570__ = new_new_n49293__ & new_new_n49532__;
  assign new_new_n49571__ = ~new_new_n49569__ & ~new_new_n49570__;
  assign new_new_n49572__ = new_new_n49568__ & new_new_n49571__;
  assign new_new_n49573__ = ~new_new_n49534__ & ~new_new_n49572__;
  assign ys__n33039 = new_new_n49565__ | new_new_n49573__;
  assign new_new_n49575__ = new_new_n10605__ & new_new_n49534__;
  assign new_new_n49576__ = new_new_n12161__ & new_new_n49306__;
  assign new_new_n49577__ = new_new_n12163__ & new_new_n49308__;
  assign new_new_n49578__ = ~new_new_n49576__ & ~new_new_n49577__;
  assign new_new_n49579__ = new_new_n12167__ & new_new_n49311__;
  assign new_new_n49580__ = new_new_n49306__ & new_new_n49532__;
  assign new_new_n49581__ = ~new_new_n49579__ & ~new_new_n49580__;
  assign new_new_n49582__ = new_new_n49578__ & new_new_n49581__;
  assign new_new_n49583__ = ~new_new_n49534__ & ~new_new_n49582__;
  assign ys__n33040 = new_new_n49575__ | new_new_n49583__;
  assign new_new_n49585__ = new_new_n44241__ & new_new_n49534__;
  assign new_new_n49586__ = new_new_n12161__ & new_new_n49319__;
  assign new_new_n49587__ = new_new_n12163__ & new_new_n49321__;
  assign new_new_n49588__ = ~new_new_n49586__ & ~new_new_n49587__;
  assign new_new_n49589__ = new_new_n12167__ & new_new_n49324__;
  assign new_new_n49590__ = new_new_n49319__ & new_new_n49532__;
  assign new_new_n49591__ = ~new_new_n49589__ & ~new_new_n49590__;
  assign new_new_n49592__ = new_new_n49588__ & new_new_n49591__;
  assign new_new_n49593__ = ~new_new_n49534__ & ~new_new_n49592__;
  assign ys__n33041 = new_new_n49585__ | new_new_n49593__;
  assign new_new_n49595__ = new_new_n26170__ & new_new_n49534__;
  assign new_new_n49596__ = new_new_n12161__ & new_new_n49332__;
  assign new_new_n49597__ = new_new_n12163__ & new_new_n49334__;
  assign new_new_n49598__ = ~new_new_n49596__ & ~new_new_n49597__;
  assign new_new_n49599__ = new_new_n12167__ & new_new_n49337__;
  assign new_new_n49600__ = new_new_n49332__ & new_new_n49532__;
  assign new_new_n49601__ = ~new_new_n49599__ & ~new_new_n49600__;
  assign new_new_n49602__ = new_new_n49598__ & new_new_n49601__;
  assign new_new_n49603__ = ~new_new_n49534__ & ~new_new_n49602__;
  assign ys__n33042 = new_new_n49595__ | new_new_n49603__;
  assign new_new_n49605__ = new_new_n26181__ & new_new_n49534__;
  assign new_new_n49606__ = new_new_n12161__ & new_new_n49345__;
  assign new_new_n49607__ = new_new_n12163__ & new_new_n49347__;
  assign new_new_n49608__ = ~new_new_n49606__ & ~new_new_n49607__;
  assign new_new_n49609__ = new_new_n12167__ & new_new_n49350__;
  assign new_new_n49610__ = new_new_n49345__ & new_new_n49532__;
  assign new_new_n49611__ = ~new_new_n49609__ & ~new_new_n49610__;
  assign new_new_n49612__ = new_new_n49608__ & new_new_n49611__;
  assign new_new_n49613__ = ~new_new_n49534__ & ~new_new_n49612__;
  assign ys__n33043 = new_new_n49605__ | new_new_n49613__;
  assign new_new_n49615__ = new_new_n26192__ & new_new_n49534__;
  assign new_new_n49616__ = new_new_n12161__ & new_new_n49358__;
  assign new_new_n49617__ = new_new_n12163__ & new_new_n49360__;
  assign new_new_n49618__ = ~new_new_n49616__ & ~new_new_n49617__;
  assign new_new_n49619__ = new_new_n12167__ & new_new_n49363__;
  assign new_new_n49620__ = new_new_n49358__ & new_new_n49532__;
  assign new_new_n49621__ = ~new_new_n49619__ & ~new_new_n49620__;
  assign new_new_n49622__ = new_new_n49618__ & new_new_n49621__;
  assign new_new_n49623__ = ~new_new_n49534__ & ~new_new_n49622__;
  assign ys__n33044 = new_new_n49615__ | new_new_n49623__;
  assign new_new_n49625__ = new_new_n16892__ & new_new_n49534__;
  assign new_new_n49626__ = new_new_n12161__ & new_new_n49371__;
  assign new_new_n49627__ = new_new_n12163__ & new_new_n49373__;
  assign new_new_n49628__ = ~new_new_n49626__ & ~new_new_n49627__;
  assign new_new_n49629__ = new_new_n12167__ & new_new_n49376__;
  assign new_new_n49630__ = new_new_n49371__ & new_new_n49532__;
  assign new_new_n49631__ = ~new_new_n49629__ & ~new_new_n49630__;
  assign new_new_n49632__ = new_new_n49628__ & new_new_n49631__;
  assign new_new_n49633__ = ~new_new_n49534__ & ~new_new_n49632__;
  assign ys__n33045 = new_new_n49625__ | new_new_n49633__;
  assign new_new_n49635__ = new_new_n44252__ & new_new_n49534__;
  assign new_new_n49636__ = new_new_n12161__ & new_new_n49384__;
  assign new_new_n49637__ = new_new_n12163__ & new_new_n49386__;
  assign new_new_n49638__ = ~new_new_n49636__ & ~new_new_n49637__;
  assign new_new_n49639__ = new_new_n12167__ & new_new_n49389__;
  assign new_new_n49640__ = new_new_n49384__ & new_new_n49532__;
  assign new_new_n49641__ = ~new_new_n49639__ & ~new_new_n49640__;
  assign new_new_n49642__ = new_new_n49638__ & new_new_n49641__;
  assign new_new_n49643__ = ~new_new_n49534__ & ~new_new_n49642__;
  assign ys__n33046 = new_new_n49635__ | new_new_n49643__;
  assign new_new_n49645__ = new_new_n44263__ & new_new_n49534__;
  assign new_new_n49646__ = new_new_n12161__ & new_new_n49397__;
  assign new_new_n49647__ = new_new_n12163__ & new_new_n49399__;
  assign new_new_n49648__ = ~new_new_n49646__ & ~new_new_n49647__;
  assign new_new_n49649__ = new_new_n12167__ & new_new_n49402__;
  assign new_new_n49650__ = new_new_n49397__ & new_new_n49532__;
  assign new_new_n49651__ = ~new_new_n49649__ & ~new_new_n49650__;
  assign new_new_n49652__ = new_new_n49648__ & new_new_n49651__;
  assign new_new_n49653__ = ~new_new_n49534__ & ~new_new_n49652__;
  assign ys__n33047 = new_new_n49645__ | new_new_n49653__;
  assign new_new_n49655__ = new_new_n44274__ & new_new_n49534__;
  assign new_new_n49656__ = new_new_n12161__ & new_new_n49410__;
  assign new_new_n49657__ = new_new_n12163__ & new_new_n49412__;
  assign new_new_n49658__ = ~new_new_n49656__ & ~new_new_n49657__;
  assign new_new_n49659__ = new_new_n12167__ & new_new_n49415__;
  assign new_new_n49660__ = new_new_n49410__ & new_new_n49532__;
  assign new_new_n49661__ = ~new_new_n49659__ & ~new_new_n49660__;
  assign new_new_n49662__ = new_new_n49658__ & new_new_n49661__;
  assign new_new_n49663__ = ~new_new_n49534__ & ~new_new_n49662__;
  assign ys__n33048 = new_new_n49655__ | new_new_n49663__;
  assign new_new_n49665__ = new_new_n44285__ & new_new_n49534__;
  assign new_new_n49666__ = new_new_n12161__ & new_new_n49423__;
  assign new_new_n49667__ = new_new_n12163__ & new_new_n49425__;
  assign new_new_n49668__ = ~new_new_n49666__ & ~new_new_n49667__;
  assign new_new_n49669__ = new_new_n12167__ & new_new_n49428__;
  assign new_new_n49670__ = new_new_n49423__ & new_new_n49532__;
  assign new_new_n49671__ = ~new_new_n49669__ & ~new_new_n49670__;
  assign new_new_n49672__ = new_new_n49668__ & new_new_n49671__;
  assign new_new_n49673__ = ~new_new_n49534__ & ~new_new_n49672__;
  assign ys__n33049 = new_new_n49665__ | new_new_n49673__;
  assign new_new_n49675__ = new_new_n44298__ & new_new_n49534__;
  assign new_new_n49676__ = new_new_n12161__ & new_new_n49436__;
  assign new_new_n49677__ = new_new_n12163__ & new_new_n49438__;
  assign new_new_n49678__ = ~new_new_n49676__ & ~new_new_n49677__;
  assign new_new_n49679__ = new_new_n12167__ & new_new_n49441__;
  assign new_new_n49680__ = new_new_n49436__ & new_new_n49532__;
  assign new_new_n49681__ = ~new_new_n49679__ & ~new_new_n49680__;
  assign new_new_n49682__ = new_new_n49678__ & new_new_n49681__;
  assign new_new_n49683__ = ~new_new_n49534__ & ~new_new_n49682__;
  assign ys__n33050 = new_new_n49675__ | new_new_n49683__;
  assign new_new_n49685__ = new_new_n44309__ & new_new_n49534__;
  assign new_new_n49686__ = new_new_n12161__ & new_new_n49449__;
  assign new_new_n49687__ = new_new_n12163__ & new_new_n49451__;
  assign new_new_n49688__ = ~new_new_n49686__ & ~new_new_n49687__;
  assign new_new_n49689__ = new_new_n12167__ & new_new_n49454__;
  assign new_new_n49690__ = new_new_n49449__ & new_new_n49532__;
  assign new_new_n49691__ = ~new_new_n49689__ & ~new_new_n49690__;
  assign new_new_n49692__ = new_new_n49688__ & new_new_n49691__;
  assign new_new_n49693__ = ~new_new_n49534__ & ~new_new_n49692__;
  assign ys__n33051 = new_new_n49685__ | new_new_n49693__;
  assign new_new_n49695__ = new_new_n16907__ & new_new_n49534__;
  assign new_new_n49696__ = new_new_n12161__ & new_new_n49462__;
  assign new_new_n49697__ = new_new_n12163__ & new_new_n49464__;
  assign new_new_n49698__ = ~new_new_n49696__ & ~new_new_n49697__;
  assign new_new_n49699__ = new_new_n12167__ & new_new_n49467__;
  assign new_new_n49700__ = new_new_n49462__ & new_new_n49532__;
  assign new_new_n49701__ = ~new_new_n49699__ & ~new_new_n49700__;
  assign new_new_n49702__ = new_new_n49698__ & new_new_n49701__;
  assign new_new_n49703__ = ~new_new_n49534__ & ~new_new_n49702__;
  assign ys__n33052 = new_new_n49695__ | new_new_n49703__;
  assign new_new_n49705__ = new_new_n12133__ & new_new_n49534__;
  assign new_new_n49706__ = new_new_n12161__ & new_new_n49475__;
  assign new_new_n49707__ = new_new_n12163__ & new_new_n49477__;
  assign new_new_n49708__ = ~new_new_n49706__ & ~new_new_n49707__;
  assign new_new_n49709__ = new_new_n12167__ & new_new_n49480__;
  assign new_new_n49710__ = new_new_n49475__ & new_new_n49532__;
  assign new_new_n49711__ = ~new_new_n49709__ & ~new_new_n49710__;
  assign new_new_n49712__ = new_new_n49708__ & new_new_n49711__;
  assign new_new_n49713__ = ~new_new_n49534__ & ~new_new_n49712__;
  assign ys__n33053 = new_new_n49705__ | new_new_n49713__;
  assign new_new_n49715__ = new_new_n12115__ & new_new_n49534__;
  assign new_new_n49716__ = new_new_n12161__ & new_new_n49488__;
  assign new_new_n49717__ = new_new_n12163__ & new_new_n49490__;
  assign new_new_n49718__ = ~new_new_n49716__ & ~new_new_n49717__;
  assign new_new_n49719__ = new_new_n12167__ & new_new_n49493__;
  assign new_new_n49720__ = new_new_n49488__ & new_new_n49532__;
  assign new_new_n49721__ = ~new_new_n49719__ & ~new_new_n49720__;
  assign new_new_n49722__ = new_new_n49718__ & new_new_n49721__;
  assign new_new_n49723__ = ~new_new_n49534__ & ~new_new_n49722__;
  assign ys__n33054 = new_new_n49715__ | new_new_n49723__;
  assign new_new_n49725__ = new_new_n12057__ & new_new_n49534__;
  assign new_new_n49726__ = new_new_n12161__ & new_new_n49501__;
  assign new_new_n49727__ = new_new_n12163__ & new_new_n49503__;
  assign new_new_n49728__ = ~new_new_n49726__ & ~new_new_n49727__;
  assign new_new_n49729__ = new_new_n12167__ & new_new_n49506__;
  assign new_new_n49730__ = new_new_n49501__ & new_new_n49532__;
  assign new_new_n49731__ = ~new_new_n49729__ & ~new_new_n49730__;
  assign new_new_n49732__ = new_new_n49728__ & new_new_n49731__;
  assign new_new_n49733__ = ~new_new_n49534__ & ~new_new_n49732__;
  assign ys__n33055 = new_new_n49725__ | new_new_n49733__;
  assign new_new_n49735__ = new_new_n10620__ & new_new_n49534__;
  assign new_new_n49736__ = new_new_n12161__ & new_new_n49514__;
  assign new_new_n49737__ = new_new_n12163__ & new_new_n49516__;
  assign new_new_n49738__ = ~new_new_n49736__ & ~new_new_n49737__;
  assign new_new_n49739__ = new_new_n12167__ & new_new_n49519__;
  assign new_new_n49740__ = new_new_n49514__ & new_new_n49532__;
  assign new_new_n49741__ = ~new_new_n49739__ & ~new_new_n49740__;
  assign new_new_n49742__ = new_new_n49738__ & new_new_n49741__;
  assign new_new_n49743__ = ~new_new_n49534__ & ~new_new_n49742__;
  assign ys__n33056 = new_new_n49735__ | new_new_n49743__;
  assign new_new_n49745__ = ~ys__n740 & new_new_n12175__;
  assign new_new_n49746__ = ~ys__n23850 & new_new_n12172__;
  assign new_new_n49747__ = ~new_new_n49745__ & ~new_new_n49746__;
  assign new_new_n49748__ = ~new_new_n12179__ & ~new_new_n49747__;
  assign ys__n33058 = new_new_n12179__ | new_new_n49748__;
  assign new_new_n49750__ = ~ys__n138 & ys__n140;
  assign new_new_n49751__ = new_new_n12198__ & new_new_n49750__;
  assign new_new_n49752__ = ~new_new_n12200__ & ~new_new_n49751__;
  assign new_new_n49753__ = new_new_n12197__ & new_new_n49752__;
  assign new_new_n49754__ = new_new_n16904__ & new_new_n49753__;
  assign new_new_n49755__ = new_new_n12194__ & new_new_n49253__;
  assign new_new_n49756__ = new_new_n12196__ & new_new_n49255__;
  assign new_new_n49757__ = ~new_new_n49755__ & ~new_new_n49756__;
  assign new_new_n49758__ = new_new_n12200__ & new_new_n49259__;
  assign new_new_n49759__ = new_new_n49253__ & new_new_n49751__;
  assign new_new_n49760__ = ~new_new_n49758__ & ~new_new_n49759__;
  assign new_new_n49761__ = new_new_n49757__ & new_new_n49760__;
  assign new_new_n49762__ = ~new_new_n49753__ & ~new_new_n49761__;
  assign ys__n33059 = new_new_n49754__ | new_new_n49762__;
  assign new_new_n49764__ = new_new_n12130__ & new_new_n49753__;
  assign new_new_n49765__ = new_new_n12194__ & new_new_n49267__;
  assign new_new_n49766__ = new_new_n12196__ & new_new_n49269__;
  assign new_new_n49767__ = ~new_new_n49765__ & ~new_new_n49766__;
  assign new_new_n49768__ = new_new_n12200__ & new_new_n49272__;
  assign new_new_n49769__ = new_new_n49267__ & new_new_n49751__;
  assign new_new_n49770__ = ~new_new_n49768__ & ~new_new_n49769__;
  assign new_new_n49771__ = new_new_n49767__ & new_new_n49770__;
  assign new_new_n49772__ = ~new_new_n49753__ & ~new_new_n49771__;
  assign ys__n33060 = new_new_n49764__ | new_new_n49772__;
  assign new_new_n49774__ = new_new_n12112__ & new_new_n49753__;
  assign new_new_n49775__ = new_new_n12194__ & new_new_n49280__;
  assign new_new_n49776__ = new_new_n12196__ & new_new_n49282__;
  assign new_new_n49777__ = ~new_new_n49775__ & ~new_new_n49776__;
  assign new_new_n49778__ = new_new_n12200__ & new_new_n49285__;
  assign new_new_n49779__ = new_new_n49280__ & new_new_n49751__;
  assign new_new_n49780__ = ~new_new_n49778__ & ~new_new_n49779__;
  assign new_new_n49781__ = new_new_n49777__ & new_new_n49780__;
  assign new_new_n49782__ = ~new_new_n49753__ & ~new_new_n49781__;
  assign ys__n33061 = new_new_n49774__ | new_new_n49782__;
  assign new_new_n49784__ = new_new_n12054__ & new_new_n49753__;
  assign new_new_n49785__ = new_new_n12194__ & new_new_n49293__;
  assign new_new_n49786__ = new_new_n12196__ & new_new_n49295__;
  assign new_new_n49787__ = ~new_new_n49785__ & ~new_new_n49786__;
  assign new_new_n49788__ = new_new_n12200__ & new_new_n49298__;
  assign new_new_n49789__ = new_new_n49293__ & new_new_n49751__;
  assign new_new_n49790__ = ~new_new_n49788__ & ~new_new_n49789__;
  assign new_new_n49791__ = new_new_n49787__ & new_new_n49790__;
  assign new_new_n49792__ = ~new_new_n49753__ & ~new_new_n49791__;
  assign ys__n33062 = new_new_n49784__ | new_new_n49792__;
  assign new_new_n49794__ = new_new_n10605__ & new_new_n49753__;
  assign new_new_n49795__ = new_new_n12194__ & new_new_n49306__;
  assign new_new_n49796__ = new_new_n12196__ & new_new_n49308__;
  assign new_new_n49797__ = ~new_new_n49795__ & ~new_new_n49796__;
  assign new_new_n49798__ = new_new_n12200__ & new_new_n49311__;
  assign new_new_n49799__ = new_new_n49306__ & new_new_n49751__;
  assign new_new_n49800__ = ~new_new_n49798__ & ~new_new_n49799__;
  assign new_new_n49801__ = new_new_n49797__ & new_new_n49800__;
  assign new_new_n49802__ = ~new_new_n49753__ & ~new_new_n49801__;
  assign ys__n33063 = new_new_n49794__ | new_new_n49802__;
  assign new_new_n49804__ = new_new_n44241__ & new_new_n49753__;
  assign new_new_n49805__ = new_new_n12194__ & new_new_n49319__;
  assign new_new_n49806__ = new_new_n12196__ & new_new_n49321__;
  assign new_new_n49807__ = ~new_new_n49805__ & ~new_new_n49806__;
  assign new_new_n49808__ = new_new_n12200__ & new_new_n49324__;
  assign new_new_n49809__ = new_new_n49319__ & new_new_n49751__;
  assign new_new_n49810__ = ~new_new_n49808__ & ~new_new_n49809__;
  assign new_new_n49811__ = new_new_n49807__ & new_new_n49810__;
  assign new_new_n49812__ = ~new_new_n49753__ & ~new_new_n49811__;
  assign ys__n33064 = new_new_n49804__ | new_new_n49812__;
  assign new_new_n49814__ = new_new_n26170__ & new_new_n49753__;
  assign new_new_n49815__ = new_new_n12194__ & new_new_n49332__;
  assign new_new_n49816__ = new_new_n12196__ & new_new_n49334__;
  assign new_new_n49817__ = ~new_new_n49815__ & ~new_new_n49816__;
  assign new_new_n49818__ = new_new_n12200__ & new_new_n49337__;
  assign new_new_n49819__ = new_new_n49332__ & new_new_n49751__;
  assign new_new_n49820__ = ~new_new_n49818__ & ~new_new_n49819__;
  assign new_new_n49821__ = new_new_n49817__ & new_new_n49820__;
  assign new_new_n49822__ = ~new_new_n49753__ & ~new_new_n49821__;
  assign ys__n33065 = new_new_n49814__ | new_new_n49822__;
  assign new_new_n49824__ = new_new_n26181__ & new_new_n49753__;
  assign new_new_n49825__ = new_new_n12194__ & new_new_n49345__;
  assign new_new_n49826__ = new_new_n12196__ & new_new_n49347__;
  assign new_new_n49827__ = ~new_new_n49825__ & ~new_new_n49826__;
  assign new_new_n49828__ = new_new_n12200__ & new_new_n49350__;
  assign new_new_n49829__ = new_new_n49345__ & new_new_n49751__;
  assign new_new_n49830__ = ~new_new_n49828__ & ~new_new_n49829__;
  assign new_new_n49831__ = new_new_n49827__ & new_new_n49830__;
  assign new_new_n49832__ = ~new_new_n49753__ & ~new_new_n49831__;
  assign ys__n33066 = new_new_n49824__ | new_new_n49832__;
  assign new_new_n49834__ = new_new_n26192__ & new_new_n49753__;
  assign new_new_n49835__ = new_new_n12194__ & new_new_n49358__;
  assign new_new_n49836__ = new_new_n12196__ & new_new_n49360__;
  assign new_new_n49837__ = ~new_new_n49835__ & ~new_new_n49836__;
  assign new_new_n49838__ = new_new_n12200__ & new_new_n49363__;
  assign new_new_n49839__ = new_new_n49358__ & new_new_n49751__;
  assign new_new_n49840__ = ~new_new_n49838__ & ~new_new_n49839__;
  assign new_new_n49841__ = new_new_n49837__ & new_new_n49840__;
  assign new_new_n49842__ = ~new_new_n49753__ & ~new_new_n49841__;
  assign ys__n33067 = new_new_n49834__ | new_new_n49842__;
  assign new_new_n49844__ = new_new_n16892__ & new_new_n49753__;
  assign new_new_n49845__ = new_new_n12194__ & new_new_n49371__;
  assign new_new_n49846__ = new_new_n12196__ & new_new_n49373__;
  assign new_new_n49847__ = ~new_new_n49845__ & ~new_new_n49846__;
  assign new_new_n49848__ = new_new_n12200__ & new_new_n49376__;
  assign new_new_n49849__ = new_new_n49371__ & new_new_n49751__;
  assign new_new_n49850__ = ~new_new_n49848__ & ~new_new_n49849__;
  assign new_new_n49851__ = new_new_n49847__ & new_new_n49850__;
  assign new_new_n49852__ = ~new_new_n49753__ & ~new_new_n49851__;
  assign ys__n33068 = new_new_n49844__ | new_new_n49852__;
  assign new_new_n49854__ = new_new_n44252__ & new_new_n49753__;
  assign new_new_n49855__ = new_new_n12194__ & new_new_n49384__;
  assign new_new_n49856__ = new_new_n12196__ & new_new_n49386__;
  assign new_new_n49857__ = ~new_new_n49855__ & ~new_new_n49856__;
  assign new_new_n49858__ = new_new_n12200__ & new_new_n49389__;
  assign new_new_n49859__ = new_new_n49384__ & new_new_n49751__;
  assign new_new_n49860__ = ~new_new_n49858__ & ~new_new_n49859__;
  assign new_new_n49861__ = new_new_n49857__ & new_new_n49860__;
  assign new_new_n49862__ = ~new_new_n49753__ & ~new_new_n49861__;
  assign ys__n33069 = new_new_n49854__ | new_new_n49862__;
  assign new_new_n49864__ = new_new_n44263__ & new_new_n49753__;
  assign new_new_n49865__ = new_new_n12194__ & new_new_n49397__;
  assign new_new_n49866__ = new_new_n12196__ & new_new_n49399__;
  assign new_new_n49867__ = ~new_new_n49865__ & ~new_new_n49866__;
  assign new_new_n49868__ = new_new_n12200__ & new_new_n49402__;
  assign new_new_n49869__ = new_new_n49397__ & new_new_n49751__;
  assign new_new_n49870__ = ~new_new_n49868__ & ~new_new_n49869__;
  assign new_new_n49871__ = new_new_n49867__ & new_new_n49870__;
  assign new_new_n49872__ = ~new_new_n49753__ & ~new_new_n49871__;
  assign ys__n33070 = new_new_n49864__ | new_new_n49872__;
  assign new_new_n49874__ = new_new_n44274__ & new_new_n49753__;
  assign new_new_n49875__ = new_new_n12194__ & new_new_n49410__;
  assign new_new_n49876__ = new_new_n12196__ & new_new_n49412__;
  assign new_new_n49877__ = ~new_new_n49875__ & ~new_new_n49876__;
  assign new_new_n49878__ = new_new_n12200__ & new_new_n49415__;
  assign new_new_n49879__ = new_new_n49410__ & new_new_n49751__;
  assign new_new_n49880__ = ~new_new_n49878__ & ~new_new_n49879__;
  assign new_new_n49881__ = new_new_n49877__ & new_new_n49880__;
  assign new_new_n49882__ = ~new_new_n49753__ & ~new_new_n49881__;
  assign ys__n33071 = new_new_n49874__ | new_new_n49882__;
  assign new_new_n49884__ = new_new_n44285__ & new_new_n49753__;
  assign new_new_n49885__ = new_new_n12194__ & new_new_n49423__;
  assign new_new_n49886__ = new_new_n12196__ & new_new_n49425__;
  assign new_new_n49887__ = ~new_new_n49885__ & ~new_new_n49886__;
  assign new_new_n49888__ = new_new_n12200__ & new_new_n49428__;
  assign new_new_n49889__ = new_new_n49423__ & new_new_n49751__;
  assign new_new_n49890__ = ~new_new_n49888__ & ~new_new_n49889__;
  assign new_new_n49891__ = new_new_n49887__ & new_new_n49890__;
  assign new_new_n49892__ = ~new_new_n49753__ & ~new_new_n49891__;
  assign ys__n33072 = new_new_n49884__ | new_new_n49892__;
  assign new_new_n49894__ = new_new_n44298__ & new_new_n49753__;
  assign new_new_n49895__ = new_new_n12194__ & new_new_n49436__;
  assign new_new_n49896__ = new_new_n12196__ & new_new_n49438__;
  assign new_new_n49897__ = ~new_new_n49895__ & ~new_new_n49896__;
  assign new_new_n49898__ = new_new_n12200__ & new_new_n49441__;
  assign new_new_n49899__ = new_new_n49436__ & new_new_n49751__;
  assign new_new_n49900__ = ~new_new_n49898__ & ~new_new_n49899__;
  assign new_new_n49901__ = new_new_n49897__ & new_new_n49900__;
  assign new_new_n49902__ = ~new_new_n49753__ & ~new_new_n49901__;
  assign ys__n33073 = new_new_n49894__ | new_new_n49902__;
  assign new_new_n49904__ = new_new_n44309__ & new_new_n49753__;
  assign new_new_n49905__ = new_new_n12194__ & new_new_n49449__;
  assign new_new_n49906__ = new_new_n12196__ & new_new_n49451__;
  assign new_new_n49907__ = ~new_new_n49905__ & ~new_new_n49906__;
  assign new_new_n49908__ = new_new_n12200__ & new_new_n49454__;
  assign new_new_n49909__ = new_new_n49449__ & new_new_n49751__;
  assign new_new_n49910__ = ~new_new_n49908__ & ~new_new_n49909__;
  assign new_new_n49911__ = new_new_n49907__ & new_new_n49910__;
  assign new_new_n49912__ = ~new_new_n49753__ & ~new_new_n49911__;
  assign ys__n33074 = new_new_n49904__ | new_new_n49912__;
  assign new_new_n49914__ = new_new_n16907__ & new_new_n49753__;
  assign new_new_n49915__ = new_new_n12194__ & new_new_n49462__;
  assign new_new_n49916__ = new_new_n12196__ & new_new_n49464__;
  assign new_new_n49917__ = ~new_new_n49915__ & ~new_new_n49916__;
  assign new_new_n49918__ = new_new_n12200__ & new_new_n49467__;
  assign new_new_n49919__ = new_new_n49462__ & new_new_n49751__;
  assign new_new_n49920__ = ~new_new_n49918__ & ~new_new_n49919__;
  assign new_new_n49921__ = new_new_n49917__ & new_new_n49920__;
  assign new_new_n49922__ = ~new_new_n49753__ & ~new_new_n49921__;
  assign ys__n33075 = new_new_n49914__ | new_new_n49922__;
  assign new_new_n49924__ = new_new_n12133__ & new_new_n49753__;
  assign new_new_n49925__ = new_new_n12194__ & new_new_n49475__;
  assign new_new_n49926__ = new_new_n12196__ & new_new_n49477__;
  assign new_new_n49927__ = ~new_new_n49925__ & ~new_new_n49926__;
  assign new_new_n49928__ = new_new_n12200__ & new_new_n49480__;
  assign new_new_n49929__ = new_new_n49475__ & new_new_n49751__;
  assign new_new_n49930__ = ~new_new_n49928__ & ~new_new_n49929__;
  assign new_new_n49931__ = new_new_n49927__ & new_new_n49930__;
  assign new_new_n49932__ = ~new_new_n49753__ & ~new_new_n49931__;
  assign ys__n33076 = new_new_n49924__ | new_new_n49932__;
  assign new_new_n49934__ = new_new_n12115__ & new_new_n49753__;
  assign new_new_n49935__ = new_new_n12194__ & new_new_n49488__;
  assign new_new_n49936__ = new_new_n12196__ & new_new_n49490__;
  assign new_new_n49937__ = ~new_new_n49935__ & ~new_new_n49936__;
  assign new_new_n49938__ = new_new_n12200__ & new_new_n49493__;
  assign new_new_n49939__ = new_new_n49488__ & new_new_n49751__;
  assign new_new_n49940__ = ~new_new_n49938__ & ~new_new_n49939__;
  assign new_new_n49941__ = new_new_n49937__ & new_new_n49940__;
  assign new_new_n49942__ = ~new_new_n49753__ & ~new_new_n49941__;
  assign ys__n33077 = new_new_n49934__ | new_new_n49942__;
  assign new_new_n49944__ = new_new_n12057__ & new_new_n49753__;
  assign new_new_n49945__ = new_new_n12194__ & new_new_n49501__;
  assign new_new_n49946__ = new_new_n12196__ & new_new_n49503__;
  assign new_new_n49947__ = ~new_new_n49945__ & ~new_new_n49946__;
  assign new_new_n49948__ = new_new_n12200__ & new_new_n49506__;
  assign new_new_n49949__ = new_new_n49501__ & new_new_n49751__;
  assign new_new_n49950__ = ~new_new_n49948__ & ~new_new_n49949__;
  assign new_new_n49951__ = new_new_n49947__ & new_new_n49950__;
  assign new_new_n49952__ = ~new_new_n49753__ & ~new_new_n49951__;
  assign ys__n33078 = new_new_n49944__ | new_new_n49952__;
  assign new_new_n49954__ = new_new_n10620__ & new_new_n49753__;
  assign new_new_n49955__ = new_new_n12194__ & new_new_n49514__;
  assign new_new_n49956__ = new_new_n12196__ & new_new_n49516__;
  assign new_new_n49957__ = ~new_new_n49955__ & ~new_new_n49956__;
  assign new_new_n49958__ = new_new_n12200__ & new_new_n49519__;
  assign new_new_n49959__ = new_new_n49514__ & new_new_n49751__;
  assign new_new_n49960__ = ~new_new_n49958__ & ~new_new_n49959__;
  assign new_new_n49961__ = new_new_n49957__ & new_new_n49960__;
  assign new_new_n49962__ = ~new_new_n49753__ & ~new_new_n49961__;
  assign ys__n33079 = new_new_n49954__ | new_new_n49962__;
  assign new_new_n49964__ = ys__n17803 & new_new_n12238__;
  assign new_new_n49965__ = new_new_n12237__ & ~new_new_n24260__;
  assign new_new_n49966__ = ~new_new_n49964__ & ~new_new_n49965__;
  assign ys__n33178 = ys__n920 & ~new_new_n49966__;
  assign new_new_n49968__ = ys__n17804 & ~ys__n30553;
  assign new_new_n49969__ = ys__n30553 & ~new_new_n39641__;
  assign new_new_n49970__ = ~new_new_n49968__ & ~new_new_n49969__;
  assign new_new_n49971__ = new_new_n12238__ & ~new_new_n49970__;
  assign new_new_n49972__ = new_new_n12237__ & ~new_new_n24329__;
  assign new_new_n49973__ = ~new_new_n49971__ & ~new_new_n49972__;
  assign ys__n33179 = ys__n920 & ~new_new_n49973__;
  assign new_new_n49975__ = ys__n17806 & ~ys__n30553;
  assign new_new_n49976__ = ys__n30553 & ~new_new_n39668__;
  assign new_new_n49977__ = ~new_new_n49975__ & ~new_new_n49976__;
  assign new_new_n49978__ = new_new_n12238__ & ~new_new_n49977__;
  assign new_new_n49979__ = new_new_n12237__ & ~new_new_n24401__;
  assign new_new_n49980__ = ~new_new_n49978__ & ~new_new_n49979__;
  assign ys__n33180 = ys__n920 & ~new_new_n49980__;
  assign new_new_n49982__ = ys__n17807 & ~ys__n30553;
  assign new_new_n49983__ = ys__n30553 & ~new_new_n39695__;
  assign new_new_n49984__ = ~new_new_n49982__ & ~new_new_n49983__;
  assign new_new_n49985__ = new_new_n12238__ & ~new_new_n49984__;
  assign new_new_n49986__ = new_new_n12237__ & ~new_new_n24476__;
  assign new_new_n49987__ = ~new_new_n49985__ & ~new_new_n49986__;
  assign ys__n33181 = ys__n920 & ~new_new_n49987__;
  assign new_new_n49989__ = ys__n17809 & ~ys__n30553;
  assign new_new_n49990__ = ys__n30553 & ~new_new_n39720__;
  assign new_new_n49991__ = ~new_new_n49989__ & ~new_new_n49990__;
  assign new_new_n49992__ = new_new_n12238__ & ~new_new_n49991__;
  assign new_new_n49993__ = new_new_n12237__ & ~new_new_n24553__;
  assign new_new_n49994__ = ~new_new_n49992__ & ~new_new_n49993__;
  assign ys__n33182 = ys__n920 & ~new_new_n49994__;
  assign new_new_n49996__ = ys__n17810 & ~ys__n30553;
  assign new_new_n49997__ = ys__n30553 & ~new_new_n39746__;
  assign new_new_n49998__ = ~new_new_n49996__ & ~new_new_n49997__;
  assign new_new_n49999__ = new_new_n12238__ & ~new_new_n49998__;
  assign new_new_n50000__ = new_new_n12237__ & ~new_new_n24629__;
  assign new_new_n50001__ = ~new_new_n49999__ & ~new_new_n50000__;
  assign ys__n33183 = ys__n920 & ~new_new_n50001__;
  assign new_new_n50003__ = ys__n17812 & ~ys__n30553;
  assign new_new_n50004__ = ys__n30553 & ~new_new_n39775__;
  assign new_new_n50005__ = ~new_new_n50003__ & ~new_new_n50004__;
  assign new_new_n50006__ = new_new_n12238__ & ~new_new_n50005__;
  assign new_new_n50007__ = new_new_n12237__ & ~new_new_n24709__;
  assign new_new_n50008__ = ~new_new_n50006__ & ~new_new_n50007__;
  assign ys__n33184 = ys__n920 & ~new_new_n50008__;
  assign new_new_n50010__ = ys__n17813 & ~ys__n30553;
  assign new_new_n50011__ = ys__n30553 & ~new_new_n39804__;
  assign new_new_n50012__ = ~new_new_n50010__ & ~new_new_n50011__;
  assign new_new_n50013__ = new_new_n12238__ & ~new_new_n50012__;
  assign new_new_n50014__ = new_new_n12237__ & ~new_new_n24785__;
  assign new_new_n50015__ = ~new_new_n50013__ & ~new_new_n50014__;
  assign ys__n33185 = ys__n920 & ~new_new_n50015__;
  assign new_new_n50017__ = ys__n17815 & ~ys__n30553;
  assign new_new_n50018__ = ys__n30553 & ~new_new_n39832__;
  assign new_new_n50019__ = ~new_new_n50017__ & ~new_new_n50018__;
  assign new_new_n50020__ = new_new_n12238__ & ~new_new_n50019__;
  assign new_new_n50021__ = new_new_n12237__ & ~new_new_n24866__;
  assign new_new_n50022__ = ~new_new_n50020__ & ~new_new_n50021__;
  assign ys__n33186 = ys__n920 & ~new_new_n50022__;
  assign new_new_n50024__ = ys__n17816 & ~ys__n30553;
  assign new_new_n50025__ = ys__n30553 & ~new_new_n39858__;
  assign new_new_n50026__ = ~new_new_n50024__ & ~new_new_n50025__;
  assign new_new_n50027__ = new_new_n12238__ & ~new_new_n50026__;
  assign new_new_n50028__ = new_new_n12237__ & ~new_new_n24942__;
  assign new_new_n50029__ = ~new_new_n50027__ & ~new_new_n50028__;
  assign ys__n33187 = ys__n920 & ~new_new_n50029__;
  assign new_new_n50031__ = ys__n17818 & ~ys__n30553;
  assign new_new_n50032__ = ys__n30553 & ~new_new_n39887__;
  assign new_new_n50033__ = ~new_new_n50031__ & ~new_new_n50032__;
  assign new_new_n50034__ = new_new_n12238__ & ~new_new_n50033__;
  assign new_new_n50035__ = new_new_n12237__ & ~new_new_n25022__;
  assign new_new_n50036__ = ~new_new_n50034__ & ~new_new_n50035__;
  assign ys__n33188 = ys__n920 & ~new_new_n50036__;
  assign new_new_n50038__ = ys__n17819 & ~ys__n30553;
  assign new_new_n50039__ = ys__n30553 & ~new_new_n39916__;
  assign new_new_n50040__ = ~new_new_n50038__ & ~new_new_n50039__;
  assign new_new_n50041__ = new_new_n12238__ & ~new_new_n50040__;
  assign new_new_n50042__ = new_new_n12237__ & ~new_new_n25098__;
  assign new_new_n50043__ = ~new_new_n50041__ & ~new_new_n50042__;
  assign ys__n33189 = ys__n920 & ~new_new_n50043__;
  assign new_new_n50045__ = ys__n17821 & ~ys__n30553;
  assign new_new_n50046__ = ys__n30553 & ~new_new_n39945__;
  assign new_new_n50047__ = ~new_new_n50045__ & ~new_new_n50046__;
  assign new_new_n50048__ = new_new_n12238__ & ~new_new_n50047__;
  assign new_new_n50049__ = new_new_n12237__ & ~new_new_n25182__;
  assign new_new_n50050__ = ~new_new_n50048__ & ~new_new_n50049__;
  assign ys__n33190 = ys__n920 & ~new_new_n50050__;
  assign new_new_n50052__ = ys__n17822 & ~ys__n30553;
  assign new_new_n50053__ = ys__n30553 & ~new_new_n39974__;
  assign new_new_n50054__ = ~new_new_n50052__ & ~new_new_n50053__;
  assign new_new_n50055__ = new_new_n12238__ & ~new_new_n50054__;
  assign new_new_n50056__ = new_new_n12237__ & ~new_new_n25258__;
  assign new_new_n50057__ = ~new_new_n50055__ & ~new_new_n50056__;
  assign ys__n33191 = ys__n920 & ~new_new_n50057__;
  assign new_new_n50059__ = ys__n17824 & ~ys__n30553;
  assign new_new_n50060__ = ys__n30553 & ~new_new_n40003__;
  assign new_new_n50061__ = ~new_new_n50059__ & ~new_new_n50060__;
  assign new_new_n50062__ = new_new_n12238__ & ~new_new_n50061__;
  assign new_new_n50063__ = new_new_n12237__ & ~new_new_n25338__;
  assign new_new_n50064__ = ~new_new_n50062__ & ~new_new_n50063__;
  assign ys__n33192 = ys__n920 & ~new_new_n50064__;
  assign new_new_n50066__ = ys__n17825 & ~ys__n30553;
  assign new_new_n50067__ = ys__n30553 & ~new_new_n40032__;
  assign new_new_n50068__ = ~new_new_n50066__ & ~new_new_n50067__;
  assign new_new_n50069__ = new_new_n12238__ & ~new_new_n50068__;
  assign new_new_n50070__ = new_new_n12237__ & ~new_new_n25412__;
  assign new_new_n50071__ = ~new_new_n50069__ & ~new_new_n50070__;
  assign ys__n33193 = ys__n920 & ~new_new_n50071__;
  assign new_new_n50073__ = ys__n17827 & ~ys__n30553;
  assign new_new_n50074__ = ys__n30553 & ~new_new_n40060__;
  assign new_new_n50075__ = ~new_new_n50073__ & ~new_new_n50074__;
  assign new_new_n50076__ = new_new_n12238__ & ~new_new_n50075__;
  assign new_new_n50077__ = new_new_n12237__ & ~new_new_n24227__;
  assign new_new_n50078__ = ~new_new_n50076__ & ~new_new_n50077__;
  assign ys__n33194 = ys__n920 & ~new_new_n50078__;
  assign new_new_n50080__ = ys__n17828 & ~ys__n30553;
  assign new_new_n50081__ = ys__n30553 & ~new_new_n40086__;
  assign new_new_n50082__ = ~new_new_n50080__ & ~new_new_n50081__;
  assign new_new_n50083__ = new_new_n12238__ & ~new_new_n50082__;
  assign new_new_n50084__ = new_new_n12237__ & ~new_new_n24306__;
  assign new_new_n50085__ = ~new_new_n50083__ & ~new_new_n50084__;
  assign ys__n33195 = ys__n920 & ~new_new_n50085__;
  assign new_new_n50087__ = ys__n17830 & ~ys__n30553;
  assign new_new_n50088__ = ys__n30553 & ~new_new_n40121__;
  assign new_new_n50089__ = ~new_new_n50087__ & ~new_new_n50088__;
  assign new_new_n50090__ = new_new_n12238__ & ~new_new_n50089__;
  assign new_new_n50091__ = new_new_n12237__ & ~new_new_n24378__;
  assign new_new_n50092__ = ~new_new_n50090__ & ~new_new_n50091__;
  assign ys__n33196 = ys__n920 & ~new_new_n50092__;
  assign new_new_n50094__ = ys__n17831 & ~ys__n30553;
  assign new_new_n50095__ = ys__n30553 & ~new_new_n40156__;
  assign new_new_n50096__ = ~new_new_n50094__ & ~new_new_n50095__;
  assign new_new_n50097__ = new_new_n12238__ & ~new_new_n50096__;
  assign new_new_n50098__ = new_new_n12237__ & ~new_new_n24451__;
  assign new_new_n50099__ = ~new_new_n50097__ & ~new_new_n50098__;
  assign ys__n33197 = ys__n920 & ~new_new_n50099__;
  assign new_new_n50101__ = ys__n17833 & ~ys__n30553;
  assign new_new_n50102__ = ys__n30553 & ~new_new_n40191__;
  assign new_new_n50103__ = ~new_new_n50101__ & ~new_new_n50102__;
  assign new_new_n50104__ = new_new_n12238__ & ~new_new_n50103__;
  assign new_new_n50105__ = new_new_n12237__ & ~new_new_n24530__;
  assign new_new_n50106__ = ~new_new_n50104__ & ~new_new_n50105__;
  assign ys__n33198 = ys__n920 & ~new_new_n50106__;
  assign new_new_n50108__ = ys__n17834 & ~ys__n30553;
  assign new_new_n50109__ = ys__n30553 & ~new_new_n40226__;
  assign new_new_n50110__ = ~new_new_n50108__ & ~new_new_n50109__;
  assign new_new_n50111__ = new_new_n12238__ & ~new_new_n50110__;
  assign new_new_n50112__ = new_new_n12237__ & ~new_new_n24603__;
  assign new_new_n50113__ = ~new_new_n50111__ & ~new_new_n50112__;
  assign ys__n33199 = ys__n920 & ~new_new_n50113__;
  assign new_new_n50115__ = ys__n17836 & ~ys__n30553;
  assign new_new_n50116__ = ys__n30553 & ~new_new_n40264__;
  assign new_new_n50117__ = ~new_new_n50115__ & ~new_new_n50116__;
  assign new_new_n50118__ = new_new_n12238__ & ~new_new_n50117__;
  assign new_new_n50119__ = new_new_n12237__ & ~new_new_n24683__;
  assign new_new_n50120__ = ~new_new_n50118__ & ~new_new_n50119__;
  assign ys__n33200 = ys__n920 & ~new_new_n50120__;
  assign new_new_n50122__ = ys__n17837 & ~ys__n30553;
  assign new_new_n50123__ = ys__n30553 & ~new_new_n40302__;
  assign new_new_n50124__ = ~new_new_n50122__ & ~new_new_n50123__;
  assign new_new_n50125__ = new_new_n12238__ & ~new_new_n50124__;
  assign new_new_n50126__ = new_new_n12237__ & ~new_new_n24759__;
  assign new_new_n50127__ = ~new_new_n50125__ & ~new_new_n50126__;
  assign ys__n33201 = ys__n920 & ~new_new_n50127__;
  assign new_new_n50129__ = ys__n17839 & ~ys__n30553;
  assign new_new_n50130__ = ys__n30553 & ~new_new_n40340__;
  assign new_new_n50131__ = ~new_new_n50129__ & ~new_new_n50130__;
  assign new_new_n50132__ = new_new_n12238__ & ~new_new_n50131__;
  assign new_new_n50133__ = new_new_n12237__ & ~new_new_n24843__;
  assign new_new_n50134__ = ~new_new_n50132__ & ~new_new_n50133__;
  assign ys__n33202 = ys__n920 & ~new_new_n50134__;
  assign new_new_n50136__ = ys__n17840 & ~ys__n30553;
  assign new_new_n50137__ = ys__n30553 & ~new_new_n40375__;
  assign new_new_n50138__ = ~new_new_n50136__ & ~new_new_n50137__;
  assign new_new_n50139__ = new_new_n12238__ & ~new_new_n50138__;
  assign new_new_n50140__ = new_new_n12237__ & ~new_new_n24916__;
  assign new_new_n50141__ = ~new_new_n50139__ & ~new_new_n50140__;
  assign ys__n33203 = ys__n920 & ~new_new_n50141__;
  assign new_new_n50143__ = ys__n17842 & ~ys__n30553;
  assign new_new_n50144__ = ys__n30553 & ~new_new_n40413__;
  assign new_new_n50145__ = ~new_new_n50143__ & ~new_new_n50144__;
  assign new_new_n50146__ = new_new_n12238__ & ~new_new_n50145__;
  assign new_new_n50147__ = new_new_n12237__ & ~new_new_n24996__;
  assign new_new_n50148__ = ~new_new_n50146__ & ~new_new_n50147__;
  assign ys__n33204 = ys__n920 & ~new_new_n50148__;
  assign new_new_n50150__ = ys__n17843 & ~ys__n30553;
  assign new_new_n50151__ = ys__n30553 & ~new_new_n40451__;
  assign new_new_n50152__ = ~new_new_n50150__ & ~new_new_n50151__;
  assign new_new_n50153__ = new_new_n12238__ & ~new_new_n50152__;
  assign new_new_n50154__ = new_new_n12237__ & ~new_new_n25072__;
  assign new_new_n50155__ = ~new_new_n50153__ & ~new_new_n50154__;
  assign ys__n33205 = ys__n920 & ~new_new_n50155__;
  assign new_new_n50157__ = ys__n17845 & ~ys__n30553;
  assign new_new_n50158__ = ys__n30553 & ~new_new_n40489__;
  assign new_new_n50159__ = ~new_new_n50157__ & ~new_new_n50158__;
  assign new_new_n50160__ = new_new_n12238__ & ~new_new_n50159__;
  assign new_new_n50161__ = new_new_n12237__ & ~new_new_n25156__;
  assign new_new_n50162__ = ~new_new_n50160__ & ~new_new_n50161__;
  assign ys__n33206 = ys__n920 & ~new_new_n50162__;
  assign new_new_n50164__ = ys__n17846 & ~ys__n30553;
  assign new_new_n50165__ = ys__n30553 & ~new_new_n40526__;
  assign new_new_n50166__ = ~new_new_n50164__ & ~new_new_n50165__;
  assign new_new_n50167__ = new_new_n12238__ & ~new_new_n50166__;
  assign new_new_n50168__ = new_new_n12237__ & ~new_new_n25232__;
  assign new_new_n50169__ = ~new_new_n50167__ & ~new_new_n50168__;
  assign ys__n33207 = ys__n920 & ~new_new_n50169__;
  assign new_new_n50171__ = ys__n17848 & ~ys__n30553;
  assign new_new_n50172__ = ys__n30553 & ~new_new_n40564__;
  assign new_new_n50173__ = ~new_new_n50171__ & ~new_new_n50172__;
  assign new_new_n50174__ = new_new_n12238__ & ~new_new_n50173__;
  assign new_new_n50175__ = new_new_n12237__ & ~new_new_n25312__;
  assign new_new_n50176__ = ~new_new_n50174__ & ~new_new_n50175__;
  assign ys__n33208 = ys__n920 & ~new_new_n50176__;
  assign new_new_n50178__ = ys__n17849 & ~ys__n30553;
  assign new_new_n50179__ = ys__n30553 & ~new_new_n40601__;
  assign new_new_n50180__ = ~new_new_n50178__ & ~new_new_n50179__;
  assign new_new_n50181__ = new_new_n12238__ & ~new_new_n50180__;
  assign new_new_n50182__ = new_new_n12237__ & ~new_new_n25386__;
  assign new_new_n50183__ = ~new_new_n50181__ & ~new_new_n50182__;
  assign ys__n33209 = ys__n920 & ~new_new_n50183__;
  assign new_new_n50185__ = ~ys__n740 & new_new_n12208__;
  assign new_new_n50186__ = ~ys__n23850 & new_new_n12205__;
  assign new_new_n50187__ = ~new_new_n50185__ & ~new_new_n50186__;
  assign new_new_n50188__ = ~new_new_n12212__ & ~new_new_n50187__;
  assign ys__n33211 = new_new_n12212__ | new_new_n50188__;
  assign new_new_n50190__ = new_new_n11175__ & ~new_new_n11628__;
  assign ys__n33366 = new_new_n10820__ & new_new_n50190__;
  assign ys__n33438 = ~ys__n1084 & ~new_new_n10845__;
  assign new_new_n50193__ = ~ys__n30216 & ~ys__n30219;
  assign new_new_n50194__ = new_new_n22487__ & new_new_n50193__;
  assign new_new_n50195__ = ys__n1106 & ~new_new_n50194__;
  assign new_new_n50196__ = ~ys__n24464 & ~ys__n24483;
  assign new_new_n50197__ = ~ys__n38649 & new_new_n50196__;
  assign new_new_n50198__ = ~ys__n1116 & ~ys__n1119;
  assign new_new_n50199__ = ~ys__n24461 & ~ys__n24463;
  assign new_new_n50200__ = new_new_n50198__ & new_new_n50199__;
  assign new_new_n50201__ = new_new_n13991__ & new_new_n22453__;
  assign new_new_n50202__ = new_new_n50200__ & new_new_n50201__;
  assign new_new_n50203__ = new_new_n50197__ & new_new_n50202__;
  assign ys__n33454 = ~new_new_n50195__ & new_new_n50203__;
  assign new_new_n50205__ = ys__n1153 & ys__n33515;
  assign new_new_n50206__ = new_new_n16222__ & new_new_n50193__;
  assign new_new_n50207__ = ys__n1151 & ~new_new_n50206__;
  assign new_new_n50208__ = ys__n33515 & new_new_n50207__;
  assign new_new_n50209__ = new_new_n23463__ & ~new_new_n50208__;
  assign ys__n33514 = ~new_new_n50205__ & new_new_n50209__;
  assign ys__n34952 = ~ys__n18166 & ~ys__n18165;
  assign ys__n34953 = ~ys__n2651 & ~ys__n18166;
  assign new_new_n50213__ = ys__n18317 & new_new_n12273__;
  assign ys__n34962 = new_new_n12284__ & new_new_n50213__;
  assign new_new_n50215__ = ys__n46248 & new_new_n43188__;
  assign new_new_n50216__ = ~ys__n46242 & ~ys__n46244;
  assign new_new_n50217__ = ~ys__n46245 & ~ys__n46247;
  assign new_new_n50218__ = new_new_n50216__ & new_new_n50217__;
  assign ys__n35052 = new_new_n50215__ | ~new_new_n50218__;
  assign new_new_n50220__ = ys__n33081 & ~ys__n33080;
  assign new_new_n50221__ = ~ys__n33081 & ys__n33080;
  assign ys__n35144 = new_new_n50220__ | new_new_n50221__;
  assign new_new_n50223__ = ~ys__n33081 & ~ys__n33080;
  assign new_new_n50224__ = ys__n33082 & new_new_n50223__;
  assign new_new_n50225__ = ~ys__n33082 & ~new_new_n50223__;
  assign ys__n35146 = new_new_n50224__ | new_new_n50225__;
  assign new_new_n50227__ = ~ys__n33082 & new_new_n50223__;
  assign new_new_n50228__ = ys__n33083 & new_new_n50227__;
  assign new_new_n50229__ = ~ys__n33083 & ~new_new_n50227__;
  assign ys__n35148 = new_new_n50228__ | new_new_n50229__;
  assign new_new_n50231__ = ~ys__n33082 & ~ys__n33083;
  assign new_new_n50232__ = new_new_n50223__ & new_new_n50231__;
  assign new_new_n50233__ = ys__n33084 & new_new_n50232__;
  assign new_new_n50234__ = ~ys__n33084 & ~new_new_n50232__;
  assign ys__n35150 = new_new_n50233__ | new_new_n50234__;
  assign new_new_n50236__ = ~ys__n33084 & new_new_n50232__;
  assign new_new_n50237__ = ys__n33085 & new_new_n50236__;
  assign new_new_n50238__ = ~ys__n33085 & ~new_new_n50236__;
  assign ys__n35152 = new_new_n50237__ | new_new_n50238__;
  assign new_new_n50240__ = ~ys__n33085 & ~ys__n33084;
  assign new_new_n50241__ = new_new_n50232__ & new_new_n50240__;
  assign new_new_n50242__ = ys__n33086 & new_new_n50241__;
  assign new_new_n50243__ = ~ys__n33086 & ~new_new_n50241__;
  assign ys__n35154 = new_new_n50242__ | new_new_n50243__;
  assign new_new_n50245__ = ~ys__n33086 & new_new_n50241__;
  assign new_new_n50246__ = ys__n33087 & new_new_n50245__;
  assign new_new_n50247__ = ~ys__n33087 & ~new_new_n50245__;
  assign ys__n35156 = new_new_n50246__ | new_new_n50247__;
  assign new_new_n50249__ = ~ys__n33087 & ~ys__n33086;
  assign new_new_n50250__ = new_new_n50240__ & new_new_n50249__;
  assign new_new_n50251__ = new_new_n50232__ & new_new_n50250__;
  assign new_new_n50252__ = ys__n33088 & new_new_n50251__;
  assign new_new_n50253__ = ~ys__n33088 & ~new_new_n50251__;
  assign ys__n35158 = new_new_n50252__ | new_new_n50253__;
  assign new_new_n50255__ = ~ys__n33088 & new_new_n50251__;
  assign new_new_n50256__ = ys__n33089 & new_new_n50255__;
  assign new_new_n50257__ = ~ys__n33089 & ~new_new_n50255__;
  assign ys__n35160 = new_new_n50256__ | new_new_n50257__;
  assign new_new_n50259__ = ~ys__n33089 & ~ys__n33088;
  assign new_new_n50260__ = new_new_n50251__ & new_new_n50259__;
  assign new_new_n50261__ = ys__n33090 & new_new_n50260__;
  assign new_new_n50262__ = ~ys__n33090 & ~new_new_n50260__;
  assign ys__n35162 = new_new_n50261__ | new_new_n50262__;
  assign new_new_n50264__ = ~ys__n33090 & new_new_n50260__;
  assign new_new_n50265__ = ys__n33091 & new_new_n50264__;
  assign new_new_n50266__ = ~ys__n33091 & ~new_new_n50264__;
  assign ys__n35164 = new_new_n50265__ | new_new_n50266__;
  assign new_new_n50268__ = ~ys__n33091 & ~ys__n33090;
  assign new_new_n50269__ = new_new_n50259__ & new_new_n50268__;
  assign new_new_n50270__ = new_new_n50251__ & new_new_n50269__;
  assign new_new_n50271__ = ys__n33092 & new_new_n50270__;
  assign new_new_n50272__ = ~ys__n33092 & ~new_new_n50270__;
  assign ys__n35166 = new_new_n50271__ | new_new_n50272__;
  assign new_new_n50274__ = ~ys__n33092 & new_new_n50270__;
  assign new_new_n50275__ = ys__n33093 & new_new_n50274__;
  assign new_new_n50276__ = ~ys__n33093 & ~new_new_n50274__;
  assign ys__n35168 = new_new_n50275__ | new_new_n50276__;
  assign new_new_n50278__ = ~ys__n33093 & ~ys__n33092;
  assign new_new_n50279__ = new_new_n50270__ & new_new_n50278__;
  assign new_new_n50280__ = ys__n33094 & new_new_n50279__;
  assign new_new_n50281__ = ~ys__n33094 & ~new_new_n50279__;
  assign ys__n35170 = new_new_n50280__ | new_new_n50281__;
  assign new_new_n50283__ = ~ys__n33094 & new_new_n50279__;
  assign new_new_n50284__ = ys__n33095 & new_new_n50283__;
  assign new_new_n50285__ = ~ys__n33095 & ~new_new_n50283__;
  assign ys__n35172 = new_new_n50284__ | new_new_n50285__;
  assign new_new_n50287__ = ~ys__n33095 & ~ys__n33094;
  assign new_new_n50288__ = new_new_n50278__ & new_new_n50287__;
  assign new_new_n50289__ = new_new_n50269__ & new_new_n50288__;
  assign new_new_n50290__ = new_new_n50251__ & new_new_n50289__;
  assign new_new_n50291__ = ys__n33096 & new_new_n50290__;
  assign new_new_n50292__ = ~ys__n33096 & ~new_new_n50290__;
  assign ys__n35174 = new_new_n50291__ | new_new_n50292__;
  assign new_new_n50294__ = ~ys__n33096 & new_new_n50290__;
  assign new_new_n50295__ = ys__n33097 & new_new_n50294__;
  assign new_new_n50296__ = ~ys__n33097 & ~new_new_n50294__;
  assign ys__n35176 = new_new_n50295__ | new_new_n50296__;
  assign new_new_n50298__ = ~ys__n33096 & ~ys__n33097;
  assign new_new_n50299__ = new_new_n50290__ & new_new_n50298__;
  assign new_new_n50300__ = ys__n33098 & new_new_n50299__;
  assign new_new_n50301__ = ~ys__n33098 & ~new_new_n50299__;
  assign ys__n35178 = new_new_n50300__ | new_new_n50301__;
  assign new_new_n50303__ = ~ys__n33098 & new_new_n50299__;
  assign new_new_n50304__ = ys__n33099 & new_new_n50303__;
  assign new_new_n50305__ = ~ys__n33099 & ~new_new_n50303__;
  assign ys__n35180 = new_new_n50304__ | new_new_n50305__;
  assign new_new_n50307__ = ~ys__n33098 & ~ys__n33099;
  assign new_new_n50308__ = new_new_n50298__ & new_new_n50307__;
  assign new_new_n50309__ = new_new_n50290__ & new_new_n50308__;
  assign new_new_n50310__ = ys__n33100 & new_new_n50309__;
  assign new_new_n50311__ = ~ys__n33100 & ~new_new_n50309__;
  assign ys__n35182 = new_new_n50310__ | new_new_n50311__;
  assign new_new_n50313__ = ~ys__n33100 & new_new_n50309__;
  assign new_new_n50314__ = ys__n33101 & new_new_n50313__;
  assign new_new_n50315__ = ~ys__n33101 & ~new_new_n50313__;
  assign ys__n35184 = new_new_n50314__ | new_new_n50315__;
  assign new_new_n50317__ = ~ys__n33100 & ~ys__n33101;
  assign new_new_n50318__ = new_new_n50309__ & new_new_n50317__;
  assign new_new_n50319__ = ys__n33102 & new_new_n50318__;
  assign new_new_n50320__ = ~ys__n33102 & ~new_new_n50318__;
  assign ys__n35186 = new_new_n50319__ | new_new_n50320__;
  assign new_new_n50322__ = ~ys__n33102 & new_new_n50318__;
  assign new_new_n50323__ = ys__n33103 & new_new_n50322__;
  assign new_new_n50324__ = ~ys__n33103 & ~new_new_n50322__;
  assign ys__n35188 = new_new_n50323__ | new_new_n50324__;
  assign new_new_n50326__ = ~ys__n33102 & ~ys__n33103;
  assign new_new_n50327__ = new_new_n50317__ & new_new_n50326__;
  assign new_new_n50328__ = new_new_n50308__ & new_new_n50327__;
  assign new_new_n50329__ = new_new_n50290__ & new_new_n50328__;
  assign new_new_n50330__ = ys__n33104 & new_new_n50329__;
  assign new_new_n50331__ = ~ys__n33104 & ~new_new_n50329__;
  assign ys__n35190 = new_new_n50330__ | new_new_n50331__;
  assign new_new_n50333__ = ~ys__n33104 & new_new_n50329__;
  assign new_new_n50334__ = ys__n33105 & new_new_n50333__;
  assign new_new_n50335__ = ~ys__n33105 & ~new_new_n50333__;
  assign ys__n35192 = new_new_n50334__ | new_new_n50335__;
  assign new_new_n50337__ = ~ys__n33104 & ~ys__n33105;
  assign new_new_n50338__ = new_new_n50329__ & new_new_n50337__;
  assign new_new_n50339__ = ys__n33106 & new_new_n50338__;
  assign new_new_n50340__ = ~ys__n33106 & ~new_new_n50338__;
  assign ys__n35194 = new_new_n50339__ | new_new_n50340__;
  assign new_new_n50342__ = ~ys__n33106 & new_new_n50338__;
  assign new_new_n50343__ = ys__n33107 & new_new_n50342__;
  assign new_new_n50344__ = ~ys__n33107 & ~new_new_n50342__;
  assign ys__n35196 = new_new_n50343__ | new_new_n50344__;
  assign new_new_n50346__ = ~ys__n33106 & ~ys__n33107;
  assign new_new_n50347__ = new_new_n50337__ & new_new_n50346__;
  assign new_new_n50348__ = new_new_n50329__ & new_new_n50347__;
  assign new_new_n50349__ = ys__n33108 & new_new_n50348__;
  assign new_new_n50350__ = ~ys__n33108 & ~new_new_n50348__;
  assign ys__n35198 = new_new_n50349__ | new_new_n50350__;
  assign new_new_n50352__ = ~ys__n33108 & new_new_n50348__;
  assign new_new_n50353__ = ys__n33109 & new_new_n50352__;
  assign new_new_n50354__ = ~ys__n33109 & ~new_new_n50352__;
  assign ys__n35200 = new_new_n50353__ | new_new_n50354__;
  assign new_new_n50356__ = ~ys__n33108 & ~ys__n33109;
  assign new_new_n50357__ = new_new_n50348__ & new_new_n50356__;
  assign new_new_n50358__ = ys__n33110 & new_new_n50357__;
  assign new_new_n50359__ = ~ys__n33110 & ~new_new_n50357__;
  assign ys__n35202 = new_new_n50358__ | new_new_n50359__;
  assign new_new_n50361__ = ~ys__n33110 & new_new_n50357__;
  assign new_new_n50362__ = ys__n33111 & new_new_n50361__;
  assign new_new_n50363__ = ~ys__n33111 & ~new_new_n50361__;
  assign ys__n35204 = new_new_n50362__ | new_new_n50363__;
  assign new_new_n50365__ = ~ys__n33110 & ~ys__n33111;
  assign new_new_n50366__ = new_new_n50356__ & new_new_n50365__;
  assign new_new_n50367__ = new_new_n50347__ & new_new_n50366__;
  assign new_new_n50368__ = new_new_n50290__ & new_new_n50367__;
  assign new_new_n50369__ = new_new_n50328__ & new_new_n50368__;
  assign new_new_n50370__ = ys__n30668 & new_new_n50369__;
  assign new_new_n50371__ = ~ys__n30668 & ~new_new_n50369__;
  assign ys__n35206 = new_new_n50370__ | new_new_n50371__;
  assign new_new_n50373__ = ys__n456 & ~ys__n710;
  assign new_new_n50374__ = ~ys__n456 & ys__n710;
  assign ys__n35402 = new_new_n50373__ | new_new_n50374__;
  assign new_new_n50376__ = ~ys__n708 & new_new_n16496__;
  assign new_new_n50377__ = ys__n708 & ~new_new_n16496__;
  assign ys__n35404 = new_new_n50376__ | new_new_n50377__;
  assign new_new_n50379__ = ys__n708 & new_new_n16496__;
  assign new_new_n50380__ = ~ys__n706 & new_new_n50379__;
  assign new_new_n50381__ = ys__n706 & ~new_new_n50379__;
  assign ys__n35406 = new_new_n50380__ | new_new_n50381__;
  assign new_new_n50383__ = ~ys__n702 & new_new_n16498__;
  assign new_new_n50384__ = ys__n702 & ~new_new_n16498__;
  assign ys__n35408 = new_new_n50383__ | new_new_n50384__;
  assign new_new_n50386__ = ys__n702 & new_new_n16498__;
  assign new_new_n50387__ = ~ys__n700 & new_new_n50386__;
  assign new_new_n50388__ = ys__n700 & ~new_new_n50386__;
  assign ys__n35410 = new_new_n50387__ | new_new_n50388__;
  assign new_new_n50390__ = new_new_n16498__ & new_new_n16499__;
  assign new_new_n50391__ = ~ys__n704 & new_new_n50390__;
  assign new_new_n50392__ = ys__n704 & ~new_new_n50390__;
  assign ys__n35412 = new_new_n50391__ | new_new_n50392__;
  assign new_new_n50394__ = ys__n414 & ~ys__n728;
  assign new_new_n50395__ = ~ys__n414 & ys__n728;
  assign ys__n35706 = new_new_n50394__ | new_new_n50395__;
  assign new_new_n50397__ = ~ys__n726 & new_new_n16482__;
  assign new_new_n50398__ = ys__n726 & ~new_new_n16482__;
  assign ys__n35708 = new_new_n50397__ | new_new_n50398__;
  assign new_new_n50400__ = ys__n726 & new_new_n16482__;
  assign new_new_n50401__ = ~ys__n724 & new_new_n50400__;
  assign new_new_n50402__ = ys__n724 & ~new_new_n50400__;
  assign ys__n35710 = new_new_n50401__ | new_new_n50402__;
  assign new_new_n50404__ = ~ys__n720 & new_new_n16484__;
  assign new_new_n50405__ = ys__n720 & ~new_new_n16484__;
  assign ys__n35712 = new_new_n50404__ | new_new_n50405__;
  assign new_new_n50407__ = ys__n720 & new_new_n16484__;
  assign new_new_n50408__ = ~ys__n718 & new_new_n50407__;
  assign new_new_n50409__ = ys__n718 & ~new_new_n50407__;
  assign ys__n35714 = new_new_n50408__ | new_new_n50409__;
  assign new_new_n50411__ = new_new_n16484__ & new_new_n16485__;
  assign new_new_n50412__ = ~ys__n722 & new_new_n50411__;
  assign new_new_n50413__ = ys__n722 & ~new_new_n50411__;
  assign ys__n35716 = new_new_n50412__ | new_new_n50413__;
  assign new_new_n50415__ = ys__n3214 & ys__n19159;
  assign new_new_n50416__ = ~new_new_n11791__ & ~new_new_n50415__;
  assign ys__n37687 = new_new_n11800__ | ~new_new_n50416__;
  assign ys__n37695 = ~new_new_n12097__ & new_new_n12103__;
  assign ys__n37697 = ~new_new_n12098__ & new_new_n12103__;
  assign new_new_n50420__ = ys__n33313 & ~new_new_n12103__;
  assign new_new_n50421__ = ys__n3214 & ~new_new_n50420__;
  assign ys__n37699 = new_new_n17020__ | new_new_n50421__;
  assign new_new_n50423__ = ys__n33311 & ~ys__n33313;
  assign new_new_n50424__ = ~new_new_n12103__ & new_new_n50423__;
  assign new_new_n50425__ = ys__n18070 & ~new_new_n50424__;
  assign ys__n37702 = new_new_n11125__ | new_new_n50425__;
  assign new_new_n50427__ = ys__n33309 & ~ys__n33311;
  assign new_new_n50428__ = ~ys__n33313 & new_new_n50427__;
  assign new_new_n50429__ = ~new_new_n12103__ & new_new_n50428__;
  assign new_new_n50430__ = ys__n18071 & ~new_new_n50429__;
  assign ys__n37707 = new_new_n11122__ | new_new_n50430__;
  assign new_new_n50432__ = ~ys__n844 & ~ys__n37710;
  assign new_new_n50433__ = ~ys__n37712 & ys__n37713;
  assign ys__n37714 = new_new_n50432__ & new_new_n50433__;
  assign ys__n37731 = ys__n24112 & ~ys__n33317;
  assign ys__n37732 = ys__n18380 & ys__n33317;
  assign ys__n37733 = ys__n18383 & ys__n33317;
  assign new_new_n50438__ = ~ys__n37668 & ys__n37669;
  assign new_new_n50439__ = ys__n37668 & ~ys__n37669;
  assign new_new_n50440__ = ~new_new_n50438__ & ~new_new_n50439__;
  assign new_new_n50441__ = ~ys__n18393 & ~new_new_n50440__;
  assign new_new_n50442__ = ys__n18393 & ys__n27598;
  assign new_new_n50443__ = ~new_new_n50441__ & ~new_new_n50442__;
  assign ys__n37738 = ys__n33320 & ~new_new_n50443__;
  assign new_new_n50445__ = ys__n33318 & ~ys__n33320;
  assign new_new_n50446__ = ~new_new_n50443__ & new_new_n50445__;
  assign ys__n37739 = new_new_n33596__ | new_new_n50446__;
  assign new_new_n50448__ = ~ys__n33318 & ~ys__n33320;
  assign new_new_n50449__ = ~new_new_n50443__ & new_new_n50448__;
  assign new_new_n50450__ = ys__n18208 & new_new_n33693__;
  assign ys__n37741 = new_new_n50449__ | new_new_n50450__;
  assign new_new_n50452__ = ys__n812 & ~ys__n3250;
  assign new_new_n50453__ = ys__n19171 & ys__n18287;
  assign new_new_n50454__ = ~ys__n18284 & new_new_n50453__;
  assign new_new_n50455__ = ys__n18284 & ys__n18763;
  assign new_new_n50456__ = ~new_new_n50454__ & ~new_new_n50455__;
  assign new_new_n50457__ = ~ys__n18281 & ~new_new_n50456__;
  assign new_new_n50458__ = ys__n18281 & ys__n18652;
  assign new_new_n50459__ = ~new_new_n50457__ & ~new_new_n50458__;
  assign new_new_n50460__ = ~ys__n18278 & ~new_new_n50459__;
  assign new_new_n50461__ = ~ys__n18278 & ~new_new_n50460__;
  assign new_new_n50462__ = ~ys__n3252 & ~new_new_n50461__;
  assign new_new_n50463__ = new_new_n50452__ & new_new_n50462__;
  assign new_new_n50464__ = ys__n804 & ys__n806;
  assign new_new_n50465__ = ys__n808 & ys__n810;
  assign new_new_n50466__ = new_new_n50464__ & new_new_n50465__;
  assign new_new_n50467__ = ys__n796 & ys__n798;
  assign new_new_n50468__ = ys__n800 & ys__n802;
  assign new_new_n50469__ = new_new_n50467__ & new_new_n50468__;
  assign new_new_n50470__ = new_new_n50466__ & new_new_n50469__;
  assign ys__n37742 = new_new_n50463__ & new_new_n50470__;
  assign ys__n38180 = ys__n38179 | ys__n18088;
  assign new_new_n50473__ = ~ys__n240 & new_new_n33805__;
  assign new_new_n50474__ = ~new_new_n33805__ & new_new_n50473__;
  assign new_new_n50475__ = ~ys__n1535 & ~new_new_n50474__;
  assign new_new_n50476__ = ~ys__n1535 & ~new_new_n50475__;
  assign new_new_n50477__ = ys__n28243 & ~ys__n4566;
  assign ys__n38182 = ~new_new_n50476__ & new_new_n50477__;
  assign ys__n38184 = ys__n38183 & ~ys__n4566;
  assign ys__n38205 = ~ys__n23627 | ~ys__n738;
  assign new_new_n50481__ = ys__n45704 & new_new_n12945__;
  assign new_new_n50482__ = ys__n45541 & new_new_n13255__;
  assign new_new_n50483__ = ~new_new_n50481__ & ~new_new_n50482__;
  assign new_new_n50484__ = ys__n45377 & new_new_n13566__;
  assign new_new_n50485__ = ys__n45214 & new_new_n13876__;
  assign new_new_n50486__ = ~new_new_n50484__ & ~new_new_n50485__;
  assign new_new_n50487__ = new_new_n50483__ & new_new_n50486__;
  assign new_new_n50488__ = ~new_new_n13883__ & ~new_new_n50487__;
  assign new_new_n50489__ = ~ys__n38282 & ~ys__n38283;
  assign new_new_n50490__ = ~ys__n38286 & ~ys__n38300;
  assign new_new_n50491__ = new_new_n50489__ & new_new_n50490__;
  assign new_new_n50492__ = ~new_new_n50488__ & new_new_n50491__;
  assign ys__n38207 = ~ys__n4566 & ~new_new_n50492__;
  assign new_new_n50494__ = ys__n45771 & ys__n46074;
  assign new_new_n50495__ = ~ys__n45771 & ~ys__n46074;
  assign new_new_n50496__ = ~ys__n46116 & ~new_new_n50495__;
  assign new_new_n50497__ = ~new_new_n50494__ & new_new_n50496__;
  assign new_new_n50498__ = ys__n45774 & ys__n46076;
  assign new_new_n50499__ = ~ys__n45774 & ~ys__n46076;
  assign new_new_n50500__ = ~ys__n46117 & ~new_new_n50499__;
  assign new_new_n50501__ = ~new_new_n50498__ & new_new_n50500__;
  assign new_new_n50502__ = ~new_new_n50497__ & ~new_new_n50501__;
  assign new_new_n50503__ = ys__n45777 & ys__n46078;
  assign new_new_n50504__ = ~ys__n45777 & ~ys__n46078;
  assign new_new_n50505__ = ~ys__n46118 & ~new_new_n50504__;
  assign new_new_n50506__ = ~new_new_n50503__ & new_new_n50505__;
  assign new_new_n50507__ = ys__n45780 & ys__n46080;
  assign new_new_n50508__ = ~ys__n45780 & ~ys__n46080;
  assign new_new_n50509__ = ~ys__n46119 & ~new_new_n50508__;
  assign new_new_n50510__ = ~new_new_n50507__ & new_new_n50509__;
  assign new_new_n50511__ = ~new_new_n50506__ & ~new_new_n50510__;
  assign new_new_n50512__ = new_new_n50502__ & new_new_n50511__;
  assign new_new_n50513__ = ys__n45759 & ys__n46066;
  assign new_new_n50514__ = ~ys__n45759 & ~ys__n46066;
  assign new_new_n50515__ = ~ys__n46112 & ~new_new_n50514__;
  assign new_new_n50516__ = ~new_new_n50513__ & new_new_n50515__;
  assign new_new_n50517__ = ys__n45762 & ys__n46068;
  assign new_new_n50518__ = ~ys__n45762 & ~ys__n46068;
  assign new_new_n50519__ = ~ys__n46113 & ~new_new_n50518__;
  assign new_new_n50520__ = ~new_new_n50517__ & new_new_n50519__;
  assign new_new_n50521__ = ~new_new_n50516__ & ~new_new_n50520__;
  assign new_new_n50522__ = ys__n45765 & ys__n46070;
  assign new_new_n50523__ = ~ys__n45765 & ~ys__n46070;
  assign new_new_n50524__ = ~ys__n46114 & ~new_new_n50523__;
  assign new_new_n50525__ = ~new_new_n50522__ & new_new_n50524__;
  assign new_new_n50526__ = ys__n45768 & ys__n46072;
  assign new_new_n50527__ = ~ys__n45768 & ~ys__n46072;
  assign new_new_n50528__ = ~ys__n46115 & ~new_new_n50527__;
  assign new_new_n50529__ = ~new_new_n50526__ & new_new_n50528__;
  assign new_new_n50530__ = ~new_new_n50525__ & ~new_new_n50529__;
  assign new_new_n50531__ = new_new_n50521__ & new_new_n50530__;
  assign new_new_n50532__ = new_new_n50512__ & new_new_n50531__;
  assign new_new_n50533__ = ys__n45801 & ys__n46094;
  assign new_new_n50534__ = ~ys__n45801 & ~ys__n46094;
  assign new_new_n50535__ = ~ys__n46126 & ~new_new_n50534__;
  assign new_new_n50536__ = ~new_new_n50533__ & new_new_n50535__;
  assign new_new_n50537__ = ys__n45795 & ys__n46090;
  assign new_new_n50538__ = ~ys__n45795 & ~ys__n46090;
  assign new_new_n50539__ = ~ys__n46124 & ~new_new_n50538__;
  assign new_new_n50540__ = ~new_new_n50537__ & new_new_n50539__;
  assign new_new_n50541__ = ys__n45798 & ys__n46092;
  assign new_new_n50542__ = ~ys__n45798 & ~ys__n46092;
  assign new_new_n50543__ = ~ys__n46125 & ~new_new_n50542__;
  assign new_new_n50544__ = ~new_new_n50541__ & new_new_n50543__;
  assign new_new_n50545__ = ~new_new_n50540__ & ~new_new_n50544__;
  assign new_new_n50546__ = ~new_new_n50536__ & new_new_n50545__;
  assign new_new_n50547__ = ys__n45783 & ys__n46082;
  assign new_new_n50548__ = ~ys__n45783 & ~ys__n46082;
  assign new_new_n50549__ = ~ys__n46120 & ~new_new_n50548__;
  assign new_new_n50550__ = ~new_new_n50547__ & new_new_n50549__;
  assign new_new_n50551__ = ys__n45786 & ys__n46084;
  assign new_new_n50552__ = ~ys__n45786 & ~ys__n46084;
  assign new_new_n50553__ = ~ys__n46121 & ~new_new_n50552__;
  assign new_new_n50554__ = ~new_new_n50551__ & new_new_n50553__;
  assign new_new_n50555__ = ~new_new_n50550__ & ~new_new_n50554__;
  assign new_new_n50556__ = ys__n45789 & ys__n46086;
  assign new_new_n50557__ = ~ys__n45789 & ~ys__n46086;
  assign new_new_n50558__ = ~ys__n46122 & ~new_new_n50557__;
  assign new_new_n50559__ = ~new_new_n50556__ & new_new_n50558__;
  assign new_new_n50560__ = ys__n45792 & ys__n46088;
  assign new_new_n50561__ = ~ys__n45792 & ~ys__n46088;
  assign new_new_n50562__ = ~ys__n46123 & ~new_new_n50561__;
  assign new_new_n50563__ = ~new_new_n50560__ & new_new_n50562__;
  assign new_new_n50564__ = ~new_new_n50559__ & ~new_new_n50563__;
  assign new_new_n50565__ = new_new_n50555__ & new_new_n50564__;
  assign new_new_n50566__ = new_new_n50546__ & new_new_n50565__;
  assign new_new_n50567__ = new_new_n50532__ & new_new_n50566__;
  assign new_new_n50568__ = ys__n45723 & ys__n46042;
  assign new_new_n50569__ = ~ys__n45723 & ~ys__n46042;
  assign new_new_n50570__ = ~ys__n46100 & ~new_new_n50569__;
  assign new_new_n50571__ = ~new_new_n50568__ & new_new_n50570__;
  assign new_new_n50572__ = ys__n45726 & ys__n46044;
  assign new_new_n50573__ = ~ys__n45726 & ~ys__n46044;
  assign new_new_n50574__ = ~ys__n46101 & ~new_new_n50573__;
  assign new_new_n50575__ = ~new_new_n50572__ & new_new_n50574__;
  assign new_new_n50576__ = ~new_new_n50571__ & ~new_new_n50575__;
  assign new_new_n50577__ = ys__n45729 & ys__n46046;
  assign new_new_n50578__ = ~ys__n45729 & ~ys__n46046;
  assign new_new_n50579__ = ~ys__n46102 & ~new_new_n50578__;
  assign new_new_n50580__ = ~new_new_n50577__ & new_new_n50579__;
  assign new_new_n50581__ = ys__n45732 & ys__n46048;
  assign new_new_n50582__ = ~ys__n45732 & ~ys__n46048;
  assign new_new_n50583__ = ~ys__n46103 & ~new_new_n50582__;
  assign new_new_n50584__ = ~new_new_n50581__ & new_new_n50583__;
  assign new_new_n50585__ = ~new_new_n50580__ & ~new_new_n50584__;
  assign new_new_n50586__ = new_new_n50576__ & new_new_n50585__;
  assign new_new_n50587__ = ys__n45711 & ys__n46034;
  assign new_new_n50588__ = ~ys__n45711 & ~ys__n46034;
  assign new_new_n50589__ = ~ys__n46096 & ~new_new_n50588__;
  assign new_new_n50590__ = ~new_new_n50587__ & new_new_n50589__;
  assign new_new_n50591__ = ys__n45714 & ys__n46036;
  assign new_new_n50592__ = ~ys__n45714 & ~ys__n46036;
  assign new_new_n50593__ = ~ys__n46097 & ~new_new_n50592__;
  assign new_new_n50594__ = ~new_new_n50591__ & new_new_n50593__;
  assign new_new_n50595__ = ~new_new_n50590__ & ~new_new_n50594__;
  assign new_new_n50596__ = ys__n45717 & ys__n46038;
  assign new_new_n50597__ = ~ys__n45717 & ~ys__n46038;
  assign new_new_n50598__ = ~ys__n46098 & ~new_new_n50597__;
  assign new_new_n50599__ = ~new_new_n50596__ & new_new_n50598__;
  assign new_new_n50600__ = ys__n45720 & ys__n46040;
  assign new_new_n50601__ = ~ys__n45720 & ~ys__n46040;
  assign new_new_n50602__ = ~ys__n46099 & ~new_new_n50601__;
  assign new_new_n50603__ = ~new_new_n50600__ & new_new_n50602__;
  assign new_new_n50604__ = ~new_new_n50599__ & ~new_new_n50603__;
  assign new_new_n50605__ = new_new_n50595__ & new_new_n50604__;
  assign new_new_n50606__ = new_new_n50586__ & new_new_n50605__;
  assign new_new_n50607__ = ys__n45747 & ys__n46058;
  assign new_new_n50608__ = ~ys__n45747 & ~ys__n46058;
  assign new_new_n50609__ = ~ys__n46108 & ~new_new_n50608__;
  assign new_new_n50610__ = ~new_new_n50607__ & new_new_n50609__;
  assign new_new_n50611__ = ys__n45750 & ys__n46060;
  assign new_new_n50612__ = ~ys__n45750 & ~ys__n46060;
  assign new_new_n50613__ = ~ys__n46109 & ~new_new_n50612__;
  assign new_new_n50614__ = ~new_new_n50611__ & new_new_n50613__;
  assign new_new_n50615__ = ~new_new_n50610__ & ~new_new_n50614__;
  assign new_new_n50616__ = ys__n45753 & ys__n46062;
  assign new_new_n50617__ = ~ys__n45753 & ~ys__n46062;
  assign new_new_n50618__ = ~ys__n46110 & ~new_new_n50617__;
  assign new_new_n50619__ = ~new_new_n50616__ & new_new_n50618__;
  assign new_new_n50620__ = ys__n45756 & ys__n46064;
  assign new_new_n50621__ = ~ys__n45756 & ~ys__n46064;
  assign new_new_n50622__ = ~ys__n46111 & ~new_new_n50621__;
  assign new_new_n50623__ = ~new_new_n50620__ & new_new_n50622__;
  assign new_new_n50624__ = ~new_new_n50619__ & ~new_new_n50623__;
  assign new_new_n50625__ = new_new_n50615__ & new_new_n50624__;
  assign new_new_n50626__ = ys__n45735 & ys__n46050;
  assign new_new_n50627__ = ~ys__n45735 & ~ys__n46050;
  assign new_new_n50628__ = ~ys__n46104 & ~new_new_n50627__;
  assign new_new_n50629__ = ~new_new_n50626__ & new_new_n50628__;
  assign new_new_n50630__ = ys__n45738 & ys__n46052;
  assign new_new_n50631__ = ~ys__n45738 & ~ys__n46052;
  assign new_new_n50632__ = ~ys__n46105 & ~new_new_n50631__;
  assign new_new_n50633__ = ~new_new_n50630__ & new_new_n50632__;
  assign new_new_n50634__ = ~new_new_n50629__ & ~new_new_n50633__;
  assign new_new_n50635__ = ys__n45741 & ys__n46054;
  assign new_new_n50636__ = ~ys__n45741 & ~ys__n46054;
  assign new_new_n50637__ = ~ys__n46106 & ~new_new_n50636__;
  assign new_new_n50638__ = ~new_new_n50635__ & new_new_n50637__;
  assign new_new_n50639__ = ys__n45744 & ys__n46056;
  assign new_new_n50640__ = ~ys__n45744 & ~ys__n46056;
  assign new_new_n50641__ = ~ys__n46107 & ~new_new_n50640__;
  assign new_new_n50642__ = ~new_new_n50639__ & new_new_n50641__;
  assign new_new_n50643__ = ~new_new_n50638__ & ~new_new_n50642__;
  assign new_new_n50644__ = new_new_n50634__ & new_new_n50643__;
  assign new_new_n50645__ = new_new_n50625__ & new_new_n50644__;
  assign new_new_n50646__ = new_new_n50606__ & new_new_n50645__;
  assign new_new_n50647__ = new_new_n50567__ & new_new_n50646__;
  assign new_new_n50648__ = ys__n46128 & new_new_n50647__;
  assign new_new_n50649__ = ys__n45771 & ys__n45976;
  assign new_new_n50650__ = ~ys__n45771 & ~ys__n45976;
  assign new_new_n50651__ = ~ys__n46018 & ~new_new_n50650__;
  assign new_new_n50652__ = ~new_new_n50649__ & new_new_n50651__;
  assign new_new_n50653__ = ys__n45774 & ys__n45978;
  assign new_new_n50654__ = ~ys__n45774 & ~ys__n45978;
  assign new_new_n50655__ = ~ys__n46019 & ~new_new_n50654__;
  assign new_new_n50656__ = ~new_new_n50653__ & new_new_n50655__;
  assign new_new_n50657__ = ~new_new_n50652__ & ~new_new_n50656__;
  assign new_new_n50658__ = ys__n45777 & ys__n45980;
  assign new_new_n50659__ = ~ys__n45777 & ~ys__n45980;
  assign new_new_n50660__ = ~ys__n46020 & ~new_new_n50659__;
  assign new_new_n50661__ = ~new_new_n50658__ & new_new_n50660__;
  assign new_new_n50662__ = ys__n45780 & ys__n45982;
  assign new_new_n50663__ = ~ys__n45780 & ~ys__n45982;
  assign new_new_n50664__ = ~ys__n46021 & ~new_new_n50663__;
  assign new_new_n50665__ = ~new_new_n50662__ & new_new_n50664__;
  assign new_new_n50666__ = ~new_new_n50661__ & ~new_new_n50665__;
  assign new_new_n50667__ = new_new_n50657__ & new_new_n50666__;
  assign new_new_n50668__ = ys__n45759 & ys__n45968;
  assign new_new_n50669__ = ~ys__n45759 & ~ys__n45968;
  assign new_new_n50670__ = ~ys__n46014 & ~new_new_n50669__;
  assign new_new_n50671__ = ~new_new_n50668__ & new_new_n50670__;
  assign new_new_n50672__ = ys__n45762 & ys__n45970;
  assign new_new_n50673__ = ~ys__n45762 & ~ys__n45970;
  assign new_new_n50674__ = ~ys__n46015 & ~new_new_n50673__;
  assign new_new_n50675__ = ~new_new_n50672__ & new_new_n50674__;
  assign new_new_n50676__ = ~new_new_n50671__ & ~new_new_n50675__;
  assign new_new_n50677__ = ys__n45765 & ys__n45972;
  assign new_new_n50678__ = ~ys__n45765 & ~ys__n45972;
  assign new_new_n50679__ = ~ys__n46016 & ~new_new_n50678__;
  assign new_new_n50680__ = ~new_new_n50677__ & new_new_n50679__;
  assign new_new_n50681__ = ys__n45768 & ys__n45974;
  assign new_new_n50682__ = ~ys__n45768 & ~ys__n45974;
  assign new_new_n50683__ = ~ys__n46017 & ~new_new_n50682__;
  assign new_new_n50684__ = ~new_new_n50681__ & new_new_n50683__;
  assign new_new_n50685__ = ~new_new_n50680__ & ~new_new_n50684__;
  assign new_new_n50686__ = new_new_n50676__ & new_new_n50685__;
  assign new_new_n50687__ = new_new_n50667__ & new_new_n50686__;
  assign new_new_n50688__ = ys__n45801 & ys__n45996;
  assign new_new_n50689__ = ~ys__n45801 & ~ys__n45996;
  assign new_new_n50690__ = ~ys__n46028 & ~new_new_n50689__;
  assign new_new_n50691__ = ~new_new_n50688__ & new_new_n50690__;
  assign new_new_n50692__ = ys__n45795 & ys__n45992;
  assign new_new_n50693__ = ~ys__n45795 & ~ys__n45992;
  assign new_new_n50694__ = ~ys__n46026 & ~new_new_n50693__;
  assign new_new_n50695__ = ~new_new_n50692__ & new_new_n50694__;
  assign new_new_n50696__ = ys__n45798 & ys__n45994;
  assign new_new_n50697__ = ~ys__n45798 & ~ys__n45994;
  assign new_new_n50698__ = ~ys__n46027 & ~new_new_n50697__;
  assign new_new_n50699__ = ~new_new_n50696__ & new_new_n50698__;
  assign new_new_n50700__ = ~new_new_n50695__ & ~new_new_n50699__;
  assign new_new_n50701__ = ~new_new_n50691__ & new_new_n50700__;
  assign new_new_n50702__ = ys__n45783 & ys__n45984;
  assign new_new_n50703__ = ~ys__n45783 & ~ys__n45984;
  assign new_new_n50704__ = ~ys__n46022 & ~new_new_n50703__;
  assign new_new_n50705__ = ~new_new_n50702__ & new_new_n50704__;
  assign new_new_n50706__ = ys__n45786 & ys__n45986;
  assign new_new_n50707__ = ~ys__n45786 & ~ys__n45986;
  assign new_new_n50708__ = ~ys__n46023 & ~new_new_n50707__;
  assign new_new_n50709__ = ~new_new_n50706__ & new_new_n50708__;
  assign new_new_n50710__ = ~new_new_n50705__ & ~new_new_n50709__;
  assign new_new_n50711__ = ys__n45789 & ys__n45988;
  assign new_new_n50712__ = ~ys__n45789 & ~ys__n45988;
  assign new_new_n50713__ = ~ys__n46024 & ~new_new_n50712__;
  assign new_new_n50714__ = ~new_new_n50711__ & new_new_n50713__;
  assign new_new_n50715__ = ys__n45792 & ys__n45990;
  assign new_new_n50716__ = ~ys__n45792 & ~ys__n45990;
  assign new_new_n50717__ = ~ys__n46025 & ~new_new_n50716__;
  assign new_new_n50718__ = ~new_new_n50715__ & new_new_n50717__;
  assign new_new_n50719__ = ~new_new_n50714__ & ~new_new_n50718__;
  assign new_new_n50720__ = new_new_n50710__ & new_new_n50719__;
  assign new_new_n50721__ = new_new_n50701__ & new_new_n50720__;
  assign new_new_n50722__ = new_new_n50687__ & new_new_n50721__;
  assign new_new_n50723__ = ys__n45723 & ys__n45944;
  assign new_new_n50724__ = ~ys__n45723 & ~ys__n45944;
  assign new_new_n50725__ = ~ys__n46002 & ~new_new_n50724__;
  assign new_new_n50726__ = ~new_new_n50723__ & new_new_n50725__;
  assign new_new_n50727__ = ys__n45726 & ys__n45946;
  assign new_new_n50728__ = ~ys__n45726 & ~ys__n45946;
  assign new_new_n50729__ = ~ys__n46003 & ~new_new_n50728__;
  assign new_new_n50730__ = ~new_new_n50727__ & new_new_n50729__;
  assign new_new_n50731__ = ~new_new_n50726__ & ~new_new_n50730__;
  assign new_new_n50732__ = ys__n45729 & ys__n45948;
  assign new_new_n50733__ = ~ys__n45729 & ~ys__n45948;
  assign new_new_n50734__ = ~ys__n46004 & ~new_new_n50733__;
  assign new_new_n50735__ = ~new_new_n50732__ & new_new_n50734__;
  assign new_new_n50736__ = ys__n45732 & ys__n45950;
  assign new_new_n50737__ = ~ys__n45732 & ~ys__n45950;
  assign new_new_n50738__ = ~ys__n46005 & ~new_new_n50737__;
  assign new_new_n50739__ = ~new_new_n50736__ & new_new_n50738__;
  assign new_new_n50740__ = ~new_new_n50735__ & ~new_new_n50739__;
  assign new_new_n50741__ = new_new_n50731__ & new_new_n50740__;
  assign new_new_n50742__ = ys__n45711 & ys__n45936;
  assign new_new_n50743__ = ~ys__n45711 & ~ys__n45936;
  assign new_new_n50744__ = ~ys__n45998 & ~new_new_n50743__;
  assign new_new_n50745__ = ~new_new_n50742__ & new_new_n50744__;
  assign new_new_n50746__ = ys__n45714 & ys__n45938;
  assign new_new_n50747__ = ~ys__n45714 & ~ys__n45938;
  assign new_new_n50748__ = ~ys__n45999 & ~new_new_n50747__;
  assign new_new_n50749__ = ~new_new_n50746__ & new_new_n50748__;
  assign new_new_n50750__ = ~new_new_n50745__ & ~new_new_n50749__;
  assign new_new_n50751__ = ys__n45717 & ys__n45940;
  assign new_new_n50752__ = ~ys__n45717 & ~ys__n45940;
  assign new_new_n50753__ = ~ys__n46000 & ~new_new_n50752__;
  assign new_new_n50754__ = ~new_new_n50751__ & new_new_n50753__;
  assign new_new_n50755__ = ys__n45720 & ys__n45942;
  assign new_new_n50756__ = ~ys__n45720 & ~ys__n45942;
  assign new_new_n50757__ = ~ys__n46001 & ~new_new_n50756__;
  assign new_new_n50758__ = ~new_new_n50755__ & new_new_n50757__;
  assign new_new_n50759__ = ~new_new_n50754__ & ~new_new_n50758__;
  assign new_new_n50760__ = new_new_n50750__ & new_new_n50759__;
  assign new_new_n50761__ = new_new_n50741__ & new_new_n50760__;
  assign new_new_n50762__ = ys__n45747 & ys__n45960;
  assign new_new_n50763__ = ~ys__n45747 & ~ys__n45960;
  assign new_new_n50764__ = ~ys__n46010 & ~new_new_n50763__;
  assign new_new_n50765__ = ~new_new_n50762__ & new_new_n50764__;
  assign new_new_n50766__ = ys__n45750 & ys__n45962;
  assign new_new_n50767__ = ~ys__n45750 & ~ys__n45962;
  assign new_new_n50768__ = ~ys__n46011 & ~new_new_n50767__;
  assign new_new_n50769__ = ~new_new_n50766__ & new_new_n50768__;
  assign new_new_n50770__ = ~new_new_n50765__ & ~new_new_n50769__;
  assign new_new_n50771__ = ys__n45753 & ys__n45964;
  assign new_new_n50772__ = ~ys__n45753 & ~ys__n45964;
  assign new_new_n50773__ = ~ys__n46012 & ~new_new_n50772__;
  assign new_new_n50774__ = ~new_new_n50771__ & new_new_n50773__;
  assign new_new_n50775__ = ys__n45756 & ys__n45966;
  assign new_new_n50776__ = ~ys__n45756 & ~ys__n45966;
  assign new_new_n50777__ = ~ys__n46013 & ~new_new_n50776__;
  assign new_new_n50778__ = ~new_new_n50775__ & new_new_n50777__;
  assign new_new_n50779__ = ~new_new_n50774__ & ~new_new_n50778__;
  assign new_new_n50780__ = new_new_n50770__ & new_new_n50779__;
  assign new_new_n50781__ = ys__n45735 & ys__n45952;
  assign new_new_n50782__ = ~ys__n45735 & ~ys__n45952;
  assign new_new_n50783__ = ~ys__n46006 & ~new_new_n50782__;
  assign new_new_n50784__ = ~new_new_n50781__ & new_new_n50783__;
  assign new_new_n50785__ = ys__n45738 & ys__n45954;
  assign new_new_n50786__ = ~ys__n45738 & ~ys__n45954;
  assign new_new_n50787__ = ~ys__n46007 & ~new_new_n50786__;
  assign new_new_n50788__ = ~new_new_n50785__ & new_new_n50787__;
  assign new_new_n50789__ = ~new_new_n50784__ & ~new_new_n50788__;
  assign new_new_n50790__ = ys__n45741 & ys__n45956;
  assign new_new_n50791__ = ~ys__n45741 & ~ys__n45956;
  assign new_new_n50792__ = ~ys__n46008 & ~new_new_n50791__;
  assign new_new_n50793__ = ~new_new_n50790__ & new_new_n50792__;
  assign new_new_n50794__ = ys__n45744 & ys__n45958;
  assign new_new_n50795__ = ~ys__n45744 & ~ys__n45958;
  assign new_new_n50796__ = ~ys__n46009 & ~new_new_n50795__;
  assign new_new_n50797__ = ~new_new_n50794__ & new_new_n50796__;
  assign new_new_n50798__ = ~new_new_n50793__ & ~new_new_n50797__;
  assign new_new_n50799__ = new_new_n50789__ & new_new_n50798__;
  assign new_new_n50800__ = new_new_n50780__ & new_new_n50799__;
  assign new_new_n50801__ = new_new_n50761__ & new_new_n50800__;
  assign new_new_n50802__ = new_new_n50722__ & new_new_n50801__;
  assign new_new_n50803__ = ys__n46031 & new_new_n50802__;
  assign new_new_n50804__ = ~new_new_n50648__ & ~new_new_n50803__;
  assign new_new_n50805__ = ys__n45771 & ys__n45878;
  assign new_new_n50806__ = ~ys__n45771 & ~ys__n45878;
  assign new_new_n50807__ = ~ys__n45920 & ~new_new_n50806__;
  assign new_new_n50808__ = ~new_new_n50805__ & new_new_n50807__;
  assign new_new_n50809__ = ys__n45774 & ys__n45880;
  assign new_new_n50810__ = ~ys__n45774 & ~ys__n45880;
  assign new_new_n50811__ = ~ys__n45921 & ~new_new_n50810__;
  assign new_new_n50812__ = ~new_new_n50809__ & new_new_n50811__;
  assign new_new_n50813__ = ~new_new_n50808__ & ~new_new_n50812__;
  assign new_new_n50814__ = ys__n45777 & ys__n45882;
  assign new_new_n50815__ = ~ys__n45777 & ~ys__n45882;
  assign new_new_n50816__ = ~ys__n45922 & ~new_new_n50815__;
  assign new_new_n50817__ = ~new_new_n50814__ & new_new_n50816__;
  assign new_new_n50818__ = ys__n45780 & ys__n45884;
  assign new_new_n50819__ = ~ys__n45780 & ~ys__n45884;
  assign new_new_n50820__ = ~ys__n45923 & ~new_new_n50819__;
  assign new_new_n50821__ = ~new_new_n50818__ & new_new_n50820__;
  assign new_new_n50822__ = ~new_new_n50817__ & ~new_new_n50821__;
  assign new_new_n50823__ = new_new_n50813__ & new_new_n50822__;
  assign new_new_n50824__ = ys__n45759 & ys__n45870;
  assign new_new_n50825__ = ~ys__n45759 & ~ys__n45870;
  assign new_new_n50826__ = ~ys__n45916 & ~new_new_n50825__;
  assign new_new_n50827__ = ~new_new_n50824__ & new_new_n50826__;
  assign new_new_n50828__ = ys__n45762 & ys__n45872;
  assign new_new_n50829__ = ~ys__n45762 & ~ys__n45872;
  assign new_new_n50830__ = ~ys__n45917 & ~new_new_n50829__;
  assign new_new_n50831__ = ~new_new_n50828__ & new_new_n50830__;
  assign new_new_n50832__ = ~new_new_n50827__ & ~new_new_n50831__;
  assign new_new_n50833__ = ys__n45765 & ys__n45874;
  assign new_new_n50834__ = ~ys__n45765 & ~ys__n45874;
  assign new_new_n50835__ = ~ys__n45918 & ~new_new_n50834__;
  assign new_new_n50836__ = ~new_new_n50833__ & new_new_n50835__;
  assign new_new_n50837__ = ys__n45768 & ys__n45876;
  assign new_new_n50838__ = ~ys__n45768 & ~ys__n45876;
  assign new_new_n50839__ = ~ys__n45919 & ~new_new_n50838__;
  assign new_new_n50840__ = ~new_new_n50837__ & new_new_n50839__;
  assign new_new_n50841__ = ~new_new_n50836__ & ~new_new_n50840__;
  assign new_new_n50842__ = new_new_n50832__ & new_new_n50841__;
  assign new_new_n50843__ = new_new_n50823__ & new_new_n50842__;
  assign new_new_n50844__ = ys__n45801 & ys__n45898;
  assign new_new_n50845__ = ~ys__n45801 & ~ys__n45898;
  assign new_new_n50846__ = ~ys__n45930 & ~new_new_n50845__;
  assign new_new_n50847__ = ~new_new_n50844__ & new_new_n50846__;
  assign new_new_n50848__ = ys__n45795 & ys__n45894;
  assign new_new_n50849__ = ~ys__n45795 & ~ys__n45894;
  assign new_new_n50850__ = ~ys__n45928 & ~new_new_n50849__;
  assign new_new_n50851__ = ~new_new_n50848__ & new_new_n50850__;
  assign new_new_n50852__ = ys__n45798 & ys__n45896;
  assign new_new_n50853__ = ~ys__n45798 & ~ys__n45896;
  assign new_new_n50854__ = ~ys__n45929 & ~new_new_n50853__;
  assign new_new_n50855__ = ~new_new_n50852__ & new_new_n50854__;
  assign new_new_n50856__ = ~new_new_n50851__ & ~new_new_n50855__;
  assign new_new_n50857__ = ~new_new_n50847__ & new_new_n50856__;
  assign new_new_n50858__ = ys__n45783 & ys__n45886;
  assign new_new_n50859__ = ~ys__n45783 & ~ys__n45886;
  assign new_new_n50860__ = ~ys__n45924 & ~new_new_n50859__;
  assign new_new_n50861__ = ~new_new_n50858__ & new_new_n50860__;
  assign new_new_n50862__ = ys__n45786 & ys__n45888;
  assign new_new_n50863__ = ~ys__n45786 & ~ys__n45888;
  assign new_new_n50864__ = ~ys__n45925 & ~new_new_n50863__;
  assign new_new_n50865__ = ~new_new_n50862__ & new_new_n50864__;
  assign new_new_n50866__ = ~new_new_n50861__ & ~new_new_n50865__;
  assign new_new_n50867__ = ys__n45789 & ys__n45890;
  assign new_new_n50868__ = ~ys__n45789 & ~ys__n45890;
  assign new_new_n50869__ = ~ys__n45926 & ~new_new_n50868__;
  assign new_new_n50870__ = ~new_new_n50867__ & new_new_n50869__;
  assign new_new_n50871__ = ys__n45792 & ys__n45892;
  assign new_new_n50872__ = ~ys__n45792 & ~ys__n45892;
  assign new_new_n50873__ = ~ys__n45927 & ~new_new_n50872__;
  assign new_new_n50874__ = ~new_new_n50871__ & new_new_n50873__;
  assign new_new_n50875__ = ~new_new_n50870__ & ~new_new_n50874__;
  assign new_new_n50876__ = new_new_n50866__ & new_new_n50875__;
  assign new_new_n50877__ = new_new_n50857__ & new_new_n50876__;
  assign new_new_n50878__ = new_new_n50843__ & new_new_n50877__;
  assign new_new_n50879__ = ys__n45723 & ys__n45846;
  assign new_new_n50880__ = ~ys__n45723 & ~ys__n45846;
  assign new_new_n50881__ = ~ys__n45904 & ~new_new_n50880__;
  assign new_new_n50882__ = ~new_new_n50879__ & new_new_n50881__;
  assign new_new_n50883__ = ys__n45726 & ys__n45848;
  assign new_new_n50884__ = ~ys__n45726 & ~ys__n45848;
  assign new_new_n50885__ = ~ys__n45905 & ~new_new_n50884__;
  assign new_new_n50886__ = ~new_new_n50883__ & new_new_n50885__;
  assign new_new_n50887__ = ~new_new_n50882__ & ~new_new_n50886__;
  assign new_new_n50888__ = ys__n45729 & ys__n45850;
  assign new_new_n50889__ = ~ys__n45729 & ~ys__n45850;
  assign new_new_n50890__ = ~ys__n45906 & ~new_new_n50889__;
  assign new_new_n50891__ = ~new_new_n50888__ & new_new_n50890__;
  assign new_new_n50892__ = ys__n45732 & ys__n45852;
  assign new_new_n50893__ = ~ys__n45732 & ~ys__n45852;
  assign new_new_n50894__ = ~ys__n45907 & ~new_new_n50893__;
  assign new_new_n50895__ = ~new_new_n50892__ & new_new_n50894__;
  assign new_new_n50896__ = ~new_new_n50891__ & ~new_new_n50895__;
  assign new_new_n50897__ = new_new_n50887__ & new_new_n50896__;
  assign new_new_n50898__ = ys__n45711 & ys__n45838;
  assign new_new_n50899__ = ~ys__n45711 & ~ys__n45838;
  assign new_new_n50900__ = ~ys__n45900 & ~new_new_n50899__;
  assign new_new_n50901__ = ~new_new_n50898__ & new_new_n50900__;
  assign new_new_n50902__ = ys__n45714 & ys__n45840;
  assign new_new_n50903__ = ~ys__n45714 & ~ys__n45840;
  assign new_new_n50904__ = ~ys__n45901 & ~new_new_n50903__;
  assign new_new_n50905__ = ~new_new_n50902__ & new_new_n50904__;
  assign new_new_n50906__ = ~new_new_n50901__ & ~new_new_n50905__;
  assign new_new_n50907__ = ys__n45717 & ys__n45842;
  assign new_new_n50908__ = ~ys__n45717 & ~ys__n45842;
  assign new_new_n50909__ = ~ys__n45902 & ~new_new_n50908__;
  assign new_new_n50910__ = ~new_new_n50907__ & new_new_n50909__;
  assign new_new_n50911__ = ys__n45720 & ys__n45844;
  assign new_new_n50912__ = ~ys__n45720 & ~ys__n45844;
  assign new_new_n50913__ = ~ys__n45903 & ~new_new_n50912__;
  assign new_new_n50914__ = ~new_new_n50911__ & new_new_n50913__;
  assign new_new_n50915__ = ~new_new_n50910__ & ~new_new_n50914__;
  assign new_new_n50916__ = new_new_n50906__ & new_new_n50915__;
  assign new_new_n50917__ = new_new_n50897__ & new_new_n50916__;
  assign new_new_n50918__ = ys__n45747 & ys__n45862;
  assign new_new_n50919__ = ~ys__n45747 & ~ys__n45862;
  assign new_new_n50920__ = ~ys__n45912 & ~new_new_n50919__;
  assign new_new_n50921__ = ~new_new_n50918__ & new_new_n50920__;
  assign new_new_n50922__ = ys__n45750 & ys__n45864;
  assign new_new_n50923__ = ~ys__n45750 & ~ys__n45864;
  assign new_new_n50924__ = ~ys__n45913 & ~new_new_n50923__;
  assign new_new_n50925__ = ~new_new_n50922__ & new_new_n50924__;
  assign new_new_n50926__ = ~new_new_n50921__ & ~new_new_n50925__;
  assign new_new_n50927__ = ys__n45753 & ys__n45866;
  assign new_new_n50928__ = ~ys__n45753 & ~ys__n45866;
  assign new_new_n50929__ = ~ys__n45914 & ~new_new_n50928__;
  assign new_new_n50930__ = ~new_new_n50927__ & new_new_n50929__;
  assign new_new_n50931__ = ys__n45756 & ys__n45868;
  assign new_new_n50932__ = ~ys__n45756 & ~ys__n45868;
  assign new_new_n50933__ = ~ys__n45915 & ~new_new_n50932__;
  assign new_new_n50934__ = ~new_new_n50931__ & new_new_n50933__;
  assign new_new_n50935__ = ~new_new_n50930__ & ~new_new_n50934__;
  assign new_new_n50936__ = new_new_n50926__ & new_new_n50935__;
  assign new_new_n50937__ = ys__n45735 & ys__n45854;
  assign new_new_n50938__ = ~ys__n45735 & ~ys__n45854;
  assign new_new_n50939__ = ~ys__n45908 & ~new_new_n50938__;
  assign new_new_n50940__ = ~new_new_n50937__ & new_new_n50939__;
  assign new_new_n50941__ = ys__n45738 & ys__n45856;
  assign new_new_n50942__ = ~ys__n45738 & ~ys__n45856;
  assign new_new_n50943__ = ~ys__n45909 & ~new_new_n50942__;
  assign new_new_n50944__ = ~new_new_n50941__ & new_new_n50943__;
  assign new_new_n50945__ = ~new_new_n50940__ & ~new_new_n50944__;
  assign new_new_n50946__ = ys__n45741 & ys__n45858;
  assign new_new_n50947__ = ~ys__n45741 & ~ys__n45858;
  assign new_new_n50948__ = ~ys__n45910 & ~new_new_n50947__;
  assign new_new_n50949__ = ~new_new_n50946__ & new_new_n50948__;
  assign new_new_n50950__ = ys__n45744 & ys__n45860;
  assign new_new_n50951__ = ~ys__n45744 & ~ys__n45860;
  assign new_new_n50952__ = ~ys__n45911 & ~new_new_n50951__;
  assign new_new_n50953__ = ~new_new_n50950__ & new_new_n50952__;
  assign new_new_n50954__ = ~new_new_n50949__ & ~new_new_n50953__;
  assign new_new_n50955__ = new_new_n50945__ & new_new_n50954__;
  assign new_new_n50956__ = new_new_n50936__ & new_new_n50955__;
  assign new_new_n50957__ = new_new_n50917__ & new_new_n50956__;
  assign new_new_n50958__ = new_new_n50878__ & new_new_n50957__;
  assign new_new_n50959__ = ys__n45933 & new_new_n50958__;
  assign new_new_n50960__ = ys__n45771 & ys__n45772;
  assign new_new_n50961__ = ~ys__n45771 & ~ys__n45772;
  assign new_new_n50962__ = ~ys__n45824 & ~new_new_n50961__;
  assign new_new_n50963__ = ~new_new_n50960__ & new_new_n50962__;
  assign new_new_n50964__ = ys__n45774 & ys__n45775;
  assign new_new_n50965__ = ~ys__n45774 & ~ys__n45775;
  assign new_new_n50966__ = ~ys__n45825 & ~new_new_n50965__;
  assign new_new_n50967__ = ~new_new_n50964__ & new_new_n50966__;
  assign new_new_n50968__ = ~new_new_n50963__ & ~new_new_n50967__;
  assign new_new_n50969__ = ys__n45777 & ys__n45778;
  assign new_new_n50970__ = ~ys__n45777 & ~ys__n45778;
  assign new_new_n50971__ = ~ys__n45826 & ~new_new_n50970__;
  assign new_new_n50972__ = ~new_new_n50969__ & new_new_n50971__;
  assign new_new_n50973__ = ys__n45780 & ys__n45781;
  assign new_new_n50974__ = ~ys__n45780 & ~ys__n45781;
  assign new_new_n50975__ = ~ys__n45827 & ~new_new_n50974__;
  assign new_new_n50976__ = ~new_new_n50973__ & new_new_n50975__;
  assign new_new_n50977__ = ~new_new_n50972__ & ~new_new_n50976__;
  assign new_new_n50978__ = new_new_n50968__ & new_new_n50977__;
  assign new_new_n50979__ = ys__n45759 & ys__n45760;
  assign new_new_n50980__ = ~ys__n45759 & ~ys__n45760;
  assign new_new_n50981__ = ~ys__n45820 & ~new_new_n50980__;
  assign new_new_n50982__ = ~new_new_n50979__ & new_new_n50981__;
  assign new_new_n50983__ = ys__n45762 & ys__n45763;
  assign new_new_n50984__ = ~ys__n45762 & ~ys__n45763;
  assign new_new_n50985__ = ~ys__n45821 & ~new_new_n50984__;
  assign new_new_n50986__ = ~new_new_n50983__ & new_new_n50985__;
  assign new_new_n50987__ = ~new_new_n50982__ & ~new_new_n50986__;
  assign new_new_n50988__ = ys__n45765 & ys__n45766;
  assign new_new_n50989__ = ~ys__n45765 & ~ys__n45766;
  assign new_new_n50990__ = ~ys__n45822 & ~new_new_n50989__;
  assign new_new_n50991__ = ~new_new_n50988__ & new_new_n50990__;
  assign new_new_n50992__ = ys__n45768 & ys__n45769;
  assign new_new_n50993__ = ~ys__n45768 & ~ys__n45769;
  assign new_new_n50994__ = ~ys__n45823 & ~new_new_n50993__;
  assign new_new_n50995__ = ~new_new_n50992__ & new_new_n50994__;
  assign new_new_n50996__ = ~new_new_n50991__ & ~new_new_n50995__;
  assign new_new_n50997__ = new_new_n50987__ & new_new_n50996__;
  assign new_new_n50998__ = new_new_n50978__ & new_new_n50997__;
  assign new_new_n50999__ = ys__n45801 & ys__n45802;
  assign new_new_n51000__ = ~ys__n45801 & ~ys__n45802;
  assign new_new_n51001__ = ~ys__n45834 & ~new_new_n51000__;
  assign new_new_n51002__ = ~new_new_n50999__ & new_new_n51001__;
  assign new_new_n51003__ = ys__n45795 & ys__n45796;
  assign new_new_n51004__ = ~ys__n45795 & ~ys__n45796;
  assign new_new_n51005__ = ~ys__n45832 & ~new_new_n51004__;
  assign new_new_n51006__ = ~new_new_n51003__ & new_new_n51005__;
  assign new_new_n51007__ = ys__n45798 & ys__n45799;
  assign new_new_n51008__ = ~ys__n45798 & ~ys__n45799;
  assign new_new_n51009__ = ~ys__n45833 & ~new_new_n51008__;
  assign new_new_n51010__ = ~new_new_n51007__ & new_new_n51009__;
  assign new_new_n51011__ = ~new_new_n51006__ & ~new_new_n51010__;
  assign new_new_n51012__ = ~new_new_n51002__ & new_new_n51011__;
  assign new_new_n51013__ = ys__n45783 & ys__n45784;
  assign new_new_n51014__ = ~ys__n45783 & ~ys__n45784;
  assign new_new_n51015__ = ~ys__n45828 & ~new_new_n51014__;
  assign new_new_n51016__ = ~new_new_n51013__ & new_new_n51015__;
  assign new_new_n51017__ = ys__n45786 & ys__n45787;
  assign new_new_n51018__ = ~ys__n45786 & ~ys__n45787;
  assign new_new_n51019__ = ~ys__n45829 & ~new_new_n51018__;
  assign new_new_n51020__ = ~new_new_n51017__ & new_new_n51019__;
  assign new_new_n51021__ = ~new_new_n51016__ & ~new_new_n51020__;
  assign new_new_n51022__ = ys__n45789 & ys__n45790;
  assign new_new_n51023__ = ~ys__n45789 & ~ys__n45790;
  assign new_new_n51024__ = ~ys__n45830 & ~new_new_n51023__;
  assign new_new_n51025__ = ~new_new_n51022__ & new_new_n51024__;
  assign new_new_n51026__ = ys__n45792 & ys__n45793;
  assign new_new_n51027__ = ~ys__n45792 & ~ys__n45793;
  assign new_new_n51028__ = ~ys__n45831 & ~new_new_n51027__;
  assign new_new_n51029__ = ~new_new_n51026__ & new_new_n51028__;
  assign new_new_n51030__ = ~new_new_n51025__ & ~new_new_n51029__;
  assign new_new_n51031__ = new_new_n51021__ & new_new_n51030__;
  assign new_new_n51032__ = new_new_n51012__ & new_new_n51031__;
  assign new_new_n51033__ = new_new_n50998__ & new_new_n51032__;
  assign new_new_n51034__ = ys__n45723 & ys__n45724;
  assign new_new_n51035__ = ~ys__n45723 & ~ys__n45724;
  assign new_new_n51036__ = ~ys__n45808 & ~new_new_n51035__;
  assign new_new_n51037__ = ~new_new_n51034__ & new_new_n51036__;
  assign new_new_n51038__ = ys__n45726 & ys__n45727;
  assign new_new_n51039__ = ~ys__n45726 & ~ys__n45727;
  assign new_new_n51040__ = ~ys__n45809 & ~new_new_n51039__;
  assign new_new_n51041__ = ~new_new_n51038__ & new_new_n51040__;
  assign new_new_n51042__ = ~new_new_n51037__ & ~new_new_n51041__;
  assign new_new_n51043__ = ys__n45729 & ys__n45730;
  assign new_new_n51044__ = ~ys__n45729 & ~ys__n45730;
  assign new_new_n51045__ = ~ys__n45810 & ~new_new_n51044__;
  assign new_new_n51046__ = ~new_new_n51043__ & new_new_n51045__;
  assign new_new_n51047__ = ys__n45732 & ys__n45733;
  assign new_new_n51048__ = ~ys__n45732 & ~ys__n45733;
  assign new_new_n51049__ = ~ys__n45811 & ~new_new_n51048__;
  assign new_new_n51050__ = ~new_new_n51047__ & new_new_n51049__;
  assign new_new_n51051__ = ~new_new_n51046__ & ~new_new_n51050__;
  assign new_new_n51052__ = new_new_n51042__ & new_new_n51051__;
  assign new_new_n51053__ = ys__n45711 & ys__n45712;
  assign new_new_n51054__ = ~ys__n45711 & ~ys__n45712;
  assign new_new_n51055__ = ~ys__n45804 & ~new_new_n51054__;
  assign new_new_n51056__ = ~new_new_n51053__ & new_new_n51055__;
  assign new_new_n51057__ = ys__n45714 & ys__n45715;
  assign new_new_n51058__ = ~ys__n45714 & ~ys__n45715;
  assign new_new_n51059__ = ~ys__n45805 & ~new_new_n51058__;
  assign new_new_n51060__ = ~new_new_n51057__ & new_new_n51059__;
  assign new_new_n51061__ = ~new_new_n51056__ & ~new_new_n51060__;
  assign new_new_n51062__ = ys__n45717 & ys__n45718;
  assign new_new_n51063__ = ~ys__n45717 & ~ys__n45718;
  assign new_new_n51064__ = ~ys__n45806 & ~new_new_n51063__;
  assign new_new_n51065__ = ~new_new_n51062__ & new_new_n51064__;
  assign new_new_n51066__ = ys__n45720 & ys__n45721;
  assign new_new_n51067__ = ~ys__n45720 & ~ys__n45721;
  assign new_new_n51068__ = ~ys__n45807 & ~new_new_n51067__;
  assign new_new_n51069__ = ~new_new_n51066__ & new_new_n51068__;
  assign new_new_n51070__ = ~new_new_n51065__ & ~new_new_n51069__;
  assign new_new_n51071__ = new_new_n51061__ & new_new_n51070__;
  assign new_new_n51072__ = new_new_n51052__ & new_new_n51071__;
  assign new_new_n51073__ = ys__n45747 & ys__n45748;
  assign new_new_n51074__ = ~ys__n45747 & ~ys__n45748;
  assign new_new_n51075__ = ~ys__n45816 & ~new_new_n51074__;
  assign new_new_n51076__ = ~new_new_n51073__ & new_new_n51075__;
  assign new_new_n51077__ = ys__n45750 & ys__n45751;
  assign new_new_n51078__ = ~ys__n45750 & ~ys__n45751;
  assign new_new_n51079__ = ~ys__n45817 & ~new_new_n51078__;
  assign new_new_n51080__ = ~new_new_n51077__ & new_new_n51079__;
  assign new_new_n51081__ = ~new_new_n51076__ & ~new_new_n51080__;
  assign new_new_n51082__ = ys__n45753 & ys__n45754;
  assign new_new_n51083__ = ~ys__n45753 & ~ys__n45754;
  assign new_new_n51084__ = ~ys__n45818 & ~new_new_n51083__;
  assign new_new_n51085__ = ~new_new_n51082__ & new_new_n51084__;
  assign new_new_n51086__ = ys__n45756 & ys__n45757;
  assign new_new_n51087__ = ~ys__n45756 & ~ys__n45757;
  assign new_new_n51088__ = ~ys__n45819 & ~new_new_n51087__;
  assign new_new_n51089__ = ~new_new_n51086__ & new_new_n51088__;
  assign new_new_n51090__ = ~new_new_n51085__ & ~new_new_n51089__;
  assign new_new_n51091__ = new_new_n51081__ & new_new_n51090__;
  assign new_new_n51092__ = ys__n45735 & ys__n45736;
  assign new_new_n51093__ = ~ys__n45735 & ~ys__n45736;
  assign new_new_n51094__ = ~ys__n45812 & ~new_new_n51093__;
  assign new_new_n51095__ = ~new_new_n51092__ & new_new_n51094__;
  assign new_new_n51096__ = ys__n45738 & ys__n45739;
  assign new_new_n51097__ = ~ys__n45738 & ~ys__n45739;
  assign new_new_n51098__ = ~ys__n45813 & ~new_new_n51097__;
  assign new_new_n51099__ = ~new_new_n51096__ & new_new_n51098__;
  assign new_new_n51100__ = ~new_new_n51095__ & ~new_new_n51099__;
  assign new_new_n51101__ = ys__n45741 & ys__n45742;
  assign new_new_n51102__ = ~ys__n45741 & ~ys__n45742;
  assign new_new_n51103__ = ~ys__n45814 & ~new_new_n51102__;
  assign new_new_n51104__ = ~new_new_n51101__ & new_new_n51103__;
  assign new_new_n51105__ = ys__n45744 & ys__n45745;
  assign new_new_n51106__ = ~ys__n45744 & ~ys__n45745;
  assign new_new_n51107__ = ~ys__n45815 & ~new_new_n51106__;
  assign new_new_n51108__ = ~new_new_n51105__ & new_new_n51107__;
  assign new_new_n51109__ = ~new_new_n51104__ & ~new_new_n51108__;
  assign new_new_n51110__ = new_new_n51100__ & new_new_n51109__;
  assign new_new_n51111__ = new_new_n51091__ & new_new_n51110__;
  assign new_new_n51112__ = new_new_n51072__ & new_new_n51111__;
  assign new_new_n51113__ = new_new_n51033__ & new_new_n51112__;
  assign new_new_n51114__ = ys__n45836 & new_new_n51113__;
  assign new_new_n51115__ = ~new_new_n50959__ & ~new_new_n51114__;
  assign new_new_n51116__ = new_new_n50804__ & new_new_n51115__;
  assign new_new_n51117__ = ~ys__n30225 & ys__n38910;
  assign new_new_n51118__ = ~ys__n1020 & new_new_n51117__;
  assign new_new_n51119__ = ~ys__n38908 & ~new_new_n51118__;
  assign new_new_n51120__ = ~new_new_n51116__ & ~new_new_n51119__;
  assign new_new_n51121__ = ~ys__n38288 & ~new_new_n51120__;
  assign ys__n38209 = ~ys__n4566 & ~new_new_n51121__;
  assign new_new_n51123__ = ys__n46127 & new_new_n50647__;
  assign new_new_n51124__ = ys__n46029 & new_new_n50802__;
  assign new_new_n51125__ = ~new_new_n51123__ & ~new_new_n51124__;
  assign new_new_n51126__ = ys__n45931 & new_new_n50958__;
  assign new_new_n51127__ = ys__n45835 & new_new_n51113__;
  assign new_new_n51128__ = ~new_new_n51126__ & ~new_new_n51127__;
  assign new_new_n51129__ = new_new_n51125__ & new_new_n51128__;
  assign new_new_n51130__ = ~new_new_n51119__ & ~new_new_n51129__;
  assign new_new_n51131__ = ~ys__n38290 & ~new_new_n51130__;
  assign ys__n38211 = ~ys__n4566 & ~new_new_n51131__;
  assign ys__n38213 = ys__n38212 & ~ys__n4566;
  assign new_new_n51134__ = ~ys__n18101 & ~ys__n18106;
  assign new_new_n51135__ = ~ys__n33375 & ys__n38315;
  assign new_new_n51136__ = new_new_n51134__ & new_new_n51135__;
  assign new_new_n51137__ = ys__n38311 & new_new_n51136__;
  assign new_new_n51138__ = ~new_new_n10820__ & new_new_n51137__;
  assign new_new_n51139__ = new_new_n16454__ & new_new_n51136__;
  assign new_new_n51140__ = ys__n23272 & ~ys__n23335;
  assign new_new_n51141__ = ys__n23332 & new_new_n51136__;
  assign new_new_n51142__ = ~new_new_n51140__ & ~new_new_n51141__;
  assign new_new_n51143__ = new_new_n11180__ & ~new_new_n51142__;
  assign new_new_n51144__ = ~new_new_n51139__ & ~new_new_n51143__;
  assign new_new_n51145__ = new_new_n10820__ & ~new_new_n51144__;
  assign new_new_n51146__ = ~new_new_n51138__ & ~new_new_n51145__;
  assign ys__n38214 = ~ys__n4566 & ~new_new_n51146__;
  assign ys__n38216 = ys__n38215 & ~ys__n4566;
  assign ys__n38218 = ys__n38217 & ~ys__n4566;
  assign ys__n38222 = ~ys__n33340 & ys__n478;
  assign new_new_n51151__ = ys__n22818 & ~ys__n33342;
  assign ys__n38224 = ys__n935 | new_new_n51151__;
  assign ys__n38246 = ~new_new_n13884__ & new_new_n13902__;
  assign ys__n38247 = ~new_new_n13884__ & new_new_n13898__;
  assign ys__n38248 = ~new_new_n13884__ & new_new_n13896__;
  assign new_new_n51156__ = new_new_n13884__ & new_new_n13914__;
  assign ys__n38250 = new_new_n13903__ | new_new_n51156__;
  assign new_new_n51158__ = new_new_n13884__ & new_new_n13913__;
  assign ys__n38252 = new_new_n13904__ | new_new_n51158__;
  assign new_new_n51160__ = ~ys__n33364 & ys__n38237;
  assign new_new_n51161__ = new_new_n13884__ & new_new_n51160__;
  assign new_new_n51162__ = ~ys__n33350 & ~new_new_n51161__;
  assign ys__n38263 = ~new_new_n13951__ & ~new_new_n51162__;
  assign new_new_n51164__ = ~ys__n33364 & ys__n38236;
  assign new_new_n51165__ = new_new_n13884__ & new_new_n51164__;
  assign new_new_n51166__ = ~ys__n33352 & ~new_new_n51165__;
  assign ys__n38266 = ~new_new_n13951__ & ~new_new_n51166__;
  assign ys__n38281 = ys__n738 & ~new_new_n50489__;
  assign new_new_n51169__ = ~ys__n38286 & ~new_new_n50488__;
  assign ys__n38285 = ys__n738 & ~new_new_n51169__;
  assign ys__n38287 = ys__n738 & ~new_new_n51121__;
  assign ys__n38289 = ys__n738 & ~new_new_n51131__;
  assign ys__n38292 = ys__n34959 | ys__n38291;
  assign new_new_n51174__ = ys__n422 & ys__n432;
  assign new_new_n51175__ = new_new_n11582__ & new_new_n51174__;
  assign new_new_n51176__ = new_new_n11687__ & new_new_n51175__;
  assign new_new_n51177__ = ~ys__n436 & ~ys__n34959;
  assign new_new_n51178__ = ys__n38291 & new_new_n51177__;
  assign new_new_n51179__ = new_new_n11607__ & new_new_n51178__;
  assign ys__n38294 = new_new_n51176__ & new_new_n51179__;
  assign new_new_n51181__ = ~ys__n935 & ~ys__n34959;
  assign ys__n38296 = ~ys__n33366 & ~new_new_n51181__;
  assign new_new_n51183__ = new_new_n15957__ & ~new_new_n15963__;
  assign new_new_n51184__ = ~new_new_n15965__ & ~new_new_n51183__;
  assign new_new_n51185__ = ~ys__n28243 & ~new_new_n51184__;
  assign new_new_n51186__ = ys__n28243 & ~new_new_n51185__;
  assign new_new_n51187__ = ys__n23480 & new_new_n51185__;
  assign ys__n38303 = new_new_n51186__ | new_new_n51187__;
  assign new_new_n51189__ = ys__n23339 & ~new_new_n11323__;
  assign new_new_n51190__ = ~ys__n28243 & new_new_n11323__;
  assign new_new_n51191__ = ~new_new_n51189__ & ~new_new_n51190__;
  assign new_new_n51192__ = ~new_new_n11175__ & ~new_new_n51191__;
  assign new_new_n51193__ = ~new_new_n34551__ & ~new_new_n51192__;
  assign new_new_n51194__ = ~new_new_n11180__ & ~new_new_n51193__;
  assign new_new_n51195__ = ys__n23335 & new_new_n11180__;
  assign new_new_n51196__ = ~new_new_n51194__ & ~new_new_n51195__;
  assign new_new_n51197__ = new_new_n10820__ & ~new_new_n51196__;
  assign new_new_n51198__ = ys__n23339 & ~new_new_n10820__;
  assign new_new_n51199__ = ~new_new_n51197__ & ~new_new_n51198__;
  assign ys__n38325 = ~ys__n4566 & ~new_new_n51199__;
  assign new_new_n51201__ = new_new_n11192__ & ~new_new_n11194__;
  assign new_new_n51202__ = ~ys__n516 & ~ys__n520;
  assign new_new_n51203__ = ~ys__n2024 & ~ys__n4478;
  assign new_new_n51204__ = ~ys__n4480 & new_new_n51203__;
  assign new_new_n51205__ = new_new_n51202__ & new_new_n51204__;
  assign new_new_n51206__ = new_new_n11212__ & new_new_n51205__;
  assign new_new_n51207__ = ~new_new_n51201__ & new_new_n51206__;
  assign new_new_n51208__ = new_new_n11330__ & ~new_new_n51207__;
  assign new_new_n51209__ = ~new_new_n11193__ & new_new_n11202__;
  assign new_new_n51210__ = new_new_n51201__ & new_new_n51209__;
  assign new_new_n51211__ = ~ys__n28243 & ~new_new_n51210__;
  assign new_new_n51212__ = ~new_new_n51208__ & new_new_n51211__;
  assign new_new_n51213__ = new_new_n11207__ & ~new_new_n15963__;
  assign new_new_n51214__ = new_new_n11257__ & new_new_n15960__;
  assign new_new_n51215__ = new_new_n15958__ & new_new_n51214__;
  assign new_new_n51216__ = ~new_new_n15962__ & ~new_new_n51215__;
  assign new_new_n51217__ = new_new_n15963__ & ~new_new_n51216__;
  assign new_new_n51218__ = new_new_n11207__ & ~new_new_n51217__;
  assign new_new_n51219__ = ~ys__n28243 & ~new_new_n51218__;
  assign new_new_n51220__ = ~new_new_n51213__ & new_new_n51219__;
  assign new_new_n51221__ = ~ys__n23730 & new_new_n15971__;
  assign new_new_n51222__ = ~ys__n23730 & ~new_new_n51221__;
  assign new_new_n51223__ = ys__n28243 & ~new_new_n51222__;
  assign new_new_n51224__ = ~new_new_n51220__ & ~new_new_n51223__;
  assign ys__n38326 = new_new_n51212__ | ~new_new_n51224__;
  assign ys__n38327 = ys__n33359 & ~ys__n4566;
  assign ys__n38328 = ys__n256 & ~ys__n4566;
  assign new_new_n51228__ = new_new_n10630__ & new_new_n10648__;
  assign new_new_n51229__ = new_new_n10658__ & new_new_n11184__;
  assign new_new_n51230__ = new_new_n51228__ & new_new_n51229__;
  assign ys__n38330 = ~ys__n4566 & new_new_n51230__;
  assign ys__n38331 = ys__n262 & ~ys__n4566;
  assign ys__n38332 = ys__n18105 & ~ys__n4566;
  assign new_new_n51234__ = new_new_n11184__ & new_new_n11203__;
  assign ys__n38334 = ~ys__n4566 & new_new_n51234__;
  assign new_new_n51236__ = new_new_n11184__ & new_new_n11250__;
  assign new_new_n51237__ = new_new_n11260__ & new_new_n51236__;
  assign ys__n38336 = ~ys__n4566 & new_new_n51237__;
  assign new_new_n51239__ = ys__n550 & ~ys__n23730;
  assign new_new_n51240__ = ys__n28243 & new_new_n51239__;
  assign new_new_n51241__ = new_new_n11203__ & new_new_n51240__;
  assign ys__n38337 = ~ys__n4566 & new_new_n51241__;
  assign new_new_n51243__ = ~ys__n28243 & new_new_n11200__;
  assign ys__n38339 = ~ys__n4566 & new_new_n51243__;
  assign new_new_n51245__ = ~new_new_n11222__ & ~new_new_n11229__;
  assign new_new_n51246__ = ~ys__n28243 & new_new_n11193__;
  assign new_new_n51247__ = ~new_new_n51245__ & new_new_n51246__;
  assign ys__n38340 = ~ys__n4566 & new_new_n51247__;
  assign new_new_n51249__ = ~new_new_n11217__ & ~new_new_n11228__;
  assign new_new_n51250__ = new_new_n51246__ & ~new_new_n51249__;
  assign ys__n38341 = ~ys__n4566 & new_new_n51250__;
  assign new_new_n51252__ = ~ys__n28243 & new_new_n11198__;
  assign ys__n38342 = ~ys__n4566 & new_new_n51252__;
  assign new_new_n51254__ = ~ys__n28243 & new_new_n10646__;
  assign new_new_n51255__ = ~ys__n23730 & new_new_n10635__;
  assign new_new_n51256__ = new_new_n10633__ & new_new_n51255__;
  assign new_new_n51257__ = ~ys__n23730 & new_new_n10646__;
  assign new_new_n51258__ = ~new_new_n51256__ & ~new_new_n51257__;
  assign new_new_n51259__ = ~new_new_n10633__ & ~new_new_n10646__;
  assign new_new_n51260__ = ys__n28243 & ~new_new_n51259__;
  assign new_new_n51261__ = ~new_new_n51258__ & new_new_n51260__;
  assign new_new_n51262__ = ~new_new_n51254__ & ~new_new_n51261__;
  assign ys__n38343 = ~ys__n4566 & ~new_new_n51262__;
  assign new_new_n51264__ = ~ys__n28243 & new_new_n10643__;
  assign new_new_n51265__ = ~ys__n23730 & new_new_n10637__;
  assign new_new_n51266__ = new_new_n10633__ & new_new_n51265__;
  assign new_new_n51267__ = ~ys__n23730 & new_new_n10643__;
  assign new_new_n51268__ = ~new_new_n51266__ & ~new_new_n51267__;
  assign new_new_n51269__ = ~new_new_n10633__ & ~new_new_n10643__;
  assign new_new_n51270__ = ys__n28243 & ~new_new_n51269__;
  assign new_new_n51271__ = ~new_new_n51268__ & new_new_n51270__;
  assign new_new_n51272__ = ~new_new_n51264__ & ~new_new_n51271__;
  assign ys__n38344 = ~ys__n4566 & ~new_new_n51272__;
  assign new_new_n51274__ = ~ys__n28243 & new_new_n51217__;
  assign new_new_n51275__ = ys__n28243 & new_new_n11250__;
  assign new_new_n51276__ = new_new_n11261__ & new_new_n51275__;
  assign new_new_n51277__ = ~new_new_n51274__ & ~new_new_n51276__;
  assign ys__n38345 = ~ys__n4566 & ~new_new_n51277__;
  assign ys__n38347 = ys__n38346 & ~ys__n4566;
  assign new_new_n51280__ = ys__n22648 & ys__n28432;
  assign new_new_n51281__ = ys__n22650 & ys__n28434;
  assign new_new_n51282__ = ~new_new_n51280__ & ~new_new_n51281__;
  assign new_new_n51283__ = ys__n22652 & ys__n28436;
  assign new_new_n51284__ = ys__n22654 & ys__n28438;
  assign new_new_n51285__ = ~new_new_n51283__ & ~new_new_n51284__;
  assign new_new_n51286__ = new_new_n51282__ & new_new_n51285__;
  assign new_new_n51287__ = ys__n22640 & ys__n28424;
  assign new_new_n51288__ = ys__n22642 & ys__n28426;
  assign new_new_n51289__ = ~new_new_n51287__ & ~new_new_n51288__;
  assign new_new_n51290__ = ys__n22644 & ys__n28428;
  assign new_new_n51291__ = ys__n22646 & ys__n28430;
  assign new_new_n51292__ = ~new_new_n51290__ & ~new_new_n51291__;
  assign new_new_n51293__ = new_new_n51289__ & new_new_n51292__;
  assign new_new_n51294__ = new_new_n51286__ & new_new_n51293__;
  assign new_new_n51295__ = ~ys__n33370 & ~ys__n33389;
  assign new_new_n51296__ = ys__n38427 & new_new_n51295__;
  assign new_new_n51297__ = ~new_new_n51294__ & new_new_n51296__;
  assign new_new_n51298__ = ~ys__n4566 & new_new_n51297__;
  assign ys__n38349 = ~ys__n18120 & new_new_n51298__;
  assign new_new_n51300__ = ~ys__n38420 & new_new_n44372__;
  assign new_new_n51301__ = ~new_new_n44368__ & new_new_n51300__;
  assign new_new_n51302__ = new_new_n44366__ & new_new_n51301__;
  assign ys__n38351 = ~ys__n4566 & ~new_new_n51302__;
  assign new_new_n51304__ = ~ys__n28243 & new_new_n11164__;
  assign ys__n38352 = ~ys__n4566 & new_new_n51304__;
  assign new_new_n51306__ = ys__n748 & ys__n750;
  assign new_new_n51307__ = new_new_n10662__ & new_new_n51306__;
  assign new_new_n51308__ = ys__n742 & ~ys__n744;
  assign new_new_n51309__ = new_new_n10644__ & new_new_n51308__;
  assign new_new_n51310__ = new_new_n51306__ & new_new_n51309__;
  assign new_new_n51311__ = ~new_new_n11194__ & ~new_new_n51310__;
  assign new_new_n51312__ = ~new_new_n51307__ & new_new_n51311__;
  assign ys__n38353 = new_new_n37128__ & ~new_new_n51312__;
  assign new_new_n51314__ = new_new_n10650__ & new_new_n51306__;
  assign new_new_n51315__ = new_new_n10648__ & new_new_n51308__;
  assign new_new_n51316__ = new_new_n51306__ & new_new_n51315__;
  assign new_new_n51317__ = ~new_new_n11191__ & ~new_new_n51316__;
  assign new_new_n51318__ = ~new_new_n51314__ & new_new_n51317__;
  assign ys__n38354 = new_new_n37128__ & ~new_new_n51318__;
  assign new_new_n51320__ = new_new_n10668__ & new_new_n51306__;
  assign new_new_n51321__ = new_new_n10667__ & new_new_n51308__;
  assign new_new_n51322__ = new_new_n51306__ & new_new_n51321__;
  assign new_new_n51323__ = ~new_new_n11190__ & ~new_new_n51322__;
  assign new_new_n51324__ = ~new_new_n51320__ & new_new_n51323__;
  assign ys__n38355 = new_new_n37128__ & ~new_new_n51324__;
  assign new_new_n51326__ = new_new_n10629__ & new_new_n51308__;
  assign new_new_n51327__ = new_new_n10632__ & new_new_n51326__;
  assign new_new_n51328__ = ~ys__n530 & ys__n752;
  assign new_new_n51329__ = new_new_n11259__ & new_new_n51328__;
  assign new_new_n51330__ = ys__n526 & ~ys__n528;
  assign new_new_n51331__ = new_new_n11258__ & new_new_n51328__;
  assign new_new_n51332__ = new_new_n51330__ & new_new_n51331__;
  assign new_new_n51333__ = ~new_new_n51329__ & ~new_new_n51332__;
  assign new_new_n51334__ = new_new_n15963__ & ~new_new_n51333__;
  assign new_new_n51335__ = ~new_new_n51327__ & ~new_new_n51334__;
  assign new_new_n51336__ = ~new_new_n15963__ & ~new_new_n51327__;
  assign new_new_n51337__ = ~ys__n28243 & ~new_new_n51336__;
  assign new_new_n51338__ = ~ys__n4566 & new_new_n51337__;
  assign ys__n38356 = ~new_new_n51335__ & new_new_n51338__;
  assign new_new_n51340__ = ~ys__n28243 & new_new_n11165__;
  assign new_new_n51341__ = new_new_n15958__ & new_new_n15959__;
  assign new_new_n51342__ = new_new_n51340__ & new_new_n51341__;
  assign new_new_n51343__ = new_new_n15963__ & new_new_n51342__;
  assign new_new_n51344__ = ~ys__n522 & ys__n524;
  assign new_new_n51345__ = new_new_n15959__ & new_new_n51344__;
  assign new_new_n51346__ = ~ys__n530 & ys__n28243;
  assign new_new_n51347__ = new_new_n51345__ & new_new_n51346__;
  assign new_new_n51348__ = new_new_n11250__ & new_new_n51347__;
  assign new_new_n51349__ = ~new_new_n51343__ & ~new_new_n51348__;
  assign ys__n38357 = ~ys__n4566 & ~new_new_n51349__;
  assign new_new_n51351__ = new_new_n11257__ & new_new_n15958__;
  assign new_new_n51352__ = new_new_n51340__ & new_new_n51351__;
  assign new_new_n51353__ = new_new_n15963__ & new_new_n51352__;
  assign ys__n38359 = ~ys__n4566 & new_new_n51353__;
  assign new_new_n51355__ = new_new_n11258__ & new_new_n15959__;
  assign new_new_n51356__ = new_new_n15958__ & new_new_n51355__;
  assign new_new_n51357__ = new_new_n11165__ & new_new_n51328__;
  assign new_new_n51358__ = ys__n530 & ys__n752;
  assign new_new_n51359__ = ~new_new_n11169__ & ~new_new_n51358__;
  assign new_new_n51360__ = ~new_new_n51357__ & new_new_n51359__;
  assign new_new_n51361__ = ~new_new_n51356__ & new_new_n51360__;
  assign new_new_n51362__ = new_new_n15958__ & new_new_n51345__;
  assign new_new_n51363__ = ys__n522 & ~ys__n530;
  assign new_new_n51364__ = ~ys__n524 & ys__n526;
  assign new_new_n51365__ = ~ys__n752 & new_new_n51364__;
  assign new_new_n51366__ = new_new_n51363__ & new_new_n51365__;
  assign new_new_n51367__ = ~new_new_n51362__ & ~new_new_n51366__;
  assign new_new_n51368__ = ys__n524 & ys__n526;
  assign new_new_n51369__ = ~ys__n752 & new_new_n51368__;
  assign new_new_n51370__ = new_new_n51363__ & new_new_n51369__;
  assign new_new_n51371__ = ~ys__n524 & ~ys__n526;
  assign new_new_n51372__ = ys__n752 & new_new_n51371__;
  assign new_new_n51373__ = new_new_n51363__ & new_new_n51372__;
  assign new_new_n51374__ = ~new_new_n51370__ & ~new_new_n51373__;
  assign new_new_n51375__ = new_new_n51367__ & new_new_n51374__;
  assign new_new_n51376__ = new_new_n51361__ & new_new_n51375__;
  assign new_new_n51377__ = new_new_n15963__ & ~new_new_n51376__;
  assign new_new_n51378__ = ys__n744 & ys__n746;
  assign new_new_n51379__ = ys__n742 & ys__n750;
  assign new_new_n51380__ = new_new_n51378__ & new_new_n51379__;
  assign new_new_n51381__ = ys__n748 & new_new_n51380__;
  assign new_new_n51382__ = new_new_n10631__ & new_new_n51306__;
  assign new_new_n51383__ = new_new_n11204__ & new_new_n51306__;
  assign new_new_n51384__ = ~new_new_n51382__ & ~new_new_n51383__;
  assign new_new_n51385__ = ~new_new_n51381__ & new_new_n51384__;
  assign new_new_n51386__ = ~ys__n742 & ys__n748;
  assign new_new_n51387__ = ~ys__n750 & new_new_n51386__;
  assign new_new_n51388__ = new_new_n51378__ & new_new_n51387__;
  assign new_new_n51389__ = new_new_n10658__ & new_new_n51315__;
  assign new_new_n51390__ = ~new_new_n51388__ & ~new_new_n51389__;
  assign new_new_n51391__ = new_new_n10657__ & new_new_n51306__;
  assign new_new_n51392__ = new_new_n51306__ & new_new_n51326__;
  assign new_new_n51393__ = ~new_new_n51391__ & ~new_new_n51392__;
  assign new_new_n51394__ = new_new_n51390__ & new_new_n51393__;
  assign new_new_n51395__ = new_new_n10641__ & new_new_n11163__;
  assign new_new_n51396__ = new_new_n11163__ & new_new_n51308__;
  assign new_new_n51397__ = ~new_new_n51395__ & ~new_new_n51396__;
  assign new_new_n51398__ = new_new_n10630__ & new_new_n10658__;
  assign new_new_n51399__ = new_new_n10641__ & new_new_n51306__;
  assign new_new_n51400__ = ~new_new_n51398__ & ~new_new_n51399__;
  assign new_new_n51401__ = new_new_n51397__ & new_new_n51400__;
  assign new_new_n51402__ = ~ys__n748 & new_new_n51380__;
  assign new_new_n51403__ = ~new_new_n10670__ & ~new_new_n51402__;
  assign new_new_n51404__ = new_new_n51401__ & new_new_n51403__;
  assign new_new_n51405__ = new_new_n51394__ & new_new_n51404__;
  assign new_new_n51406__ = new_new_n51385__ & new_new_n51405__;
  assign new_new_n51407__ = new_new_n11167__ & new_new_n51358__;
  assign new_new_n51408__ = new_new_n10631__ & new_new_n11163__;
  assign new_new_n51409__ = ~new_new_n51407__ & new_new_n51408__;
  assign new_new_n51410__ = new_new_n11169__ & new_new_n51214__;
  assign new_new_n51411__ = new_new_n11164__ & new_new_n51410__;
  assign new_new_n51412__ = ~new_new_n51409__ & ~new_new_n51411__;
  assign new_new_n51413__ = new_new_n51406__ & new_new_n51412__;
  assign new_new_n51414__ = ~new_new_n51377__ & new_new_n51413__;
  assign new_new_n51415__ = ~new_new_n11164__ & ~new_new_n15963__;
  assign new_new_n51416__ = ~new_new_n51408__ & new_new_n51415__;
  assign new_new_n51417__ = new_new_n51406__ & new_new_n51416__;
  assign new_new_n51418__ = ~ys__n28243 & ~new_new_n51417__;
  assign new_new_n51419__ = ~new_new_n51414__ & new_new_n51418__;
  assign new_new_n51420__ = new_new_n10630__ & new_new_n10667__;
  assign new_new_n51421__ = new_new_n10632__ & new_new_n51420__;
  assign new_new_n51422__ = ~new_new_n11200__ & ~new_new_n51421__;
  assign new_new_n51423__ = new_new_n10658__ & new_new_n11199__;
  assign new_new_n51424__ = new_new_n10658__ & new_new_n51420__;
  assign new_new_n51425__ = ~new_new_n51423__ & ~new_new_n51424__;
  assign new_new_n51426__ = new_new_n51422__ & new_new_n51425__;
  assign new_new_n51427__ = ~new_new_n10633__ & ~new_new_n11198__;
  assign new_new_n51428__ = new_new_n10631__ & new_new_n10658__;
  assign new_new_n51429__ = ~new_new_n11250__ & ~new_new_n51327__;
  assign new_new_n51430__ = ~new_new_n51428__ & new_new_n51429__;
  assign new_new_n51431__ = new_new_n51427__ & new_new_n51430__;
  assign new_new_n51432__ = new_new_n51426__ & new_new_n51431__;
  assign new_new_n51433__ = ys__n47659 & new_new_n11250__;
  assign new_new_n51434__ = ys__n530 & new_new_n51327__;
  assign new_new_n51435__ = ~new_new_n11257__ & ~new_new_n51330__;
  assign new_new_n51436__ = new_new_n51428__ & ~new_new_n51435__;
  assign new_new_n51437__ = ~new_new_n51434__ & ~new_new_n51436__;
  assign new_new_n51438__ = ~new_new_n51433__ & new_new_n51437__;
  assign new_new_n51439__ = ys__n550 & new_new_n10636__;
  assign new_new_n51440__ = ~ys__n518 & ys__n548;
  assign new_new_n51441__ = ys__n550 & new_new_n51440__;
  assign new_new_n51442__ = ~new_new_n51439__ & ~new_new_n51441__;
  assign new_new_n51443__ = new_new_n10633__ & ~new_new_n51442__;
  assign new_new_n51444__ = new_new_n11198__ & new_new_n15959__;
  assign new_new_n51445__ = ~new_new_n51443__ & ~new_new_n51444__;
  assign new_new_n51446__ = new_new_n51426__ & new_new_n51445__;
  assign new_new_n51447__ = new_new_n51438__ & new_new_n51446__;
  assign new_new_n51448__ = ys__n28243 & ~new_new_n51447__;
  assign new_new_n51449__ = ~new_new_n51432__ & new_new_n51448__;
  assign new_new_n51450__ = ~new_new_n51419__ & ~new_new_n51449__;
  assign ys__n38360 = ~ys__n4566 & ~new_new_n51450__;
  assign ys__n38362 = ys__n38361 & ~ys__n4566;
  assign new_new_n51453__ = ys__n520 & new_new_n51358__;
  assign new_new_n51454__ = new_new_n51214__ & new_new_n51453__;
  assign new_new_n51455__ = new_new_n51304__ & new_new_n51454__;
  assign ys__n38364 = ~ys__n4566 & new_new_n51455__;
  assign new_new_n51457__ = ~ys__n512 & ~ys__n520;
  assign new_new_n51458__ = ~ys__n632 & new_new_n51457__;
  assign new_new_n51459__ = new_new_n11210__ & new_new_n51458__;
  assign new_new_n51460__ = ys__n23705 & ~ys__n28243;
  assign new_new_n51461__ = new_new_n11164__ & new_new_n51460__;
  assign new_new_n51462__ = new_new_n51459__ & new_new_n51461__;
  assign ys__n38365 = ~ys__n4566 & new_new_n51462__;
  assign new_new_n51464__ = ys__n23706 & ~ys__n28243;
  assign new_new_n51465__ = new_new_n11164__ & new_new_n51464__;
  assign new_new_n51466__ = new_new_n51459__ & new_new_n51465__;
  assign ys__n38366 = ~ys__n4566 & new_new_n51466__;
  assign new_new_n51468__ = ys__n23707 & ~ys__n28243;
  assign new_new_n51469__ = new_new_n11164__ & new_new_n51468__;
  assign new_new_n51470__ = new_new_n51459__ & new_new_n51469__;
  assign ys__n38367 = ~ys__n4566 & new_new_n51470__;
  assign new_new_n51472__ = ys__n23708 & ~ys__n28243;
  assign new_new_n51473__ = new_new_n11164__ & new_new_n51472__;
  assign new_new_n51474__ = new_new_n51459__ & new_new_n51473__;
  assign ys__n38368 = ~ys__n4566 & new_new_n51474__;
  assign new_new_n51476__ = ys__n23709 & ~ys__n28243;
  assign new_new_n51477__ = new_new_n11164__ & new_new_n51476__;
  assign new_new_n51478__ = new_new_n51459__ & new_new_n51477__;
  assign ys__n38369 = ~ys__n4566 & new_new_n51478__;
  assign new_new_n51480__ = ys__n23710 & ~ys__n28243;
  assign new_new_n51481__ = new_new_n11164__ & new_new_n51480__;
  assign new_new_n51482__ = new_new_n51459__ & new_new_n51481__;
  assign ys__n38370 = ~ys__n4566 & new_new_n51482__;
  assign new_new_n51484__ = ys__n23711 & ~ys__n28243;
  assign new_new_n51485__ = new_new_n11164__ & new_new_n51484__;
  assign new_new_n51486__ = new_new_n51459__ & new_new_n51485__;
  assign ys__n38371 = ~ys__n4566 & new_new_n51486__;
  assign new_new_n51488__ = ys__n23712 & ~ys__n28243;
  assign new_new_n51489__ = new_new_n11164__ & new_new_n51488__;
  assign new_new_n51490__ = new_new_n51459__ & new_new_n51489__;
  assign ys__n38372 = ~ys__n4566 & new_new_n51490__;
  assign new_new_n51492__ = ys__n23713 & ~ys__n28243;
  assign new_new_n51493__ = new_new_n11164__ & new_new_n51492__;
  assign new_new_n51494__ = new_new_n51459__ & new_new_n51493__;
  assign ys__n38373 = ~ys__n4566 & new_new_n51494__;
  assign new_new_n51496__ = ys__n23714 & ~ys__n28243;
  assign new_new_n51497__ = new_new_n11164__ & new_new_n51496__;
  assign new_new_n51498__ = new_new_n51459__ & new_new_n51497__;
  assign ys__n38374 = ~ys__n4566 & new_new_n51498__;
  assign new_new_n51500__ = ys__n23715 & ~ys__n28243;
  assign new_new_n51501__ = new_new_n11164__ & new_new_n51500__;
  assign new_new_n51502__ = new_new_n51459__ & new_new_n51501__;
  assign ys__n38375 = ~ys__n4566 & new_new_n51502__;
  assign ys__n38377 = ys__n38376 & ~ys__n4566;
  assign ys__n38379 = ys__n38378 & ~ys__n4566;
  assign ys__n38381 = ys__n38380 & ~ys__n4566;
  assign ys__n38383 = ys__n38382 & ~ys__n4566;
  assign ys__n38385 = ys__n38384 & ~ys__n4566;
  assign ys__n38387 = ys__n38386 & ~ys__n4566;
  assign new_new_n51510__ = ys__n632 & new_new_n51457__;
  assign new_new_n51511__ = new_new_n11210__ & new_new_n51510__;
  assign new_new_n51512__ = ys__n634 & ys__n636;
  assign new_new_n51513__ = ~ys__n638 & ~ys__n640;
  assign new_new_n51514__ = ~ys__n642 & ~ys__n28243;
  assign new_new_n51515__ = new_new_n51513__ & new_new_n51514__;
  assign new_new_n51516__ = new_new_n51512__ & new_new_n51515__;
  assign new_new_n51517__ = new_new_n11164__ & new_new_n51516__;
  assign new_new_n51518__ = new_new_n51511__ & new_new_n51517__;
  assign ys__n38388 = ~ys__n4566 & new_new_n51518__;
  assign new_new_n51520__ = ~ys__n638 & ys__n640;
  assign new_new_n51521__ = new_new_n51512__ & new_new_n51514__;
  assign new_new_n51522__ = new_new_n51520__ & new_new_n51521__;
  assign new_new_n51523__ = new_new_n11164__ & new_new_n51522__;
  assign new_new_n51524__ = new_new_n51511__ & new_new_n51523__;
  assign ys__n38389 = ~ys__n4566 & new_new_n51524__;
  assign new_new_n51526__ = ~ys__n634 & ys__n636;
  assign new_new_n51527__ = new_new_n11565__ & new_new_n51526__;
  assign new_new_n51528__ = new_new_n51513__ & new_new_n51527__;
  assign new_new_n51529__ = new_new_n11164__ & new_new_n51528__;
  assign new_new_n51530__ = new_new_n51511__ & new_new_n51529__;
  assign ys__n38390 = ~ys__n4566 & new_new_n51530__;
  assign new_new_n51532__ = ~ys__n634 & ~ys__n636;
  assign new_new_n51533__ = new_new_n11565__ & new_new_n51513__;
  assign new_new_n51534__ = new_new_n51532__ & new_new_n51533__;
  assign new_new_n51535__ = new_new_n11164__ & new_new_n51534__;
  assign new_new_n51536__ = new_new_n51511__ & new_new_n51535__;
  assign ys__n38391 = ~ys__n4566 & new_new_n51536__;
  assign new_new_n51538__ = new_new_n11565__ & new_new_n51520__;
  assign new_new_n51539__ = new_new_n51532__ & new_new_n51538__;
  assign new_new_n51540__ = new_new_n11164__ & new_new_n51539__;
  assign new_new_n51541__ = new_new_n51511__ & new_new_n51540__;
  assign ys__n38392 = ~ys__n4566 & new_new_n51541__;
  assign new_new_n51543__ = ys__n640 & ys__n642;
  assign new_new_n51544__ = new_new_n11466__ & new_new_n51543__;
  assign new_new_n51545__ = new_new_n51512__ & new_new_n51544__;
  assign new_new_n51546__ = new_new_n11164__ & new_new_n51545__;
  assign new_new_n51547__ = new_new_n51511__ & new_new_n51546__;
  assign ys__n38393 = ~ys__n4566 & new_new_n51547__;
  assign new_new_n51549__ = ~ys__n4458 & ~ys__n4461;
  assign new_new_n51550__ = ~ys__n4465 & new_new_n51549__;
  assign new_new_n51551__ = ~ys__n4454 & ~ys__n4455;
  assign new_new_n51552__ = new_new_n34089__ & new_new_n51551__;
  assign new_new_n51553__ = new_new_n33965__ & new_new_n34127__;
  assign new_new_n51554__ = new_new_n51552__ & new_new_n51553__;
  assign new_new_n51555__ = new_new_n51550__ & new_new_n51554__;
  assign ys__n38394 = ~ys__n4566 & ~new_new_n51555__;
  assign new_new_n51557__ = ~ys__n28243 & new_new_n11210__;
  assign new_new_n51558__ = new_new_n11216__ & new_new_n51557__;
  assign new_new_n51559__ = new_new_n11259__ & new_new_n51558__;
  assign new_new_n51560__ = ~ys__n516 & ~ys__n550;
  assign new_new_n51561__ = new_new_n10636__ & new_new_n51560__;
  assign new_new_n51562__ = new_new_n11170__ & new_new_n51561__;
  assign new_new_n51563__ = ~ys__n640 & ~ys__n642;
  assign new_new_n51564__ = ~ys__n736 & ~ys__n4488;
  assign new_new_n51565__ = new_new_n51563__ & new_new_n51564__;
  assign new_new_n51566__ = ~ys__n632 & ~ys__n634;
  assign new_new_n51567__ = ~ys__n636 & ~ys__n638;
  assign new_new_n51568__ = new_new_n51566__ & new_new_n51567__;
  assign new_new_n51569__ = new_new_n51565__ & new_new_n51568__;
  assign new_new_n51570__ = new_new_n51562__ & new_new_n51569__;
  assign new_new_n51571__ = new_new_n11164__ & new_new_n51570__;
  assign new_new_n51572__ = new_new_n51559__ & new_new_n51571__;
  assign ys__n38396 = ~ys__n4566 & new_new_n51572__;
  assign new_new_n51574__ = ~ys__n28243 & new_new_n51407__;
  assign new_new_n51575__ = new_new_n51408__ & new_new_n51574__;
  assign new_new_n51576__ = ~ys__n23730 & new_new_n51346__;
  assign new_new_n51577__ = new_new_n51355__ & new_new_n51576__;
  assign new_new_n51578__ = new_new_n11250__ & new_new_n51577__;
  assign new_new_n51579__ = ~new_new_n51575__ & ~new_new_n51578__;
  assign ys__n38397 = ~ys__n4566 & ~new_new_n51579__;
  assign new_new_n51581__ = new_new_n18424__ & ~new_new_n20775__;
  assign new_new_n51582__ = ~new_new_n18424__ & new_new_n20775__;
  assign new_new_n51583__ = ~new_new_n51581__ & ~new_new_n51582__;
  assign new_new_n51584__ = ys__n38418 & ~ys__n4566;
  assign ys__n38417 = ~new_new_n51583__ & new_new_n51584__;
  assign new_new_n51586__ = new_new_n10990__ & new_new_n11003__;
  assign new_new_n51587__ = ys__n23717 & ys__n33403;
  assign new_new_n51588__ = ~new_new_n51586__ & new_new_n51587__;
  assign new_new_n51589__ = new_new_n11006__ & new_new_n51588__;
  assign new_new_n51590__ = ~ys__n935 & ~ys__n38473;
  assign new_new_n51591__ = ys__n33403 & new_new_n10993__;
  assign new_new_n51592__ = new_new_n51590__ & ~new_new_n51591__;
  assign new_new_n51593__ = ~new_new_n10990__ & ~new_new_n51592__;
  assign new_new_n51594__ = ys__n738 & new_new_n51593__;
  assign new_new_n51595__ = ys__n935 & ~new_new_n10990__;
  assign new_new_n51596__ = new_new_n12583__ & new_new_n51595__;
  assign new_new_n51597__ = ~new_new_n51594__ & ~new_new_n51596__;
  assign new_new_n51598__ = ~new_new_n51589__ & new_new_n51597__;
  assign new_new_n51599__ = ~new_new_n44177__ & ~new_new_n51598__;
  assign new_new_n51600__ = ~new_new_n12555__ & ~new_new_n12629__;
  assign new_new_n51601__ = ~new_new_n41468__ & ~new_new_n41483__;
  assign new_new_n51602__ = new_new_n12629__ & ~new_new_n51601__;
  assign new_new_n51603__ = ~new_new_n51600__ & ~new_new_n51602__;
  assign new_new_n51604__ = ~ys__n33396 & ~ys__n33398;
  assign new_new_n51605__ = ys__n33403 & new_new_n51604__;
  assign new_new_n51606__ = ~ys__n4566 & new_new_n51605__;
  assign new_new_n51607__ = new_new_n11006__ & new_new_n51606__;
  assign new_new_n51608__ = ~new_new_n51603__ & new_new_n51607__;
  assign new_new_n51609__ = new_new_n51590__ & ~new_new_n51606__;
  assign new_new_n51610__ = ys__n738 & ~new_new_n51609__;
  assign new_new_n51611__ = ~new_new_n51603__ & new_new_n51610__;
  assign new_new_n51612__ = ys__n935 & new_new_n12555__;
  assign new_new_n51613__ = ys__n935 & ~new_new_n51612__;
  assign new_new_n51614__ = new_new_n12583__ & new_new_n51613__;
  assign new_new_n51615__ = ~new_new_n51611__ & ~new_new_n51614__;
  assign new_new_n51616__ = ~new_new_n51608__ & new_new_n51615__;
  assign new_new_n51617__ = ~new_new_n44177__ & ~new_new_n51616__;
  assign new_new_n51618__ = ~new_new_n51599__ & ~new_new_n51617__;
  assign ys__n38456 = ys__n30863 & ~new_new_n51618__;
  assign new_new_n51620__ = ~ys__n626 & ys__n664;
  assign new_new_n51621__ = new_new_n21880__ & new_new_n51620__;
  assign new_new_n51622__ = ~ys__n662 & ~ys__n668;
  assign new_new_n51623__ = new_new_n21879__ & new_new_n51622__;
  assign new_new_n51624__ = new_new_n51620__ & new_new_n51623__;
  assign new_new_n51625__ = ys__n662 & ~ys__n668;
  assign new_new_n51626__ = new_new_n21879__ & new_new_n51620__;
  assign new_new_n51627__ = new_new_n51625__ & new_new_n51626__;
  assign new_new_n51628__ = ~new_new_n51624__ & ~new_new_n51627__;
  assign new_new_n51629__ = ~new_new_n51621__ & new_new_n51628__;
  assign ys__n38508 = ys__n33414 & ~new_new_n51629__;
  assign new_new_n51631__ = new_new_n21852__ & new_new_n51622__;
  assign new_new_n51632__ = new_new_n51620__ & new_new_n51631__;
  assign new_new_n51633__ = ys__n660 & ~ys__n666;
  assign new_new_n51634__ = new_new_n51620__ & new_new_n51622__;
  assign new_new_n51635__ = new_new_n51633__ & new_new_n51634__;
  assign new_new_n51636__ = ~new_new_n51632__ & ~new_new_n51635__;
  assign new_new_n51637__ = new_new_n21853__ & new_new_n51620__;
  assign new_new_n51638__ = new_new_n21852__ & new_new_n51620__;
  assign new_new_n51639__ = new_new_n51625__ & new_new_n51638__;
  assign new_new_n51640__ = new_new_n51620__ & new_new_n51625__;
  assign new_new_n51641__ = new_new_n51633__ & new_new_n51640__;
  assign new_new_n51642__ = ~new_new_n51639__ & ~new_new_n51641__;
  assign new_new_n51643__ = ~new_new_n51637__ & new_new_n51642__;
  assign new_new_n51644__ = new_new_n51636__ & new_new_n51643__;
  assign ys__n38509 = ys__n33414 & ~new_new_n51644__;
  assign ys__n38510 = ys__n846 | ~new_new_n22618__;
  assign ys__n38515 = ~ys__n18120 & new_new_n22060__;
  assign new_new_n51648__ = ~ys__n33431 & ys__n38553;
  assign new_new_n51649__ = ~ys__n24131 & ~new_new_n51648__;
  assign ys__n38518 = ~ys__n1036 & ~new_new_n51649__;
  assign new_new_n51651__ = ys__n24145 & ys__n38518;
  assign ys__n38520 = ~ys__n24145 | new_new_n51651__;
  assign new_new_n51653__ = ~ys__n4185 & new_new_n22014__;
  assign ys__n38523 = ys__n38522 | new_new_n51653__;
  assign ys__n38525 = ys__n1029 | ys__n1036;
  assign new_new_n51656__ = ys__n33442 & ~ys__n18120;
  assign ys__n38552 = new_new_n22387__ & ~new_new_n51656__;
  assign new_new_n51658__ = ~ys__n24228 & ~new_new_n51648__;
  assign ys__n38555 = ~ys__n1076 & ~new_new_n51658__;
  assign new_new_n51660__ = ys__n24236 & ys__n38555;
  assign ys__n38563 = ~ys__n24236 | new_new_n51660__;
  assign new_new_n51662__ = ys__n33491 & ys__n33497;
  assign new_new_n51663__ = ~ys__n33495 & ~new_new_n51662__;
  assign new_new_n51664__ = ~ys__n4566 & new_new_n51663__;
  assign ys__n38615 = ys__n24271 & new_new_n51664__;
  assign new_new_n51666__ = ~ys__n33451 & ys__n38620;
  assign new_new_n51667__ = ~ys__n33499 & ~new_new_n51666__;
  assign ys__n38623 = ~ys__n1094 & ~new_new_n51667__;
  assign ys__n38650 = ~ys__n33455 & ys__n33454;
  assign new_new_n51670__ = ~ys__n33457 & ys__n24268;
  assign new_new_n51671__ = ys__n24502 & new_new_n51670__;
  assign ys__n38662 = ys__n24255 | new_new_n51671__;
  assign new_new_n51673__ = ~ys__n24447 & ~ys__n24541;
  assign new_new_n51674__ = ~ys__n24502 & new_new_n51673__;
  assign new_new_n51675__ = new_new_n16582__ & ys__n38623;
  assign new_new_n51676__ = ~ys__n4566 & new_new_n51675__;
  assign new_new_n51677__ = ~ys__n24259 & new_new_n51676__;
  assign new_new_n51678__ = ~ys__n24262 & new_new_n51677__;
  assign new_new_n51679__ = ys__n24502 & new_new_n51678__;
  assign ys__n38668 = new_new_n51674__ | new_new_n51679__;
  assign ys__n38669 = ys__n38662 | ys__n38668;
  assign new_new_n51682__ = ys__n18214 & ~ys__n18216;
  assign ys__n38672 = ys__n18218 & new_new_n51682__;
  assign new_new_n51684__ = ys__n1511 & ys__n30216;
  assign ys__n38674 = ~ys__n4566 & new_new_n51684__;
  assign new_new_n51686__ = ys__n1110 & ys__n33488;
  assign ys__n38689 = new_new_n23427__ | new_new_n51686__;
  assign new_new_n51688__ = ys__n33552 & new_new_n12472__;
  assign new_new_n51689__ = ~new_new_n23364__ & ~new_new_n51688__;
  assign new_new_n51690__ = ~ys__n33491 & ~new_new_n51689__;
  assign new_new_n51691__ = ~ys__n33491 & ys__n33552;
  assign new_new_n51692__ = new_new_n12472__ & ~new_new_n51691__;
  assign new_new_n51693__ = ~new_new_n22467__ & new_new_n51692__;
  assign new_new_n51694__ = ~new_new_n51690__ & ~new_new_n51693__;
  assign new_new_n51695__ = ~ys__n4566 & new_new_n22447__;
  assign new_new_n51696__ = ~new_new_n51694__ & new_new_n51695__;
  assign ys__n38742 = ~ys__n4696 & new_new_n51696__;
  assign new_new_n51698__ = ys__n1106 & new_new_n12472__;
  assign new_new_n51699__ = ~new_new_n51691__ & new_new_n51698__;
  assign new_new_n51700__ = new_new_n16582__ & new_new_n51699__;
  assign new_new_n51701__ = ~new_new_n22467__ & new_new_n51700__;
  assign new_new_n51702__ = new_new_n22446__ & new_new_n51701__;
  assign new_new_n51703__ = ~ys__n4566 & new_new_n51702__;
  assign ys__n38768 = ~ys__n4696 & new_new_n51703__;
  assign ys__n38795 = ys__n33515 & ys__n33514;
  assign new_new_n51706__ = ~ys__n24581 & ~ys__n24604;
  assign new_new_n51707__ = new_new_n16608__ & new_new_n51706__;
  assign ys__n38799 = ys__n18136 | new_new_n51707__;
  assign ys__n38884 = ~ys__n29117 & ys__n38883;
  assign ys__n38886 = ~ys__n29117 & ys__n38885;
  assign new_new_n51711__ = ys__n48 & ~ys__n50;
  assign new_new_n51712__ = ys__n52 & new_new_n51711__;
  assign new_new_n51713__ = ys__n56 & ys__n58;
  assign new_new_n51714__ = ys__n60 & ys__n62;
  assign new_new_n51715__ = new_new_n51713__ & new_new_n51714__;
  assign new_new_n51716__ = ys__n48 & ys__n50;
  assign new_new_n51717__ = ys__n52 & ys__n54;
  assign new_new_n51718__ = new_new_n51716__ & new_new_n51717__;
  assign new_new_n51719__ = new_new_n51715__ & new_new_n51718__;
  assign ys__n38887 = new_new_n51712__ | new_new_n51719__;
  assign ys__n38900 = ~ys__n33558 & ys__n740;
  assign new_new_n51722__ = ys__n30214 & ~ys__n3039;
  assign ys__n38912 = ys__n23850 | new_new_n51722__;
  assign ys__n38913 = ys__n30217 & ~ys__n4566;
  assign new_new_n51725__ = ys__n30216 & ~ys__n740;
  assign new_new_n51726__ = ys__n30217 & ys__n740;
  assign new_new_n51727__ = ~new_new_n51725__ & ~new_new_n51726__;
  assign ys__n38914 = ~ys__n4566 & ~new_new_n51727__;
  assign new_new_n51729__ = ys__n30219 & ~ys__n740;
  assign new_new_n51730__ = ys__n30220 & ys__n740;
  assign new_new_n51731__ = ~new_new_n51729__ & ~new_new_n51730__;
  assign ys__n38915 = ~ys__n4566 & ~new_new_n51731__;
  assign new_new_n51733__ = ys__n30225 & ~ys__n30223;
  assign ys__n38917 = ys__n1020 | new_new_n51733__;
  assign new_new_n51735__ = ys__n28438 & ~ys__n33574;
  assign new_new_n51736__ = ys__n28434 & ~ys__n33570;
  assign new_new_n51737__ = ys__n28436 & ~ys__n33572;
  assign new_new_n51738__ = ~new_new_n51736__ & ~new_new_n51737__;
  assign new_new_n51739__ = ~new_new_n51735__ & new_new_n51738__;
  assign new_new_n51740__ = ys__n28428 & ~ys__n33564;
  assign new_new_n51741__ = ~ys__n38277 & ~new_new_n51740__;
  assign new_new_n51742__ = ys__n28430 & ~ys__n33566;
  assign new_new_n51743__ = ys__n28432 & ~ys__n33568;
  assign new_new_n51744__ = ~new_new_n51742__ & ~new_new_n51743__;
  assign new_new_n51745__ = new_new_n51741__ & new_new_n51744__;
  assign ys__n38923 = ~new_new_n51739__ | ~new_new_n51745__;
  assign new_new_n51747__ = ~ys__n33576 & ys__n38927;
  assign new_new_n51748__ = ys__n38928 & ys__n38929;
  assign ys__n38925 = new_new_n51747__ & new_new_n51748__;
  assign ys__n38930 = ~ys__n398 & ~new_new_n14002__;
  assign new_new_n51751__ = ys__n196 & ys__n198;
  assign new_new_n51752__ = ~ys__n2830 & new_new_n51751__;
  assign new_new_n51753__ = ys__n196 & ys__n2830;
  assign new_new_n51754__ = ~ys__n196 & ~ys__n2830;
  assign new_new_n51755__ = ~new_new_n51753__ & ~new_new_n51754__;
  assign new_new_n51756__ = ~new_new_n51752__ & new_new_n51755__;
  assign new_new_n51757__ = ~ys__n196 & new_new_n40638__;
  assign new_new_n51758__ = ys__n196 & ~ys__n198;
  assign new_new_n51759__ = ~ys__n2830 & new_new_n51758__;
  assign new_new_n51760__ = ~ys__n196 & new_new_n51753__;
  assign new_new_n51761__ = ~new_new_n51759__ & ~new_new_n51760__;
  assign new_new_n51762__ = ~new_new_n51757__ & new_new_n51761__;
  assign new_new_n51763__ = new_new_n51756__ & new_new_n51762__;
  assign new_new_n51764__ = ys__n48259 & new_new_n51759__;
  assign new_new_n51765__ = ys__n48259 & new_new_n51753__;
  assign ys__n44968 = ys__n352 & ys__n27855;
  assign new_new_n51767__ = new_new_n51754__ & ys__n44968;
  assign new_new_n51768__ = ~new_new_n51765__ & ~new_new_n51767__;
  assign new_new_n51769__ = ~new_new_n51764__ & new_new_n51768__;
  assign new_new_n51770__ = new_new_n51757__ & ys__n44968;
  assign new_new_n51771__ = ys__n48259 & new_new_n51752__;
  assign ys__n44952 = ys__n352 & ys__n28015;
  assign new_new_n51773__ = new_new_n51760__ & ys__n44952;
  assign new_new_n51774__ = ~new_new_n51771__ & ~new_new_n51773__;
  assign new_new_n51775__ = ~new_new_n51770__ & new_new_n51774__;
  assign new_new_n51776__ = new_new_n51769__ & new_new_n51775__;
  assign new_new_n51777__ = ~new_new_n51763__ & ~new_new_n51776__;
  assign new_new_n51778__ = ys__n48275 & new_new_n51752__;
  assign new_new_n51779__ = ~new_new_n51763__ & new_new_n51778__;
  assign new_new_n51780__ = new_new_n51777__ & ~new_new_n51779__;
  assign new_new_n51781__ = new_new_n51777__ & ~new_new_n51780__;
  assign new_new_n51782__ = ys__n48260 & new_new_n51759__;
  assign new_new_n51783__ = ys__n48260 & new_new_n51753__;
  assign ys__n44969 = ys__n352 & ys__n27857;
  assign new_new_n51785__ = new_new_n51754__ & ys__n44969;
  assign new_new_n51786__ = ~new_new_n51783__ & ~new_new_n51785__;
  assign new_new_n51787__ = ~new_new_n51782__ & new_new_n51786__;
  assign new_new_n51788__ = new_new_n51757__ & ys__n44969;
  assign new_new_n51789__ = ys__n48260 & new_new_n51752__;
  assign ys__n44953 = ys__n352 & ys__n28016;
  assign new_new_n51791__ = new_new_n51760__ & ys__n44953;
  assign new_new_n51792__ = ~new_new_n51789__ & ~new_new_n51791__;
  assign new_new_n51793__ = ~new_new_n51788__ & new_new_n51792__;
  assign new_new_n51794__ = new_new_n51787__ & new_new_n51793__;
  assign new_new_n51795__ = ~new_new_n51763__ & ~new_new_n51794__;
  assign new_new_n51796__ = ~new_new_n51781__ & ~new_new_n51795__;
  assign new_new_n51797__ = ys__n48261 & new_new_n51759__;
  assign new_new_n51798__ = ys__n48261 & new_new_n51753__;
  assign ys__n44970 = ys__n352 & ys__n27859;
  assign new_new_n51800__ = new_new_n51754__ & ys__n44970;
  assign new_new_n51801__ = ~new_new_n51798__ & ~new_new_n51800__;
  assign new_new_n51802__ = ~new_new_n51797__ & new_new_n51801__;
  assign new_new_n51803__ = new_new_n51757__ & ys__n44970;
  assign new_new_n51804__ = ys__n48261 & new_new_n51752__;
  assign ys__n44954 = ys__n352 & ys__n28017;
  assign new_new_n51806__ = new_new_n51760__ & ys__n44954;
  assign new_new_n51807__ = ~new_new_n51804__ & ~new_new_n51806__;
  assign new_new_n51808__ = ~new_new_n51803__ & new_new_n51807__;
  assign new_new_n51809__ = new_new_n51802__ & new_new_n51808__;
  assign new_new_n51810__ = ~new_new_n51763__ & ~new_new_n51809__;
  assign new_new_n51811__ = new_new_n51796__ & ~new_new_n51810__;
  assign new_new_n51812__ = ~new_new_n51777__ & ~new_new_n51779__;
  assign new_new_n51813__ = new_new_n51795__ & new_new_n51812__;
  assign new_new_n51814__ = new_new_n51795__ & ~new_new_n51813__;
  assign new_new_n51815__ = new_new_n51810__ & ~new_new_n51814__;
  assign new_new_n51816__ = ~new_new_n51811__ & ~new_new_n51815__;
  assign new_new_n51817__ = ys__n162 & ~ys__n346;
  assign new_new_n51818__ = new_new_n12339__ & new_new_n51817__;
  assign new_new_n51819__ = ys__n352 & new_new_n41384__;
  assign new_new_n51820__ = new_new_n51818__ & new_new_n51819__;
  assign new_new_n51821__ = ys__n352 & new_new_n41391__;
  assign new_new_n51822__ = new_new_n51818__ & new_new_n51821__;
  assign new_new_n51823__ = ~new_new_n51820__ & ~new_new_n51822__;
  assign new_new_n51824__ = new_new_n12598__ & new_new_n51818__;
  assign new_new_n51825__ = new_new_n12344__ & new_new_n12596__;
  assign new_new_n51826__ = ys__n352 & new_new_n51818__;
  assign new_new_n51827__ = new_new_n51825__ & new_new_n51826__;
  assign new_new_n51828__ = ~new_new_n51824__ & ~new_new_n51827__;
  assign new_new_n51829__ = new_new_n51823__ & new_new_n51828__;
  assign new_new_n51830__ = new_new_n41389__ & new_new_n41402__;
  assign new_new_n51831__ = new_new_n12604__ & new_new_n41393__;
  assign new_new_n51832__ = new_new_n51830__ & new_new_n51831__;
  assign new_new_n51833__ = ~ys__n196 & ys__n948;
  assign ys__n44836 = ~new_new_n51832__ & new_new_n51833__;
  assign new_new_n51835__ = ys__n1817 & ys__n44836;
  assign new_new_n51836__ = new_new_n51829__ & ~new_new_n51835__;
  assign new_new_n51837__ = ys__n948 & ~new_new_n51836__;
  assign new_new_n51838__ = ys__n196 & ys__n44833;
  assign new_new_n51839__ = ~new_new_n51837__ & ~new_new_n51838__;
  assign new_new_n51840__ = new_new_n51816__ & ~new_new_n51839__;
  assign new_new_n51841__ = ~new_new_n51816__ & new_new_n51839__;
  assign ys__n39395 = new_new_n51840__ | new_new_n51841__;
  assign new_new_n51843__ = new_new_n51777__ & new_new_n51779__;
  assign new_new_n51844__ = ~new_new_n51795__ & new_new_n51843__;
  assign new_new_n51845__ = ~new_new_n51813__ & ~new_new_n51844__;
  assign new_new_n51846__ = ~new_new_n51810__ & ~new_new_n51845__;
  assign new_new_n51847__ = ~new_new_n51777__ & new_new_n51779__;
  assign new_new_n51848__ = ~new_new_n51777__ & ~new_new_n51847__;
  assign new_new_n51849__ = new_new_n51795__ & ~new_new_n51848__;
  assign new_new_n51850__ = ~new_new_n51796__ & ~new_new_n51849__;
  assign new_new_n51851__ = new_new_n51810__ & ~new_new_n51850__;
  assign new_new_n51852__ = ~new_new_n51846__ & ~new_new_n51851__;
  assign new_new_n51853__ = ~new_new_n51839__ & new_new_n51852__;
  assign new_new_n51854__ = new_new_n51839__ & ~new_new_n51852__;
  assign ys__n39396 = new_new_n51853__ | new_new_n51854__;
  assign new_new_n51856__ = ~new_new_n51795__ & new_new_n51812__;
  assign new_new_n51857__ = ~new_new_n51780__ & ~new_new_n51847__;
  assign new_new_n51858__ = new_new_n51795__ & ~new_new_n51857__;
  assign new_new_n51859__ = ~new_new_n51856__ & ~new_new_n51858__;
  assign new_new_n51860__ = ~new_new_n51810__ & ~new_new_n51859__;
  assign new_new_n51861__ = ~new_new_n51812__ & ~new_new_n51843__;
  assign new_new_n51862__ = ~new_new_n51795__ & ~new_new_n51861__;
  assign new_new_n51863__ = ~new_new_n51781__ & new_new_n51795__;
  assign new_new_n51864__ = ~new_new_n51862__ & ~new_new_n51863__;
  assign new_new_n51865__ = new_new_n51810__ & ~new_new_n51864__;
  assign new_new_n51866__ = ~new_new_n51860__ & ~new_new_n51865__;
  assign new_new_n51867__ = ~new_new_n51839__ & new_new_n51866__;
  assign new_new_n51868__ = new_new_n51839__ & ~new_new_n51866__;
  assign ys__n39397 = new_new_n51867__ | new_new_n51868__;
  assign new_new_n51870__ = new_new_n51795__ & ~new_new_n51810__;
  assign new_new_n51871__ = new_new_n51843__ & new_new_n51870__;
  assign new_new_n51872__ = ~new_new_n51795__ & ~new_new_n51848__;
  assign new_new_n51873__ = ~new_new_n51795__ & ~new_new_n51872__;
  assign new_new_n51874__ = new_new_n51810__ & ~new_new_n51873__;
  assign new_new_n51875__ = ~new_new_n51871__ & ~new_new_n51874__;
  assign new_new_n51876__ = ~new_new_n51839__ & new_new_n51875__;
  assign new_new_n51877__ = new_new_n51839__ & ~new_new_n51875__;
  assign ys__n39398 = new_new_n51876__ | new_new_n51877__;
  assign new_new_n51879__ = ys__n48262 & new_new_n51759__;
  assign new_new_n51880__ = ys__n48262 & new_new_n51753__;
  assign ys__n44971 = ys__n352 & ys__n27861;
  assign new_new_n51882__ = new_new_n51754__ & ys__n44971;
  assign new_new_n51883__ = ~new_new_n51880__ & ~new_new_n51882__;
  assign new_new_n51884__ = ~new_new_n51879__ & new_new_n51883__;
  assign new_new_n51885__ = new_new_n51757__ & ys__n44971;
  assign new_new_n51886__ = ys__n48262 & new_new_n51752__;
  assign ys__n44955 = ys__n352 & ys__n28018;
  assign new_new_n51888__ = new_new_n51760__ & ys__n44955;
  assign new_new_n51889__ = ~new_new_n51886__ & ~new_new_n51888__;
  assign new_new_n51890__ = ~new_new_n51885__ & new_new_n51889__;
  assign new_new_n51891__ = new_new_n51884__ & new_new_n51890__;
  assign new_new_n51892__ = ~new_new_n51763__ & ~new_new_n51891__;
  assign new_new_n51893__ = ~new_new_n51810__ & new_new_n51892__;
  assign new_new_n51894__ = new_new_n51892__ & ~new_new_n51893__;
  assign new_new_n51895__ = ys__n48263 & new_new_n51759__;
  assign new_new_n51896__ = ys__n48263 & new_new_n51753__;
  assign ys__n44972 = ys__n352 & ys__n27863;
  assign new_new_n51898__ = new_new_n51754__ & ys__n44972;
  assign new_new_n51899__ = ~new_new_n51896__ & ~new_new_n51898__;
  assign new_new_n51900__ = ~new_new_n51895__ & new_new_n51899__;
  assign new_new_n51901__ = new_new_n51757__ & ys__n44972;
  assign new_new_n51902__ = ys__n48263 & new_new_n51752__;
  assign ys__n44956 = ys__n352 & ys__n28019;
  assign new_new_n51904__ = new_new_n51760__ & ys__n44956;
  assign new_new_n51905__ = ~new_new_n51902__ & ~new_new_n51904__;
  assign new_new_n51906__ = ~new_new_n51901__ & new_new_n51905__;
  assign new_new_n51907__ = new_new_n51900__ & new_new_n51906__;
  assign new_new_n51908__ = ~new_new_n51763__ & ~new_new_n51907__;
  assign new_new_n51909__ = ~new_new_n51894__ & ~new_new_n51908__;
  assign new_new_n51910__ = ys__n48264 & new_new_n51759__;
  assign new_new_n51911__ = ys__n48264 & new_new_n51753__;
  assign ys__n44973 = ys__n352 & ys__n27865;
  assign new_new_n51913__ = new_new_n51754__ & ys__n44973;
  assign new_new_n51914__ = ~new_new_n51911__ & ~new_new_n51913__;
  assign new_new_n51915__ = ~new_new_n51910__ & new_new_n51914__;
  assign new_new_n51916__ = new_new_n51757__ & ys__n44973;
  assign new_new_n51917__ = ys__n48264 & new_new_n51752__;
  assign ys__n44957 = ys__n352 & ys__n28020;
  assign new_new_n51919__ = new_new_n51760__ & ys__n44957;
  assign new_new_n51920__ = ~new_new_n51917__ & ~new_new_n51919__;
  assign new_new_n51921__ = ~new_new_n51916__ & new_new_n51920__;
  assign new_new_n51922__ = new_new_n51915__ & new_new_n51921__;
  assign new_new_n51923__ = ~new_new_n51763__ & ~new_new_n51922__;
  assign new_new_n51924__ = new_new_n51909__ & ~new_new_n51923__;
  assign new_new_n51925__ = ~new_new_n51810__ & ~new_new_n51892__;
  assign new_new_n51926__ = new_new_n51908__ & new_new_n51925__;
  assign new_new_n51927__ = new_new_n51908__ & ~new_new_n51926__;
  assign new_new_n51928__ = new_new_n51923__ & ~new_new_n51927__;
  assign new_new_n51929__ = ~new_new_n51924__ & ~new_new_n51928__;
  assign new_new_n51930__ = ~new_new_n51839__ & new_new_n51929__;
  assign new_new_n51931__ = new_new_n51839__ & ~new_new_n51929__;
  assign ys__n39399 = new_new_n51930__ | new_new_n51931__;
  assign new_new_n51933__ = new_new_n51810__ & new_new_n51892__;
  assign new_new_n51934__ = ~new_new_n51908__ & new_new_n51933__;
  assign new_new_n51935__ = ~new_new_n51926__ & ~new_new_n51934__;
  assign new_new_n51936__ = ~new_new_n51923__ & ~new_new_n51935__;
  assign new_new_n51937__ = new_new_n51810__ & ~new_new_n51892__;
  assign new_new_n51938__ = ~new_new_n51892__ & ~new_new_n51937__;
  assign new_new_n51939__ = new_new_n51908__ & ~new_new_n51938__;
  assign new_new_n51940__ = ~new_new_n51909__ & ~new_new_n51939__;
  assign new_new_n51941__ = new_new_n51923__ & ~new_new_n51940__;
  assign new_new_n51942__ = ~new_new_n51936__ & ~new_new_n51941__;
  assign new_new_n51943__ = ~new_new_n51839__ & new_new_n51942__;
  assign new_new_n51944__ = new_new_n51839__ & ~new_new_n51942__;
  assign ys__n39400 = new_new_n51943__ | new_new_n51944__;
  assign new_new_n51946__ = ~new_new_n51908__ & new_new_n51925__;
  assign new_new_n51947__ = ~new_new_n51893__ & ~new_new_n51937__;
  assign new_new_n51948__ = new_new_n51908__ & ~new_new_n51947__;
  assign new_new_n51949__ = ~new_new_n51946__ & ~new_new_n51948__;
  assign new_new_n51950__ = ~new_new_n51923__ & ~new_new_n51949__;
  assign new_new_n51951__ = ~new_new_n51925__ & ~new_new_n51933__;
  assign new_new_n51952__ = ~new_new_n51908__ & ~new_new_n51951__;
  assign new_new_n51953__ = ~new_new_n51894__ & new_new_n51908__;
  assign new_new_n51954__ = ~new_new_n51952__ & ~new_new_n51953__;
  assign new_new_n51955__ = new_new_n51923__ & ~new_new_n51954__;
  assign new_new_n51956__ = ~new_new_n51950__ & ~new_new_n51955__;
  assign new_new_n51957__ = ~new_new_n51839__ & new_new_n51956__;
  assign new_new_n51958__ = new_new_n51839__ & ~new_new_n51956__;
  assign ys__n39401 = new_new_n51957__ | new_new_n51958__;
  assign new_new_n51960__ = new_new_n51908__ & ~new_new_n51923__;
  assign new_new_n51961__ = new_new_n51933__ & new_new_n51960__;
  assign new_new_n51962__ = ~new_new_n51908__ & ~new_new_n51938__;
  assign new_new_n51963__ = ~new_new_n51908__ & ~new_new_n51962__;
  assign new_new_n51964__ = new_new_n51923__ & ~new_new_n51963__;
  assign new_new_n51965__ = ~new_new_n51961__ & ~new_new_n51964__;
  assign new_new_n51966__ = ~new_new_n51839__ & new_new_n51965__;
  assign new_new_n51967__ = new_new_n51839__ & ~new_new_n51965__;
  assign ys__n39402 = new_new_n51966__ | new_new_n51967__;
  assign new_new_n51969__ = ys__n48265 & new_new_n51759__;
  assign new_new_n51970__ = ys__n48265 & new_new_n51753__;
  assign ys__n44974 = ys__n352 & ys__n27867;
  assign new_new_n51972__ = new_new_n51754__ & ys__n44974;
  assign new_new_n51973__ = ~new_new_n51970__ & ~new_new_n51972__;
  assign new_new_n51974__ = ~new_new_n51969__ & new_new_n51973__;
  assign new_new_n51975__ = new_new_n51757__ & ys__n44974;
  assign new_new_n51976__ = ys__n48265 & new_new_n51752__;
  assign ys__n44958 = ys__n352 & ys__n28021;
  assign new_new_n51978__ = new_new_n51760__ & ys__n44958;
  assign new_new_n51979__ = ~new_new_n51976__ & ~new_new_n51978__;
  assign new_new_n51980__ = ~new_new_n51975__ & new_new_n51979__;
  assign new_new_n51981__ = new_new_n51974__ & new_new_n51980__;
  assign new_new_n51982__ = ~new_new_n51763__ & ~new_new_n51981__;
  assign new_new_n51983__ = ~new_new_n51923__ & new_new_n51982__;
  assign new_new_n51984__ = new_new_n51982__ & ~new_new_n51983__;
  assign new_new_n51985__ = ys__n48266 & new_new_n51759__;
  assign new_new_n51986__ = ys__n48266 & new_new_n51753__;
  assign ys__n44975 = ys__n352 & ys__n27869;
  assign new_new_n51988__ = new_new_n51754__ & ys__n44975;
  assign new_new_n51989__ = ~new_new_n51986__ & ~new_new_n51988__;
  assign new_new_n51990__ = ~new_new_n51985__ & new_new_n51989__;
  assign new_new_n51991__ = new_new_n51757__ & ys__n44975;
  assign new_new_n51992__ = ys__n48266 & new_new_n51752__;
  assign ys__n44959 = ys__n352 & ys__n28022;
  assign new_new_n51994__ = new_new_n51760__ & ys__n44959;
  assign new_new_n51995__ = ~new_new_n51992__ & ~new_new_n51994__;
  assign new_new_n51996__ = ~new_new_n51991__ & new_new_n51995__;
  assign new_new_n51997__ = new_new_n51990__ & new_new_n51996__;
  assign new_new_n51998__ = ~new_new_n51763__ & ~new_new_n51997__;
  assign new_new_n51999__ = ~new_new_n51984__ & ~new_new_n51998__;
  assign new_new_n52000__ = ys__n48267 & new_new_n51759__;
  assign new_new_n52001__ = ys__n48267 & new_new_n51753__;
  assign ys__n44976 = ys__n352 & ys__n27871;
  assign new_new_n52003__ = new_new_n51754__ & ys__n44976;
  assign new_new_n52004__ = ~new_new_n52001__ & ~new_new_n52003__;
  assign new_new_n52005__ = ~new_new_n52000__ & new_new_n52004__;
  assign new_new_n52006__ = new_new_n51757__ & ys__n44976;
  assign new_new_n52007__ = ys__n48267 & new_new_n51752__;
  assign ys__n44960 = ys__n352 & ys__n28023;
  assign new_new_n52009__ = new_new_n51760__ & ys__n44960;
  assign new_new_n52010__ = ~new_new_n52007__ & ~new_new_n52009__;
  assign new_new_n52011__ = ~new_new_n52006__ & new_new_n52010__;
  assign new_new_n52012__ = new_new_n52005__ & new_new_n52011__;
  assign new_new_n52013__ = ~new_new_n51763__ & ~new_new_n52012__;
  assign new_new_n52014__ = new_new_n51999__ & ~new_new_n52013__;
  assign new_new_n52015__ = ~new_new_n51923__ & ~new_new_n51982__;
  assign new_new_n52016__ = new_new_n51998__ & new_new_n52015__;
  assign new_new_n52017__ = new_new_n51998__ & ~new_new_n52016__;
  assign new_new_n52018__ = new_new_n52013__ & ~new_new_n52017__;
  assign new_new_n52019__ = ~new_new_n52014__ & ~new_new_n52018__;
  assign new_new_n52020__ = ~new_new_n51839__ & new_new_n52019__;
  assign new_new_n52021__ = new_new_n51839__ & ~new_new_n52019__;
  assign ys__n39403 = new_new_n52020__ | new_new_n52021__;
  assign new_new_n52023__ = new_new_n51923__ & new_new_n51982__;
  assign new_new_n52024__ = ~new_new_n51998__ & new_new_n52023__;
  assign new_new_n52025__ = ~new_new_n52016__ & ~new_new_n52024__;
  assign new_new_n52026__ = ~new_new_n52013__ & ~new_new_n52025__;
  assign new_new_n52027__ = new_new_n51923__ & ~new_new_n51982__;
  assign new_new_n52028__ = ~new_new_n51982__ & ~new_new_n52027__;
  assign new_new_n52029__ = new_new_n51998__ & ~new_new_n52028__;
  assign new_new_n52030__ = ~new_new_n51999__ & ~new_new_n52029__;
  assign new_new_n52031__ = new_new_n52013__ & ~new_new_n52030__;
  assign new_new_n52032__ = ~new_new_n52026__ & ~new_new_n52031__;
  assign new_new_n52033__ = ~new_new_n51839__ & new_new_n52032__;
  assign new_new_n52034__ = new_new_n51839__ & ~new_new_n52032__;
  assign ys__n39404 = new_new_n52033__ | new_new_n52034__;
  assign new_new_n52036__ = ~new_new_n51998__ & new_new_n52015__;
  assign new_new_n52037__ = ~new_new_n51983__ & ~new_new_n52027__;
  assign new_new_n52038__ = new_new_n51998__ & ~new_new_n52037__;
  assign new_new_n52039__ = ~new_new_n52036__ & ~new_new_n52038__;
  assign new_new_n52040__ = ~new_new_n52013__ & ~new_new_n52039__;
  assign new_new_n52041__ = ~new_new_n52015__ & ~new_new_n52023__;
  assign new_new_n52042__ = ~new_new_n51998__ & ~new_new_n52041__;
  assign new_new_n52043__ = ~new_new_n51984__ & new_new_n51998__;
  assign new_new_n52044__ = ~new_new_n52042__ & ~new_new_n52043__;
  assign new_new_n52045__ = new_new_n52013__ & ~new_new_n52044__;
  assign new_new_n52046__ = ~new_new_n52040__ & ~new_new_n52045__;
  assign new_new_n52047__ = ~new_new_n51839__ & new_new_n52046__;
  assign new_new_n52048__ = new_new_n51839__ & ~new_new_n52046__;
  assign ys__n39405 = new_new_n52047__ | new_new_n52048__;
  assign new_new_n52050__ = new_new_n51998__ & ~new_new_n52013__;
  assign new_new_n52051__ = new_new_n52023__ & new_new_n52050__;
  assign new_new_n52052__ = ~new_new_n51998__ & ~new_new_n52028__;
  assign new_new_n52053__ = ~new_new_n51998__ & ~new_new_n52052__;
  assign new_new_n52054__ = new_new_n52013__ & ~new_new_n52053__;
  assign new_new_n52055__ = ~new_new_n52051__ & ~new_new_n52054__;
  assign new_new_n52056__ = ~new_new_n51839__ & new_new_n52055__;
  assign new_new_n52057__ = new_new_n51839__ & ~new_new_n52055__;
  assign ys__n39406 = new_new_n52056__ | new_new_n52057__;
  assign new_new_n52059__ = ys__n48268 & new_new_n51759__;
  assign new_new_n52060__ = ys__n48268 & new_new_n51753__;
  assign ys__n44977 = ys__n352 & ys__n27873;
  assign new_new_n52062__ = new_new_n51754__ & ys__n44977;
  assign new_new_n52063__ = ~new_new_n52060__ & ~new_new_n52062__;
  assign new_new_n52064__ = ~new_new_n52059__ & new_new_n52063__;
  assign new_new_n52065__ = new_new_n51757__ & ys__n44977;
  assign new_new_n52066__ = ys__n48268 & new_new_n51752__;
  assign ys__n44961 = ys__n352 & ys__n28024;
  assign new_new_n52068__ = new_new_n51760__ & ys__n44961;
  assign new_new_n52069__ = ~new_new_n52066__ & ~new_new_n52068__;
  assign new_new_n52070__ = ~new_new_n52065__ & new_new_n52069__;
  assign new_new_n52071__ = new_new_n52064__ & new_new_n52070__;
  assign new_new_n52072__ = ~new_new_n51763__ & ~new_new_n52071__;
  assign new_new_n52073__ = ~new_new_n52013__ & new_new_n52072__;
  assign new_new_n52074__ = new_new_n52072__ & ~new_new_n52073__;
  assign new_new_n52075__ = ys__n48269 & new_new_n51759__;
  assign new_new_n52076__ = ys__n48269 & new_new_n51753__;
  assign ys__n44978 = ys__n352 & ys__n27875;
  assign new_new_n52078__ = new_new_n51754__ & ys__n44978;
  assign new_new_n52079__ = ~new_new_n52076__ & ~new_new_n52078__;
  assign new_new_n52080__ = ~new_new_n52075__ & new_new_n52079__;
  assign new_new_n52081__ = new_new_n51757__ & ys__n44978;
  assign new_new_n52082__ = ys__n48269 & new_new_n51752__;
  assign ys__n44962 = ys__n352 & ys__n28025;
  assign new_new_n52084__ = new_new_n51760__ & ys__n44962;
  assign new_new_n52085__ = ~new_new_n52082__ & ~new_new_n52084__;
  assign new_new_n52086__ = ~new_new_n52081__ & new_new_n52085__;
  assign new_new_n52087__ = new_new_n52080__ & new_new_n52086__;
  assign new_new_n52088__ = ~new_new_n51763__ & ~new_new_n52087__;
  assign new_new_n52089__ = ~new_new_n52074__ & ~new_new_n52088__;
  assign new_new_n52090__ = ys__n48270 & new_new_n51759__;
  assign new_new_n52091__ = ys__n48270 & new_new_n51753__;
  assign ys__n44979 = ys__n352 & ys__n27877;
  assign new_new_n52093__ = new_new_n51754__ & ys__n44979;
  assign new_new_n52094__ = ~new_new_n52091__ & ~new_new_n52093__;
  assign new_new_n52095__ = ~new_new_n52090__ & new_new_n52094__;
  assign new_new_n52096__ = new_new_n51757__ & ys__n44979;
  assign new_new_n52097__ = ys__n48270 & new_new_n51752__;
  assign ys__n44963 = ys__n352 & ys__n28026;
  assign new_new_n52099__ = new_new_n51760__ & ys__n44963;
  assign new_new_n52100__ = ~new_new_n52097__ & ~new_new_n52099__;
  assign new_new_n52101__ = ~new_new_n52096__ & new_new_n52100__;
  assign new_new_n52102__ = new_new_n52095__ & new_new_n52101__;
  assign new_new_n52103__ = ~new_new_n51763__ & ~new_new_n52102__;
  assign new_new_n52104__ = new_new_n52089__ & ~new_new_n52103__;
  assign new_new_n52105__ = ~new_new_n52013__ & ~new_new_n52072__;
  assign new_new_n52106__ = new_new_n52088__ & new_new_n52105__;
  assign new_new_n52107__ = new_new_n52088__ & ~new_new_n52106__;
  assign new_new_n52108__ = new_new_n52103__ & ~new_new_n52107__;
  assign new_new_n52109__ = ~new_new_n52104__ & ~new_new_n52108__;
  assign new_new_n52110__ = ~new_new_n51839__ & new_new_n52109__;
  assign new_new_n52111__ = new_new_n51839__ & ~new_new_n52109__;
  assign ys__n39407 = new_new_n52110__ | new_new_n52111__;
  assign new_new_n52113__ = new_new_n52013__ & new_new_n52072__;
  assign new_new_n52114__ = ~new_new_n52088__ & new_new_n52113__;
  assign new_new_n52115__ = ~new_new_n52106__ & ~new_new_n52114__;
  assign new_new_n52116__ = ~new_new_n52103__ & ~new_new_n52115__;
  assign new_new_n52117__ = new_new_n52013__ & ~new_new_n52072__;
  assign new_new_n52118__ = ~new_new_n52072__ & ~new_new_n52117__;
  assign new_new_n52119__ = new_new_n52088__ & ~new_new_n52118__;
  assign new_new_n52120__ = ~new_new_n52089__ & ~new_new_n52119__;
  assign new_new_n52121__ = new_new_n52103__ & ~new_new_n52120__;
  assign new_new_n52122__ = ~new_new_n52116__ & ~new_new_n52121__;
  assign new_new_n52123__ = ~new_new_n51839__ & new_new_n52122__;
  assign new_new_n52124__ = new_new_n51839__ & ~new_new_n52122__;
  assign ys__n39408 = new_new_n52123__ | new_new_n52124__;
  assign new_new_n52126__ = ~new_new_n52088__ & new_new_n52105__;
  assign new_new_n52127__ = ~new_new_n52073__ & ~new_new_n52117__;
  assign new_new_n52128__ = new_new_n52088__ & ~new_new_n52127__;
  assign new_new_n52129__ = ~new_new_n52126__ & ~new_new_n52128__;
  assign new_new_n52130__ = ~new_new_n52103__ & ~new_new_n52129__;
  assign new_new_n52131__ = ~new_new_n52105__ & ~new_new_n52113__;
  assign new_new_n52132__ = ~new_new_n52088__ & ~new_new_n52131__;
  assign new_new_n52133__ = ~new_new_n52074__ & new_new_n52088__;
  assign new_new_n52134__ = ~new_new_n52132__ & ~new_new_n52133__;
  assign new_new_n52135__ = new_new_n52103__ & ~new_new_n52134__;
  assign new_new_n52136__ = ~new_new_n52130__ & ~new_new_n52135__;
  assign new_new_n52137__ = ~new_new_n51839__ & new_new_n52136__;
  assign new_new_n52138__ = new_new_n51839__ & ~new_new_n52136__;
  assign ys__n39409 = new_new_n52137__ | new_new_n52138__;
  assign new_new_n52140__ = new_new_n52088__ & ~new_new_n52103__;
  assign new_new_n52141__ = new_new_n52113__ & new_new_n52140__;
  assign new_new_n52142__ = ~new_new_n52088__ & ~new_new_n52118__;
  assign new_new_n52143__ = ~new_new_n52088__ & ~new_new_n52142__;
  assign new_new_n52144__ = new_new_n52103__ & ~new_new_n52143__;
  assign new_new_n52145__ = ~new_new_n52141__ & ~new_new_n52144__;
  assign new_new_n52146__ = ~new_new_n51839__ & new_new_n52145__;
  assign new_new_n52147__ = new_new_n51839__ & ~new_new_n52145__;
  assign ys__n39410 = new_new_n52146__ | new_new_n52147__;
  assign new_new_n52149__ = ys__n48271 & new_new_n51759__;
  assign new_new_n52150__ = ys__n48271 & new_new_n51753__;
  assign ys__n44980 = ys__n352 & ys__n27879;
  assign new_new_n52152__ = new_new_n51754__ & ys__n44980;
  assign new_new_n52153__ = ~new_new_n52150__ & ~new_new_n52152__;
  assign new_new_n52154__ = ~new_new_n52149__ & new_new_n52153__;
  assign new_new_n52155__ = new_new_n51757__ & ys__n44980;
  assign new_new_n52156__ = ys__n48271 & new_new_n51752__;
  assign ys__n44964 = ys__n352 & ys__n28027;
  assign new_new_n52158__ = new_new_n51760__ & ys__n44964;
  assign new_new_n52159__ = ~new_new_n52156__ & ~new_new_n52158__;
  assign new_new_n52160__ = ~new_new_n52155__ & new_new_n52159__;
  assign new_new_n52161__ = new_new_n52154__ & new_new_n52160__;
  assign new_new_n52162__ = ~new_new_n51763__ & ~new_new_n52161__;
  assign new_new_n52163__ = ~new_new_n52103__ & new_new_n52162__;
  assign new_new_n52164__ = new_new_n52162__ & ~new_new_n52163__;
  assign new_new_n52165__ = ys__n48272 & new_new_n51759__;
  assign new_new_n52166__ = ys__n48272 & new_new_n51753__;
  assign ys__n44981 = ys__n352 & ys__n27881;
  assign new_new_n52168__ = new_new_n51754__ & ys__n44981;
  assign new_new_n52169__ = ~new_new_n52166__ & ~new_new_n52168__;
  assign new_new_n52170__ = ~new_new_n52165__ & new_new_n52169__;
  assign new_new_n52171__ = new_new_n51757__ & ys__n44981;
  assign new_new_n52172__ = ys__n48272 & new_new_n51752__;
  assign ys__n44965 = ys__n352 & ys__n28028;
  assign new_new_n52174__ = new_new_n51760__ & ys__n44965;
  assign new_new_n52175__ = ~new_new_n52172__ & ~new_new_n52174__;
  assign new_new_n52176__ = ~new_new_n52171__ & new_new_n52175__;
  assign new_new_n52177__ = new_new_n52170__ & new_new_n52176__;
  assign new_new_n52178__ = ~new_new_n51763__ & ~new_new_n52177__;
  assign new_new_n52179__ = ~new_new_n52164__ & ~new_new_n52178__;
  assign new_new_n52180__ = ys__n48273 & new_new_n51759__;
  assign new_new_n52181__ = ys__n48273 & new_new_n51753__;
  assign ys__n44982 = ys__n352 & ys__n27883;
  assign new_new_n52183__ = new_new_n51754__ & ys__n44982;
  assign new_new_n52184__ = ~new_new_n52181__ & ~new_new_n52183__;
  assign new_new_n52185__ = ~new_new_n52180__ & new_new_n52184__;
  assign new_new_n52186__ = new_new_n51757__ & ys__n44982;
  assign new_new_n52187__ = ys__n48273 & new_new_n51752__;
  assign ys__n44966 = ys__n352 & ys__n28029;
  assign new_new_n52189__ = new_new_n51760__ & ys__n44966;
  assign new_new_n52190__ = ~new_new_n52187__ & ~new_new_n52189__;
  assign new_new_n52191__ = ~new_new_n52186__ & new_new_n52190__;
  assign new_new_n52192__ = new_new_n52185__ & new_new_n52191__;
  assign new_new_n52193__ = ~new_new_n51763__ & ~new_new_n52192__;
  assign new_new_n52194__ = new_new_n52179__ & ~new_new_n52193__;
  assign new_new_n52195__ = ~new_new_n52103__ & ~new_new_n52162__;
  assign new_new_n52196__ = new_new_n52178__ & new_new_n52195__;
  assign new_new_n52197__ = new_new_n52178__ & ~new_new_n52196__;
  assign new_new_n52198__ = new_new_n52193__ & ~new_new_n52197__;
  assign new_new_n52199__ = ~new_new_n52194__ & ~new_new_n52198__;
  assign new_new_n52200__ = ~new_new_n51839__ & new_new_n52199__;
  assign new_new_n52201__ = new_new_n51839__ & ~new_new_n52199__;
  assign ys__n39411 = new_new_n52200__ | new_new_n52201__;
  assign new_new_n52203__ = new_new_n52103__ & new_new_n52162__;
  assign new_new_n52204__ = ~new_new_n52178__ & new_new_n52203__;
  assign new_new_n52205__ = ~new_new_n52196__ & ~new_new_n52204__;
  assign new_new_n52206__ = ~new_new_n52193__ & ~new_new_n52205__;
  assign new_new_n52207__ = new_new_n52103__ & ~new_new_n52162__;
  assign new_new_n52208__ = ~new_new_n52162__ & ~new_new_n52207__;
  assign new_new_n52209__ = new_new_n52178__ & ~new_new_n52208__;
  assign new_new_n52210__ = ~new_new_n52179__ & ~new_new_n52209__;
  assign new_new_n52211__ = new_new_n52193__ & ~new_new_n52210__;
  assign new_new_n52212__ = ~new_new_n52206__ & ~new_new_n52211__;
  assign new_new_n52213__ = ~new_new_n51839__ & new_new_n52212__;
  assign new_new_n52214__ = new_new_n51839__ & ~new_new_n52212__;
  assign ys__n39412 = new_new_n52213__ | new_new_n52214__;
  assign new_new_n52216__ = ~new_new_n52178__ & new_new_n52195__;
  assign new_new_n52217__ = ~new_new_n52163__ & ~new_new_n52207__;
  assign new_new_n52218__ = new_new_n52178__ & ~new_new_n52217__;
  assign new_new_n52219__ = ~new_new_n52216__ & ~new_new_n52218__;
  assign new_new_n52220__ = ~new_new_n52193__ & ~new_new_n52219__;
  assign new_new_n52221__ = ~new_new_n52195__ & ~new_new_n52203__;
  assign new_new_n52222__ = ~new_new_n52178__ & ~new_new_n52221__;
  assign new_new_n52223__ = ~new_new_n52164__ & new_new_n52178__;
  assign new_new_n52224__ = ~new_new_n52222__ & ~new_new_n52223__;
  assign new_new_n52225__ = new_new_n52193__ & ~new_new_n52224__;
  assign new_new_n52226__ = ~new_new_n52220__ & ~new_new_n52225__;
  assign new_new_n52227__ = ~new_new_n51839__ & new_new_n52226__;
  assign new_new_n52228__ = new_new_n51839__ & ~new_new_n52226__;
  assign ys__n39413 = new_new_n52227__ | new_new_n52228__;
  assign new_new_n52230__ = new_new_n52178__ & ~new_new_n52193__;
  assign new_new_n52231__ = new_new_n52203__ & new_new_n52230__;
  assign new_new_n52232__ = ~new_new_n52178__ & ~new_new_n52208__;
  assign new_new_n52233__ = ~new_new_n52178__ & ~new_new_n52232__;
  assign new_new_n52234__ = new_new_n52193__ & ~new_new_n52233__;
  assign new_new_n52235__ = ~new_new_n52231__ & ~new_new_n52234__;
  assign new_new_n52236__ = ~new_new_n51839__ & new_new_n52235__;
  assign new_new_n52237__ = new_new_n51839__ & ~new_new_n52235__;
  assign ys__n39414 = new_new_n52236__ | new_new_n52237__;
  assign ys__n44983 = ys__n352 & ys__n27885;
  assign new_new_n52240__ = new_new_n51754__ & ys__n44983;
  assign new_new_n52241__ = ys__n48274 & new_new_n51759__;
  assign new_new_n52242__ = ys__n48274 & new_new_n51752__;
  assign new_new_n52243__ = ~new_new_n52241__ & ~new_new_n52242__;
  assign new_new_n52244__ = ~new_new_n52240__ & new_new_n52243__;
  assign new_new_n52245__ = ~new_new_n51763__ & ~new_new_n52244__;
  assign new_new_n52246__ = new_new_n51757__ & ys__n44983;
  assign ys__n44967 = ys__n352 & ys__n28030;
  assign new_new_n52248__ = new_new_n51760__ & ys__n44967;
  assign new_new_n52249__ = ys__n48274 & new_new_n51753__;
  assign new_new_n52250__ = ~new_new_n52240__ & ~new_new_n52249__;
  assign new_new_n52251__ = ~new_new_n52248__ & new_new_n52250__;
  assign new_new_n52252__ = ~new_new_n52246__ & new_new_n52251__;
  assign new_new_n52253__ = new_new_n52243__ & new_new_n52252__;
  assign new_new_n52254__ = ~new_new_n51763__ & ~new_new_n52253__;
  assign new_new_n52255__ = ~new_new_n52193__ & new_new_n52254__;
  assign new_new_n52256__ = new_new_n52254__ & ~new_new_n52255__;
  assign new_new_n52257__ = ~new_new_n52245__ & ~new_new_n52256__;
  assign new_new_n52258__ = ~new_new_n52245__ & new_new_n52257__;
  assign new_new_n52259__ = ~new_new_n52193__ & ~new_new_n52254__;
  assign new_new_n52260__ = new_new_n52245__ & new_new_n52259__;
  assign new_new_n52261__ = new_new_n52245__ & ~new_new_n52260__;
  assign new_new_n52262__ = new_new_n52245__ & ~new_new_n52261__;
  assign new_new_n52263__ = ~new_new_n52258__ & ~new_new_n52262__;
  assign new_new_n52264__ = ~new_new_n51839__ & new_new_n52263__;
  assign new_new_n52265__ = new_new_n51839__ & ~new_new_n52263__;
  assign ys__n39415 = new_new_n52264__ | new_new_n52265__;
  assign new_new_n52267__ = new_new_n52193__ & new_new_n52254__;
  assign new_new_n52268__ = ~new_new_n52245__ & new_new_n52267__;
  assign new_new_n52269__ = ~new_new_n52260__ & ~new_new_n52268__;
  assign new_new_n52270__ = ~new_new_n52245__ & ~new_new_n52269__;
  assign new_new_n52271__ = new_new_n52193__ & ~new_new_n52254__;
  assign new_new_n52272__ = ~new_new_n52254__ & ~new_new_n52271__;
  assign new_new_n52273__ = new_new_n52245__ & ~new_new_n52272__;
  assign new_new_n52274__ = ~new_new_n52257__ & ~new_new_n52273__;
  assign new_new_n52275__ = new_new_n52245__ & ~new_new_n52274__;
  assign new_new_n52276__ = ~new_new_n52270__ & ~new_new_n52275__;
  assign new_new_n52277__ = ~new_new_n51839__ & new_new_n52276__;
  assign new_new_n52278__ = new_new_n51839__ & ~new_new_n52276__;
  assign ys__n39416 = new_new_n52277__ | new_new_n52278__;
  assign new_new_n52280__ = ~new_new_n52245__ & new_new_n52259__;
  assign new_new_n52281__ = ~new_new_n52255__ & ~new_new_n52271__;
  assign new_new_n52282__ = new_new_n52245__ & ~new_new_n52281__;
  assign new_new_n52283__ = ~new_new_n52280__ & ~new_new_n52282__;
  assign new_new_n52284__ = ~new_new_n52245__ & ~new_new_n52283__;
  assign new_new_n52285__ = ~new_new_n52259__ & ~new_new_n52267__;
  assign new_new_n52286__ = ~new_new_n52245__ & ~new_new_n52285__;
  assign new_new_n52287__ = new_new_n52245__ & ~new_new_n52256__;
  assign new_new_n52288__ = ~new_new_n52286__ & ~new_new_n52287__;
  assign new_new_n52289__ = new_new_n52245__ & ~new_new_n52288__;
  assign new_new_n52290__ = ~new_new_n52284__ & ~new_new_n52289__;
  assign new_new_n52291__ = ~new_new_n51839__ & new_new_n52290__;
  assign new_new_n52292__ = new_new_n51839__ & ~new_new_n52290__;
  assign ys__n39417 = new_new_n52291__ | new_new_n52292__;
  assign new_new_n52294__ = ~new_new_n52245__ & ~new_new_n52272__;
  assign new_new_n52295__ = ~new_new_n52245__ & ~new_new_n52294__;
  assign new_new_n52296__ = new_new_n52245__ & ~new_new_n52295__;
  assign new_new_n52297__ = ~new_new_n51839__ & ~new_new_n52296__;
  assign new_new_n52298__ = new_new_n51839__ & new_new_n52296__;
  assign ys__n39418 = new_new_n52297__ | new_new_n52298__;
  assign new_new_n52300__ = ys__n33634 & ys__n33636;
  assign new_new_n52301__ = ys__n33632 & new_new_n52300__;
  assign new_new_n52302__ = ys__n39718 & new_new_n52301__;
  assign new_new_n52303__ = ys__n33632 & ys__n33636;
  assign new_new_n52304__ = ys__n33638 & new_new_n52303__;
  assign new_new_n52305__ = ys__n24741 & new_new_n52304__;
  assign new_new_n52306__ = ~new_new_n52302__ & ~new_new_n52305__;
  assign new_new_n52307__ = ~ys__n33632 & ~ys__n33634;
  assign new_new_n52308__ = ~ys__n33638 & new_new_n52307__;
  assign new_new_n52309__ = ys__n33683 & new_new_n52308__;
  assign new_new_n52310__ = ys__n33632 & ys__n33634;
  assign new_new_n52311__ = ys__n33638 & new_new_n52310__;
  assign new_new_n52312__ = ~ys__n33683 & new_new_n52311__;
  assign new_new_n52313__ = ~new_new_n52309__ & ~new_new_n52312__;
  assign new_new_n52314__ = new_new_n52306__ & new_new_n52313__;
  assign new_new_n52315__ = ~ys__n33634 & ~ys__n33636;
  assign new_new_n52316__ = ~ys__n33638 & new_new_n52315__;
  assign new_new_n52317__ = ys__n24747 & new_new_n52316__;
  assign new_new_n52318__ = ~ys__n33632 & new_new_n52315__;
  assign new_new_n52319__ = ys__n24744 & new_new_n52318__;
  assign new_new_n52320__ = ~new_new_n52317__ & ~new_new_n52319__;
  assign new_new_n52321__ = ~ys__n33632 & ~ys__n33636;
  assign new_new_n52322__ = ~ys__n33638 & new_new_n52321__;
  assign new_new_n52323__ = ys__n24741 & new_new_n52322__;
  assign new_new_n52324__ = ys__n33638 & new_new_n52300__;
  assign new_new_n52325__ = ys__n39720 & new_new_n52324__;
  assign new_new_n52326__ = ~new_new_n52323__ & ~new_new_n52325__;
  assign new_new_n52327__ = new_new_n52320__ & new_new_n52326__;
  assign ys__n40052 = ~new_new_n52314__ | ~new_new_n52327__;
  assign ys__n42129 = new_new_n25452__ & new_new_n25490__;
  assign new_new_n52330__ = ys__n33658 & ys__n33660;
  assign new_new_n52331__ = ys__n33662 & new_new_n52330__;
  assign new_new_n52332__ = ys__n33656 & ys__n33660;
  assign new_new_n52333__ = ys__n33662 & new_new_n52332__;
  assign new_new_n52334__ = ys__n33656 & new_new_n52330__;
  assign new_new_n52335__ = ~new_new_n52333__ & ~new_new_n52334__;
  assign new_new_n52336__ = ~new_new_n52331__ & new_new_n52335__;
  assign new_new_n52337__ = ys__n39520 & ~new_new_n52336__;
  assign new_new_n52338__ = ~ys__n33658 & ~ys__n33660;
  assign new_new_n52339__ = ~ys__n33662 & new_new_n52338__;
  assign new_new_n52340__ = ~ys__n33656 & ~ys__n33660;
  assign new_new_n52341__ = ~ys__n33662 & new_new_n52340__;
  assign new_new_n52342__ = ~ys__n33656 & new_new_n52338__;
  assign new_new_n52343__ = ~new_new_n52341__ & ~new_new_n52342__;
  assign new_new_n52344__ = ~new_new_n52339__ & new_new_n52343__;
  assign new_new_n52345__ = ys__n39518 & ~new_new_n52344__;
  assign new_new_n52346__ = ~ys__n33656 & ~ys__n33658;
  assign new_new_n52347__ = ~ys__n33662 & new_new_n52346__;
  assign new_new_n52348__ = ys__n33747 & new_new_n52347__;
  assign new_new_n52349__ = ys__n33656 & ys__n33658;
  assign new_new_n52350__ = ys__n33662 & new_new_n52349__;
  assign new_new_n52351__ = ~ys__n33747 & new_new_n52350__;
  assign new_new_n52352__ = ~new_new_n52348__ & ~new_new_n52351__;
  assign new_new_n52353__ = ~new_new_n52345__ & new_new_n52352__;
  assign new_new_n52354__ = ~new_new_n52337__ & new_new_n52353__;
  assign new_new_n52355__ = ys__n33666 & ys__n33668;
  assign new_new_n52356__ = ys__n33670 & new_new_n52355__;
  assign new_new_n52357__ = ys__n33664 & ys__n33668;
  assign new_new_n52358__ = ys__n33670 & new_new_n52357__;
  assign new_new_n52359__ = ys__n33664 & new_new_n52355__;
  assign new_new_n52360__ = ~new_new_n52358__ & ~new_new_n52359__;
  assign new_new_n52361__ = ~new_new_n52356__ & new_new_n52360__;
  assign new_new_n52362__ = ys__n39520 & ~new_new_n52361__;
  assign new_new_n52363__ = ~ys__n33666 & ~ys__n33668;
  assign new_new_n52364__ = ~ys__n33670 & new_new_n52363__;
  assign new_new_n52365__ = ~ys__n33664 & ~ys__n33668;
  assign new_new_n52366__ = ~ys__n33670 & new_new_n52365__;
  assign new_new_n52367__ = ~ys__n33664 & new_new_n52363__;
  assign new_new_n52368__ = ~new_new_n52366__ & ~new_new_n52367__;
  assign new_new_n52369__ = ~new_new_n52364__ & new_new_n52368__;
  assign new_new_n52370__ = ys__n39518 & ~new_new_n52369__;
  assign new_new_n52371__ = ~ys__n33664 & ~ys__n33666;
  assign new_new_n52372__ = ~ys__n33670 & new_new_n52371__;
  assign new_new_n52373__ = ys__n33747 & new_new_n52372__;
  assign new_new_n52374__ = ys__n33664 & ys__n33666;
  assign new_new_n52375__ = ys__n33670 & new_new_n52374__;
  assign new_new_n52376__ = ~ys__n33747 & new_new_n52375__;
  assign new_new_n52377__ = ~new_new_n52373__ & ~new_new_n52376__;
  assign new_new_n52378__ = ~new_new_n52370__ & new_new_n52377__;
  assign new_new_n52379__ = ~new_new_n52362__ & new_new_n52378__;
  assign new_new_n52380__ = ~ys__n33672 & ~ys__n33676;
  assign new_new_n52381__ = ~ys__n33678 & new_new_n52380__;
  assign new_new_n52382__ = ~ys__n33674 & ~ys__n33676;
  assign new_new_n52383__ = ~ys__n33678 & new_new_n52382__;
  assign new_new_n52384__ = ~ys__n33672 & new_new_n52382__;
  assign new_new_n52385__ = ~new_new_n52383__ & ~new_new_n52384__;
  assign new_new_n52386__ = ~new_new_n52381__ & new_new_n52385__;
  assign new_new_n52387__ = ys__n39518 & ~new_new_n52386__;
  assign new_new_n52388__ = ys__n33672 & ys__n33676;
  assign new_new_n52389__ = ys__n33678 & new_new_n52388__;
  assign new_new_n52390__ = ys__n33674 & ys__n33676;
  assign new_new_n52391__ = ys__n33678 & new_new_n52390__;
  assign new_new_n52392__ = ys__n33672 & new_new_n52390__;
  assign new_new_n52393__ = ~new_new_n52391__ & ~new_new_n52392__;
  assign new_new_n52394__ = ~new_new_n52389__ & new_new_n52393__;
  assign new_new_n52395__ = ys__n39520 & ~new_new_n52394__;
  assign new_new_n52396__ = ~new_new_n52387__ & ~new_new_n52395__;
  assign new_new_n52397__ = ~new_new_n52379__ & ~new_new_n52396__;
  assign new_new_n52398__ = ~new_new_n52354__ & new_new_n52397__;
  assign new_new_n52399__ = new_new_n52379__ & new_new_n52396__;
  assign new_new_n52400__ = ~new_new_n52354__ & new_new_n52399__;
  assign new_new_n52401__ = ~new_new_n52398__ & ~new_new_n52400__;
  assign new_new_n52402__ = ~new_new_n52379__ & new_new_n52396__;
  assign new_new_n52403__ = new_new_n52354__ & new_new_n52402__;
  assign new_new_n52404__ = new_new_n52379__ & ~new_new_n52396__;
  assign new_new_n52405__ = new_new_n52354__ & new_new_n52404__;
  assign new_new_n52406__ = ~new_new_n52403__ & ~new_new_n52405__;
  assign new_new_n52407__ = new_new_n52401__ & new_new_n52406__;
  assign new_new_n52408__ = ys__n33642 & ys__n33644;
  assign new_new_n52409__ = ys__n33646 & new_new_n52408__;
  assign new_new_n52410__ = ys__n33640 & ys__n33644;
  assign new_new_n52411__ = ys__n33646 & new_new_n52410__;
  assign new_new_n52412__ = ys__n33640 & new_new_n52408__;
  assign new_new_n52413__ = ~new_new_n52411__ & ~new_new_n52412__;
  assign new_new_n52414__ = ~new_new_n52409__ & new_new_n52413__;
  assign new_new_n52415__ = ys__n39520 & ~new_new_n52414__;
  assign new_new_n52416__ = ~ys__n33642 & ~ys__n33644;
  assign new_new_n52417__ = ~ys__n33646 & new_new_n52416__;
  assign new_new_n52418__ = ~ys__n33640 & ~ys__n33644;
  assign new_new_n52419__ = ~ys__n33646 & new_new_n52418__;
  assign new_new_n52420__ = ~ys__n33640 & new_new_n52416__;
  assign new_new_n52421__ = ~new_new_n52419__ & ~new_new_n52420__;
  assign new_new_n52422__ = ~new_new_n52417__ & new_new_n52421__;
  assign new_new_n52423__ = ys__n39518 & ~new_new_n52422__;
  assign new_new_n52424__ = ~ys__n33640 & ~ys__n33642;
  assign new_new_n52425__ = ~ys__n33646 & new_new_n52424__;
  assign new_new_n52426__ = ys__n33747 & new_new_n52425__;
  assign new_new_n52427__ = ys__n33640 & ys__n33642;
  assign new_new_n52428__ = ys__n33646 & new_new_n52427__;
  assign new_new_n52429__ = ~ys__n33747 & new_new_n52428__;
  assign new_new_n52430__ = ~new_new_n52426__ & ~new_new_n52429__;
  assign new_new_n52431__ = ~new_new_n52423__ & new_new_n52430__;
  assign new_new_n52432__ = ~new_new_n52415__ & new_new_n52431__;
  assign new_new_n52433__ = ~new_new_n52301__ & ~new_new_n52324__;
  assign new_new_n52434__ = ~new_new_n52304__ & new_new_n52433__;
  assign new_new_n52435__ = ys__n39520 & ~new_new_n52434__;
  assign new_new_n52436__ = ~new_new_n52316__ & ~new_new_n52318__;
  assign new_new_n52437__ = ~new_new_n52322__ & new_new_n52436__;
  assign new_new_n52438__ = ys__n39518 & ~new_new_n52437__;
  assign new_new_n52439__ = ys__n33747 & new_new_n52308__;
  assign new_new_n52440__ = ~ys__n33747 & new_new_n52311__;
  assign new_new_n52441__ = ~new_new_n52439__ & ~new_new_n52440__;
  assign new_new_n52442__ = ~new_new_n52438__ & new_new_n52441__;
  assign new_new_n52443__ = ~new_new_n52435__ & new_new_n52442__;
  assign new_new_n52444__ = ~new_new_n52432__ & ~new_new_n52443__;
  assign new_new_n52445__ = ys__n33650 & ys__n33652;
  assign new_new_n52446__ = ys__n33654 & new_new_n52445__;
  assign new_new_n52447__ = ys__n33648 & ys__n33652;
  assign new_new_n52448__ = ys__n33654 & new_new_n52447__;
  assign new_new_n52449__ = ys__n33648 & new_new_n52445__;
  assign new_new_n52450__ = ~new_new_n52448__ & ~new_new_n52449__;
  assign new_new_n52451__ = ~new_new_n52446__ & new_new_n52450__;
  assign new_new_n52452__ = ys__n39520 & ~new_new_n52451__;
  assign new_new_n52453__ = ~ys__n33650 & ~ys__n33652;
  assign new_new_n52454__ = ~ys__n33654 & new_new_n52453__;
  assign new_new_n52455__ = ~ys__n33648 & ~ys__n33652;
  assign new_new_n52456__ = ~ys__n33654 & new_new_n52455__;
  assign new_new_n52457__ = ~ys__n33648 & new_new_n52453__;
  assign new_new_n52458__ = ~new_new_n52456__ & ~new_new_n52457__;
  assign new_new_n52459__ = ~new_new_n52454__ & new_new_n52458__;
  assign new_new_n52460__ = ys__n39518 & ~new_new_n52459__;
  assign new_new_n52461__ = ~ys__n33648 & ~ys__n33650;
  assign new_new_n52462__ = ~ys__n33654 & new_new_n52461__;
  assign new_new_n52463__ = ys__n33747 & new_new_n52462__;
  assign new_new_n52464__ = ys__n33648 & ys__n33650;
  assign new_new_n52465__ = ys__n33654 & new_new_n52464__;
  assign new_new_n52466__ = ~ys__n33747 & new_new_n52465__;
  assign new_new_n52467__ = ~new_new_n52463__ & ~new_new_n52466__;
  assign new_new_n52468__ = ~new_new_n52460__ & new_new_n52467__;
  assign new_new_n52469__ = ~new_new_n52452__ & new_new_n52468__;
  assign new_new_n52470__ = ~new_new_n52432__ & ~new_new_n52469__;
  assign new_new_n52471__ = ~new_new_n52443__ & ~new_new_n52469__;
  assign new_new_n52472__ = ~new_new_n52470__ & ~new_new_n52471__;
  assign new_new_n52473__ = ~new_new_n52444__ & new_new_n52472__;
  assign new_new_n52474__ = ys__n39518 & new_new_n52383__;
  assign new_new_n52475__ = ys__n39520 & new_new_n52391__;
  assign new_new_n52476__ = ~new_new_n52474__ & ~new_new_n52475__;
  assign new_new_n52477__ = ys__n39518 & new_new_n52384__;
  assign new_new_n52478__ = ys__n39520 & new_new_n52392__;
  assign new_new_n52479__ = ~new_new_n52477__ & ~new_new_n52478__;
  assign new_new_n52480__ = new_new_n52476__ & new_new_n52479__;
  assign new_new_n52481__ = ~new_new_n52354__ & ~new_new_n52480__;
  assign new_new_n52482__ = ~new_new_n52354__ & ~new_new_n52379__;
  assign new_new_n52483__ = ~new_new_n52379__ & ~new_new_n52480__;
  assign new_new_n52484__ = ~new_new_n52482__ & ~new_new_n52483__;
  assign new_new_n52485__ = ~new_new_n52481__ & new_new_n52484__;
  assign new_new_n52486__ = ~new_new_n52473__ & ~new_new_n52485__;
  assign new_new_n52487__ = ~new_new_n52407__ & new_new_n52486__;
  assign new_new_n52488__ = ~new_new_n52473__ & new_new_n52485__;
  assign new_new_n52489__ = new_new_n52407__ & new_new_n52488__;
  assign new_new_n52490__ = ~new_new_n52487__ & ~new_new_n52489__;
  assign new_new_n52491__ = new_new_n52473__ & new_new_n52485__;
  assign new_new_n52492__ = ~new_new_n52407__ & new_new_n52491__;
  assign new_new_n52493__ = new_new_n52473__ & ~new_new_n52485__;
  assign new_new_n52494__ = new_new_n52407__ & new_new_n52493__;
  assign new_new_n52495__ = ~new_new_n52492__ & ~new_new_n52494__;
  assign new_new_n52496__ = new_new_n52490__ & new_new_n52495__;
  assign new_new_n52497__ = ~new_new_n52354__ & new_new_n52483__;
  assign new_new_n52498__ = new_new_n52379__ & new_new_n52480__;
  assign new_new_n52499__ = ~new_new_n52354__ & new_new_n52498__;
  assign new_new_n52500__ = ~new_new_n52497__ & ~new_new_n52499__;
  assign new_new_n52501__ = ~new_new_n52379__ & new_new_n52480__;
  assign new_new_n52502__ = new_new_n52354__ & new_new_n52501__;
  assign new_new_n52503__ = new_new_n52379__ & ~new_new_n52480__;
  assign new_new_n52504__ = new_new_n52354__ & new_new_n52503__;
  assign new_new_n52505__ = ~new_new_n52502__ & ~new_new_n52504__;
  assign new_new_n52506__ = new_new_n52500__ & new_new_n52505__;
  assign new_new_n52507__ = ~new_new_n52473__ & ~new_new_n52506__;
  assign new_new_n52508__ = ys__n24834 & new_new_n52384__;
  assign new_new_n52509__ = ~new_new_n52474__ & ~new_new_n52508__;
  assign new_new_n52510__ = ys__n39778 & new_new_n52392__;
  assign new_new_n52511__ = ~new_new_n52475__ & ~new_new_n52510__;
  assign new_new_n52512__ = new_new_n52509__ & new_new_n52511__;
  assign new_new_n52513__ = ~new_new_n52379__ & ~new_new_n52512__;
  assign new_new_n52514__ = ~new_new_n52354__ & ~new_new_n52512__;
  assign new_new_n52515__ = ~new_new_n52513__ & ~new_new_n52514__;
  assign new_new_n52516__ = ~new_new_n52482__ & new_new_n52515__;
  assign new_new_n52517__ = ~new_new_n52506__ & ~new_new_n52516__;
  assign new_new_n52518__ = ~new_new_n52473__ & ~new_new_n52516__;
  assign new_new_n52519__ = ~new_new_n52517__ & ~new_new_n52518__;
  assign new_new_n52520__ = ~new_new_n52507__ & new_new_n52519__;
  assign new_new_n52521__ = ~new_new_n52443__ & new_new_n52470__;
  assign new_new_n52522__ = new_new_n52432__ & new_new_n52469__;
  assign new_new_n52523__ = ~new_new_n52443__ & new_new_n52522__;
  assign new_new_n52524__ = ~new_new_n52521__ & ~new_new_n52523__;
  assign new_new_n52525__ = ~new_new_n52432__ & new_new_n52469__;
  assign new_new_n52526__ = new_new_n52443__ & new_new_n52525__;
  assign new_new_n52527__ = new_new_n52432__ & ~new_new_n52469__;
  assign new_new_n52528__ = new_new_n52443__ & new_new_n52527__;
  assign new_new_n52529__ = ~new_new_n52526__ & ~new_new_n52528__;
  assign new_new_n52530__ = new_new_n52524__ & new_new_n52529__;
  assign new_new_n52531__ = ~new_new_n52520__ & ~new_new_n52530__;
  assign new_new_n52532__ = ~new_new_n52496__ & new_new_n52531__;
  assign new_new_n52533__ = new_new_n52520__ & ~new_new_n52530__;
  assign new_new_n52534__ = new_new_n52496__ & new_new_n52533__;
  assign new_new_n52535__ = ~new_new_n52532__ & ~new_new_n52534__;
  assign new_new_n52536__ = new_new_n52520__ & new_new_n52530__;
  assign new_new_n52537__ = ~new_new_n52496__ & new_new_n52536__;
  assign new_new_n52538__ = ~new_new_n52520__ & new_new_n52530__;
  assign new_new_n52539__ = new_new_n52496__ & new_new_n52538__;
  assign new_new_n52540__ = ~new_new_n52537__ & ~new_new_n52539__;
  assign ys__n42153 = ~new_new_n52535__ | ~new_new_n52540__;
  assign new_new_n52542__ = ~new_new_n52473__ & new_new_n52517__;
  assign new_new_n52543__ = new_new_n52473__ & ~new_new_n52516__;
  assign new_new_n52544__ = new_new_n52506__ & new_new_n52543__;
  assign new_new_n52545__ = ~new_new_n52473__ & new_new_n52516__;
  assign new_new_n52546__ = new_new_n52506__ & new_new_n52545__;
  assign new_new_n52547__ = new_new_n52473__ & new_new_n52516__;
  assign new_new_n52548__ = ~new_new_n52506__ & new_new_n52547__;
  assign new_new_n52549__ = ~new_new_n52546__ & ~new_new_n52548__;
  assign new_new_n52550__ = ~new_new_n52544__ & new_new_n52549__;
  assign new_new_n52551__ = ~new_new_n52542__ & new_new_n52550__;
  assign new_new_n52552__ = ~new_new_n52530__ & ~new_new_n52551__;
  assign new_new_n52553__ = ~new_new_n52354__ & new_new_n52513__;
  assign new_new_n52554__ = new_new_n52379__ & new_new_n52512__;
  assign new_new_n52555__ = ~new_new_n52354__ & new_new_n52554__;
  assign new_new_n52556__ = ~new_new_n52553__ & ~new_new_n52555__;
  assign new_new_n52557__ = ~new_new_n52379__ & new_new_n52512__;
  assign new_new_n52558__ = new_new_n52354__ & new_new_n52557__;
  assign new_new_n52559__ = new_new_n52379__ & ~new_new_n52512__;
  assign new_new_n52560__ = new_new_n52354__ & new_new_n52559__;
  assign new_new_n52561__ = ~new_new_n52558__ & ~new_new_n52560__;
  assign new_new_n52562__ = new_new_n52556__ & new_new_n52561__;
  assign new_new_n52563__ = ~new_new_n52473__ & ~new_new_n52562__;
  assign new_new_n52564__ = ys__n39518 & new_new_n52366__;
  assign new_new_n52565__ = ys__n39520 & new_new_n52356__;
  assign new_new_n52566__ = ~new_new_n52564__ & ~new_new_n52565__;
  assign new_new_n52567__ = ys__n39520 & new_new_n52359__;
  assign new_new_n52568__ = ys__n39520 & new_new_n52358__;
  assign new_new_n52569__ = ~new_new_n52567__ & ~new_new_n52568__;
  assign new_new_n52570__ = new_new_n52566__ & new_new_n52569__;
  assign new_new_n52571__ = ys__n39518 & new_new_n52364__;
  assign new_new_n52572__ = ys__n39518 & new_new_n52367__;
  assign new_new_n52573__ = ~new_new_n52571__ & ~new_new_n52572__;
  assign new_new_n52574__ = new_new_n52377__ & new_new_n52573__;
  assign new_new_n52575__ = new_new_n52570__ & new_new_n52574__;
  assign new_new_n52576__ = ~new_new_n52354__ & ~new_new_n52575__;
  assign new_new_n52577__ = ys__n24834 & new_new_n52383__;
  assign new_new_n52578__ = ys__n24831 & new_new_n52384__;
  assign new_new_n52579__ = ~new_new_n52577__ & ~new_new_n52578__;
  assign new_new_n52580__ = ys__n39778 & new_new_n52391__;
  assign new_new_n52581__ = ys__n39776 & new_new_n52392__;
  assign new_new_n52582__ = ~new_new_n52580__ & ~new_new_n52581__;
  assign new_new_n52583__ = new_new_n52579__ & new_new_n52582__;
  assign new_new_n52584__ = ~new_new_n52575__ & ~new_new_n52583__;
  assign new_new_n52585__ = ~new_new_n52354__ & ~new_new_n52583__;
  assign new_new_n52586__ = ~new_new_n52584__ & ~new_new_n52585__;
  assign new_new_n52587__ = ~new_new_n52576__ & new_new_n52586__;
  assign new_new_n52588__ = ~new_new_n52562__ & ~new_new_n52587__;
  assign new_new_n52589__ = ~new_new_n52473__ & ~new_new_n52587__;
  assign new_new_n52590__ = ~new_new_n52588__ & ~new_new_n52589__;
  assign new_new_n52591__ = ~new_new_n52563__ & new_new_n52590__;
  assign new_new_n52592__ = ~new_new_n52551__ & ~new_new_n52591__;
  assign new_new_n52593__ = ~new_new_n52530__ & ~new_new_n52591__;
  assign new_new_n52594__ = ~new_new_n52592__ & ~new_new_n52593__;
  assign ys__n42189 = new_new_n52552__ | ~new_new_n52594__;
  assign new_new_n52596__ = ~new_new_n52530__ & new_new_n52592__;
  assign new_new_n52597__ = new_new_n52530__ & ~new_new_n52591__;
  assign new_new_n52598__ = new_new_n52551__ & new_new_n52597__;
  assign new_new_n52599__ = ~new_new_n52530__ & new_new_n52591__;
  assign new_new_n52600__ = new_new_n52551__ & new_new_n52599__;
  assign new_new_n52601__ = new_new_n52530__ & new_new_n52591__;
  assign new_new_n52602__ = ~new_new_n52551__ & new_new_n52601__;
  assign new_new_n52603__ = ~new_new_n52600__ & ~new_new_n52602__;
  assign new_new_n52604__ = ~new_new_n52598__ & new_new_n52603__;
  assign ys__n42194 = new_new_n52596__ | ~new_new_n52604__;
  assign new_new_n52606__ = ~new_new_n52473__ & new_new_n52588__;
  assign new_new_n52607__ = new_new_n52473__ & ~new_new_n52587__;
  assign new_new_n52608__ = new_new_n52562__ & new_new_n52607__;
  assign new_new_n52609__ = ~new_new_n52473__ & new_new_n52587__;
  assign new_new_n52610__ = new_new_n52562__ & new_new_n52609__;
  assign new_new_n52611__ = new_new_n52473__ & new_new_n52587__;
  assign new_new_n52612__ = ~new_new_n52562__ & new_new_n52611__;
  assign new_new_n52613__ = ~new_new_n52610__ & ~new_new_n52612__;
  assign new_new_n52614__ = ~new_new_n52608__ & new_new_n52613__;
  assign new_new_n52615__ = ~new_new_n52606__ & new_new_n52614__;
  assign new_new_n52616__ = ~new_new_n52530__ & ~new_new_n52615__;
  assign new_new_n52617__ = ~new_new_n52354__ & new_new_n52584__;
  assign new_new_n52618__ = new_new_n52575__ & new_new_n52583__;
  assign new_new_n52619__ = ~new_new_n52354__ & new_new_n52618__;
  assign new_new_n52620__ = ~new_new_n52617__ & ~new_new_n52619__;
  assign new_new_n52621__ = ~new_new_n52575__ & new_new_n52583__;
  assign new_new_n52622__ = new_new_n52354__ & new_new_n52621__;
  assign new_new_n52623__ = new_new_n52575__ & ~new_new_n52583__;
  assign new_new_n52624__ = new_new_n52354__ & new_new_n52623__;
  assign new_new_n52625__ = ~new_new_n52622__ & ~new_new_n52624__;
  assign new_new_n52626__ = new_new_n52620__ & new_new_n52625__;
  assign new_new_n52627__ = ~new_new_n52473__ & ~new_new_n52626__;
  assign new_new_n52628__ = ys__n24834 & new_new_n52366__;
  assign new_new_n52629__ = ys__n39778 & new_new_n52358__;
  assign new_new_n52630__ = ~new_new_n52628__ & ~new_new_n52629__;
  assign new_new_n52631__ = ys__n33745 & new_new_n52372__;
  assign new_new_n52632__ = ~ys__n33745 & new_new_n52375__;
  assign new_new_n52633__ = ~new_new_n52631__ & ~new_new_n52632__;
  assign new_new_n52634__ = new_new_n52630__ & new_new_n52633__;
  assign new_new_n52635__ = ~new_new_n52565__ & ~new_new_n52567__;
  assign new_new_n52636__ = new_new_n52573__ & new_new_n52635__;
  assign new_new_n52637__ = new_new_n52634__ & new_new_n52636__;
  assign new_new_n52638__ = ~new_new_n52354__ & ~new_new_n52637__;
  assign new_new_n52639__ = ys__n24831 & new_new_n52383__;
  assign new_new_n52640__ = ys__n24828 & new_new_n52384__;
  assign new_new_n52641__ = ~new_new_n52639__ & ~new_new_n52640__;
  assign new_new_n52642__ = ys__n39776 & new_new_n52391__;
  assign new_new_n52643__ = ys__n39774 & new_new_n52392__;
  assign new_new_n52644__ = ~new_new_n52642__ & ~new_new_n52643__;
  assign new_new_n52645__ = new_new_n52641__ & new_new_n52644__;
  assign new_new_n52646__ = ~new_new_n52637__ & ~new_new_n52645__;
  assign new_new_n52647__ = ~new_new_n52354__ & ~new_new_n52645__;
  assign new_new_n52648__ = ~new_new_n52646__ & ~new_new_n52647__;
  assign new_new_n52649__ = ~new_new_n52638__ & new_new_n52648__;
  assign new_new_n52650__ = ~new_new_n52626__ & ~new_new_n52649__;
  assign new_new_n52651__ = ~new_new_n52473__ & ~new_new_n52649__;
  assign new_new_n52652__ = ~new_new_n52650__ & ~new_new_n52651__;
  assign new_new_n52653__ = ~new_new_n52627__ & new_new_n52652__;
  assign new_new_n52654__ = ~new_new_n52615__ & ~new_new_n52653__;
  assign new_new_n52655__ = ~new_new_n52530__ & ~new_new_n52653__;
  assign new_new_n52656__ = ~new_new_n52654__ & ~new_new_n52655__;
  assign ys__n42229 = new_new_n52616__ | ~new_new_n52656__;
  assign new_new_n52658__ = ~new_new_n52530__ & new_new_n52654__;
  assign new_new_n52659__ = new_new_n52530__ & ~new_new_n52653__;
  assign new_new_n52660__ = new_new_n52615__ & new_new_n52659__;
  assign new_new_n52661__ = ~new_new_n52530__ & new_new_n52653__;
  assign new_new_n52662__ = new_new_n52615__ & new_new_n52661__;
  assign new_new_n52663__ = new_new_n52530__ & new_new_n52653__;
  assign new_new_n52664__ = ~new_new_n52615__ & new_new_n52663__;
  assign new_new_n52665__ = ~new_new_n52662__ & ~new_new_n52664__;
  assign new_new_n52666__ = ~new_new_n52660__ & new_new_n52665__;
  assign ys__n42234 = new_new_n52658__ | ~new_new_n52666__;
  assign new_new_n52668__ = ~new_new_n52473__ & new_new_n52650__;
  assign new_new_n52669__ = ~new_new_n52473__ & new_new_n52649__;
  assign new_new_n52670__ = new_new_n52626__ & new_new_n52669__;
  assign new_new_n52671__ = ~new_new_n52668__ & ~new_new_n52670__;
  assign new_new_n52672__ = new_new_n52473__ & new_new_n52649__;
  assign new_new_n52673__ = ~new_new_n52626__ & new_new_n52672__;
  assign new_new_n52674__ = new_new_n52473__ & ~new_new_n52649__;
  assign new_new_n52675__ = new_new_n52626__ & new_new_n52674__;
  assign new_new_n52676__ = ~new_new_n52673__ & ~new_new_n52675__;
  assign new_new_n52677__ = new_new_n52671__ & new_new_n52676__;
  assign new_new_n52678__ = ~new_new_n52530__ & ~new_new_n52677__;
  assign new_new_n52679__ = ~new_new_n52354__ & new_new_n52646__;
  assign new_new_n52680__ = new_new_n52637__ & new_new_n52645__;
  assign new_new_n52681__ = ~new_new_n52354__ & new_new_n52680__;
  assign new_new_n52682__ = ~new_new_n52679__ & ~new_new_n52681__;
  assign new_new_n52683__ = ~new_new_n52637__ & new_new_n52645__;
  assign new_new_n52684__ = new_new_n52354__ & new_new_n52683__;
  assign new_new_n52685__ = new_new_n52637__ & ~new_new_n52645__;
  assign new_new_n52686__ = new_new_n52354__ & new_new_n52685__;
  assign new_new_n52687__ = ~new_new_n52684__ & ~new_new_n52686__;
  assign new_new_n52688__ = new_new_n52682__ & new_new_n52687__;
  assign new_new_n52689__ = ~new_new_n52473__ & ~new_new_n52688__;
  assign new_new_n52690__ = ys__n39778 & new_new_n52359__;
  assign new_new_n52691__ = ys__n39776 & new_new_n52358__;
  assign new_new_n52692__ = ~new_new_n52690__ & ~new_new_n52691__;
  assign new_new_n52693__ = ys__n33743 & new_new_n52372__;
  assign new_new_n52694__ = ~ys__n33743 & new_new_n52375__;
  assign new_new_n52695__ = ~new_new_n52693__ & ~new_new_n52694__;
  assign new_new_n52696__ = new_new_n52692__ & new_new_n52695__;
  assign new_new_n52697__ = ~new_new_n52565__ & ~new_new_n52571__;
  assign new_new_n52698__ = ys__n24834 & new_new_n52367__;
  assign new_new_n52699__ = ys__n24831 & new_new_n52366__;
  assign new_new_n52700__ = ~new_new_n52698__ & ~new_new_n52699__;
  assign new_new_n52701__ = new_new_n52697__ & new_new_n52700__;
  assign new_new_n52702__ = new_new_n52696__ & new_new_n52701__;
  assign new_new_n52703__ = ~new_new_n52354__ & ~new_new_n52702__;
  assign new_new_n52704__ = ys__n24828 & new_new_n52383__;
  assign new_new_n52705__ = ys__n24825 & new_new_n52384__;
  assign new_new_n52706__ = ~new_new_n52704__ & ~new_new_n52705__;
  assign new_new_n52707__ = ys__n39774 & new_new_n52391__;
  assign new_new_n52708__ = ys__n39772 & new_new_n52392__;
  assign new_new_n52709__ = ~new_new_n52707__ & ~new_new_n52708__;
  assign new_new_n52710__ = new_new_n52706__ & new_new_n52709__;
  assign new_new_n52711__ = ~new_new_n52702__ & ~new_new_n52710__;
  assign new_new_n52712__ = ~new_new_n52354__ & ~new_new_n52710__;
  assign new_new_n52713__ = ~new_new_n52711__ & ~new_new_n52712__;
  assign new_new_n52714__ = ~new_new_n52703__ & new_new_n52713__;
  assign new_new_n52715__ = ~new_new_n52688__ & ~new_new_n52714__;
  assign new_new_n52716__ = ~new_new_n52473__ & ~new_new_n52714__;
  assign new_new_n52717__ = ~new_new_n52715__ & ~new_new_n52716__;
  assign new_new_n52718__ = ~new_new_n52689__ & new_new_n52717__;
  assign new_new_n52719__ = ~new_new_n52677__ & ~new_new_n52718__;
  assign new_new_n52720__ = ~new_new_n52530__ & ~new_new_n52718__;
  assign new_new_n52721__ = ~new_new_n52719__ & ~new_new_n52720__;
  assign ys__n42270 = new_new_n52678__ | ~new_new_n52721__;
  assign new_new_n52723__ = ~new_new_n52530__ & new_new_n52719__;
  assign new_new_n52724__ = new_new_n52530__ & ~new_new_n52718__;
  assign new_new_n52725__ = new_new_n52677__ & new_new_n52724__;
  assign new_new_n52726__ = ~new_new_n52530__ & new_new_n52718__;
  assign new_new_n52727__ = new_new_n52677__ & new_new_n52726__;
  assign new_new_n52728__ = new_new_n52530__ & new_new_n52718__;
  assign new_new_n52729__ = ~new_new_n52677__ & new_new_n52728__;
  assign new_new_n52730__ = ~new_new_n52727__ & ~new_new_n52729__;
  assign new_new_n52731__ = ~new_new_n52725__ & new_new_n52730__;
  assign ys__n42275 = new_new_n52723__ | ~new_new_n52731__;
  assign new_new_n52733__ = ~new_new_n52473__ & new_new_n52715__;
  assign new_new_n52734__ = ~new_new_n52473__ & new_new_n52714__;
  assign new_new_n52735__ = new_new_n52688__ & new_new_n52734__;
  assign new_new_n52736__ = ~new_new_n52733__ & ~new_new_n52735__;
  assign new_new_n52737__ = new_new_n52473__ & new_new_n52714__;
  assign new_new_n52738__ = ~new_new_n52688__ & new_new_n52737__;
  assign new_new_n52739__ = new_new_n52473__ & ~new_new_n52714__;
  assign new_new_n52740__ = new_new_n52688__ & new_new_n52739__;
  assign new_new_n52741__ = ~new_new_n52738__ & ~new_new_n52740__;
  assign new_new_n52742__ = new_new_n52736__ & new_new_n52741__;
  assign new_new_n52743__ = ~new_new_n52530__ & ~new_new_n52742__;
  assign new_new_n52744__ = ~new_new_n52354__ & new_new_n52711__;
  assign new_new_n52745__ = new_new_n52702__ & new_new_n52710__;
  assign new_new_n52746__ = ~new_new_n52354__ & new_new_n52745__;
  assign new_new_n52747__ = ~new_new_n52744__ & ~new_new_n52746__;
  assign new_new_n52748__ = ~new_new_n52702__ & new_new_n52710__;
  assign new_new_n52749__ = new_new_n52354__ & new_new_n52748__;
  assign new_new_n52750__ = new_new_n52702__ & ~new_new_n52710__;
  assign new_new_n52751__ = new_new_n52354__ & new_new_n52750__;
  assign new_new_n52752__ = ~new_new_n52749__ & ~new_new_n52751__;
  assign new_new_n52753__ = new_new_n52747__ & new_new_n52752__;
  assign new_new_n52754__ = ~new_new_n52473__ & ~new_new_n52753__;
  assign new_new_n52755__ = ys__n39776 & new_new_n52359__;
  assign new_new_n52756__ = ys__n39774 & new_new_n52358__;
  assign new_new_n52757__ = ~new_new_n52755__ & ~new_new_n52756__;
  assign new_new_n52758__ = ys__n33741 & new_new_n52372__;
  assign new_new_n52759__ = ~ys__n33741 & new_new_n52375__;
  assign new_new_n52760__ = ~new_new_n52758__ & ~new_new_n52759__;
  assign new_new_n52761__ = new_new_n52757__ & new_new_n52760__;
  assign new_new_n52762__ = ys__n24834 & new_new_n52364__;
  assign new_new_n52763__ = ys__n24831 & new_new_n52367__;
  assign new_new_n52764__ = ~new_new_n52762__ & ~new_new_n52763__;
  assign new_new_n52765__ = ys__n24828 & new_new_n52366__;
  assign new_new_n52766__ = ys__n39778 & new_new_n52356__;
  assign new_new_n52767__ = ~new_new_n52765__ & ~new_new_n52766__;
  assign new_new_n52768__ = new_new_n52764__ & new_new_n52767__;
  assign new_new_n52769__ = new_new_n52761__ & new_new_n52768__;
  assign new_new_n52770__ = ys__n39518 & new_new_n52341__;
  assign new_new_n52771__ = ys__n39520 & new_new_n52331__;
  assign new_new_n52772__ = ~new_new_n52770__ & ~new_new_n52771__;
  assign new_new_n52773__ = ys__n39520 & new_new_n52334__;
  assign new_new_n52774__ = ys__n39520 & new_new_n52333__;
  assign new_new_n52775__ = ~new_new_n52773__ & ~new_new_n52774__;
  assign new_new_n52776__ = new_new_n52772__ & new_new_n52775__;
  assign new_new_n52777__ = ys__n39518 & new_new_n52339__;
  assign new_new_n52778__ = ys__n39518 & new_new_n52342__;
  assign new_new_n52779__ = ~new_new_n52777__ & ~new_new_n52778__;
  assign new_new_n52780__ = new_new_n52352__ & new_new_n52779__;
  assign new_new_n52781__ = new_new_n52776__ & new_new_n52780__;
  assign new_new_n52782__ = ~new_new_n52769__ & ~new_new_n52781__;
  assign new_new_n52783__ = ys__n24825 & new_new_n52383__;
  assign new_new_n52784__ = ys__n24822 & new_new_n52384__;
  assign new_new_n52785__ = ~new_new_n52783__ & ~new_new_n52784__;
  assign new_new_n52786__ = ys__n39772 & new_new_n52391__;
  assign new_new_n52787__ = ys__n39770 & new_new_n52392__;
  assign new_new_n52788__ = ~new_new_n52786__ & ~new_new_n52787__;
  assign new_new_n52789__ = new_new_n52785__ & new_new_n52788__;
  assign new_new_n52790__ = ~new_new_n52769__ & ~new_new_n52789__;
  assign new_new_n52791__ = ~new_new_n52781__ & ~new_new_n52789__;
  assign new_new_n52792__ = ~new_new_n52790__ & ~new_new_n52791__;
  assign new_new_n52793__ = ~new_new_n52782__ & new_new_n52792__;
  assign new_new_n52794__ = ~new_new_n52753__ & ~new_new_n52793__;
  assign new_new_n52795__ = ~new_new_n52473__ & ~new_new_n52793__;
  assign new_new_n52796__ = ~new_new_n52794__ & ~new_new_n52795__;
  assign new_new_n52797__ = ~new_new_n52754__ & new_new_n52796__;
  assign new_new_n52798__ = ~new_new_n52742__ & ~new_new_n52797__;
  assign new_new_n52799__ = ~new_new_n52530__ & ~new_new_n52797__;
  assign new_new_n52800__ = ~new_new_n52798__ & ~new_new_n52799__;
  assign ys__n42311 = new_new_n52743__ | ~new_new_n52800__;
  assign new_new_n52802__ = ~new_new_n52530__ & new_new_n52798__;
  assign new_new_n52803__ = new_new_n52530__ & ~new_new_n52797__;
  assign new_new_n52804__ = new_new_n52742__ & new_new_n52803__;
  assign new_new_n52805__ = ~new_new_n52530__ & new_new_n52797__;
  assign new_new_n52806__ = new_new_n52742__ & new_new_n52805__;
  assign new_new_n52807__ = new_new_n52530__ & new_new_n52797__;
  assign new_new_n52808__ = ~new_new_n52742__ & new_new_n52807__;
  assign new_new_n52809__ = ~new_new_n52806__ & ~new_new_n52808__;
  assign new_new_n52810__ = ~new_new_n52804__ & new_new_n52809__;
  assign ys__n42316 = new_new_n52802__ | ~new_new_n52810__;
  assign new_new_n52812__ = ~new_new_n52473__ & new_new_n52794__;
  assign new_new_n52813__ = ~new_new_n52473__ & new_new_n52793__;
  assign new_new_n52814__ = new_new_n52753__ & new_new_n52813__;
  assign new_new_n52815__ = ~new_new_n52812__ & ~new_new_n52814__;
  assign new_new_n52816__ = new_new_n52473__ & new_new_n52793__;
  assign new_new_n52817__ = ~new_new_n52753__ & new_new_n52816__;
  assign new_new_n52818__ = new_new_n52473__ & ~new_new_n52793__;
  assign new_new_n52819__ = new_new_n52753__ & new_new_n52818__;
  assign new_new_n52820__ = ~new_new_n52817__ & ~new_new_n52819__;
  assign new_new_n52821__ = new_new_n52815__ & new_new_n52820__;
  assign new_new_n52822__ = ~new_new_n52530__ & ~new_new_n52821__;
  assign new_new_n52823__ = ~new_new_n52781__ & new_new_n52790__;
  assign new_new_n52824__ = new_new_n52769__ & new_new_n52789__;
  assign new_new_n52825__ = ~new_new_n52781__ & new_new_n52824__;
  assign new_new_n52826__ = ~new_new_n52823__ & ~new_new_n52825__;
  assign new_new_n52827__ = ~new_new_n52769__ & new_new_n52789__;
  assign new_new_n52828__ = new_new_n52781__ & new_new_n52827__;
  assign new_new_n52829__ = new_new_n52769__ & ~new_new_n52789__;
  assign new_new_n52830__ = new_new_n52781__ & new_new_n52829__;
  assign new_new_n52831__ = ~new_new_n52828__ & ~new_new_n52830__;
  assign new_new_n52832__ = new_new_n52826__ & new_new_n52831__;
  assign new_new_n52833__ = ~new_new_n52473__ & ~new_new_n52832__;
  assign new_new_n52834__ = ys__n39774 & new_new_n52359__;
  assign new_new_n52835__ = ys__n39772 & new_new_n52358__;
  assign new_new_n52836__ = ~new_new_n52834__ & ~new_new_n52835__;
  assign new_new_n52837__ = ys__n33739 & new_new_n52372__;
  assign new_new_n52838__ = ~ys__n33739 & new_new_n52375__;
  assign new_new_n52839__ = ~new_new_n52837__ & ~new_new_n52838__;
  assign new_new_n52840__ = new_new_n52836__ & new_new_n52839__;
  assign new_new_n52841__ = ys__n24831 & new_new_n52364__;
  assign new_new_n52842__ = ys__n24828 & new_new_n52367__;
  assign new_new_n52843__ = ~new_new_n52841__ & ~new_new_n52842__;
  assign new_new_n52844__ = ys__n24825 & new_new_n52366__;
  assign new_new_n52845__ = ys__n39776 & new_new_n52356__;
  assign new_new_n52846__ = ~new_new_n52844__ & ~new_new_n52845__;
  assign new_new_n52847__ = new_new_n52843__ & new_new_n52846__;
  assign new_new_n52848__ = new_new_n52840__ & new_new_n52847__;
  assign new_new_n52849__ = ys__n24834 & new_new_n52341__;
  assign new_new_n52850__ = ys__n39778 & new_new_n52333__;
  assign new_new_n52851__ = ~new_new_n52849__ & ~new_new_n52850__;
  assign new_new_n52852__ = ys__n33745 & new_new_n52347__;
  assign new_new_n52853__ = ~ys__n33745 & new_new_n52350__;
  assign new_new_n52854__ = ~new_new_n52852__ & ~new_new_n52853__;
  assign new_new_n52855__ = new_new_n52851__ & new_new_n52854__;
  assign new_new_n52856__ = ~new_new_n52771__ & ~new_new_n52773__;
  assign new_new_n52857__ = new_new_n52779__ & new_new_n52856__;
  assign new_new_n52858__ = new_new_n52855__ & new_new_n52857__;
  assign new_new_n52859__ = ~new_new_n52848__ & ~new_new_n52858__;
  assign new_new_n52860__ = ys__n24822 & new_new_n52383__;
  assign new_new_n52861__ = ys__n24819 & new_new_n52384__;
  assign new_new_n52862__ = ~new_new_n52860__ & ~new_new_n52861__;
  assign new_new_n52863__ = ys__n39770 & new_new_n52391__;
  assign new_new_n52864__ = ys__n39768 & new_new_n52392__;
  assign new_new_n52865__ = ~new_new_n52863__ & ~new_new_n52864__;
  assign new_new_n52866__ = new_new_n52862__ & new_new_n52865__;
  assign new_new_n52867__ = ~new_new_n52848__ & ~new_new_n52866__;
  assign new_new_n52868__ = ~new_new_n52858__ & ~new_new_n52866__;
  assign new_new_n52869__ = ~new_new_n52867__ & ~new_new_n52868__;
  assign new_new_n52870__ = ~new_new_n52859__ & new_new_n52869__;
  assign new_new_n52871__ = ~new_new_n52832__ & ~new_new_n52870__;
  assign new_new_n52872__ = ~new_new_n52473__ & ~new_new_n52870__;
  assign new_new_n52873__ = ~new_new_n52871__ & ~new_new_n52872__;
  assign new_new_n52874__ = ~new_new_n52833__ & new_new_n52873__;
  assign new_new_n52875__ = ~new_new_n52821__ & ~new_new_n52874__;
  assign new_new_n52876__ = ~new_new_n52530__ & ~new_new_n52874__;
  assign new_new_n52877__ = ~new_new_n52875__ & ~new_new_n52876__;
  assign ys__n42352 = new_new_n52822__ | ~new_new_n52877__;
  assign new_new_n52879__ = ~new_new_n52530__ & new_new_n52875__;
  assign new_new_n52880__ = new_new_n52530__ & ~new_new_n52874__;
  assign new_new_n52881__ = new_new_n52821__ & new_new_n52880__;
  assign new_new_n52882__ = ~new_new_n52530__ & new_new_n52874__;
  assign new_new_n52883__ = new_new_n52821__ & new_new_n52882__;
  assign new_new_n52884__ = new_new_n52530__ & new_new_n52874__;
  assign new_new_n52885__ = ~new_new_n52821__ & new_new_n52884__;
  assign new_new_n52886__ = ~new_new_n52883__ & ~new_new_n52885__;
  assign new_new_n52887__ = ~new_new_n52881__ & new_new_n52886__;
  assign ys__n42357 = new_new_n52879__ | ~new_new_n52887__;
  assign new_new_n52889__ = ~new_new_n52473__ & new_new_n52871__;
  assign new_new_n52890__ = ~new_new_n52473__ & new_new_n52870__;
  assign new_new_n52891__ = new_new_n52832__ & new_new_n52890__;
  assign new_new_n52892__ = ~new_new_n52889__ & ~new_new_n52891__;
  assign new_new_n52893__ = new_new_n52473__ & new_new_n52870__;
  assign new_new_n52894__ = ~new_new_n52832__ & new_new_n52893__;
  assign new_new_n52895__ = new_new_n52473__ & ~new_new_n52870__;
  assign new_new_n52896__ = new_new_n52832__ & new_new_n52895__;
  assign new_new_n52897__ = ~new_new_n52894__ & ~new_new_n52896__;
  assign new_new_n52898__ = new_new_n52892__ & new_new_n52897__;
  assign new_new_n52899__ = ~new_new_n52530__ & ~new_new_n52898__;
  assign new_new_n52900__ = ~new_new_n52858__ & new_new_n52867__;
  assign new_new_n52901__ = new_new_n52848__ & new_new_n52866__;
  assign new_new_n52902__ = ~new_new_n52858__ & new_new_n52901__;
  assign new_new_n52903__ = ~new_new_n52900__ & ~new_new_n52902__;
  assign new_new_n52904__ = ~new_new_n52848__ & new_new_n52866__;
  assign new_new_n52905__ = new_new_n52858__ & new_new_n52904__;
  assign new_new_n52906__ = new_new_n52848__ & ~new_new_n52866__;
  assign new_new_n52907__ = new_new_n52858__ & new_new_n52906__;
  assign new_new_n52908__ = ~new_new_n52905__ & ~new_new_n52907__;
  assign new_new_n52909__ = new_new_n52903__ & new_new_n52908__;
  assign new_new_n52910__ = ~new_new_n52473__ & ~new_new_n52909__;
  assign new_new_n52911__ = ys__n39772 & new_new_n52359__;
  assign new_new_n52912__ = ys__n39770 & new_new_n52358__;
  assign new_new_n52913__ = ~new_new_n52911__ & ~new_new_n52912__;
  assign new_new_n52914__ = ys__n33737 & new_new_n52372__;
  assign new_new_n52915__ = ~ys__n33737 & new_new_n52375__;
  assign new_new_n52916__ = ~new_new_n52914__ & ~new_new_n52915__;
  assign new_new_n52917__ = new_new_n52913__ & new_new_n52916__;
  assign new_new_n52918__ = ys__n24828 & new_new_n52364__;
  assign new_new_n52919__ = ys__n24825 & new_new_n52367__;
  assign new_new_n52920__ = ~new_new_n52918__ & ~new_new_n52919__;
  assign new_new_n52921__ = ys__n24822 & new_new_n52366__;
  assign new_new_n52922__ = ys__n39774 & new_new_n52356__;
  assign new_new_n52923__ = ~new_new_n52921__ & ~new_new_n52922__;
  assign new_new_n52924__ = new_new_n52920__ & new_new_n52923__;
  assign new_new_n52925__ = new_new_n52917__ & new_new_n52924__;
  assign new_new_n52926__ = ys__n39778 & new_new_n52334__;
  assign new_new_n52927__ = ys__n39776 & new_new_n52333__;
  assign new_new_n52928__ = ~new_new_n52926__ & ~new_new_n52927__;
  assign new_new_n52929__ = ys__n33743 & new_new_n52347__;
  assign new_new_n52930__ = ~ys__n33743 & new_new_n52350__;
  assign new_new_n52931__ = ~new_new_n52929__ & ~new_new_n52930__;
  assign new_new_n52932__ = new_new_n52928__ & new_new_n52931__;
  assign new_new_n52933__ = ~new_new_n52771__ & ~new_new_n52777__;
  assign new_new_n52934__ = ys__n24834 & new_new_n52342__;
  assign new_new_n52935__ = ys__n24831 & new_new_n52341__;
  assign new_new_n52936__ = ~new_new_n52934__ & ~new_new_n52935__;
  assign new_new_n52937__ = new_new_n52933__ & new_new_n52936__;
  assign new_new_n52938__ = new_new_n52932__ & new_new_n52937__;
  assign new_new_n52939__ = ~new_new_n52925__ & ~new_new_n52938__;
  assign new_new_n52940__ = ys__n24819 & new_new_n52383__;
  assign new_new_n52941__ = ys__n24816 & new_new_n52384__;
  assign new_new_n52942__ = ~new_new_n52940__ & ~new_new_n52941__;
  assign new_new_n52943__ = ys__n39768 & new_new_n52391__;
  assign new_new_n52944__ = ys__n39766 & new_new_n52392__;
  assign new_new_n52945__ = ~new_new_n52943__ & ~new_new_n52944__;
  assign new_new_n52946__ = new_new_n52942__ & new_new_n52945__;
  assign new_new_n52947__ = ~new_new_n52925__ & ~new_new_n52946__;
  assign new_new_n52948__ = ~new_new_n52938__ & ~new_new_n52946__;
  assign new_new_n52949__ = ~new_new_n52947__ & ~new_new_n52948__;
  assign new_new_n52950__ = ~new_new_n52939__ & new_new_n52949__;
  assign new_new_n52951__ = ~new_new_n52909__ & ~new_new_n52950__;
  assign new_new_n52952__ = ~new_new_n52473__ & ~new_new_n52950__;
  assign new_new_n52953__ = ~new_new_n52951__ & ~new_new_n52952__;
  assign new_new_n52954__ = ~new_new_n52910__ & new_new_n52953__;
  assign new_new_n52955__ = ~new_new_n52898__ & ~new_new_n52954__;
  assign new_new_n52956__ = ~new_new_n52530__ & ~new_new_n52954__;
  assign new_new_n52957__ = ~new_new_n52955__ & ~new_new_n52956__;
  assign ys__n42393 = new_new_n52899__ | ~new_new_n52957__;
  assign new_new_n52959__ = ~new_new_n52530__ & new_new_n52955__;
  assign new_new_n52960__ = new_new_n52530__ & ~new_new_n52954__;
  assign new_new_n52961__ = new_new_n52898__ & new_new_n52960__;
  assign new_new_n52962__ = ~new_new_n52530__ & new_new_n52954__;
  assign new_new_n52963__ = new_new_n52898__ & new_new_n52962__;
  assign new_new_n52964__ = new_new_n52530__ & new_new_n52954__;
  assign new_new_n52965__ = ~new_new_n52898__ & new_new_n52964__;
  assign new_new_n52966__ = ~new_new_n52963__ & ~new_new_n52965__;
  assign new_new_n52967__ = ~new_new_n52961__ & new_new_n52966__;
  assign ys__n42398 = new_new_n52959__ | ~new_new_n52967__;
  assign new_new_n52969__ = ~new_new_n52473__ & new_new_n52951__;
  assign new_new_n52970__ = ~new_new_n52473__ & new_new_n52950__;
  assign new_new_n52971__ = new_new_n52909__ & new_new_n52970__;
  assign new_new_n52972__ = ~new_new_n52969__ & ~new_new_n52971__;
  assign new_new_n52973__ = new_new_n52473__ & new_new_n52950__;
  assign new_new_n52974__ = ~new_new_n52909__ & new_new_n52973__;
  assign new_new_n52975__ = new_new_n52473__ & ~new_new_n52950__;
  assign new_new_n52976__ = new_new_n52909__ & new_new_n52975__;
  assign new_new_n52977__ = ~new_new_n52974__ & ~new_new_n52976__;
  assign new_new_n52978__ = new_new_n52972__ & new_new_n52977__;
  assign new_new_n52979__ = ~new_new_n52530__ & ~new_new_n52978__;
  assign new_new_n52980__ = ~new_new_n52938__ & new_new_n52947__;
  assign new_new_n52981__ = new_new_n52925__ & new_new_n52946__;
  assign new_new_n52982__ = ~new_new_n52938__ & new_new_n52981__;
  assign new_new_n52983__ = ~new_new_n52980__ & ~new_new_n52982__;
  assign new_new_n52984__ = ~new_new_n52925__ & new_new_n52946__;
  assign new_new_n52985__ = new_new_n52938__ & new_new_n52984__;
  assign new_new_n52986__ = new_new_n52925__ & ~new_new_n52946__;
  assign new_new_n52987__ = new_new_n52938__ & new_new_n52986__;
  assign new_new_n52988__ = ~new_new_n52985__ & ~new_new_n52987__;
  assign new_new_n52989__ = new_new_n52983__ & new_new_n52988__;
  assign new_new_n52990__ = ys__n39518 & new_new_n52456__;
  assign new_new_n52991__ = ys__n39520 & new_new_n52446__;
  assign new_new_n52992__ = ~new_new_n52990__ & ~new_new_n52991__;
  assign new_new_n52993__ = ys__n39520 & new_new_n52449__;
  assign new_new_n52994__ = ys__n39520 & new_new_n52448__;
  assign new_new_n52995__ = ~new_new_n52993__ & ~new_new_n52994__;
  assign new_new_n52996__ = new_new_n52992__ & new_new_n52995__;
  assign new_new_n52997__ = ys__n39518 & new_new_n52454__;
  assign new_new_n52998__ = ys__n39518 & new_new_n52457__;
  assign new_new_n52999__ = ~new_new_n52997__ & ~new_new_n52998__;
  assign new_new_n53000__ = new_new_n52467__ & new_new_n52999__;
  assign new_new_n53001__ = new_new_n52996__ & new_new_n53000__;
  assign new_new_n53002__ = ~new_new_n52443__ & ~new_new_n53001__;
  assign new_new_n53003__ = ~new_new_n52432__ & ~new_new_n53001__;
  assign new_new_n53004__ = ~new_new_n52444__ & ~new_new_n53003__;
  assign new_new_n53005__ = ~new_new_n53002__ & new_new_n53004__;
  assign new_new_n53006__ = ~new_new_n52989__ & ~new_new_n53005__;
  assign new_new_n53007__ = ys__n39770 & new_new_n52359__;
  assign new_new_n53008__ = ys__n39768 & new_new_n52358__;
  assign new_new_n53009__ = ~new_new_n53007__ & ~new_new_n53008__;
  assign new_new_n53010__ = ys__n33735 & new_new_n52372__;
  assign new_new_n53011__ = ~ys__n33735 & new_new_n52375__;
  assign new_new_n53012__ = ~new_new_n53010__ & ~new_new_n53011__;
  assign new_new_n53013__ = new_new_n53009__ & new_new_n53012__;
  assign new_new_n53014__ = ys__n24825 & new_new_n52364__;
  assign new_new_n53015__ = ys__n24822 & new_new_n52367__;
  assign new_new_n53016__ = ~new_new_n53014__ & ~new_new_n53015__;
  assign new_new_n53017__ = ys__n24819 & new_new_n52366__;
  assign new_new_n53018__ = ys__n39772 & new_new_n52356__;
  assign new_new_n53019__ = ~new_new_n53017__ & ~new_new_n53018__;
  assign new_new_n53020__ = new_new_n53016__ & new_new_n53019__;
  assign new_new_n53021__ = new_new_n53013__ & new_new_n53020__;
  assign new_new_n53022__ = ys__n39776 & new_new_n52334__;
  assign new_new_n53023__ = ys__n39774 & new_new_n52333__;
  assign new_new_n53024__ = ~new_new_n53022__ & ~new_new_n53023__;
  assign new_new_n53025__ = ys__n33741 & new_new_n52347__;
  assign new_new_n53026__ = ~ys__n33741 & new_new_n52350__;
  assign new_new_n53027__ = ~new_new_n53025__ & ~new_new_n53026__;
  assign new_new_n53028__ = new_new_n53024__ & new_new_n53027__;
  assign new_new_n53029__ = ys__n24834 & new_new_n52339__;
  assign new_new_n53030__ = ys__n24831 & new_new_n52342__;
  assign new_new_n53031__ = ~new_new_n53029__ & ~new_new_n53030__;
  assign new_new_n53032__ = ys__n24828 & new_new_n52341__;
  assign new_new_n53033__ = ys__n39778 & new_new_n52331__;
  assign new_new_n53034__ = ~new_new_n53032__ & ~new_new_n53033__;
  assign new_new_n53035__ = new_new_n53031__ & new_new_n53034__;
  assign new_new_n53036__ = new_new_n53028__ & new_new_n53035__;
  assign new_new_n53037__ = ~new_new_n53021__ & ~new_new_n53036__;
  assign new_new_n53038__ = ys__n24816 & new_new_n52383__;
  assign new_new_n53039__ = ys__n24813 & new_new_n52384__;
  assign new_new_n53040__ = ~new_new_n53038__ & ~new_new_n53039__;
  assign new_new_n53041__ = ys__n39766 & new_new_n52391__;
  assign new_new_n53042__ = ys__n39764 & new_new_n52392__;
  assign new_new_n53043__ = ~new_new_n53041__ & ~new_new_n53042__;
  assign new_new_n53044__ = new_new_n53040__ & new_new_n53043__;
  assign new_new_n53045__ = ~new_new_n53021__ & ~new_new_n53044__;
  assign new_new_n53046__ = ~new_new_n53036__ & ~new_new_n53044__;
  assign new_new_n53047__ = ~new_new_n53045__ & ~new_new_n53046__;
  assign new_new_n53048__ = ~new_new_n53037__ & new_new_n53047__;
  assign new_new_n53049__ = ~new_new_n52989__ & ~new_new_n53048__;
  assign new_new_n53050__ = ~new_new_n53005__ & ~new_new_n53048__;
  assign new_new_n53051__ = ~new_new_n53049__ & ~new_new_n53050__;
  assign new_new_n53052__ = ~new_new_n53006__ & new_new_n53051__;
  assign new_new_n53053__ = ~new_new_n52978__ & ~new_new_n53052__;
  assign new_new_n53054__ = ~new_new_n52530__ & ~new_new_n53052__;
  assign new_new_n53055__ = ~new_new_n53053__ & ~new_new_n53054__;
  assign ys__n42434 = new_new_n52979__ | ~new_new_n53055__;
  assign new_new_n53057__ = ~new_new_n52530__ & new_new_n53053__;
  assign new_new_n53058__ = new_new_n52530__ & ~new_new_n53052__;
  assign new_new_n53059__ = new_new_n52978__ & new_new_n53058__;
  assign new_new_n53060__ = ~new_new_n52530__ & new_new_n53052__;
  assign new_new_n53061__ = new_new_n52978__ & new_new_n53060__;
  assign new_new_n53062__ = new_new_n52530__ & new_new_n53052__;
  assign new_new_n53063__ = ~new_new_n52978__ & new_new_n53062__;
  assign new_new_n53064__ = ~new_new_n53061__ & ~new_new_n53063__;
  assign new_new_n53065__ = ~new_new_n53059__ & new_new_n53064__;
  assign ys__n42439 = new_new_n53057__ | ~new_new_n53065__;
  assign new_new_n53067__ = ~new_new_n53005__ & new_new_n53049__;
  assign new_new_n53068__ = new_new_n52989__ & new_new_n53048__;
  assign new_new_n53069__ = ~new_new_n53005__ & new_new_n53068__;
  assign new_new_n53070__ = ~new_new_n53067__ & ~new_new_n53069__;
  assign new_new_n53071__ = ~new_new_n52989__ & new_new_n53048__;
  assign new_new_n53072__ = new_new_n53005__ & new_new_n53071__;
  assign new_new_n53073__ = new_new_n52989__ & ~new_new_n53048__;
  assign new_new_n53074__ = new_new_n53005__ & new_new_n53073__;
  assign new_new_n53075__ = ~new_new_n53072__ & ~new_new_n53074__;
  assign new_new_n53076__ = new_new_n53070__ & new_new_n53075__;
  assign new_new_n53077__ = ~new_new_n52530__ & ~new_new_n53076__;
  assign new_new_n53078__ = ~new_new_n53036__ & new_new_n53045__;
  assign new_new_n53079__ = new_new_n53021__ & new_new_n53044__;
  assign new_new_n53080__ = ~new_new_n53036__ & new_new_n53079__;
  assign new_new_n53081__ = ~new_new_n53078__ & ~new_new_n53080__;
  assign new_new_n53082__ = ~new_new_n53021__ & new_new_n53044__;
  assign new_new_n53083__ = new_new_n53036__ & new_new_n53082__;
  assign new_new_n53084__ = new_new_n53021__ & ~new_new_n53044__;
  assign new_new_n53085__ = new_new_n53036__ & new_new_n53084__;
  assign new_new_n53086__ = ~new_new_n53083__ & ~new_new_n53085__;
  assign new_new_n53087__ = new_new_n53081__ & new_new_n53086__;
  assign new_new_n53088__ = ys__n24834 & new_new_n52456__;
  assign new_new_n53089__ = ys__n39778 & new_new_n52448__;
  assign new_new_n53090__ = ~new_new_n53088__ & ~new_new_n53089__;
  assign new_new_n53091__ = ys__n33745 & new_new_n52462__;
  assign new_new_n53092__ = ~ys__n33745 & new_new_n52465__;
  assign new_new_n53093__ = ~new_new_n53091__ & ~new_new_n53092__;
  assign new_new_n53094__ = new_new_n53090__ & new_new_n53093__;
  assign new_new_n53095__ = ~new_new_n52991__ & ~new_new_n52993__;
  assign new_new_n53096__ = new_new_n52999__ & new_new_n53095__;
  assign new_new_n53097__ = new_new_n53094__ & new_new_n53096__;
  assign new_new_n53098__ = ~new_new_n52443__ & ~new_new_n53097__;
  assign new_new_n53099__ = ~new_new_n52432__ & ~new_new_n53097__;
  assign new_new_n53100__ = ~new_new_n52444__ & ~new_new_n53099__;
  assign new_new_n53101__ = ~new_new_n53098__ & new_new_n53100__;
  assign new_new_n53102__ = ~new_new_n53087__ & ~new_new_n53101__;
  assign new_new_n53103__ = ys__n39768 & new_new_n52359__;
  assign new_new_n53104__ = ys__n39766 & new_new_n52358__;
  assign new_new_n53105__ = ~new_new_n53103__ & ~new_new_n53104__;
  assign new_new_n53106__ = ys__n33733 & new_new_n52372__;
  assign new_new_n53107__ = ~ys__n33733 & new_new_n52375__;
  assign new_new_n53108__ = ~new_new_n53106__ & ~new_new_n53107__;
  assign new_new_n53109__ = new_new_n53105__ & new_new_n53108__;
  assign new_new_n53110__ = ys__n24822 & new_new_n52364__;
  assign new_new_n53111__ = ys__n24819 & new_new_n52367__;
  assign new_new_n53112__ = ~new_new_n53110__ & ~new_new_n53111__;
  assign new_new_n53113__ = ys__n24816 & new_new_n52366__;
  assign new_new_n53114__ = ys__n39770 & new_new_n52356__;
  assign new_new_n53115__ = ~new_new_n53113__ & ~new_new_n53114__;
  assign new_new_n53116__ = new_new_n53112__ & new_new_n53115__;
  assign new_new_n53117__ = new_new_n53109__ & new_new_n53116__;
  assign new_new_n53118__ = ys__n39774 & new_new_n52334__;
  assign new_new_n53119__ = ys__n39772 & new_new_n52333__;
  assign new_new_n53120__ = ~new_new_n53118__ & ~new_new_n53119__;
  assign new_new_n53121__ = ys__n33739 & new_new_n52347__;
  assign new_new_n53122__ = ~ys__n33739 & new_new_n52350__;
  assign new_new_n53123__ = ~new_new_n53121__ & ~new_new_n53122__;
  assign new_new_n53124__ = new_new_n53120__ & new_new_n53123__;
  assign new_new_n53125__ = ys__n24831 & new_new_n52339__;
  assign new_new_n53126__ = ys__n24828 & new_new_n52342__;
  assign new_new_n53127__ = ~new_new_n53125__ & ~new_new_n53126__;
  assign new_new_n53128__ = ys__n24825 & new_new_n52341__;
  assign new_new_n53129__ = ys__n39776 & new_new_n52331__;
  assign new_new_n53130__ = ~new_new_n53128__ & ~new_new_n53129__;
  assign new_new_n53131__ = new_new_n53127__ & new_new_n53130__;
  assign new_new_n53132__ = new_new_n53124__ & new_new_n53131__;
  assign new_new_n53133__ = ~new_new_n53117__ & ~new_new_n53132__;
  assign new_new_n53134__ = ys__n24813 & new_new_n52383__;
  assign new_new_n53135__ = ys__n24810 & new_new_n52384__;
  assign new_new_n53136__ = ~new_new_n53134__ & ~new_new_n53135__;
  assign new_new_n53137__ = ys__n39764 & new_new_n52391__;
  assign new_new_n53138__ = ys__n39762 & new_new_n52392__;
  assign new_new_n53139__ = ~new_new_n53137__ & ~new_new_n53138__;
  assign new_new_n53140__ = new_new_n53136__ & new_new_n53139__;
  assign new_new_n53141__ = ~new_new_n53117__ & ~new_new_n53140__;
  assign new_new_n53142__ = ~new_new_n53132__ & ~new_new_n53140__;
  assign new_new_n53143__ = ~new_new_n53141__ & ~new_new_n53142__;
  assign new_new_n53144__ = ~new_new_n53133__ & new_new_n53143__;
  assign new_new_n53145__ = ~new_new_n53087__ & ~new_new_n53144__;
  assign new_new_n53146__ = ~new_new_n53101__ & ~new_new_n53144__;
  assign new_new_n53147__ = ~new_new_n53145__ & ~new_new_n53146__;
  assign new_new_n53148__ = ~new_new_n53102__ & new_new_n53147__;
  assign new_new_n53149__ = ~new_new_n53076__ & ~new_new_n53148__;
  assign new_new_n53150__ = ~new_new_n52530__ & ~new_new_n53148__;
  assign new_new_n53151__ = ~new_new_n53149__ & ~new_new_n53150__;
  assign ys__n42488 = new_new_n53077__ | ~new_new_n53151__;
  assign new_new_n53153__ = ~new_new_n52530__ & new_new_n53149__;
  assign new_new_n53154__ = new_new_n52530__ & ~new_new_n53148__;
  assign new_new_n53155__ = new_new_n53076__ & new_new_n53154__;
  assign new_new_n53156__ = ~new_new_n52530__ & new_new_n53148__;
  assign new_new_n53157__ = new_new_n53076__ & new_new_n53156__;
  assign new_new_n53158__ = new_new_n52530__ & new_new_n53148__;
  assign new_new_n53159__ = ~new_new_n53076__ & new_new_n53158__;
  assign new_new_n53160__ = ~new_new_n53157__ & ~new_new_n53159__;
  assign new_new_n53161__ = ~new_new_n53155__ & new_new_n53160__;
  assign ys__n42493 = new_new_n53153__ | ~new_new_n53161__;
  assign new_new_n53163__ = ~new_new_n53101__ & new_new_n53145__;
  assign new_new_n53164__ = new_new_n53087__ & new_new_n53144__;
  assign new_new_n53165__ = ~new_new_n53101__ & new_new_n53164__;
  assign new_new_n53166__ = ~new_new_n53163__ & ~new_new_n53165__;
  assign new_new_n53167__ = ~new_new_n53087__ & new_new_n53144__;
  assign new_new_n53168__ = new_new_n53101__ & new_new_n53167__;
  assign new_new_n53169__ = new_new_n53087__ & ~new_new_n53144__;
  assign new_new_n53170__ = new_new_n53101__ & new_new_n53169__;
  assign new_new_n53171__ = ~new_new_n53168__ & ~new_new_n53170__;
  assign new_new_n53172__ = new_new_n53166__ & new_new_n53171__;
  assign new_new_n53173__ = ~new_new_n52443__ & new_new_n53003__;
  assign new_new_n53174__ = new_new_n52432__ & new_new_n53001__;
  assign new_new_n53175__ = ~new_new_n52443__ & new_new_n53174__;
  assign new_new_n53176__ = ~new_new_n53173__ & ~new_new_n53175__;
  assign new_new_n53177__ = ~new_new_n52432__ & new_new_n53001__;
  assign new_new_n53178__ = new_new_n52443__ & new_new_n53177__;
  assign new_new_n53179__ = new_new_n52432__ & ~new_new_n53001__;
  assign new_new_n53180__ = new_new_n52443__ & new_new_n53179__;
  assign new_new_n53181__ = ~new_new_n53178__ & ~new_new_n53180__;
  assign new_new_n53182__ = new_new_n53176__ & new_new_n53181__;
  assign new_new_n53183__ = ~new_new_n53172__ & ~new_new_n53182__;
  assign new_new_n53184__ = ~new_new_n53132__ & new_new_n53141__;
  assign new_new_n53185__ = new_new_n53117__ & new_new_n53140__;
  assign new_new_n53186__ = ~new_new_n53132__ & new_new_n53185__;
  assign new_new_n53187__ = ~new_new_n53184__ & ~new_new_n53186__;
  assign new_new_n53188__ = ~new_new_n53117__ & new_new_n53140__;
  assign new_new_n53189__ = new_new_n53132__ & new_new_n53188__;
  assign new_new_n53190__ = new_new_n53117__ & ~new_new_n53140__;
  assign new_new_n53191__ = new_new_n53132__ & new_new_n53190__;
  assign new_new_n53192__ = ~new_new_n53189__ & ~new_new_n53191__;
  assign new_new_n53193__ = new_new_n53187__ & new_new_n53192__;
  assign new_new_n53194__ = ys__n39778 & new_new_n52449__;
  assign new_new_n53195__ = ys__n39776 & new_new_n52448__;
  assign new_new_n53196__ = ~new_new_n53194__ & ~new_new_n53195__;
  assign new_new_n53197__ = ys__n33743 & new_new_n52462__;
  assign new_new_n53198__ = ~ys__n33743 & new_new_n52465__;
  assign new_new_n53199__ = ~new_new_n53197__ & ~new_new_n53198__;
  assign new_new_n53200__ = new_new_n53196__ & new_new_n53199__;
  assign new_new_n53201__ = ~new_new_n52991__ & ~new_new_n52997__;
  assign new_new_n53202__ = ys__n24834 & new_new_n52457__;
  assign new_new_n53203__ = ys__n24831 & new_new_n52456__;
  assign new_new_n53204__ = ~new_new_n53202__ & ~new_new_n53203__;
  assign new_new_n53205__ = new_new_n53201__ & new_new_n53204__;
  assign new_new_n53206__ = new_new_n53200__ & new_new_n53205__;
  assign new_new_n53207__ = ~new_new_n52443__ & ~new_new_n53206__;
  assign new_new_n53208__ = ~new_new_n52432__ & ~new_new_n53206__;
  assign new_new_n53209__ = ~new_new_n52444__ & ~new_new_n53208__;
  assign new_new_n53210__ = ~new_new_n53207__ & new_new_n53209__;
  assign new_new_n53211__ = ~new_new_n53193__ & ~new_new_n53210__;
  assign new_new_n53212__ = ys__n39766 & new_new_n52359__;
  assign new_new_n53213__ = ys__n39764 & new_new_n52358__;
  assign new_new_n53214__ = ~new_new_n53212__ & ~new_new_n53213__;
  assign new_new_n53215__ = ys__n33731 & new_new_n52372__;
  assign new_new_n53216__ = ~ys__n33731 & new_new_n52375__;
  assign new_new_n53217__ = ~new_new_n53215__ & ~new_new_n53216__;
  assign new_new_n53218__ = new_new_n53214__ & new_new_n53217__;
  assign new_new_n53219__ = ys__n24819 & new_new_n52364__;
  assign new_new_n53220__ = ys__n24816 & new_new_n52367__;
  assign new_new_n53221__ = ~new_new_n53219__ & ~new_new_n53220__;
  assign new_new_n53222__ = ys__n24813 & new_new_n52366__;
  assign new_new_n53223__ = ys__n39768 & new_new_n52356__;
  assign new_new_n53224__ = ~new_new_n53222__ & ~new_new_n53223__;
  assign new_new_n53225__ = new_new_n53221__ & new_new_n53224__;
  assign new_new_n53226__ = new_new_n53218__ & new_new_n53225__;
  assign new_new_n53227__ = ys__n39772 & new_new_n52334__;
  assign new_new_n53228__ = ys__n39770 & new_new_n52333__;
  assign new_new_n53229__ = ~new_new_n53227__ & ~new_new_n53228__;
  assign new_new_n53230__ = ys__n33737 & new_new_n52347__;
  assign new_new_n53231__ = ~ys__n33737 & new_new_n52350__;
  assign new_new_n53232__ = ~new_new_n53230__ & ~new_new_n53231__;
  assign new_new_n53233__ = new_new_n53229__ & new_new_n53232__;
  assign new_new_n53234__ = ys__n24828 & new_new_n52339__;
  assign new_new_n53235__ = ys__n24825 & new_new_n52342__;
  assign new_new_n53236__ = ~new_new_n53234__ & ~new_new_n53235__;
  assign new_new_n53237__ = ys__n24822 & new_new_n52341__;
  assign new_new_n53238__ = ys__n39774 & new_new_n52331__;
  assign new_new_n53239__ = ~new_new_n53237__ & ~new_new_n53238__;
  assign new_new_n53240__ = new_new_n53236__ & new_new_n53239__;
  assign new_new_n53241__ = new_new_n53233__ & new_new_n53240__;
  assign new_new_n53242__ = ~new_new_n53226__ & ~new_new_n53241__;
  assign new_new_n53243__ = ys__n24810 & new_new_n52383__;
  assign new_new_n53244__ = ys__n24807 & new_new_n52384__;
  assign new_new_n53245__ = ~new_new_n53243__ & ~new_new_n53244__;
  assign new_new_n53246__ = ys__n39762 & new_new_n52391__;
  assign new_new_n53247__ = ys__n39760 & new_new_n52392__;
  assign new_new_n53248__ = ~new_new_n53246__ & ~new_new_n53247__;
  assign new_new_n53249__ = new_new_n53245__ & new_new_n53248__;
  assign new_new_n53250__ = ~new_new_n53226__ & ~new_new_n53249__;
  assign new_new_n53251__ = ~new_new_n53241__ & ~new_new_n53249__;
  assign new_new_n53252__ = ~new_new_n53250__ & ~new_new_n53251__;
  assign new_new_n53253__ = ~new_new_n53242__ & new_new_n53252__;
  assign new_new_n53254__ = ~new_new_n53193__ & ~new_new_n53253__;
  assign new_new_n53255__ = ~new_new_n53210__ & ~new_new_n53253__;
  assign new_new_n53256__ = ~new_new_n53254__ & ~new_new_n53255__;
  assign new_new_n53257__ = ~new_new_n53211__ & new_new_n53256__;
  assign new_new_n53258__ = ~new_new_n53172__ & ~new_new_n53257__;
  assign new_new_n53259__ = ~new_new_n53182__ & ~new_new_n53257__;
  assign new_new_n53260__ = ~new_new_n53258__ & ~new_new_n53259__;
  assign ys__n42541 = new_new_n53183__ | ~new_new_n53260__;
  assign new_new_n53262__ = ~new_new_n53182__ & new_new_n53258__;
  assign new_new_n53263__ = new_new_n53182__ & ~new_new_n53257__;
  assign new_new_n53264__ = new_new_n53172__ & new_new_n53263__;
  assign new_new_n53265__ = ~new_new_n53182__ & new_new_n53257__;
  assign new_new_n53266__ = new_new_n53172__ & new_new_n53265__;
  assign new_new_n53267__ = new_new_n53182__ & new_new_n53257__;
  assign new_new_n53268__ = ~new_new_n53172__ & new_new_n53267__;
  assign new_new_n53269__ = ~new_new_n53266__ & ~new_new_n53268__;
  assign new_new_n53270__ = ~new_new_n53264__ & new_new_n53269__;
  assign ys__n42546 = new_new_n53262__ | ~new_new_n53270__;
  assign new_new_n53272__ = ~new_new_n53210__ & new_new_n53254__;
  assign new_new_n53273__ = new_new_n53193__ & new_new_n53253__;
  assign new_new_n53274__ = ~new_new_n53210__ & new_new_n53273__;
  assign new_new_n53275__ = ~new_new_n53272__ & ~new_new_n53274__;
  assign new_new_n53276__ = ~new_new_n53193__ & new_new_n53253__;
  assign new_new_n53277__ = new_new_n53210__ & new_new_n53276__;
  assign new_new_n53278__ = new_new_n53193__ & ~new_new_n53253__;
  assign new_new_n53279__ = new_new_n53210__ & new_new_n53278__;
  assign new_new_n53280__ = ~new_new_n53277__ & ~new_new_n53279__;
  assign new_new_n53281__ = new_new_n53275__ & new_new_n53280__;
  assign new_new_n53282__ = ~new_new_n52443__ & new_new_n53099__;
  assign new_new_n53283__ = new_new_n52432__ & new_new_n53097__;
  assign new_new_n53284__ = ~new_new_n52443__ & new_new_n53283__;
  assign new_new_n53285__ = ~new_new_n53282__ & ~new_new_n53284__;
  assign new_new_n53286__ = ~new_new_n52432__ & new_new_n53097__;
  assign new_new_n53287__ = new_new_n52443__ & new_new_n53286__;
  assign new_new_n53288__ = new_new_n52432__ & ~new_new_n53097__;
  assign new_new_n53289__ = new_new_n52443__ & new_new_n53288__;
  assign new_new_n53290__ = ~new_new_n53287__ & ~new_new_n53289__;
  assign new_new_n53291__ = new_new_n53285__ & new_new_n53290__;
  assign new_new_n53292__ = ~new_new_n53281__ & ~new_new_n53291__;
  assign new_new_n53293__ = ~new_new_n53241__ & new_new_n53250__;
  assign new_new_n53294__ = new_new_n53226__ & new_new_n53249__;
  assign new_new_n53295__ = ~new_new_n53241__ & new_new_n53294__;
  assign new_new_n53296__ = ~new_new_n53293__ & ~new_new_n53295__;
  assign new_new_n53297__ = ~new_new_n53226__ & new_new_n53249__;
  assign new_new_n53298__ = new_new_n53241__ & new_new_n53297__;
  assign new_new_n53299__ = new_new_n53226__ & ~new_new_n53249__;
  assign new_new_n53300__ = new_new_n53241__ & new_new_n53299__;
  assign new_new_n53301__ = ~new_new_n53298__ & ~new_new_n53300__;
  assign new_new_n53302__ = new_new_n53296__ & new_new_n53301__;
  assign new_new_n53303__ = ys__n39518 & new_new_n52419__;
  assign new_new_n53304__ = ys__n39520 & new_new_n52409__;
  assign new_new_n53305__ = ~new_new_n53303__ & ~new_new_n53304__;
  assign new_new_n53306__ = ys__n39520 & new_new_n52412__;
  assign new_new_n53307__ = ys__n39520 & new_new_n52411__;
  assign new_new_n53308__ = ~new_new_n53306__ & ~new_new_n53307__;
  assign new_new_n53309__ = new_new_n53305__ & new_new_n53308__;
  assign new_new_n53310__ = ys__n39518 & new_new_n52417__;
  assign new_new_n53311__ = ys__n39518 & new_new_n52420__;
  assign new_new_n53312__ = ~new_new_n53310__ & ~new_new_n53311__;
  assign new_new_n53313__ = new_new_n52430__ & new_new_n53312__;
  assign new_new_n53314__ = new_new_n53309__ & new_new_n53313__;
  assign new_new_n53315__ = ~new_new_n52443__ & ~new_new_n53314__;
  assign new_new_n53316__ = ys__n39776 & new_new_n52449__;
  assign new_new_n53317__ = ys__n39774 & new_new_n52448__;
  assign new_new_n53318__ = ~new_new_n53316__ & ~new_new_n53317__;
  assign new_new_n53319__ = ys__n33741 & new_new_n52462__;
  assign new_new_n53320__ = ~ys__n33741 & new_new_n52465__;
  assign new_new_n53321__ = ~new_new_n53319__ & ~new_new_n53320__;
  assign new_new_n53322__ = new_new_n53318__ & new_new_n53321__;
  assign new_new_n53323__ = ys__n24834 & new_new_n52454__;
  assign new_new_n53324__ = ys__n24831 & new_new_n52457__;
  assign new_new_n53325__ = ~new_new_n53323__ & ~new_new_n53324__;
  assign new_new_n53326__ = ys__n24828 & new_new_n52456__;
  assign new_new_n53327__ = ys__n39778 & new_new_n52446__;
  assign new_new_n53328__ = ~new_new_n53326__ & ~new_new_n53327__;
  assign new_new_n53329__ = new_new_n53325__ & new_new_n53328__;
  assign new_new_n53330__ = new_new_n53322__ & new_new_n53329__;
  assign new_new_n53331__ = ~new_new_n53314__ & ~new_new_n53330__;
  assign new_new_n53332__ = ~new_new_n52443__ & ~new_new_n53330__;
  assign new_new_n53333__ = ~new_new_n53331__ & ~new_new_n53332__;
  assign new_new_n53334__ = ~new_new_n53315__ & new_new_n53333__;
  assign new_new_n53335__ = ~new_new_n53302__ & ~new_new_n53334__;
  assign new_new_n53336__ = ys__n39764 & new_new_n52359__;
  assign new_new_n53337__ = ys__n39762 & new_new_n52358__;
  assign new_new_n53338__ = ~new_new_n53336__ & ~new_new_n53337__;
  assign new_new_n53339__ = ys__n33729 & new_new_n52372__;
  assign new_new_n53340__ = ~ys__n33729 & new_new_n52375__;
  assign new_new_n53341__ = ~new_new_n53339__ & ~new_new_n53340__;
  assign new_new_n53342__ = new_new_n53338__ & new_new_n53341__;
  assign new_new_n53343__ = ys__n24816 & new_new_n52364__;
  assign new_new_n53344__ = ys__n24813 & new_new_n52367__;
  assign new_new_n53345__ = ~new_new_n53343__ & ~new_new_n53344__;
  assign new_new_n53346__ = ys__n24810 & new_new_n52366__;
  assign new_new_n53347__ = ys__n39766 & new_new_n52356__;
  assign new_new_n53348__ = ~new_new_n53346__ & ~new_new_n53347__;
  assign new_new_n53349__ = new_new_n53345__ & new_new_n53348__;
  assign new_new_n53350__ = new_new_n53342__ & new_new_n53349__;
  assign new_new_n53351__ = ys__n39770 & new_new_n52334__;
  assign new_new_n53352__ = ys__n39768 & new_new_n52333__;
  assign new_new_n53353__ = ~new_new_n53351__ & ~new_new_n53352__;
  assign new_new_n53354__ = ys__n33735 & new_new_n52347__;
  assign new_new_n53355__ = ~ys__n33735 & new_new_n52350__;
  assign new_new_n53356__ = ~new_new_n53354__ & ~new_new_n53355__;
  assign new_new_n53357__ = new_new_n53353__ & new_new_n53356__;
  assign new_new_n53358__ = ys__n24825 & new_new_n52339__;
  assign new_new_n53359__ = ys__n24822 & new_new_n52342__;
  assign new_new_n53360__ = ~new_new_n53358__ & ~new_new_n53359__;
  assign new_new_n53361__ = ys__n24819 & new_new_n52341__;
  assign new_new_n53362__ = ys__n39772 & new_new_n52331__;
  assign new_new_n53363__ = ~new_new_n53361__ & ~new_new_n53362__;
  assign new_new_n53364__ = new_new_n53360__ & new_new_n53363__;
  assign new_new_n53365__ = new_new_n53357__ & new_new_n53364__;
  assign new_new_n53366__ = ~new_new_n53350__ & ~new_new_n53365__;
  assign new_new_n53367__ = ys__n24807 & new_new_n52383__;
  assign new_new_n53368__ = ys__n24804 & new_new_n52384__;
  assign new_new_n53369__ = ~new_new_n53367__ & ~new_new_n53368__;
  assign new_new_n53370__ = ys__n39760 & new_new_n52391__;
  assign new_new_n53371__ = ys__n39758 & new_new_n52392__;
  assign new_new_n53372__ = ~new_new_n53370__ & ~new_new_n53371__;
  assign new_new_n53373__ = new_new_n53369__ & new_new_n53372__;
  assign new_new_n53374__ = ~new_new_n53350__ & ~new_new_n53373__;
  assign new_new_n53375__ = ~new_new_n53365__ & ~new_new_n53373__;
  assign new_new_n53376__ = ~new_new_n53374__ & ~new_new_n53375__;
  assign new_new_n53377__ = ~new_new_n53366__ & new_new_n53376__;
  assign new_new_n53378__ = ~new_new_n53302__ & ~new_new_n53377__;
  assign new_new_n53379__ = ~new_new_n53334__ & ~new_new_n53377__;
  assign new_new_n53380__ = ~new_new_n53378__ & ~new_new_n53379__;
  assign new_new_n53381__ = ~new_new_n53335__ & new_new_n53380__;
  assign new_new_n53382__ = ~new_new_n53281__ & ~new_new_n53381__;
  assign new_new_n53383__ = ~new_new_n53291__ & ~new_new_n53381__;
  assign new_new_n53384__ = ~new_new_n53382__ & ~new_new_n53383__;
  assign ys__n42594 = new_new_n53292__ | ~new_new_n53384__;
  assign new_new_n53386__ = ~new_new_n53291__ & new_new_n53382__;
  assign new_new_n53387__ = new_new_n53291__ & ~new_new_n53381__;
  assign new_new_n53388__ = new_new_n53281__ & new_new_n53387__;
  assign new_new_n53389__ = ~new_new_n53291__ & new_new_n53381__;
  assign new_new_n53390__ = new_new_n53281__ & new_new_n53389__;
  assign new_new_n53391__ = new_new_n53291__ & new_new_n53381__;
  assign new_new_n53392__ = ~new_new_n53281__ & new_new_n53391__;
  assign new_new_n53393__ = ~new_new_n53390__ & ~new_new_n53392__;
  assign new_new_n53394__ = ~new_new_n53388__ & new_new_n53393__;
  assign ys__n42599 = new_new_n53386__ | ~new_new_n53394__;
  assign new_new_n53396__ = ~new_new_n53334__ & new_new_n53378__;
  assign new_new_n53397__ = new_new_n53302__ & new_new_n53377__;
  assign new_new_n53398__ = ~new_new_n53334__ & new_new_n53397__;
  assign new_new_n53399__ = ~new_new_n53396__ & ~new_new_n53398__;
  assign new_new_n53400__ = ~new_new_n53302__ & new_new_n53377__;
  assign new_new_n53401__ = new_new_n53334__ & new_new_n53400__;
  assign new_new_n53402__ = new_new_n53302__ & ~new_new_n53377__;
  assign new_new_n53403__ = new_new_n53334__ & new_new_n53402__;
  assign new_new_n53404__ = ~new_new_n53401__ & ~new_new_n53403__;
  assign new_new_n53405__ = new_new_n53399__ & new_new_n53404__;
  assign new_new_n53406__ = ~new_new_n52443__ & new_new_n53208__;
  assign new_new_n53407__ = new_new_n52432__ & new_new_n53206__;
  assign new_new_n53408__ = ~new_new_n52443__ & new_new_n53407__;
  assign new_new_n53409__ = ~new_new_n53406__ & ~new_new_n53408__;
  assign new_new_n53410__ = ~new_new_n52432__ & new_new_n53206__;
  assign new_new_n53411__ = new_new_n52443__ & new_new_n53410__;
  assign new_new_n53412__ = new_new_n52432__ & ~new_new_n53206__;
  assign new_new_n53413__ = new_new_n52443__ & new_new_n53412__;
  assign new_new_n53414__ = ~new_new_n53411__ & ~new_new_n53413__;
  assign new_new_n53415__ = new_new_n53409__ & new_new_n53414__;
  assign new_new_n53416__ = ~new_new_n53405__ & ~new_new_n53415__;
  assign new_new_n53417__ = ~new_new_n53365__ & new_new_n53374__;
  assign new_new_n53418__ = new_new_n53350__ & new_new_n53373__;
  assign new_new_n53419__ = ~new_new_n53365__ & new_new_n53418__;
  assign new_new_n53420__ = ~new_new_n53417__ & ~new_new_n53419__;
  assign new_new_n53421__ = ~new_new_n53350__ & new_new_n53373__;
  assign new_new_n53422__ = new_new_n53365__ & new_new_n53421__;
  assign new_new_n53423__ = new_new_n53350__ & ~new_new_n53373__;
  assign new_new_n53424__ = new_new_n53365__ & new_new_n53423__;
  assign new_new_n53425__ = ~new_new_n53422__ & ~new_new_n53424__;
  assign new_new_n53426__ = new_new_n53420__ & new_new_n53425__;
  assign new_new_n53427__ = ys__n24834 & new_new_n52419__;
  assign new_new_n53428__ = ys__n39778 & new_new_n52411__;
  assign new_new_n53429__ = ~new_new_n53427__ & ~new_new_n53428__;
  assign new_new_n53430__ = ys__n33745 & new_new_n52425__;
  assign new_new_n53431__ = ~ys__n33745 & new_new_n52428__;
  assign new_new_n53432__ = ~new_new_n53430__ & ~new_new_n53431__;
  assign new_new_n53433__ = new_new_n53429__ & new_new_n53432__;
  assign new_new_n53434__ = ~new_new_n53304__ & ~new_new_n53306__;
  assign new_new_n53435__ = new_new_n53312__ & new_new_n53434__;
  assign new_new_n53436__ = new_new_n53433__ & new_new_n53435__;
  assign new_new_n53437__ = ~new_new_n52443__ & ~new_new_n53436__;
  assign new_new_n53438__ = ys__n39774 & new_new_n52449__;
  assign new_new_n53439__ = ys__n39772 & new_new_n52448__;
  assign new_new_n53440__ = ~new_new_n53438__ & ~new_new_n53439__;
  assign new_new_n53441__ = ys__n33739 & new_new_n52462__;
  assign new_new_n53442__ = ~ys__n33739 & new_new_n52465__;
  assign new_new_n53443__ = ~new_new_n53441__ & ~new_new_n53442__;
  assign new_new_n53444__ = new_new_n53440__ & new_new_n53443__;
  assign new_new_n53445__ = ys__n24831 & new_new_n52454__;
  assign new_new_n53446__ = ys__n24828 & new_new_n52457__;
  assign new_new_n53447__ = ~new_new_n53445__ & ~new_new_n53446__;
  assign new_new_n53448__ = ys__n24825 & new_new_n52456__;
  assign new_new_n53449__ = ys__n39776 & new_new_n52446__;
  assign new_new_n53450__ = ~new_new_n53448__ & ~new_new_n53449__;
  assign new_new_n53451__ = new_new_n53447__ & new_new_n53450__;
  assign new_new_n53452__ = new_new_n53444__ & new_new_n53451__;
  assign new_new_n53453__ = ~new_new_n53436__ & ~new_new_n53452__;
  assign new_new_n53454__ = ~new_new_n52443__ & ~new_new_n53452__;
  assign new_new_n53455__ = ~new_new_n53453__ & ~new_new_n53454__;
  assign new_new_n53456__ = ~new_new_n53437__ & new_new_n53455__;
  assign new_new_n53457__ = ~new_new_n53426__ & ~new_new_n53456__;
  assign new_new_n53458__ = ys__n39762 & new_new_n52359__;
  assign new_new_n53459__ = ys__n39760 & new_new_n52358__;
  assign new_new_n53460__ = ~new_new_n53458__ & ~new_new_n53459__;
  assign new_new_n53461__ = ys__n33727 & new_new_n52372__;
  assign new_new_n53462__ = ~ys__n33727 & new_new_n52375__;
  assign new_new_n53463__ = ~new_new_n53461__ & ~new_new_n53462__;
  assign new_new_n53464__ = new_new_n53460__ & new_new_n53463__;
  assign new_new_n53465__ = ys__n24813 & new_new_n52364__;
  assign new_new_n53466__ = ys__n24810 & new_new_n52367__;
  assign new_new_n53467__ = ~new_new_n53465__ & ~new_new_n53466__;
  assign new_new_n53468__ = ys__n24807 & new_new_n52366__;
  assign new_new_n53469__ = ys__n39764 & new_new_n52356__;
  assign new_new_n53470__ = ~new_new_n53468__ & ~new_new_n53469__;
  assign new_new_n53471__ = new_new_n53467__ & new_new_n53470__;
  assign new_new_n53472__ = new_new_n53464__ & new_new_n53471__;
  assign new_new_n53473__ = ys__n39768 & new_new_n52334__;
  assign new_new_n53474__ = ys__n39766 & new_new_n52333__;
  assign new_new_n53475__ = ~new_new_n53473__ & ~new_new_n53474__;
  assign new_new_n53476__ = ys__n33733 & new_new_n52347__;
  assign new_new_n53477__ = ~ys__n33733 & new_new_n52350__;
  assign new_new_n53478__ = ~new_new_n53476__ & ~new_new_n53477__;
  assign new_new_n53479__ = new_new_n53475__ & new_new_n53478__;
  assign new_new_n53480__ = ys__n24822 & new_new_n52339__;
  assign new_new_n53481__ = ys__n24819 & new_new_n52342__;
  assign new_new_n53482__ = ~new_new_n53480__ & ~new_new_n53481__;
  assign new_new_n53483__ = ys__n24816 & new_new_n52341__;
  assign new_new_n53484__ = ys__n39770 & new_new_n52331__;
  assign new_new_n53485__ = ~new_new_n53483__ & ~new_new_n53484__;
  assign new_new_n53486__ = new_new_n53482__ & new_new_n53485__;
  assign new_new_n53487__ = new_new_n53479__ & new_new_n53486__;
  assign new_new_n53488__ = ~new_new_n53472__ & ~new_new_n53487__;
  assign new_new_n53489__ = ys__n24804 & new_new_n52383__;
  assign new_new_n53490__ = ys__n24801 & new_new_n52384__;
  assign new_new_n53491__ = ~new_new_n53489__ & ~new_new_n53490__;
  assign new_new_n53492__ = ys__n39758 & new_new_n52391__;
  assign new_new_n53493__ = ys__n39756 & new_new_n52392__;
  assign new_new_n53494__ = ~new_new_n53492__ & ~new_new_n53493__;
  assign new_new_n53495__ = new_new_n53491__ & new_new_n53494__;
  assign new_new_n53496__ = ~new_new_n53472__ & ~new_new_n53495__;
  assign new_new_n53497__ = ~new_new_n53487__ & ~new_new_n53495__;
  assign new_new_n53498__ = ~new_new_n53496__ & ~new_new_n53497__;
  assign new_new_n53499__ = ~new_new_n53488__ & new_new_n53498__;
  assign new_new_n53500__ = ~new_new_n53426__ & ~new_new_n53499__;
  assign new_new_n53501__ = ~new_new_n53456__ & ~new_new_n53499__;
  assign new_new_n53502__ = ~new_new_n53500__ & ~new_new_n53501__;
  assign new_new_n53503__ = ~new_new_n53457__ & new_new_n53502__;
  assign new_new_n53504__ = ~new_new_n53405__ & ~new_new_n53503__;
  assign new_new_n53505__ = ~new_new_n53415__ & ~new_new_n53503__;
  assign new_new_n53506__ = ~new_new_n53504__ & ~new_new_n53505__;
  assign ys__n42647 = new_new_n53416__ | ~new_new_n53506__;
  assign new_new_n53508__ = ~new_new_n53415__ & new_new_n53504__;
  assign new_new_n53509__ = new_new_n53415__ & ~new_new_n53503__;
  assign new_new_n53510__ = new_new_n53405__ & new_new_n53509__;
  assign new_new_n53511__ = ~new_new_n53415__ & new_new_n53503__;
  assign new_new_n53512__ = new_new_n53405__ & new_new_n53511__;
  assign new_new_n53513__ = new_new_n53415__ & new_new_n53503__;
  assign new_new_n53514__ = ~new_new_n53405__ & new_new_n53513__;
  assign new_new_n53515__ = ~new_new_n53512__ & ~new_new_n53514__;
  assign new_new_n53516__ = ~new_new_n53510__ & new_new_n53515__;
  assign ys__n42652 = new_new_n53508__ | ~new_new_n53516__;
  assign new_new_n53518__ = ~new_new_n53456__ & new_new_n53500__;
  assign new_new_n53519__ = new_new_n53426__ & new_new_n53499__;
  assign new_new_n53520__ = ~new_new_n53456__ & new_new_n53519__;
  assign new_new_n53521__ = ~new_new_n53518__ & ~new_new_n53520__;
  assign new_new_n53522__ = ~new_new_n53426__ & new_new_n53499__;
  assign new_new_n53523__ = new_new_n53456__ & new_new_n53522__;
  assign new_new_n53524__ = new_new_n53426__ & ~new_new_n53499__;
  assign new_new_n53525__ = new_new_n53456__ & new_new_n53524__;
  assign new_new_n53526__ = ~new_new_n53523__ & ~new_new_n53525__;
  assign new_new_n53527__ = new_new_n53521__ & new_new_n53526__;
  assign new_new_n53528__ = ~new_new_n52443__ & new_new_n53331__;
  assign new_new_n53529__ = new_new_n53314__ & new_new_n53330__;
  assign new_new_n53530__ = ~new_new_n52443__ & new_new_n53529__;
  assign new_new_n53531__ = ~new_new_n53528__ & ~new_new_n53530__;
  assign new_new_n53532__ = ~new_new_n53314__ & new_new_n53330__;
  assign new_new_n53533__ = new_new_n52443__ & new_new_n53532__;
  assign new_new_n53534__ = new_new_n53314__ & ~new_new_n53330__;
  assign new_new_n53535__ = new_new_n52443__ & new_new_n53534__;
  assign new_new_n53536__ = ~new_new_n53533__ & ~new_new_n53535__;
  assign new_new_n53537__ = new_new_n53531__ & new_new_n53536__;
  assign new_new_n53538__ = ~new_new_n53527__ & ~new_new_n53537__;
  assign new_new_n53539__ = ~new_new_n53487__ & new_new_n53496__;
  assign new_new_n53540__ = new_new_n53472__ & new_new_n53495__;
  assign new_new_n53541__ = ~new_new_n53487__ & new_new_n53540__;
  assign new_new_n53542__ = ~new_new_n53539__ & ~new_new_n53541__;
  assign new_new_n53543__ = ~new_new_n53472__ & new_new_n53495__;
  assign new_new_n53544__ = new_new_n53487__ & new_new_n53543__;
  assign new_new_n53545__ = new_new_n53472__ & ~new_new_n53495__;
  assign new_new_n53546__ = new_new_n53487__ & new_new_n53545__;
  assign new_new_n53547__ = ~new_new_n53544__ & ~new_new_n53546__;
  assign new_new_n53548__ = new_new_n53542__ & new_new_n53547__;
  assign new_new_n53549__ = ys__n39778 & new_new_n52412__;
  assign new_new_n53550__ = ys__n39776 & new_new_n52411__;
  assign new_new_n53551__ = ~new_new_n53549__ & ~new_new_n53550__;
  assign new_new_n53552__ = ys__n33743 & new_new_n52425__;
  assign new_new_n53553__ = ~ys__n33743 & new_new_n52428__;
  assign new_new_n53554__ = ~new_new_n53552__ & ~new_new_n53553__;
  assign new_new_n53555__ = new_new_n53551__ & new_new_n53554__;
  assign new_new_n53556__ = ~new_new_n53304__ & ~new_new_n53310__;
  assign new_new_n53557__ = ys__n24834 & new_new_n52420__;
  assign new_new_n53558__ = ys__n24831 & new_new_n52419__;
  assign new_new_n53559__ = ~new_new_n53557__ & ~new_new_n53558__;
  assign new_new_n53560__ = new_new_n53556__ & new_new_n53559__;
  assign new_new_n53561__ = new_new_n53555__ & new_new_n53560__;
  assign new_new_n53562__ = ~new_new_n52443__ & ~new_new_n53561__;
  assign new_new_n53563__ = ys__n39772 & new_new_n52449__;
  assign new_new_n53564__ = ys__n39770 & new_new_n52448__;
  assign new_new_n53565__ = ~new_new_n53563__ & ~new_new_n53564__;
  assign new_new_n53566__ = ys__n33737 & new_new_n52462__;
  assign new_new_n53567__ = ~ys__n33737 & new_new_n52465__;
  assign new_new_n53568__ = ~new_new_n53566__ & ~new_new_n53567__;
  assign new_new_n53569__ = new_new_n53565__ & new_new_n53568__;
  assign new_new_n53570__ = ys__n24828 & new_new_n52454__;
  assign new_new_n53571__ = ys__n24825 & new_new_n52457__;
  assign new_new_n53572__ = ~new_new_n53570__ & ~new_new_n53571__;
  assign new_new_n53573__ = ys__n24822 & new_new_n52456__;
  assign new_new_n53574__ = ys__n39774 & new_new_n52446__;
  assign new_new_n53575__ = ~new_new_n53573__ & ~new_new_n53574__;
  assign new_new_n53576__ = new_new_n53572__ & new_new_n53575__;
  assign new_new_n53577__ = new_new_n53569__ & new_new_n53576__;
  assign new_new_n53578__ = ~new_new_n53561__ & ~new_new_n53577__;
  assign new_new_n53579__ = ~new_new_n52443__ & ~new_new_n53577__;
  assign new_new_n53580__ = ~new_new_n53578__ & ~new_new_n53579__;
  assign new_new_n53581__ = ~new_new_n53562__ & new_new_n53580__;
  assign new_new_n53582__ = ~new_new_n53548__ & ~new_new_n53581__;
  assign new_new_n53583__ = ys__n39760 & new_new_n52359__;
  assign new_new_n53584__ = ys__n39758 & new_new_n52358__;
  assign new_new_n53585__ = ~new_new_n53583__ & ~new_new_n53584__;
  assign new_new_n53586__ = ys__n33725 & new_new_n52372__;
  assign new_new_n53587__ = ~ys__n33725 & new_new_n52375__;
  assign new_new_n53588__ = ~new_new_n53586__ & ~new_new_n53587__;
  assign new_new_n53589__ = new_new_n53585__ & new_new_n53588__;
  assign new_new_n53590__ = ys__n24810 & new_new_n52364__;
  assign new_new_n53591__ = ys__n24807 & new_new_n52367__;
  assign new_new_n53592__ = ~new_new_n53590__ & ~new_new_n53591__;
  assign new_new_n53593__ = ys__n24804 & new_new_n52366__;
  assign new_new_n53594__ = ys__n39762 & new_new_n52356__;
  assign new_new_n53595__ = ~new_new_n53593__ & ~new_new_n53594__;
  assign new_new_n53596__ = new_new_n53592__ & new_new_n53595__;
  assign new_new_n53597__ = new_new_n53589__ & new_new_n53596__;
  assign new_new_n53598__ = ys__n39766 & new_new_n52334__;
  assign new_new_n53599__ = ys__n39764 & new_new_n52333__;
  assign new_new_n53600__ = ~new_new_n53598__ & ~new_new_n53599__;
  assign new_new_n53601__ = ys__n33731 & new_new_n52347__;
  assign new_new_n53602__ = ~ys__n33731 & new_new_n52350__;
  assign new_new_n53603__ = ~new_new_n53601__ & ~new_new_n53602__;
  assign new_new_n53604__ = new_new_n53600__ & new_new_n53603__;
  assign new_new_n53605__ = ys__n24819 & new_new_n52339__;
  assign new_new_n53606__ = ys__n24816 & new_new_n52342__;
  assign new_new_n53607__ = ~new_new_n53605__ & ~new_new_n53606__;
  assign new_new_n53608__ = ys__n24813 & new_new_n52341__;
  assign new_new_n53609__ = ys__n39768 & new_new_n52331__;
  assign new_new_n53610__ = ~new_new_n53608__ & ~new_new_n53609__;
  assign new_new_n53611__ = new_new_n53607__ & new_new_n53610__;
  assign new_new_n53612__ = new_new_n53604__ & new_new_n53611__;
  assign new_new_n53613__ = ~new_new_n53597__ & ~new_new_n53612__;
  assign new_new_n53614__ = ys__n24801 & new_new_n52383__;
  assign new_new_n53615__ = ys__n24798 & new_new_n52384__;
  assign new_new_n53616__ = ~new_new_n53614__ & ~new_new_n53615__;
  assign new_new_n53617__ = ys__n39756 & new_new_n52391__;
  assign new_new_n53618__ = ys__n39754 & new_new_n52392__;
  assign new_new_n53619__ = ~new_new_n53617__ & ~new_new_n53618__;
  assign new_new_n53620__ = new_new_n53616__ & new_new_n53619__;
  assign new_new_n53621__ = ~new_new_n53597__ & ~new_new_n53620__;
  assign new_new_n53622__ = ~new_new_n53612__ & ~new_new_n53620__;
  assign new_new_n53623__ = ~new_new_n53621__ & ~new_new_n53622__;
  assign new_new_n53624__ = ~new_new_n53613__ & new_new_n53623__;
  assign new_new_n53625__ = ~new_new_n53548__ & ~new_new_n53624__;
  assign new_new_n53626__ = ~new_new_n53581__ & ~new_new_n53624__;
  assign new_new_n53627__ = ~new_new_n53625__ & ~new_new_n53626__;
  assign new_new_n53628__ = ~new_new_n53582__ & new_new_n53627__;
  assign new_new_n53629__ = ~new_new_n53527__ & ~new_new_n53628__;
  assign new_new_n53630__ = ~new_new_n53537__ & ~new_new_n53628__;
  assign new_new_n53631__ = ~new_new_n53629__ & ~new_new_n53630__;
  assign ys__n42701 = new_new_n53538__ | ~new_new_n53631__;
  assign new_new_n53633__ = ~new_new_n53537__ & new_new_n53629__;
  assign new_new_n53634__ = new_new_n53537__ & ~new_new_n53628__;
  assign new_new_n53635__ = new_new_n53527__ & new_new_n53634__;
  assign new_new_n53636__ = ~new_new_n53537__ & new_new_n53628__;
  assign new_new_n53637__ = new_new_n53527__ & new_new_n53636__;
  assign new_new_n53638__ = new_new_n53537__ & new_new_n53628__;
  assign new_new_n53639__ = ~new_new_n53527__ & new_new_n53638__;
  assign new_new_n53640__ = ~new_new_n53637__ & ~new_new_n53639__;
  assign new_new_n53641__ = ~new_new_n53635__ & new_new_n53640__;
  assign ys__n42706 = new_new_n53633__ | ~new_new_n53641__;
  assign new_new_n53643__ = ~new_new_n53581__ & new_new_n53625__;
  assign new_new_n53644__ = new_new_n53548__ & new_new_n53624__;
  assign new_new_n53645__ = ~new_new_n53581__ & new_new_n53644__;
  assign new_new_n53646__ = ~new_new_n53643__ & ~new_new_n53645__;
  assign new_new_n53647__ = ~new_new_n53548__ & new_new_n53624__;
  assign new_new_n53648__ = new_new_n53581__ & new_new_n53647__;
  assign new_new_n53649__ = new_new_n53548__ & ~new_new_n53624__;
  assign new_new_n53650__ = new_new_n53581__ & new_new_n53649__;
  assign new_new_n53651__ = ~new_new_n53648__ & ~new_new_n53650__;
  assign new_new_n53652__ = new_new_n53646__ & new_new_n53651__;
  assign new_new_n53653__ = ~new_new_n52443__ & new_new_n53453__;
  assign new_new_n53654__ = new_new_n53436__ & new_new_n53452__;
  assign new_new_n53655__ = ~new_new_n52443__ & new_new_n53654__;
  assign new_new_n53656__ = ~new_new_n53653__ & ~new_new_n53655__;
  assign new_new_n53657__ = ~new_new_n53436__ & new_new_n53452__;
  assign new_new_n53658__ = new_new_n52443__ & new_new_n53657__;
  assign new_new_n53659__ = new_new_n53436__ & ~new_new_n53452__;
  assign new_new_n53660__ = new_new_n52443__ & new_new_n53659__;
  assign new_new_n53661__ = ~new_new_n53658__ & ~new_new_n53660__;
  assign new_new_n53662__ = new_new_n53656__ & new_new_n53661__;
  assign new_new_n53663__ = ~new_new_n53652__ & ~new_new_n53662__;
  assign new_new_n53664__ = ~new_new_n53612__ & new_new_n53621__;
  assign new_new_n53665__ = new_new_n53597__ & new_new_n53620__;
  assign new_new_n53666__ = ~new_new_n53612__ & new_new_n53665__;
  assign new_new_n53667__ = ~new_new_n53664__ & ~new_new_n53666__;
  assign new_new_n53668__ = ~new_new_n53597__ & new_new_n53620__;
  assign new_new_n53669__ = new_new_n53612__ & new_new_n53668__;
  assign new_new_n53670__ = new_new_n53597__ & ~new_new_n53620__;
  assign new_new_n53671__ = new_new_n53612__ & new_new_n53670__;
  assign new_new_n53672__ = ~new_new_n53669__ & ~new_new_n53671__;
  assign new_new_n53673__ = new_new_n53667__ & new_new_n53672__;
  assign new_new_n53674__ = ys__n39776 & new_new_n52412__;
  assign new_new_n53675__ = ys__n39774 & new_new_n52411__;
  assign new_new_n53676__ = ~new_new_n53674__ & ~new_new_n53675__;
  assign new_new_n53677__ = ys__n33741 & new_new_n52425__;
  assign new_new_n53678__ = ~ys__n33741 & new_new_n52428__;
  assign new_new_n53679__ = ~new_new_n53677__ & ~new_new_n53678__;
  assign new_new_n53680__ = new_new_n53676__ & new_new_n53679__;
  assign new_new_n53681__ = ys__n24834 & new_new_n52417__;
  assign new_new_n53682__ = ys__n24831 & new_new_n52420__;
  assign new_new_n53683__ = ~new_new_n53681__ & ~new_new_n53682__;
  assign new_new_n53684__ = ys__n24828 & new_new_n52419__;
  assign new_new_n53685__ = ys__n39778 & new_new_n52409__;
  assign new_new_n53686__ = ~new_new_n53684__ & ~new_new_n53685__;
  assign new_new_n53687__ = new_new_n53683__ & new_new_n53686__;
  assign new_new_n53688__ = new_new_n53680__ & new_new_n53687__;
  assign new_new_n53689__ = ys__n39518 & new_new_n52322__;
  assign new_new_n53690__ = ys__n39520 & new_new_n52324__;
  assign new_new_n53691__ = ~new_new_n53689__ & ~new_new_n53690__;
  assign new_new_n53692__ = ys__n39520 & new_new_n52301__;
  assign new_new_n53693__ = ys__n39520 & new_new_n52304__;
  assign new_new_n53694__ = ~new_new_n53692__ & ~new_new_n53693__;
  assign new_new_n53695__ = new_new_n53691__ & new_new_n53694__;
  assign new_new_n53696__ = ys__n39518 & new_new_n52316__;
  assign new_new_n53697__ = ys__n39518 & new_new_n52318__;
  assign new_new_n53698__ = ~new_new_n53696__ & ~new_new_n53697__;
  assign new_new_n53699__ = new_new_n52441__ & new_new_n53698__;
  assign new_new_n53700__ = new_new_n53695__ & new_new_n53699__;
  assign new_new_n53701__ = ~new_new_n53688__ & ~new_new_n53700__;
  assign new_new_n53702__ = ys__n39770 & new_new_n52449__;
  assign new_new_n53703__ = ys__n39768 & new_new_n52448__;
  assign new_new_n53704__ = ~new_new_n53702__ & ~new_new_n53703__;
  assign new_new_n53705__ = ys__n33735 & new_new_n52462__;
  assign new_new_n53706__ = ~ys__n33735 & new_new_n52465__;
  assign new_new_n53707__ = ~new_new_n53705__ & ~new_new_n53706__;
  assign new_new_n53708__ = new_new_n53704__ & new_new_n53707__;
  assign new_new_n53709__ = ys__n24825 & new_new_n52454__;
  assign new_new_n53710__ = ys__n24822 & new_new_n52457__;
  assign new_new_n53711__ = ~new_new_n53709__ & ~new_new_n53710__;
  assign new_new_n53712__ = ys__n24819 & new_new_n52456__;
  assign new_new_n53713__ = ys__n39772 & new_new_n52446__;
  assign new_new_n53714__ = ~new_new_n53712__ & ~new_new_n53713__;
  assign new_new_n53715__ = new_new_n53711__ & new_new_n53714__;
  assign new_new_n53716__ = new_new_n53708__ & new_new_n53715__;
  assign new_new_n53717__ = ~new_new_n53688__ & ~new_new_n53716__;
  assign new_new_n53718__ = ~new_new_n53700__ & ~new_new_n53716__;
  assign new_new_n53719__ = ~new_new_n53717__ & ~new_new_n53718__;
  assign new_new_n53720__ = ~new_new_n53701__ & new_new_n53719__;
  assign new_new_n53721__ = ~new_new_n53673__ & ~new_new_n53720__;
  assign new_new_n53722__ = ys__n39758 & new_new_n52359__;
  assign new_new_n53723__ = ys__n39756 & new_new_n52358__;
  assign new_new_n53724__ = ~new_new_n53722__ & ~new_new_n53723__;
  assign new_new_n53725__ = ys__n33723 & new_new_n52372__;
  assign new_new_n53726__ = ~ys__n33723 & new_new_n52375__;
  assign new_new_n53727__ = ~new_new_n53725__ & ~new_new_n53726__;
  assign new_new_n53728__ = new_new_n53724__ & new_new_n53727__;
  assign new_new_n53729__ = ys__n24807 & new_new_n52364__;
  assign new_new_n53730__ = ys__n24804 & new_new_n52367__;
  assign new_new_n53731__ = ~new_new_n53729__ & ~new_new_n53730__;
  assign new_new_n53732__ = ys__n24801 & new_new_n52366__;
  assign new_new_n53733__ = ys__n39760 & new_new_n52356__;
  assign new_new_n53734__ = ~new_new_n53732__ & ~new_new_n53733__;
  assign new_new_n53735__ = new_new_n53731__ & new_new_n53734__;
  assign new_new_n53736__ = new_new_n53728__ & new_new_n53735__;
  assign new_new_n53737__ = ys__n39764 & new_new_n52334__;
  assign new_new_n53738__ = ys__n39762 & new_new_n52333__;
  assign new_new_n53739__ = ~new_new_n53737__ & ~new_new_n53738__;
  assign new_new_n53740__ = ys__n33729 & new_new_n52347__;
  assign new_new_n53741__ = ~ys__n33729 & new_new_n52350__;
  assign new_new_n53742__ = ~new_new_n53740__ & ~new_new_n53741__;
  assign new_new_n53743__ = new_new_n53739__ & new_new_n53742__;
  assign new_new_n53744__ = ys__n24816 & new_new_n52339__;
  assign new_new_n53745__ = ys__n24813 & new_new_n52342__;
  assign new_new_n53746__ = ~new_new_n53744__ & ~new_new_n53745__;
  assign new_new_n53747__ = ys__n24810 & new_new_n52341__;
  assign new_new_n53748__ = ys__n39766 & new_new_n52331__;
  assign new_new_n53749__ = ~new_new_n53747__ & ~new_new_n53748__;
  assign new_new_n53750__ = new_new_n53746__ & new_new_n53749__;
  assign new_new_n53751__ = new_new_n53743__ & new_new_n53750__;
  assign new_new_n53752__ = ~new_new_n53736__ & ~new_new_n53751__;
  assign new_new_n53753__ = ys__n24798 & new_new_n52383__;
  assign new_new_n53754__ = ys__n24795 & new_new_n52384__;
  assign new_new_n53755__ = ~new_new_n53753__ & ~new_new_n53754__;
  assign new_new_n53756__ = ys__n39754 & new_new_n52391__;
  assign new_new_n53757__ = ys__n39752 & new_new_n52392__;
  assign new_new_n53758__ = ~new_new_n53756__ & ~new_new_n53757__;
  assign new_new_n53759__ = new_new_n53755__ & new_new_n53758__;
  assign new_new_n53760__ = ~new_new_n53736__ & ~new_new_n53759__;
  assign new_new_n53761__ = ~new_new_n53751__ & ~new_new_n53759__;
  assign new_new_n53762__ = ~new_new_n53760__ & ~new_new_n53761__;
  assign new_new_n53763__ = ~new_new_n53752__ & new_new_n53762__;
  assign new_new_n53764__ = ~new_new_n53673__ & ~new_new_n53763__;
  assign new_new_n53765__ = ~new_new_n53720__ & ~new_new_n53763__;
  assign new_new_n53766__ = ~new_new_n53764__ & ~new_new_n53765__;
  assign new_new_n53767__ = ~new_new_n53721__ & new_new_n53766__;
  assign new_new_n53768__ = ~new_new_n53652__ & ~new_new_n53767__;
  assign new_new_n53769__ = ~new_new_n53662__ & ~new_new_n53767__;
  assign new_new_n53770__ = ~new_new_n53768__ & ~new_new_n53769__;
  assign ys__n42755 = new_new_n53663__ | ~new_new_n53770__;
  assign new_new_n53772__ = ~new_new_n53662__ & new_new_n53768__;
  assign new_new_n53773__ = new_new_n53662__ & ~new_new_n53767__;
  assign new_new_n53774__ = new_new_n53652__ & new_new_n53773__;
  assign new_new_n53775__ = ~new_new_n53662__ & new_new_n53767__;
  assign new_new_n53776__ = new_new_n53652__ & new_new_n53775__;
  assign new_new_n53777__ = new_new_n53662__ & new_new_n53767__;
  assign new_new_n53778__ = ~new_new_n53652__ & new_new_n53777__;
  assign new_new_n53779__ = ~new_new_n53776__ & ~new_new_n53778__;
  assign new_new_n53780__ = ~new_new_n53774__ & new_new_n53779__;
  assign ys__n42760 = new_new_n53772__ | ~new_new_n53780__;
  assign new_new_n53782__ = ~new_new_n53720__ & new_new_n53764__;
  assign new_new_n53783__ = new_new_n53720__ & ~new_new_n53763__;
  assign new_new_n53784__ = new_new_n53673__ & new_new_n53783__;
  assign new_new_n53785__ = ~new_new_n53720__ & new_new_n53763__;
  assign new_new_n53786__ = new_new_n53673__ & new_new_n53785__;
  assign new_new_n53787__ = new_new_n53720__ & new_new_n53763__;
  assign new_new_n53788__ = ~new_new_n53673__ & new_new_n53787__;
  assign new_new_n53789__ = ~new_new_n53786__ & ~new_new_n53788__;
  assign new_new_n53790__ = ~new_new_n53784__ & new_new_n53789__;
  assign new_new_n53791__ = ~new_new_n53782__ & new_new_n53790__;
  assign new_new_n53792__ = ~new_new_n52443__ & new_new_n53578__;
  assign new_new_n53793__ = new_new_n53561__ & new_new_n53577__;
  assign new_new_n53794__ = ~new_new_n52443__ & new_new_n53793__;
  assign new_new_n53795__ = ~new_new_n53792__ & ~new_new_n53794__;
  assign new_new_n53796__ = ~new_new_n53561__ & new_new_n53577__;
  assign new_new_n53797__ = new_new_n52443__ & new_new_n53796__;
  assign new_new_n53798__ = new_new_n53561__ & ~new_new_n53577__;
  assign new_new_n53799__ = new_new_n52443__ & new_new_n53798__;
  assign new_new_n53800__ = ~new_new_n53797__ & ~new_new_n53799__;
  assign new_new_n53801__ = new_new_n53795__ & new_new_n53800__;
  assign new_new_n53802__ = ~new_new_n53791__ & ~new_new_n53801__;
  assign new_new_n53803__ = ~new_new_n53751__ & new_new_n53760__;
  assign new_new_n53804__ = new_new_n53736__ & new_new_n53759__;
  assign new_new_n53805__ = ~new_new_n53751__ & new_new_n53804__;
  assign new_new_n53806__ = ~new_new_n53803__ & ~new_new_n53805__;
  assign new_new_n53807__ = ~new_new_n53736__ & new_new_n53759__;
  assign new_new_n53808__ = new_new_n53751__ & new_new_n53807__;
  assign new_new_n53809__ = new_new_n53736__ & ~new_new_n53759__;
  assign new_new_n53810__ = new_new_n53751__ & new_new_n53809__;
  assign new_new_n53811__ = ~new_new_n53808__ & ~new_new_n53810__;
  assign new_new_n53812__ = new_new_n53806__ & new_new_n53811__;
  assign new_new_n53813__ = ys__n39774 & new_new_n52412__;
  assign new_new_n53814__ = ys__n39772 & new_new_n52411__;
  assign new_new_n53815__ = ~new_new_n53813__ & ~new_new_n53814__;
  assign new_new_n53816__ = ys__n33739 & new_new_n52425__;
  assign new_new_n53817__ = ~ys__n33739 & new_new_n52428__;
  assign new_new_n53818__ = ~new_new_n53816__ & ~new_new_n53817__;
  assign new_new_n53819__ = new_new_n53815__ & new_new_n53818__;
  assign new_new_n53820__ = ys__n24831 & new_new_n52417__;
  assign new_new_n53821__ = ys__n24828 & new_new_n52420__;
  assign new_new_n53822__ = ~new_new_n53820__ & ~new_new_n53821__;
  assign new_new_n53823__ = ys__n24825 & new_new_n52419__;
  assign new_new_n53824__ = ys__n39776 & new_new_n52409__;
  assign new_new_n53825__ = ~new_new_n53823__ & ~new_new_n53824__;
  assign new_new_n53826__ = new_new_n53822__ & new_new_n53825__;
  assign new_new_n53827__ = new_new_n53819__ & new_new_n53826__;
  assign new_new_n53828__ = ys__n24834 & new_new_n52322__;
  assign new_new_n53829__ = ys__n39778 & new_new_n52304__;
  assign new_new_n53830__ = ~new_new_n53828__ & ~new_new_n53829__;
  assign new_new_n53831__ = ys__n33745 & new_new_n52308__;
  assign new_new_n53832__ = ~ys__n33745 & new_new_n52311__;
  assign new_new_n53833__ = ~new_new_n53831__ & ~new_new_n53832__;
  assign new_new_n53834__ = new_new_n53830__ & new_new_n53833__;
  assign new_new_n53835__ = ~new_new_n53690__ & ~new_new_n53692__;
  assign new_new_n53836__ = new_new_n53698__ & new_new_n53835__;
  assign new_new_n53837__ = new_new_n53834__ & new_new_n53836__;
  assign new_new_n53838__ = ~new_new_n53827__ & ~new_new_n53837__;
  assign new_new_n53839__ = ys__n39768 & new_new_n52449__;
  assign new_new_n53840__ = ys__n39766 & new_new_n52448__;
  assign new_new_n53841__ = ~new_new_n53839__ & ~new_new_n53840__;
  assign new_new_n53842__ = ys__n33733 & new_new_n52462__;
  assign new_new_n53843__ = ~ys__n33733 & new_new_n52465__;
  assign new_new_n53844__ = ~new_new_n53842__ & ~new_new_n53843__;
  assign new_new_n53845__ = new_new_n53841__ & new_new_n53844__;
  assign new_new_n53846__ = ys__n24822 & new_new_n52454__;
  assign new_new_n53847__ = ys__n24819 & new_new_n52457__;
  assign new_new_n53848__ = ~new_new_n53846__ & ~new_new_n53847__;
  assign new_new_n53849__ = ys__n24816 & new_new_n52456__;
  assign new_new_n53850__ = ys__n39770 & new_new_n52446__;
  assign new_new_n53851__ = ~new_new_n53849__ & ~new_new_n53850__;
  assign new_new_n53852__ = new_new_n53848__ & new_new_n53851__;
  assign new_new_n53853__ = new_new_n53845__ & new_new_n53852__;
  assign new_new_n53854__ = ~new_new_n53827__ & ~new_new_n53853__;
  assign new_new_n53855__ = ~new_new_n53837__ & ~new_new_n53853__;
  assign new_new_n53856__ = ~new_new_n53854__ & ~new_new_n53855__;
  assign new_new_n53857__ = ~new_new_n53838__ & new_new_n53856__;
  assign new_new_n53858__ = ~new_new_n53812__ & ~new_new_n53857__;
  assign new_new_n53859__ = ys__n39756 & new_new_n52359__;
  assign new_new_n53860__ = ys__n39754 & new_new_n52358__;
  assign new_new_n53861__ = ~new_new_n53859__ & ~new_new_n53860__;
  assign new_new_n53862__ = ys__n33721 & new_new_n52372__;
  assign new_new_n53863__ = ~ys__n33721 & new_new_n52375__;
  assign new_new_n53864__ = ~new_new_n53862__ & ~new_new_n53863__;
  assign new_new_n53865__ = new_new_n53861__ & new_new_n53864__;
  assign new_new_n53866__ = ys__n24804 & new_new_n52364__;
  assign new_new_n53867__ = ys__n24801 & new_new_n52367__;
  assign new_new_n53868__ = ~new_new_n53866__ & ~new_new_n53867__;
  assign new_new_n53869__ = ys__n24798 & new_new_n52366__;
  assign new_new_n53870__ = ys__n39758 & new_new_n52356__;
  assign new_new_n53871__ = ~new_new_n53869__ & ~new_new_n53870__;
  assign new_new_n53872__ = new_new_n53868__ & new_new_n53871__;
  assign new_new_n53873__ = new_new_n53865__ & new_new_n53872__;
  assign new_new_n53874__ = ys__n39762 & new_new_n52334__;
  assign new_new_n53875__ = ys__n39760 & new_new_n52333__;
  assign new_new_n53876__ = ~new_new_n53874__ & ~new_new_n53875__;
  assign new_new_n53877__ = ys__n33727 & new_new_n52347__;
  assign new_new_n53878__ = ~ys__n33727 & new_new_n52350__;
  assign new_new_n53879__ = ~new_new_n53877__ & ~new_new_n53878__;
  assign new_new_n53880__ = new_new_n53876__ & new_new_n53879__;
  assign new_new_n53881__ = ys__n24813 & new_new_n52339__;
  assign new_new_n53882__ = ys__n24810 & new_new_n52342__;
  assign new_new_n53883__ = ~new_new_n53881__ & ~new_new_n53882__;
  assign new_new_n53884__ = ys__n24807 & new_new_n52341__;
  assign new_new_n53885__ = ys__n39764 & new_new_n52331__;
  assign new_new_n53886__ = ~new_new_n53884__ & ~new_new_n53885__;
  assign new_new_n53887__ = new_new_n53883__ & new_new_n53886__;
  assign new_new_n53888__ = new_new_n53880__ & new_new_n53887__;
  assign new_new_n53889__ = ~new_new_n53873__ & ~new_new_n53888__;
  assign new_new_n53890__ = ys__n24795 & new_new_n52383__;
  assign new_new_n53891__ = ys__n24792 & new_new_n52384__;
  assign new_new_n53892__ = ~new_new_n53890__ & ~new_new_n53891__;
  assign new_new_n53893__ = ys__n39752 & new_new_n52391__;
  assign new_new_n53894__ = ys__n39750 & new_new_n52392__;
  assign new_new_n53895__ = ~new_new_n53893__ & ~new_new_n53894__;
  assign new_new_n53896__ = new_new_n53892__ & new_new_n53895__;
  assign new_new_n53897__ = ~new_new_n53873__ & ~new_new_n53896__;
  assign new_new_n53898__ = ~new_new_n53888__ & ~new_new_n53896__;
  assign new_new_n53899__ = ~new_new_n53897__ & ~new_new_n53898__;
  assign new_new_n53900__ = ~new_new_n53889__ & new_new_n53899__;
  assign new_new_n53901__ = ~new_new_n53812__ & ~new_new_n53900__;
  assign new_new_n53902__ = ~new_new_n53857__ & ~new_new_n53900__;
  assign new_new_n53903__ = ~new_new_n53901__ & ~new_new_n53902__;
  assign new_new_n53904__ = ~new_new_n53858__ & new_new_n53903__;
  assign new_new_n53905__ = ~new_new_n53791__ & ~new_new_n53904__;
  assign new_new_n53906__ = ~new_new_n53801__ & ~new_new_n53904__;
  assign new_new_n53907__ = ~new_new_n53905__ & ~new_new_n53906__;
  assign ys__n42809 = new_new_n53802__ | ~new_new_n53907__;
  assign new_new_n53909__ = ~new_new_n53801__ & new_new_n53905__;
  assign new_new_n53910__ = new_new_n53801__ & ~new_new_n53904__;
  assign new_new_n53911__ = new_new_n53791__ & new_new_n53910__;
  assign new_new_n53912__ = ~new_new_n53801__ & new_new_n53904__;
  assign new_new_n53913__ = new_new_n53791__ & new_new_n53912__;
  assign new_new_n53914__ = new_new_n53801__ & new_new_n53904__;
  assign new_new_n53915__ = ~new_new_n53791__ & new_new_n53914__;
  assign new_new_n53916__ = ~new_new_n53913__ & ~new_new_n53915__;
  assign new_new_n53917__ = ~new_new_n53911__ & new_new_n53916__;
  assign ys__n42814 = new_new_n53909__ | ~new_new_n53917__;
  assign new_new_n53919__ = ~new_new_n53857__ & new_new_n53901__;
  assign new_new_n53920__ = new_new_n53857__ & ~new_new_n53900__;
  assign new_new_n53921__ = new_new_n53812__ & new_new_n53920__;
  assign new_new_n53922__ = ~new_new_n53857__ & new_new_n53900__;
  assign new_new_n53923__ = new_new_n53812__ & new_new_n53922__;
  assign new_new_n53924__ = new_new_n53857__ & new_new_n53900__;
  assign new_new_n53925__ = ~new_new_n53812__ & new_new_n53924__;
  assign new_new_n53926__ = ~new_new_n53923__ & ~new_new_n53925__;
  assign new_new_n53927__ = ~new_new_n53921__ & new_new_n53926__;
  assign new_new_n53928__ = ~new_new_n53919__ & new_new_n53927__;
  assign new_new_n53929__ = ~new_new_n53700__ & new_new_n53717__;
  assign new_new_n53930__ = new_new_n53688__ & new_new_n53716__;
  assign new_new_n53931__ = ~new_new_n53700__ & new_new_n53930__;
  assign new_new_n53932__ = ~new_new_n53929__ & ~new_new_n53931__;
  assign new_new_n53933__ = ~new_new_n53688__ & new_new_n53716__;
  assign new_new_n53934__ = new_new_n53700__ & new_new_n53933__;
  assign new_new_n53935__ = new_new_n53688__ & ~new_new_n53716__;
  assign new_new_n53936__ = new_new_n53700__ & new_new_n53935__;
  assign new_new_n53937__ = ~new_new_n53934__ & ~new_new_n53936__;
  assign new_new_n53938__ = new_new_n53932__ & new_new_n53937__;
  assign new_new_n53939__ = ~new_new_n53928__ & ~new_new_n53938__;
  assign new_new_n53940__ = ~new_new_n53888__ & new_new_n53897__;
  assign new_new_n53941__ = new_new_n53873__ & new_new_n53896__;
  assign new_new_n53942__ = ~new_new_n53888__ & new_new_n53941__;
  assign new_new_n53943__ = ~new_new_n53940__ & ~new_new_n53942__;
  assign new_new_n53944__ = ~new_new_n53873__ & new_new_n53896__;
  assign new_new_n53945__ = new_new_n53888__ & new_new_n53944__;
  assign new_new_n53946__ = new_new_n53873__ & ~new_new_n53896__;
  assign new_new_n53947__ = new_new_n53888__ & new_new_n53946__;
  assign new_new_n53948__ = ~new_new_n53945__ & ~new_new_n53947__;
  assign new_new_n53949__ = new_new_n53943__ & new_new_n53948__;
  assign new_new_n53950__ = ys__n39772 & new_new_n52412__;
  assign new_new_n53951__ = ys__n39770 & new_new_n52411__;
  assign new_new_n53952__ = ~new_new_n53950__ & ~new_new_n53951__;
  assign new_new_n53953__ = ys__n33737 & new_new_n52425__;
  assign new_new_n53954__ = ~ys__n33737 & new_new_n52428__;
  assign new_new_n53955__ = ~new_new_n53953__ & ~new_new_n53954__;
  assign new_new_n53956__ = new_new_n53952__ & new_new_n53955__;
  assign new_new_n53957__ = ys__n24828 & new_new_n52417__;
  assign new_new_n53958__ = ys__n24825 & new_new_n52420__;
  assign new_new_n53959__ = ~new_new_n53957__ & ~new_new_n53958__;
  assign new_new_n53960__ = ys__n24822 & new_new_n52419__;
  assign new_new_n53961__ = ys__n39774 & new_new_n52409__;
  assign new_new_n53962__ = ~new_new_n53960__ & ~new_new_n53961__;
  assign new_new_n53963__ = new_new_n53959__ & new_new_n53962__;
  assign new_new_n53964__ = new_new_n53956__ & new_new_n53963__;
  assign new_new_n53965__ = ys__n39778 & new_new_n52301__;
  assign new_new_n53966__ = ys__n39776 & new_new_n52304__;
  assign new_new_n53967__ = ~new_new_n53965__ & ~new_new_n53966__;
  assign new_new_n53968__ = ys__n33743 & new_new_n52308__;
  assign new_new_n53969__ = ~ys__n33743 & new_new_n52311__;
  assign new_new_n53970__ = ~new_new_n53968__ & ~new_new_n53969__;
  assign new_new_n53971__ = new_new_n53967__ & new_new_n53970__;
  assign new_new_n53972__ = ~new_new_n53690__ & ~new_new_n53696__;
  assign new_new_n53973__ = ys__n24834 & new_new_n52318__;
  assign new_new_n53974__ = ys__n24831 & new_new_n52322__;
  assign new_new_n53975__ = ~new_new_n53973__ & ~new_new_n53974__;
  assign new_new_n53976__ = new_new_n53972__ & new_new_n53975__;
  assign new_new_n53977__ = new_new_n53971__ & new_new_n53976__;
  assign new_new_n53978__ = ~new_new_n53964__ & ~new_new_n53977__;
  assign new_new_n53979__ = ys__n39766 & new_new_n52449__;
  assign new_new_n53980__ = ys__n39764 & new_new_n52448__;
  assign new_new_n53981__ = ~new_new_n53979__ & ~new_new_n53980__;
  assign new_new_n53982__ = ys__n33731 & new_new_n52462__;
  assign new_new_n53983__ = ~ys__n33731 & new_new_n52465__;
  assign new_new_n53984__ = ~new_new_n53982__ & ~new_new_n53983__;
  assign new_new_n53985__ = new_new_n53981__ & new_new_n53984__;
  assign new_new_n53986__ = ys__n24819 & new_new_n52454__;
  assign new_new_n53987__ = ys__n24816 & new_new_n52457__;
  assign new_new_n53988__ = ~new_new_n53986__ & ~new_new_n53987__;
  assign new_new_n53989__ = ys__n24813 & new_new_n52456__;
  assign new_new_n53990__ = ys__n39768 & new_new_n52446__;
  assign new_new_n53991__ = ~new_new_n53989__ & ~new_new_n53990__;
  assign new_new_n53992__ = new_new_n53988__ & new_new_n53991__;
  assign new_new_n53993__ = new_new_n53985__ & new_new_n53992__;
  assign new_new_n53994__ = ~new_new_n53964__ & ~new_new_n53993__;
  assign new_new_n53995__ = ~new_new_n53977__ & ~new_new_n53993__;
  assign new_new_n53996__ = ~new_new_n53994__ & ~new_new_n53995__;
  assign new_new_n53997__ = ~new_new_n53978__ & new_new_n53996__;
  assign new_new_n53998__ = ~new_new_n53949__ & ~new_new_n53997__;
  assign new_new_n53999__ = ys__n39754 & new_new_n52359__;
  assign new_new_n54000__ = ys__n39752 & new_new_n52358__;
  assign new_new_n54001__ = ~new_new_n53999__ & ~new_new_n54000__;
  assign new_new_n54002__ = ys__n33719 & new_new_n52372__;
  assign new_new_n54003__ = ~ys__n33719 & new_new_n52375__;
  assign new_new_n54004__ = ~new_new_n54002__ & ~new_new_n54003__;
  assign new_new_n54005__ = new_new_n54001__ & new_new_n54004__;
  assign new_new_n54006__ = ys__n24801 & new_new_n52364__;
  assign new_new_n54007__ = ys__n24798 & new_new_n52367__;
  assign new_new_n54008__ = ~new_new_n54006__ & ~new_new_n54007__;
  assign new_new_n54009__ = ys__n24795 & new_new_n52366__;
  assign new_new_n54010__ = ys__n39756 & new_new_n52356__;
  assign new_new_n54011__ = ~new_new_n54009__ & ~new_new_n54010__;
  assign new_new_n54012__ = new_new_n54008__ & new_new_n54011__;
  assign new_new_n54013__ = new_new_n54005__ & new_new_n54012__;
  assign new_new_n54014__ = ys__n39760 & new_new_n52334__;
  assign new_new_n54015__ = ys__n39758 & new_new_n52333__;
  assign new_new_n54016__ = ~new_new_n54014__ & ~new_new_n54015__;
  assign new_new_n54017__ = ys__n33725 & new_new_n52347__;
  assign new_new_n54018__ = ~ys__n33725 & new_new_n52350__;
  assign new_new_n54019__ = ~new_new_n54017__ & ~new_new_n54018__;
  assign new_new_n54020__ = new_new_n54016__ & new_new_n54019__;
  assign new_new_n54021__ = ys__n24810 & new_new_n52339__;
  assign new_new_n54022__ = ys__n24807 & new_new_n52342__;
  assign new_new_n54023__ = ~new_new_n54021__ & ~new_new_n54022__;
  assign new_new_n54024__ = ys__n24804 & new_new_n52341__;
  assign new_new_n54025__ = ys__n39762 & new_new_n52331__;
  assign new_new_n54026__ = ~new_new_n54024__ & ~new_new_n54025__;
  assign new_new_n54027__ = new_new_n54023__ & new_new_n54026__;
  assign new_new_n54028__ = new_new_n54020__ & new_new_n54027__;
  assign new_new_n54029__ = ~new_new_n54013__ & ~new_new_n54028__;
  assign new_new_n54030__ = ys__n24792 & new_new_n52383__;
  assign new_new_n54031__ = ys__n24789 & new_new_n52384__;
  assign new_new_n54032__ = ~new_new_n54030__ & ~new_new_n54031__;
  assign new_new_n54033__ = ys__n39750 & new_new_n52391__;
  assign new_new_n54034__ = ys__n39748 & new_new_n52392__;
  assign new_new_n54035__ = ~new_new_n54033__ & ~new_new_n54034__;
  assign new_new_n54036__ = new_new_n54032__ & new_new_n54035__;
  assign new_new_n54037__ = ~new_new_n54013__ & ~new_new_n54036__;
  assign new_new_n54038__ = ~new_new_n54028__ & ~new_new_n54036__;
  assign new_new_n54039__ = ~new_new_n54037__ & ~new_new_n54038__;
  assign new_new_n54040__ = ~new_new_n54029__ & new_new_n54039__;
  assign new_new_n54041__ = ~new_new_n53949__ & ~new_new_n54040__;
  assign new_new_n54042__ = ~new_new_n53997__ & ~new_new_n54040__;
  assign new_new_n54043__ = ~new_new_n54041__ & ~new_new_n54042__;
  assign new_new_n54044__ = ~new_new_n53998__ & new_new_n54043__;
  assign new_new_n54045__ = ~new_new_n53928__ & ~new_new_n54044__;
  assign new_new_n54046__ = ~new_new_n53938__ & ~new_new_n54044__;
  assign new_new_n54047__ = ~new_new_n54045__ & ~new_new_n54046__;
  assign ys__n42863 = new_new_n53939__ | ~new_new_n54047__;
  assign new_new_n54049__ = ~new_new_n53938__ & new_new_n54045__;
  assign new_new_n54050__ = new_new_n53938__ & ~new_new_n54044__;
  assign new_new_n54051__ = new_new_n53928__ & new_new_n54050__;
  assign new_new_n54052__ = ~new_new_n53938__ & new_new_n54044__;
  assign new_new_n54053__ = new_new_n53928__ & new_new_n54052__;
  assign new_new_n54054__ = new_new_n53938__ & new_new_n54044__;
  assign new_new_n54055__ = ~new_new_n53928__ & new_new_n54054__;
  assign new_new_n54056__ = ~new_new_n54053__ & ~new_new_n54055__;
  assign new_new_n54057__ = ~new_new_n54051__ & new_new_n54056__;
  assign ys__n42868 = new_new_n54049__ | ~new_new_n54057__;
  assign new_new_n54059__ = ~new_new_n53997__ & new_new_n54041__;
  assign new_new_n54060__ = new_new_n53997__ & ~new_new_n54040__;
  assign new_new_n54061__ = new_new_n53949__ & new_new_n54060__;
  assign new_new_n54062__ = ~new_new_n53997__ & new_new_n54040__;
  assign new_new_n54063__ = new_new_n53949__ & new_new_n54062__;
  assign new_new_n54064__ = new_new_n53997__ & new_new_n54040__;
  assign new_new_n54065__ = ~new_new_n53949__ & new_new_n54064__;
  assign new_new_n54066__ = ~new_new_n54063__ & ~new_new_n54065__;
  assign new_new_n54067__ = ~new_new_n54061__ & new_new_n54066__;
  assign new_new_n54068__ = ~new_new_n54059__ & new_new_n54067__;
  assign new_new_n54069__ = ~new_new_n53837__ & new_new_n53854__;
  assign new_new_n54070__ = new_new_n53827__ & new_new_n53853__;
  assign new_new_n54071__ = ~new_new_n53837__ & new_new_n54070__;
  assign new_new_n54072__ = ~new_new_n54069__ & ~new_new_n54071__;
  assign new_new_n54073__ = ~new_new_n53827__ & new_new_n53853__;
  assign new_new_n54074__ = new_new_n53837__ & new_new_n54073__;
  assign new_new_n54075__ = new_new_n53827__ & ~new_new_n53853__;
  assign new_new_n54076__ = new_new_n53837__ & new_new_n54075__;
  assign new_new_n54077__ = ~new_new_n54074__ & ~new_new_n54076__;
  assign new_new_n54078__ = new_new_n54072__ & new_new_n54077__;
  assign new_new_n54079__ = ~new_new_n54068__ & ~new_new_n54078__;
  assign new_new_n54080__ = ~new_new_n54028__ & new_new_n54037__;
  assign new_new_n54081__ = new_new_n54013__ & new_new_n54036__;
  assign new_new_n54082__ = ~new_new_n54028__ & new_new_n54081__;
  assign new_new_n54083__ = ~new_new_n54080__ & ~new_new_n54082__;
  assign new_new_n54084__ = ~new_new_n54013__ & new_new_n54036__;
  assign new_new_n54085__ = new_new_n54028__ & new_new_n54084__;
  assign new_new_n54086__ = new_new_n54013__ & ~new_new_n54036__;
  assign new_new_n54087__ = new_new_n54028__ & new_new_n54086__;
  assign new_new_n54088__ = ~new_new_n54085__ & ~new_new_n54087__;
  assign new_new_n54089__ = new_new_n54083__ & new_new_n54088__;
  assign new_new_n54090__ = ys__n39770 & new_new_n52412__;
  assign new_new_n54091__ = ys__n39768 & new_new_n52411__;
  assign new_new_n54092__ = ~new_new_n54090__ & ~new_new_n54091__;
  assign new_new_n54093__ = ys__n33735 & new_new_n52425__;
  assign new_new_n54094__ = ~ys__n33735 & new_new_n52428__;
  assign new_new_n54095__ = ~new_new_n54093__ & ~new_new_n54094__;
  assign new_new_n54096__ = new_new_n54092__ & new_new_n54095__;
  assign new_new_n54097__ = ys__n24825 & new_new_n52417__;
  assign new_new_n54098__ = ys__n24822 & new_new_n52420__;
  assign new_new_n54099__ = ~new_new_n54097__ & ~new_new_n54098__;
  assign new_new_n54100__ = ys__n24819 & new_new_n52419__;
  assign new_new_n54101__ = ys__n39772 & new_new_n52409__;
  assign new_new_n54102__ = ~new_new_n54100__ & ~new_new_n54101__;
  assign new_new_n54103__ = new_new_n54099__ & new_new_n54102__;
  assign new_new_n54104__ = new_new_n54096__ & new_new_n54103__;
  assign new_new_n54105__ = ys__n39776 & new_new_n52301__;
  assign new_new_n54106__ = ys__n39774 & new_new_n52304__;
  assign new_new_n54107__ = ~new_new_n54105__ & ~new_new_n54106__;
  assign new_new_n54108__ = ys__n33741 & new_new_n52308__;
  assign new_new_n54109__ = ~ys__n33741 & new_new_n52311__;
  assign new_new_n54110__ = ~new_new_n54108__ & ~new_new_n54109__;
  assign new_new_n54111__ = new_new_n54107__ & new_new_n54110__;
  assign new_new_n54112__ = ys__n24834 & new_new_n52316__;
  assign new_new_n54113__ = ys__n24831 & new_new_n52318__;
  assign new_new_n54114__ = ~new_new_n54112__ & ~new_new_n54113__;
  assign new_new_n54115__ = ys__n24828 & new_new_n52322__;
  assign new_new_n54116__ = ys__n39778 & new_new_n52324__;
  assign new_new_n54117__ = ~new_new_n54115__ & ~new_new_n54116__;
  assign new_new_n54118__ = new_new_n54114__ & new_new_n54117__;
  assign new_new_n54119__ = new_new_n54111__ & new_new_n54118__;
  assign new_new_n54120__ = ~new_new_n54104__ & ~new_new_n54119__;
  assign new_new_n54121__ = ys__n39764 & new_new_n52449__;
  assign new_new_n54122__ = ys__n39762 & new_new_n52448__;
  assign new_new_n54123__ = ~new_new_n54121__ & ~new_new_n54122__;
  assign new_new_n54124__ = ys__n33729 & new_new_n52462__;
  assign new_new_n54125__ = ~ys__n33729 & new_new_n52465__;
  assign new_new_n54126__ = ~new_new_n54124__ & ~new_new_n54125__;
  assign new_new_n54127__ = new_new_n54123__ & new_new_n54126__;
  assign new_new_n54128__ = ys__n24816 & new_new_n52454__;
  assign new_new_n54129__ = ys__n24813 & new_new_n52457__;
  assign new_new_n54130__ = ~new_new_n54128__ & ~new_new_n54129__;
  assign new_new_n54131__ = ys__n24810 & new_new_n52456__;
  assign new_new_n54132__ = ys__n39766 & new_new_n52446__;
  assign new_new_n54133__ = ~new_new_n54131__ & ~new_new_n54132__;
  assign new_new_n54134__ = new_new_n54130__ & new_new_n54133__;
  assign new_new_n54135__ = new_new_n54127__ & new_new_n54134__;
  assign new_new_n54136__ = ~new_new_n54104__ & ~new_new_n54135__;
  assign new_new_n54137__ = ~new_new_n54119__ & ~new_new_n54135__;
  assign new_new_n54138__ = ~new_new_n54136__ & ~new_new_n54137__;
  assign new_new_n54139__ = ~new_new_n54120__ & new_new_n54138__;
  assign new_new_n54140__ = ~new_new_n54089__ & ~new_new_n54139__;
  assign new_new_n54141__ = ys__n39752 & new_new_n52359__;
  assign new_new_n54142__ = ys__n39750 & new_new_n52358__;
  assign new_new_n54143__ = ~new_new_n54141__ & ~new_new_n54142__;
  assign new_new_n54144__ = ys__n33717 & new_new_n52372__;
  assign new_new_n54145__ = ~ys__n33717 & new_new_n52375__;
  assign new_new_n54146__ = ~new_new_n54144__ & ~new_new_n54145__;
  assign new_new_n54147__ = new_new_n54143__ & new_new_n54146__;
  assign new_new_n54148__ = ys__n24798 & new_new_n52364__;
  assign new_new_n54149__ = ys__n24795 & new_new_n52367__;
  assign new_new_n54150__ = ~new_new_n54148__ & ~new_new_n54149__;
  assign new_new_n54151__ = ys__n24792 & new_new_n52366__;
  assign new_new_n54152__ = ys__n39754 & new_new_n52356__;
  assign new_new_n54153__ = ~new_new_n54151__ & ~new_new_n54152__;
  assign new_new_n54154__ = new_new_n54150__ & new_new_n54153__;
  assign new_new_n54155__ = new_new_n54147__ & new_new_n54154__;
  assign new_new_n54156__ = ys__n39758 & new_new_n52334__;
  assign new_new_n54157__ = ys__n39756 & new_new_n52333__;
  assign new_new_n54158__ = ~new_new_n54156__ & ~new_new_n54157__;
  assign new_new_n54159__ = ys__n33723 & new_new_n52347__;
  assign new_new_n54160__ = ~ys__n33723 & new_new_n52350__;
  assign new_new_n54161__ = ~new_new_n54159__ & ~new_new_n54160__;
  assign new_new_n54162__ = new_new_n54158__ & new_new_n54161__;
  assign new_new_n54163__ = ys__n24807 & new_new_n52339__;
  assign new_new_n54164__ = ys__n24804 & new_new_n52342__;
  assign new_new_n54165__ = ~new_new_n54163__ & ~new_new_n54164__;
  assign new_new_n54166__ = ys__n24801 & new_new_n52341__;
  assign new_new_n54167__ = ys__n39760 & new_new_n52331__;
  assign new_new_n54168__ = ~new_new_n54166__ & ~new_new_n54167__;
  assign new_new_n54169__ = new_new_n54165__ & new_new_n54168__;
  assign new_new_n54170__ = new_new_n54162__ & new_new_n54169__;
  assign new_new_n54171__ = ~new_new_n54155__ & ~new_new_n54170__;
  assign new_new_n54172__ = ys__n24789 & new_new_n52383__;
  assign new_new_n54173__ = ys__n24786 & new_new_n52384__;
  assign new_new_n54174__ = ~new_new_n54172__ & ~new_new_n54173__;
  assign new_new_n54175__ = ys__n39748 & new_new_n52391__;
  assign new_new_n54176__ = ys__n39746 & new_new_n52392__;
  assign new_new_n54177__ = ~new_new_n54175__ & ~new_new_n54176__;
  assign new_new_n54178__ = new_new_n54174__ & new_new_n54177__;
  assign new_new_n54179__ = ~new_new_n54155__ & ~new_new_n54178__;
  assign new_new_n54180__ = ~new_new_n54170__ & ~new_new_n54178__;
  assign new_new_n54181__ = ~new_new_n54179__ & ~new_new_n54180__;
  assign new_new_n54182__ = ~new_new_n54171__ & new_new_n54181__;
  assign new_new_n54183__ = ~new_new_n54089__ & ~new_new_n54182__;
  assign new_new_n54184__ = ~new_new_n54139__ & ~new_new_n54182__;
  assign new_new_n54185__ = ~new_new_n54183__ & ~new_new_n54184__;
  assign new_new_n54186__ = ~new_new_n54140__ & new_new_n54185__;
  assign new_new_n54187__ = ~new_new_n54068__ & ~new_new_n54186__;
  assign new_new_n54188__ = ~new_new_n54078__ & ~new_new_n54186__;
  assign new_new_n54189__ = ~new_new_n54187__ & ~new_new_n54188__;
  assign ys__n42917 = new_new_n54079__ | ~new_new_n54189__;
  assign new_new_n54191__ = ~new_new_n54078__ & new_new_n54187__;
  assign new_new_n54192__ = new_new_n54078__ & ~new_new_n54186__;
  assign new_new_n54193__ = new_new_n54068__ & new_new_n54192__;
  assign new_new_n54194__ = ~new_new_n54078__ & new_new_n54186__;
  assign new_new_n54195__ = new_new_n54068__ & new_new_n54194__;
  assign new_new_n54196__ = new_new_n54078__ & new_new_n54186__;
  assign new_new_n54197__ = ~new_new_n54068__ & new_new_n54196__;
  assign new_new_n54198__ = ~new_new_n54195__ & ~new_new_n54197__;
  assign new_new_n54199__ = ~new_new_n54193__ & new_new_n54198__;
  assign ys__n42922 = new_new_n54191__ | ~new_new_n54199__;
  assign new_new_n54201__ = ~new_new_n54139__ & new_new_n54183__;
  assign new_new_n54202__ = new_new_n54139__ & ~new_new_n54182__;
  assign new_new_n54203__ = new_new_n54089__ & new_new_n54202__;
  assign new_new_n54204__ = ~new_new_n54139__ & new_new_n54182__;
  assign new_new_n54205__ = new_new_n54089__ & new_new_n54204__;
  assign new_new_n54206__ = new_new_n54139__ & new_new_n54182__;
  assign new_new_n54207__ = ~new_new_n54089__ & new_new_n54206__;
  assign new_new_n54208__ = ~new_new_n54205__ & ~new_new_n54207__;
  assign new_new_n54209__ = ~new_new_n54203__ & new_new_n54208__;
  assign new_new_n54210__ = ~new_new_n54201__ & new_new_n54209__;
  assign new_new_n54211__ = ~new_new_n53977__ & new_new_n53994__;
  assign new_new_n54212__ = new_new_n53964__ & new_new_n53993__;
  assign new_new_n54213__ = ~new_new_n53977__ & new_new_n54212__;
  assign new_new_n54214__ = ~new_new_n54211__ & ~new_new_n54213__;
  assign new_new_n54215__ = ~new_new_n53964__ & new_new_n53993__;
  assign new_new_n54216__ = new_new_n53977__ & new_new_n54215__;
  assign new_new_n54217__ = new_new_n53964__ & ~new_new_n53993__;
  assign new_new_n54218__ = new_new_n53977__ & new_new_n54217__;
  assign new_new_n54219__ = ~new_new_n54216__ & ~new_new_n54218__;
  assign new_new_n54220__ = new_new_n54214__ & new_new_n54219__;
  assign new_new_n54221__ = ~new_new_n54210__ & ~new_new_n54220__;
  assign new_new_n54222__ = ~new_new_n54170__ & new_new_n54179__;
  assign new_new_n54223__ = new_new_n54155__ & new_new_n54178__;
  assign new_new_n54224__ = ~new_new_n54170__ & new_new_n54223__;
  assign new_new_n54225__ = ~new_new_n54222__ & ~new_new_n54224__;
  assign new_new_n54226__ = ~new_new_n54155__ & new_new_n54178__;
  assign new_new_n54227__ = new_new_n54170__ & new_new_n54226__;
  assign new_new_n54228__ = new_new_n54155__ & ~new_new_n54178__;
  assign new_new_n54229__ = new_new_n54170__ & new_new_n54228__;
  assign new_new_n54230__ = ~new_new_n54227__ & ~new_new_n54229__;
  assign new_new_n54231__ = new_new_n54225__ & new_new_n54230__;
  assign new_new_n54232__ = ys__n39768 & new_new_n52412__;
  assign new_new_n54233__ = ys__n39766 & new_new_n52411__;
  assign new_new_n54234__ = ~new_new_n54232__ & ~new_new_n54233__;
  assign new_new_n54235__ = ys__n33733 & new_new_n52425__;
  assign new_new_n54236__ = ~ys__n33733 & new_new_n52428__;
  assign new_new_n54237__ = ~new_new_n54235__ & ~new_new_n54236__;
  assign new_new_n54238__ = new_new_n54234__ & new_new_n54237__;
  assign new_new_n54239__ = ys__n24822 & new_new_n52417__;
  assign new_new_n54240__ = ys__n24819 & new_new_n52420__;
  assign new_new_n54241__ = ~new_new_n54239__ & ~new_new_n54240__;
  assign new_new_n54242__ = ys__n24816 & new_new_n52419__;
  assign new_new_n54243__ = ys__n39770 & new_new_n52409__;
  assign new_new_n54244__ = ~new_new_n54242__ & ~new_new_n54243__;
  assign new_new_n54245__ = new_new_n54241__ & new_new_n54244__;
  assign new_new_n54246__ = new_new_n54238__ & new_new_n54245__;
  assign new_new_n54247__ = ys__n39774 & new_new_n52301__;
  assign new_new_n54248__ = ys__n39772 & new_new_n52304__;
  assign new_new_n54249__ = ~new_new_n54247__ & ~new_new_n54248__;
  assign new_new_n54250__ = ys__n33739 & new_new_n52308__;
  assign new_new_n54251__ = ~ys__n33739 & new_new_n52311__;
  assign new_new_n54252__ = ~new_new_n54250__ & ~new_new_n54251__;
  assign new_new_n54253__ = new_new_n54249__ & new_new_n54252__;
  assign new_new_n54254__ = ys__n24831 & new_new_n52316__;
  assign new_new_n54255__ = ys__n24828 & new_new_n52318__;
  assign new_new_n54256__ = ~new_new_n54254__ & ~new_new_n54255__;
  assign new_new_n54257__ = ys__n24825 & new_new_n52322__;
  assign new_new_n54258__ = ys__n39776 & new_new_n52324__;
  assign new_new_n54259__ = ~new_new_n54257__ & ~new_new_n54258__;
  assign new_new_n54260__ = new_new_n54256__ & new_new_n54259__;
  assign new_new_n54261__ = new_new_n54253__ & new_new_n54260__;
  assign new_new_n54262__ = ~new_new_n54246__ & ~new_new_n54261__;
  assign new_new_n54263__ = ys__n39762 & new_new_n52449__;
  assign new_new_n54264__ = ys__n39760 & new_new_n52448__;
  assign new_new_n54265__ = ~new_new_n54263__ & ~new_new_n54264__;
  assign new_new_n54266__ = ys__n33727 & new_new_n52462__;
  assign new_new_n54267__ = ~ys__n33727 & new_new_n52465__;
  assign new_new_n54268__ = ~new_new_n54266__ & ~new_new_n54267__;
  assign new_new_n54269__ = new_new_n54265__ & new_new_n54268__;
  assign new_new_n54270__ = ys__n24813 & new_new_n52454__;
  assign new_new_n54271__ = ys__n24810 & new_new_n52457__;
  assign new_new_n54272__ = ~new_new_n54270__ & ~new_new_n54271__;
  assign new_new_n54273__ = ys__n24807 & new_new_n52456__;
  assign new_new_n54274__ = ys__n39764 & new_new_n52446__;
  assign new_new_n54275__ = ~new_new_n54273__ & ~new_new_n54274__;
  assign new_new_n54276__ = new_new_n54272__ & new_new_n54275__;
  assign new_new_n54277__ = new_new_n54269__ & new_new_n54276__;
  assign new_new_n54278__ = ~new_new_n54246__ & ~new_new_n54277__;
  assign new_new_n54279__ = ~new_new_n54261__ & ~new_new_n54277__;
  assign new_new_n54280__ = ~new_new_n54278__ & ~new_new_n54279__;
  assign new_new_n54281__ = ~new_new_n54262__ & new_new_n54280__;
  assign new_new_n54282__ = ~new_new_n54231__ & ~new_new_n54281__;
  assign new_new_n54283__ = ys__n39750 & new_new_n52359__;
  assign new_new_n54284__ = ys__n39748 & new_new_n52358__;
  assign new_new_n54285__ = ~new_new_n54283__ & ~new_new_n54284__;
  assign new_new_n54286__ = ys__n33715 & new_new_n52372__;
  assign new_new_n54287__ = ~ys__n33715 & new_new_n52375__;
  assign new_new_n54288__ = ~new_new_n54286__ & ~new_new_n54287__;
  assign new_new_n54289__ = new_new_n54285__ & new_new_n54288__;
  assign new_new_n54290__ = ys__n24795 & new_new_n52364__;
  assign new_new_n54291__ = ys__n24792 & new_new_n52367__;
  assign new_new_n54292__ = ~new_new_n54290__ & ~new_new_n54291__;
  assign new_new_n54293__ = ys__n24789 & new_new_n52366__;
  assign new_new_n54294__ = ys__n39752 & new_new_n52356__;
  assign new_new_n54295__ = ~new_new_n54293__ & ~new_new_n54294__;
  assign new_new_n54296__ = new_new_n54292__ & new_new_n54295__;
  assign new_new_n54297__ = new_new_n54289__ & new_new_n54296__;
  assign new_new_n54298__ = ys__n39756 & new_new_n52334__;
  assign new_new_n54299__ = ys__n39754 & new_new_n52333__;
  assign new_new_n54300__ = ~new_new_n54298__ & ~new_new_n54299__;
  assign new_new_n54301__ = ys__n33721 & new_new_n52347__;
  assign new_new_n54302__ = ~ys__n33721 & new_new_n52350__;
  assign new_new_n54303__ = ~new_new_n54301__ & ~new_new_n54302__;
  assign new_new_n54304__ = new_new_n54300__ & new_new_n54303__;
  assign new_new_n54305__ = ys__n24804 & new_new_n52339__;
  assign new_new_n54306__ = ys__n24801 & new_new_n52342__;
  assign new_new_n54307__ = ~new_new_n54305__ & ~new_new_n54306__;
  assign new_new_n54308__ = ys__n24798 & new_new_n52341__;
  assign new_new_n54309__ = ys__n39758 & new_new_n52331__;
  assign new_new_n54310__ = ~new_new_n54308__ & ~new_new_n54309__;
  assign new_new_n54311__ = new_new_n54307__ & new_new_n54310__;
  assign new_new_n54312__ = new_new_n54304__ & new_new_n54311__;
  assign new_new_n54313__ = ~new_new_n54297__ & ~new_new_n54312__;
  assign new_new_n54314__ = ys__n24786 & new_new_n52383__;
  assign new_new_n54315__ = ys__n24783 & new_new_n52384__;
  assign new_new_n54316__ = ~new_new_n54314__ & ~new_new_n54315__;
  assign new_new_n54317__ = ys__n39746 & new_new_n52391__;
  assign new_new_n54318__ = ys__n39744 & new_new_n52392__;
  assign new_new_n54319__ = ~new_new_n54317__ & ~new_new_n54318__;
  assign new_new_n54320__ = new_new_n54316__ & new_new_n54319__;
  assign new_new_n54321__ = ~new_new_n54297__ & ~new_new_n54320__;
  assign new_new_n54322__ = ~new_new_n54312__ & ~new_new_n54320__;
  assign new_new_n54323__ = ~new_new_n54321__ & ~new_new_n54322__;
  assign new_new_n54324__ = ~new_new_n54313__ & new_new_n54323__;
  assign new_new_n54325__ = ~new_new_n54231__ & ~new_new_n54324__;
  assign new_new_n54326__ = ~new_new_n54281__ & ~new_new_n54324__;
  assign new_new_n54327__ = ~new_new_n54325__ & ~new_new_n54326__;
  assign new_new_n54328__ = ~new_new_n54282__ & new_new_n54327__;
  assign new_new_n54329__ = ~new_new_n54210__ & ~new_new_n54328__;
  assign new_new_n54330__ = ~new_new_n54220__ & ~new_new_n54328__;
  assign new_new_n54331__ = ~new_new_n54329__ & ~new_new_n54330__;
  assign ys__n42971 = new_new_n54221__ | ~new_new_n54331__;
  assign new_new_n54333__ = ~new_new_n54220__ & new_new_n54329__;
  assign new_new_n54334__ = new_new_n54220__ & ~new_new_n54328__;
  assign new_new_n54335__ = new_new_n54210__ & new_new_n54334__;
  assign new_new_n54336__ = ~new_new_n54220__ & new_new_n54328__;
  assign new_new_n54337__ = new_new_n54210__ & new_new_n54336__;
  assign new_new_n54338__ = new_new_n54220__ & new_new_n54328__;
  assign new_new_n54339__ = ~new_new_n54210__ & new_new_n54338__;
  assign new_new_n54340__ = ~new_new_n54337__ & ~new_new_n54339__;
  assign new_new_n54341__ = ~new_new_n54335__ & new_new_n54340__;
  assign ys__n42976 = new_new_n54333__ | ~new_new_n54341__;
  assign new_new_n54343__ = ~new_new_n54281__ & new_new_n54325__;
  assign new_new_n54344__ = new_new_n54281__ & ~new_new_n54324__;
  assign new_new_n54345__ = new_new_n54231__ & new_new_n54344__;
  assign new_new_n54346__ = ~new_new_n54281__ & new_new_n54324__;
  assign new_new_n54347__ = new_new_n54231__ & new_new_n54346__;
  assign new_new_n54348__ = new_new_n54281__ & new_new_n54324__;
  assign new_new_n54349__ = ~new_new_n54231__ & new_new_n54348__;
  assign new_new_n54350__ = ~new_new_n54347__ & ~new_new_n54349__;
  assign new_new_n54351__ = ~new_new_n54345__ & new_new_n54350__;
  assign new_new_n54352__ = ~new_new_n54343__ & new_new_n54351__;
  assign new_new_n54353__ = ~new_new_n54119__ & new_new_n54136__;
  assign new_new_n54354__ = new_new_n54104__ & new_new_n54135__;
  assign new_new_n54355__ = ~new_new_n54119__ & new_new_n54354__;
  assign new_new_n54356__ = ~new_new_n54353__ & ~new_new_n54355__;
  assign new_new_n54357__ = ~new_new_n54104__ & new_new_n54135__;
  assign new_new_n54358__ = new_new_n54119__ & new_new_n54357__;
  assign new_new_n54359__ = new_new_n54104__ & ~new_new_n54135__;
  assign new_new_n54360__ = new_new_n54119__ & new_new_n54359__;
  assign new_new_n54361__ = ~new_new_n54358__ & ~new_new_n54360__;
  assign new_new_n54362__ = new_new_n54356__ & new_new_n54361__;
  assign new_new_n54363__ = ~new_new_n54352__ & ~new_new_n54362__;
  assign new_new_n54364__ = ~new_new_n54312__ & new_new_n54321__;
  assign new_new_n54365__ = new_new_n54297__ & new_new_n54320__;
  assign new_new_n54366__ = ~new_new_n54312__ & new_new_n54365__;
  assign new_new_n54367__ = ~new_new_n54364__ & ~new_new_n54366__;
  assign new_new_n54368__ = ~new_new_n54297__ & new_new_n54320__;
  assign new_new_n54369__ = new_new_n54312__ & new_new_n54368__;
  assign new_new_n54370__ = new_new_n54297__ & ~new_new_n54320__;
  assign new_new_n54371__ = new_new_n54312__ & new_new_n54370__;
  assign new_new_n54372__ = ~new_new_n54369__ & ~new_new_n54371__;
  assign new_new_n54373__ = new_new_n54367__ & new_new_n54372__;
  assign new_new_n54374__ = ys__n39766 & new_new_n52412__;
  assign new_new_n54375__ = ys__n39764 & new_new_n52411__;
  assign new_new_n54376__ = ~new_new_n54374__ & ~new_new_n54375__;
  assign new_new_n54377__ = ys__n33731 & new_new_n52425__;
  assign new_new_n54378__ = ~ys__n33731 & new_new_n52428__;
  assign new_new_n54379__ = ~new_new_n54377__ & ~new_new_n54378__;
  assign new_new_n54380__ = new_new_n54376__ & new_new_n54379__;
  assign new_new_n54381__ = ys__n24819 & new_new_n52417__;
  assign new_new_n54382__ = ys__n24816 & new_new_n52420__;
  assign new_new_n54383__ = ~new_new_n54381__ & ~new_new_n54382__;
  assign new_new_n54384__ = ys__n24813 & new_new_n52419__;
  assign new_new_n54385__ = ys__n39768 & new_new_n52409__;
  assign new_new_n54386__ = ~new_new_n54384__ & ~new_new_n54385__;
  assign new_new_n54387__ = new_new_n54383__ & new_new_n54386__;
  assign new_new_n54388__ = new_new_n54380__ & new_new_n54387__;
  assign new_new_n54389__ = ys__n39772 & new_new_n52301__;
  assign new_new_n54390__ = ys__n39770 & new_new_n52304__;
  assign new_new_n54391__ = ~new_new_n54389__ & ~new_new_n54390__;
  assign new_new_n54392__ = ys__n33737 & new_new_n52308__;
  assign new_new_n54393__ = ~ys__n33737 & new_new_n52311__;
  assign new_new_n54394__ = ~new_new_n54392__ & ~new_new_n54393__;
  assign new_new_n54395__ = new_new_n54391__ & new_new_n54394__;
  assign new_new_n54396__ = ys__n24828 & new_new_n52316__;
  assign new_new_n54397__ = ys__n24825 & new_new_n52318__;
  assign new_new_n54398__ = ~new_new_n54396__ & ~new_new_n54397__;
  assign new_new_n54399__ = ys__n24822 & new_new_n52322__;
  assign new_new_n54400__ = ys__n39774 & new_new_n52324__;
  assign new_new_n54401__ = ~new_new_n54399__ & ~new_new_n54400__;
  assign new_new_n54402__ = new_new_n54398__ & new_new_n54401__;
  assign new_new_n54403__ = new_new_n54395__ & new_new_n54402__;
  assign new_new_n54404__ = ~new_new_n54388__ & ~new_new_n54403__;
  assign new_new_n54405__ = ys__n39760 & new_new_n52449__;
  assign new_new_n54406__ = ys__n39758 & new_new_n52448__;
  assign new_new_n54407__ = ~new_new_n54405__ & ~new_new_n54406__;
  assign new_new_n54408__ = ys__n33725 & new_new_n52462__;
  assign new_new_n54409__ = ~ys__n33725 & new_new_n52465__;
  assign new_new_n54410__ = ~new_new_n54408__ & ~new_new_n54409__;
  assign new_new_n54411__ = new_new_n54407__ & new_new_n54410__;
  assign new_new_n54412__ = ys__n24810 & new_new_n52454__;
  assign new_new_n54413__ = ys__n24807 & new_new_n52457__;
  assign new_new_n54414__ = ~new_new_n54412__ & ~new_new_n54413__;
  assign new_new_n54415__ = ys__n24804 & new_new_n52456__;
  assign new_new_n54416__ = ys__n39762 & new_new_n52446__;
  assign new_new_n54417__ = ~new_new_n54415__ & ~new_new_n54416__;
  assign new_new_n54418__ = new_new_n54414__ & new_new_n54417__;
  assign new_new_n54419__ = new_new_n54411__ & new_new_n54418__;
  assign new_new_n54420__ = ~new_new_n54388__ & ~new_new_n54419__;
  assign new_new_n54421__ = ~new_new_n54403__ & ~new_new_n54419__;
  assign new_new_n54422__ = ~new_new_n54420__ & ~new_new_n54421__;
  assign new_new_n54423__ = ~new_new_n54404__ & new_new_n54422__;
  assign new_new_n54424__ = ~new_new_n54373__ & ~new_new_n54423__;
  assign new_new_n54425__ = ys__n39748 & new_new_n52359__;
  assign new_new_n54426__ = ys__n39746 & new_new_n52358__;
  assign new_new_n54427__ = ~new_new_n54425__ & ~new_new_n54426__;
  assign new_new_n54428__ = ys__n33713 & new_new_n52372__;
  assign new_new_n54429__ = ~ys__n33713 & new_new_n52375__;
  assign new_new_n54430__ = ~new_new_n54428__ & ~new_new_n54429__;
  assign new_new_n54431__ = new_new_n54427__ & new_new_n54430__;
  assign new_new_n54432__ = ys__n24792 & new_new_n52364__;
  assign new_new_n54433__ = ys__n24789 & new_new_n52367__;
  assign new_new_n54434__ = ~new_new_n54432__ & ~new_new_n54433__;
  assign new_new_n54435__ = ys__n24786 & new_new_n52366__;
  assign new_new_n54436__ = ys__n39750 & new_new_n52356__;
  assign new_new_n54437__ = ~new_new_n54435__ & ~new_new_n54436__;
  assign new_new_n54438__ = new_new_n54434__ & new_new_n54437__;
  assign new_new_n54439__ = new_new_n54431__ & new_new_n54438__;
  assign new_new_n54440__ = ys__n39754 & new_new_n52334__;
  assign new_new_n54441__ = ys__n39752 & new_new_n52333__;
  assign new_new_n54442__ = ~new_new_n54440__ & ~new_new_n54441__;
  assign new_new_n54443__ = ys__n33719 & new_new_n52347__;
  assign new_new_n54444__ = ~ys__n33719 & new_new_n52350__;
  assign new_new_n54445__ = ~new_new_n54443__ & ~new_new_n54444__;
  assign new_new_n54446__ = new_new_n54442__ & new_new_n54445__;
  assign new_new_n54447__ = ys__n24801 & new_new_n52339__;
  assign new_new_n54448__ = ys__n24798 & new_new_n52342__;
  assign new_new_n54449__ = ~new_new_n54447__ & ~new_new_n54448__;
  assign new_new_n54450__ = ys__n24795 & new_new_n52341__;
  assign new_new_n54451__ = ys__n39756 & new_new_n52331__;
  assign new_new_n54452__ = ~new_new_n54450__ & ~new_new_n54451__;
  assign new_new_n54453__ = new_new_n54449__ & new_new_n54452__;
  assign new_new_n54454__ = new_new_n54446__ & new_new_n54453__;
  assign new_new_n54455__ = ~new_new_n54439__ & ~new_new_n54454__;
  assign new_new_n54456__ = ys__n24783 & new_new_n52383__;
  assign new_new_n54457__ = ys__n24780 & new_new_n52384__;
  assign new_new_n54458__ = ~new_new_n54456__ & ~new_new_n54457__;
  assign new_new_n54459__ = ys__n39744 & new_new_n52391__;
  assign new_new_n54460__ = ys__n39742 & new_new_n52392__;
  assign new_new_n54461__ = ~new_new_n54459__ & ~new_new_n54460__;
  assign new_new_n54462__ = new_new_n54458__ & new_new_n54461__;
  assign new_new_n54463__ = ~new_new_n54439__ & ~new_new_n54462__;
  assign new_new_n54464__ = ~new_new_n54454__ & ~new_new_n54462__;
  assign new_new_n54465__ = ~new_new_n54463__ & ~new_new_n54464__;
  assign new_new_n54466__ = ~new_new_n54455__ & new_new_n54465__;
  assign new_new_n54467__ = ~new_new_n54373__ & ~new_new_n54466__;
  assign new_new_n54468__ = ~new_new_n54423__ & ~new_new_n54466__;
  assign new_new_n54469__ = ~new_new_n54467__ & ~new_new_n54468__;
  assign new_new_n54470__ = ~new_new_n54424__ & new_new_n54469__;
  assign new_new_n54471__ = ~new_new_n54352__ & ~new_new_n54470__;
  assign new_new_n54472__ = ~new_new_n54362__ & ~new_new_n54470__;
  assign new_new_n54473__ = ~new_new_n54471__ & ~new_new_n54472__;
  assign ys__n43025 = new_new_n54363__ | ~new_new_n54473__;
  assign new_new_n54475__ = ~new_new_n54362__ & new_new_n54471__;
  assign new_new_n54476__ = new_new_n54362__ & ~new_new_n54470__;
  assign new_new_n54477__ = new_new_n54352__ & new_new_n54476__;
  assign new_new_n54478__ = ~new_new_n54362__ & new_new_n54470__;
  assign new_new_n54479__ = new_new_n54352__ & new_new_n54478__;
  assign new_new_n54480__ = new_new_n54362__ & new_new_n54470__;
  assign new_new_n54481__ = ~new_new_n54352__ & new_new_n54480__;
  assign new_new_n54482__ = ~new_new_n54479__ & ~new_new_n54481__;
  assign new_new_n54483__ = ~new_new_n54477__ & new_new_n54482__;
  assign ys__n43030 = new_new_n54475__ | ~new_new_n54483__;
  assign new_new_n54485__ = ~new_new_n54423__ & new_new_n54467__;
  assign new_new_n54486__ = new_new_n54423__ & ~new_new_n54466__;
  assign new_new_n54487__ = new_new_n54373__ & new_new_n54486__;
  assign new_new_n54488__ = ~new_new_n54423__ & new_new_n54466__;
  assign new_new_n54489__ = new_new_n54373__ & new_new_n54488__;
  assign new_new_n54490__ = new_new_n54423__ & new_new_n54466__;
  assign new_new_n54491__ = ~new_new_n54373__ & new_new_n54490__;
  assign new_new_n54492__ = ~new_new_n54489__ & ~new_new_n54491__;
  assign new_new_n54493__ = ~new_new_n54487__ & new_new_n54492__;
  assign new_new_n54494__ = ~new_new_n54485__ & new_new_n54493__;
  assign new_new_n54495__ = ~new_new_n54261__ & new_new_n54278__;
  assign new_new_n54496__ = new_new_n54246__ & new_new_n54277__;
  assign new_new_n54497__ = ~new_new_n54261__ & new_new_n54496__;
  assign new_new_n54498__ = ~new_new_n54495__ & ~new_new_n54497__;
  assign new_new_n54499__ = ~new_new_n54246__ & new_new_n54277__;
  assign new_new_n54500__ = new_new_n54261__ & new_new_n54499__;
  assign new_new_n54501__ = new_new_n54246__ & ~new_new_n54277__;
  assign new_new_n54502__ = new_new_n54261__ & new_new_n54501__;
  assign new_new_n54503__ = ~new_new_n54500__ & ~new_new_n54502__;
  assign new_new_n54504__ = new_new_n54498__ & new_new_n54503__;
  assign new_new_n54505__ = ~new_new_n54494__ & ~new_new_n54504__;
  assign new_new_n54506__ = ~new_new_n54454__ & new_new_n54463__;
  assign new_new_n54507__ = new_new_n54439__ & new_new_n54462__;
  assign new_new_n54508__ = ~new_new_n54454__ & new_new_n54507__;
  assign new_new_n54509__ = ~new_new_n54506__ & ~new_new_n54508__;
  assign new_new_n54510__ = ~new_new_n54439__ & new_new_n54462__;
  assign new_new_n54511__ = new_new_n54454__ & new_new_n54510__;
  assign new_new_n54512__ = new_new_n54439__ & ~new_new_n54462__;
  assign new_new_n54513__ = new_new_n54454__ & new_new_n54512__;
  assign new_new_n54514__ = ~new_new_n54511__ & ~new_new_n54513__;
  assign new_new_n54515__ = new_new_n54509__ & new_new_n54514__;
  assign new_new_n54516__ = ys__n39764 & new_new_n52412__;
  assign new_new_n54517__ = ys__n39762 & new_new_n52411__;
  assign new_new_n54518__ = ~new_new_n54516__ & ~new_new_n54517__;
  assign new_new_n54519__ = ys__n33729 & new_new_n52425__;
  assign new_new_n54520__ = ~ys__n33729 & new_new_n52428__;
  assign new_new_n54521__ = ~new_new_n54519__ & ~new_new_n54520__;
  assign new_new_n54522__ = new_new_n54518__ & new_new_n54521__;
  assign new_new_n54523__ = ys__n24816 & new_new_n52417__;
  assign new_new_n54524__ = ys__n24813 & new_new_n52420__;
  assign new_new_n54525__ = ~new_new_n54523__ & ~new_new_n54524__;
  assign new_new_n54526__ = ys__n24810 & new_new_n52419__;
  assign new_new_n54527__ = ys__n39766 & new_new_n52409__;
  assign new_new_n54528__ = ~new_new_n54526__ & ~new_new_n54527__;
  assign new_new_n54529__ = new_new_n54525__ & new_new_n54528__;
  assign new_new_n54530__ = new_new_n54522__ & new_new_n54529__;
  assign new_new_n54531__ = ys__n39770 & new_new_n52301__;
  assign new_new_n54532__ = ys__n39768 & new_new_n52304__;
  assign new_new_n54533__ = ~new_new_n54531__ & ~new_new_n54532__;
  assign new_new_n54534__ = ys__n33735 & new_new_n52308__;
  assign new_new_n54535__ = ~ys__n33735 & new_new_n52311__;
  assign new_new_n54536__ = ~new_new_n54534__ & ~new_new_n54535__;
  assign new_new_n54537__ = new_new_n54533__ & new_new_n54536__;
  assign new_new_n54538__ = ys__n24825 & new_new_n52316__;
  assign new_new_n54539__ = ys__n24822 & new_new_n52318__;
  assign new_new_n54540__ = ~new_new_n54538__ & ~new_new_n54539__;
  assign new_new_n54541__ = ys__n24819 & new_new_n52322__;
  assign new_new_n54542__ = ys__n39772 & new_new_n52324__;
  assign new_new_n54543__ = ~new_new_n54541__ & ~new_new_n54542__;
  assign new_new_n54544__ = new_new_n54540__ & new_new_n54543__;
  assign new_new_n54545__ = new_new_n54537__ & new_new_n54544__;
  assign new_new_n54546__ = ~new_new_n54530__ & ~new_new_n54545__;
  assign new_new_n54547__ = ys__n39758 & new_new_n52449__;
  assign new_new_n54548__ = ys__n39756 & new_new_n52448__;
  assign new_new_n54549__ = ~new_new_n54547__ & ~new_new_n54548__;
  assign new_new_n54550__ = ys__n33723 & new_new_n52462__;
  assign new_new_n54551__ = ~ys__n33723 & new_new_n52465__;
  assign new_new_n54552__ = ~new_new_n54550__ & ~new_new_n54551__;
  assign new_new_n54553__ = new_new_n54549__ & new_new_n54552__;
  assign new_new_n54554__ = ys__n24807 & new_new_n52454__;
  assign new_new_n54555__ = ys__n24804 & new_new_n52457__;
  assign new_new_n54556__ = ~new_new_n54554__ & ~new_new_n54555__;
  assign new_new_n54557__ = ys__n24801 & new_new_n52456__;
  assign new_new_n54558__ = ys__n39760 & new_new_n52446__;
  assign new_new_n54559__ = ~new_new_n54557__ & ~new_new_n54558__;
  assign new_new_n54560__ = new_new_n54556__ & new_new_n54559__;
  assign new_new_n54561__ = new_new_n54553__ & new_new_n54560__;
  assign new_new_n54562__ = ~new_new_n54530__ & ~new_new_n54561__;
  assign new_new_n54563__ = ~new_new_n54545__ & ~new_new_n54561__;
  assign new_new_n54564__ = ~new_new_n54562__ & ~new_new_n54563__;
  assign new_new_n54565__ = ~new_new_n54546__ & new_new_n54564__;
  assign new_new_n54566__ = ~new_new_n54515__ & ~new_new_n54565__;
  assign new_new_n54567__ = ys__n39746 & new_new_n52359__;
  assign new_new_n54568__ = ys__n39744 & new_new_n52358__;
  assign new_new_n54569__ = ~new_new_n54567__ & ~new_new_n54568__;
  assign new_new_n54570__ = ys__n33711 & new_new_n52372__;
  assign new_new_n54571__ = ~ys__n33711 & new_new_n52375__;
  assign new_new_n54572__ = ~new_new_n54570__ & ~new_new_n54571__;
  assign new_new_n54573__ = new_new_n54569__ & new_new_n54572__;
  assign new_new_n54574__ = ys__n24789 & new_new_n52364__;
  assign new_new_n54575__ = ys__n24786 & new_new_n52367__;
  assign new_new_n54576__ = ~new_new_n54574__ & ~new_new_n54575__;
  assign new_new_n54577__ = ys__n24783 & new_new_n52366__;
  assign new_new_n54578__ = ys__n39748 & new_new_n52356__;
  assign new_new_n54579__ = ~new_new_n54577__ & ~new_new_n54578__;
  assign new_new_n54580__ = new_new_n54576__ & new_new_n54579__;
  assign new_new_n54581__ = new_new_n54573__ & new_new_n54580__;
  assign new_new_n54582__ = ys__n39752 & new_new_n52334__;
  assign new_new_n54583__ = ys__n39750 & new_new_n52333__;
  assign new_new_n54584__ = ~new_new_n54582__ & ~new_new_n54583__;
  assign new_new_n54585__ = ys__n33717 & new_new_n52347__;
  assign new_new_n54586__ = ~ys__n33717 & new_new_n52350__;
  assign new_new_n54587__ = ~new_new_n54585__ & ~new_new_n54586__;
  assign new_new_n54588__ = new_new_n54584__ & new_new_n54587__;
  assign new_new_n54589__ = ys__n24798 & new_new_n52339__;
  assign new_new_n54590__ = ys__n24795 & new_new_n52342__;
  assign new_new_n54591__ = ~new_new_n54589__ & ~new_new_n54590__;
  assign new_new_n54592__ = ys__n24792 & new_new_n52341__;
  assign new_new_n54593__ = ys__n39754 & new_new_n52331__;
  assign new_new_n54594__ = ~new_new_n54592__ & ~new_new_n54593__;
  assign new_new_n54595__ = new_new_n54591__ & new_new_n54594__;
  assign new_new_n54596__ = new_new_n54588__ & new_new_n54595__;
  assign new_new_n54597__ = ~new_new_n54581__ & ~new_new_n54596__;
  assign new_new_n54598__ = ys__n24780 & new_new_n52383__;
  assign new_new_n54599__ = ys__n24777 & new_new_n52384__;
  assign new_new_n54600__ = ~new_new_n54598__ & ~new_new_n54599__;
  assign new_new_n54601__ = ys__n39742 & new_new_n52391__;
  assign new_new_n54602__ = ys__n39740 & new_new_n52392__;
  assign new_new_n54603__ = ~new_new_n54601__ & ~new_new_n54602__;
  assign new_new_n54604__ = new_new_n54600__ & new_new_n54603__;
  assign new_new_n54605__ = ~new_new_n54581__ & ~new_new_n54604__;
  assign new_new_n54606__ = ~new_new_n54596__ & ~new_new_n54604__;
  assign new_new_n54607__ = ~new_new_n54605__ & ~new_new_n54606__;
  assign new_new_n54608__ = ~new_new_n54597__ & new_new_n54607__;
  assign new_new_n54609__ = ~new_new_n54515__ & ~new_new_n54608__;
  assign new_new_n54610__ = ~new_new_n54565__ & ~new_new_n54608__;
  assign new_new_n54611__ = ~new_new_n54609__ & ~new_new_n54610__;
  assign new_new_n54612__ = ~new_new_n54566__ & new_new_n54611__;
  assign new_new_n54613__ = ~new_new_n54494__ & ~new_new_n54612__;
  assign new_new_n54614__ = ~new_new_n54504__ & ~new_new_n54612__;
  assign new_new_n54615__ = ~new_new_n54613__ & ~new_new_n54614__;
  assign ys__n43079 = new_new_n54505__ | ~new_new_n54615__;
  assign new_new_n54617__ = ~new_new_n54504__ & new_new_n54613__;
  assign new_new_n54618__ = new_new_n54504__ & ~new_new_n54612__;
  assign new_new_n54619__ = new_new_n54494__ & new_new_n54618__;
  assign new_new_n54620__ = ~new_new_n54504__ & new_new_n54612__;
  assign new_new_n54621__ = new_new_n54494__ & new_new_n54620__;
  assign new_new_n54622__ = new_new_n54504__ & new_new_n54612__;
  assign new_new_n54623__ = ~new_new_n54494__ & new_new_n54622__;
  assign new_new_n54624__ = ~new_new_n54621__ & ~new_new_n54623__;
  assign new_new_n54625__ = ~new_new_n54619__ & new_new_n54624__;
  assign ys__n43084 = new_new_n54617__ | ~new_new_n54625__;
  assign new_new_n54627__ = ~new_new_n54565__ & new_new_n54609__;
  assign new_new_n54628__ = new_new_n54565__ & ~new_new_n54608__;
  assign new_new_n54629__ = new_new_n54515__ & new_new_n54628__;
  assign new_new_n54630__ = ~new_new_n54565__ & new_new_n54608__;
  assign new_new_n54631__ = new_new_n54515__ & new_new_n54630__;
  assign new_new_n54632__ = new_new_n54565__ & new_new_n54608__;
  assign new_new_n54633__ = ~new_new_n54515__ & new_new_n54632__;
  assign new_new_n54634__ = ~new_new_n54631__ & ~new_new_n54633__;
  assign new_new_n54635__ = ~new_new_n54629__ & new_new_n54634__;
  assign new_new_n54636__ = ~new_new_n54627__ & new_new_n54635__;
  assign new_new_n54637__ = ~new_new_n54403__ & new_new_n54420__;
  assign new_new_n54638__ = new_new_n54388__ & new_new_n54419__;
  assign new_new_n54639__ = ~new_new_n54403__ & new_new_n54638__;
  assign new_new_n54640__ = ~new_new_n54637__ & ~new_new_n54639__;
  assign new_new_n54641__ = ~new_new_n54388__ & new_new_n54419__;
  assign new_new_n54642__ = new_new_n54403__ & new_new_n54641__;
  assign new_new_n54643__ = new_new_n54388__ & ~new_new_n54419__;
  assign new_new_n54644__ = new_new_n54403__ & new_new_n54643__;
  assign new_new_n54645__ = ~new_new_n54642__ & ~new_new_n54644__;
  assign new_new_n54646__ = new_new_n54640__ & new_new_n54645__;
  assign new_new_n54647__ = ~new_new_n54636__ & ~new_new_n54646__;
  assign new_new_n54648__ = ~new_new_n54596__ & new_new_n54605__;
  assign new_new_n54649__ = new_new_n54581__ & new_new_n54604__;
  assign new_new_n54650__ = ~new_new_n54596__ & new_new_n54649__;
  assign new_new_n54651__ = ~new_new_n54648__ & ~new_new_n54650__;
  assign new_new_n54652__ = ~new_new_n54581__ & new_new_n54604__;
  assign new_new_n54653__ = new_new_n54596__ & new_new_n54652__;
  assign new_new_n54654__ = new_new_n54581__ & ~new_new_n54604__;
  assign new_new_n54655__ = new_new_n54596__ & new_new_n54654__;
  assign new_new_n54656__ = ~new_new_n54653__ & ~new_new_n54655__;
  assign new_new_n54657__ = new_new_n54651__ & new_new_n54656__;
  assign new_new_n54658__ = ys__n39762 & new_new_n52412__;
  assign new_new_n54659__ = ys__n39760 & new_new_n52411__;
  assign new_new_n54660__ = ~new_new_n54658__ & ~new_new_n54659__;
  assign new_new_n54661__ = ys__n33727 & new_new_n52425__;
  assign new_new_n54662__ = ~ys__n33727 & new_new_n52428__;
  assign new_new_n54663__ = ~new_new_n54661__ & ~new_new_n54662__;
  assign new_new_n54664__ = new_new_n54660__ & new_new_n54663__;
  assign new_new_n54665__ = ys__n24813 & new_new_n52417__;
  assign new_new_n54666__ = ys__n24810 & new_new_n52420__;
  assign new_new_n54667__ = ~new_new_n54665__ & ~new_new_n54666__;
  assign new_new_n54668__ = ys__n24807 & new_new_n52419__;
  assign new_new_n54669__ = ys__n39764 & new_new_n52409__;
  assign new_new_n54670__ = ~new_new_n54668__ & ~new_new_n54669__;
  assign new_new_n54671__ = new_new_n54667__ & new_new_n54670__;
  assign new_new_n54672__ = new_new_n54664__ & new_new_n54671__;
  assign new_new_n54673__ = ys__n39768 & new_new_n52301__;
  assign new_new_n54674__ = ys__n39766 & new_new_n52304__;
  assign new_new_n54675__ = ~new_new_n54673__ & ~new_new_n54674__;
  assign new_new_n54676__ = ys__n33733 & new_new_n52308__;
  assign new_new_n54677__ = ~ys__n33733 & new_new_n52311__;
  assign new_new_n54678__ = ~new_new_n54676__ & ~new_new_n54677__;
  assign new_new_n54679__ = new_new_n54675__ & new_new_n54678__;
  assign new_new_n54680__ = ys__n24822 & new_new_n52316__;
  assign new_new_n54681__ = ys__n24819 & new_new_n52318__;
  assign new_new_n54682__ = ~new_new_n54680__ & ~new_new_n54681__;
  assign new_new_n54683__ = ys__n24816 & new_new_n52322__;
  assign new_new_n54684__ = ys__n39770 & new_new_n52324__;
  assign new_new_n54685__ = ~new_new_n54683__ & ~new_new_n54684__;
  assign new_new_n54686__ = new_new_n54682__ & new_new_n54685__;
  assign new_new_n54687__ = new_new_n54679__ & new_new_n54686__;
  assign new_new_n54688__ = ~new_new_n54672__ & ~new_new_n54687__;
  assign new_new_n54689__ = ys__n39756 & new_new_n52449__;
  assign new_new_n54690__ = ys__n39754 & new_new_n52448__;
  assign new_new_n54691__ = ~new_new_n54689__ & ~new_new_n54690__;
  assign new_new_n54692__ = ys__n33721 & new_new_n52462__;
  assign new_new_n54693__ = ~ys__n33721 & new_new_n52465__;
  assign new_new_n54694__ = ~new_new_n54692__ & ~new_new_n54693__;
  assign new_new_n54695__ = new_new_n54691__ & new_new_n54694__;
  assign new_new_n54696__ = ys__n24804 & new_new_n52454__;
  assign new_new_n54697__ = ys__n24801 & new_new_n52457__;
  assign new_new_n54698__ = ~new_new_n54696__ & ~new_new_n54697__;
  assign new_new_n54699__ = ys__n24798 & new_new_n52456__;
  assign new_new_n54700__ = ys__n39758 & new_new_n52446__;
  assign new_new_n54701__ = ~new_new_n54699__ & ~new_new_n54700__;
  assign new_new_n54702__ = new_new_n54698__ & new_new_n54701__;
  assign new_new_n54703__ = new_new_n54695__ & new_new_n54702__;
  assign new_new_n54704__ = ~new_new_n54672__ & ~new_new_n54703__;
  assign new_new_n54705__ = ~new_new_n54687__ & ~new_new_n54703__;
  assign new_new_n54706__ = ~new_new_n54704__ & ~new_new_n54705__;
  assign new_new_n54707__ = ~new_new_n54688__ & new_new_n54706__;
  assign new_new_n54708__ = ~new_new_n54657__ & ~new_new_n54707__;
  assign new_new_n54709__ = ys__n39744 & new_new_n52359__;
  assign new_new_n54710__ = ys__n39742 & new_new_n52358__;
  assign new_new_n54711__ = ~new_new_n54709__ & ~new_new_n54710__;
  assign new_new_n54712__ = ys__n33709 & new_new_n52372__;
  assign new_new_n54713__ = ~ys__n33709 & new_new_n52375__;
  assign new_new_n54714__ = ~new_new_n54712__ & ~new_new_n54713__;
  assign new_new_n54715__ = new_new_n54711__ & new_new_n54714__;
  assign new_new_n54716__ = ys__n24786 & new_new_n52364__;
  assign new_new_n54717__ = ys__n24783 & new_new_n52367__;
  assign new_new_n54718__ = ~new_new_n54716__ & ~new_new_n54717__;
  assign new_new_n54719__ = ys__n24780 & new_new_n52366__;
  assign new_new_n54720__ = ys__n39746 & new_new_n52356__;
  assign new_new_n54721__ = ~new_new_n54719__ & ~new_new_n54720__;
  assign new_new_n54722__ = new_new_n54718__ & new_new_n54721__;
  assign new_new_n54723__ = new_new_n54715__ & new_new_n54722__;
  assign new_new_n54724__ = ys__n39750 & new_new_n52334__;
  assign new_new_n54725__ = ys__n39748 & new_new_n52333__;
  assign new_new_n54726__ = ~new_new_n54724__ & ~new_new_n54725__;
  assign new_new_n54727__ = ys__n33715 & new_new_n52347__;
  assign new_new_n54728__ = ~ys__n33715 & new_new_n52350__;
  assign new_new_n54729__ = ~new_new_n54727__ & ~new_new_n54728__;
  assign new_new_n54730__ = new_new_n54726__ & new_new_n54729__;
  assign new_new_n54731__ = ys__n24795 & new_new_n52339__;
  assign new_new_n54732__ = ys__n24792 & new_new_n52342__;
  assign new_new_n54733__ = ~new_new_n54731__ & ~new_new_n54732__;
  assign new_new_n54734__ = ys__n24789 & new_new_n52341__;
  assign new_new_n54735__ = ys__n39752 & new_new_n52331__;
  assign new_new_n54736__ = ~new_new_n54734__ & ~new_new_n54735__;
  assign new_new_n54737__ = new_new_n54733__ & new_new_n54736__;
  assign new_new_n54738__ = new_new_n54730__ & new_new_n54737__;
  assign new_new_n54739__ = ~new_new_n54723__ & ~new_new_n54738__;
  assign new_new_n54740__ = ys__n24777 & new_new_n52383__;
  assign new_new_n54741__ = ys__n24774 & new_new_n52384__;
  assign new_new_n54742__ = ~new_new_n54740__ & ~new_new_n54741__;
  assign new_new_n54743__ = ys__n39740 & new_new_n52391__;
  assign new_new_n54744__ = ys__n39738 & new_new_n52392__;
  assign new_new_n54745__ = ~new_new_n54743__ & ~new_new_n54744__;
  assign new_new_n54746__ = new_new_n54742__ & new_new_n54745__;
  assign new_new_n54747__ = ~new_new_n54723__ & ~new_new_n54746__;
  assign new_new_n54748__ = ~new_new_n54738__ & ~new_new_n54746__;
  assign new_new_n54749__ = ~new_new_n54747__ & ~new_new_n54748__;
  assign new_new_n54750__ = ~new_new_n54739__ & new_new_n54749__;
  assign new_new_n54751__ = ~new_new_n54657__ & ~new_new_n54750__;
  assign new_new_n54752__ = ~new_new_n54707__ & ~new_new_n54750__;
  assign new_new_n54753__ = ~new_new_n54751__ & ~new_new_n54752__;
  assign new_new_n54754__ = ~new_new_n54708__ & new_new_n54753__;
  assign new_new_n54755__ = ~new_new_n54636__ & ~new_new_n54754__;
  assign new_new_n54756__ = ~new_new_n54646__ & ~new_new_n54754__;
  assign new_new_n54757__ = ~new_new_n54755__ & ~new_new_n54756__;
  assign ys__n43133 = new_new_n54647__ | ~new_new_n54757__;
  assign new_new_n54759__ = ~new_new_n54646__ & new_new_n54755__;
  assign new_new_n54760__ = new_new_n54646__ & ~new_new_n54754__;
  assign new_new_n54761__ = new_new_n54636__ & new_new_n54760__;
  assign new_new_n54762__ = ~new_new_n54646__ & new_new_n54754__;
  assign new_new_n54763__ = new_new_n54636__ & new_new_n54762__;
  assign new_new_n54764__ = new_new_n54646__ & new_new_n54754__;
  assign new_new_n54765__ = ~new_new_n54636__ & new_new_n54764__;
  assign new_new_n54766__ = ~new_new_n54763__ & ~new_new_n54765__;
  assign new_new_n54767__ = ~new_new_n54761__ & new_new_n54766__;
  assign ys__n43138 = new_new_n54759__ | ~new_new_n54767__;
  assign new_new_n54769__ = ~new_new_n54707__ & new_new_n54751__;
  assign new_new_n54770__ = new_new_n54707__ & ~new_new_n54750__;
  assign new_new_n54771__ = new_new_n54657__ & new_new_n54770__;
  assign new_new_n54772__ = ~new_new_n54707__ & new_new_n54750__;
  assign new_new_n54773__ = new_new_n54657__ & new_new_n54772__;
  assign new_new_n54774__ = new_new_n54707__ & new_new_n54750__;
  assign new_new_n54775__ = ~new_new_n54657__ & new_new_n54774__;
  assign new_new_n54776__ = ~new_new_n54773__ & ~new_new_n54775__;
  assign new_new_n54777__ = ~new_new_n54771__ & new_new_n54776__;
  assign new_new_n54778__ = ~new_new_n54769__ & new_new_n54777__;
  assign new_new_n54779__ = ~new_new_n54545__ & new_new_n54562__;
  assign new_new_n54780__ = new_new_n54530__ & new_new_n54561__;
  assign new_new_n54781__ = ~new_new_n54545__ & new_new_n54780__;
  assign new_new_n54782__ = ~new_new_n54779__ & ~new_new_n54781__;
  assign new_new_n54783__ = ~new_new_n54530__ & new_new_n54561__;
  assign new_new_n54784__ = new_new_n54545__ & new_new_n54783__;
  assign new_new_n54785__ = new_new_n54530__ & ~new_new_n54561__;
  assign new_new_n54786__ = new_new_n54545__ & new_new_n54785__;
  assign new_new_n54787__ = ~new_new_n54784__ & ~new_new_n54786__;
  assign new_new_n54788__ = new_new_n54782__ & new_new_n54787__;
  assign new_new_n54789__ = ~new_new_n54778__ & ~new_new_n54788__;
  assign new_new_n54790__ = ~new_new_n54738__ & new_new_n54747__;
  assign new_new_n54791__ = new_new_n54723__ & new_new_n54746__;
  assign new_new_n54792__ = ~new_new_n54738__ & new_new_n54791__;
  assign new_new_n54793__ = ~new_new_n54790__ & ~new_new_n54792__;
  assign new_new_n54794__ = ~new_new_n54723__ & new_new_n54746__;
  assign new_new_n54795__ = new_new_n54738__ & new_new_n54794__;
  assign new_new_n54796__ = new_new_n54723__ & ~new_new_n54746__;
  assign new_new_n54797__ = new_new_n54738__ & new_new_n54796__;
  assign new_new_n54798__ = ~new_new_n54795__ & ~new_new_n54797__;
  assign new_new_n54799__ = new_new_n54793__ & new_new_n54798__;
  assign new_new_n54800__ = ys__n39760 & new_new_n52412__;
  assign new_new_n54801__ = ys__n39758 & new_new_n52411__;
  assign new_new_n54802__ = ~new_new_n54800__ & ~new_new_n54801__;
  assign new_new_n54803__ = ys__n33725 & new_new_n52425__;
  assign new_new_n54804__ = ~ys__n33725 & new_new_n52428__;
  assign new_new_n54805__ = ~new_new_n54803__ & ~new_new_n54804__;
  assign new_new_n54806__ = new_new_n54802__ & new_new_n54805__;
  assign new_new_n54807__ = ys__n24810 & new_new_n52417__;
  assign new_new_n54808__ = ys__n24807 & new_new_n52420__;
  assign new_new_n54809__ = ~new_new_n54807__ & ~new_new_n54808__;
  assign new_new_n54810__ = ys__n24804 & new_new_n52419__;
  assign new_new_n54811__ = ys__n39762 & new_new_n52409__;
  assign new_new_n54812__ = ~new_new_n54810__ & ~new_new_n54811__;
  assign new_new_n54813__ = new_new_n54809__ & new_new_n54812__;
  assign new_new_n54814__ = new_new_n54806__ & new_new_n54813__;
  assign new_new_n54815__ = ys__n39766 & new_new_n52301__;
  assign new_new_n54816__ = ys__n39764 & new_new_n52304__;
  assign new_new_n54817__ = ~new_new_n54815__ & ~new_new_n54816__;
  assign new_new_n54818__ = ys__n33731 & new_new_n52308__;
  assign new_new_n54819__ = ~ys__n33731 & new_new_n52311__;
  assign new_new_n54820__ = ~new_new_n54818__ & ~new_new_n54819__;
  assign new_new_n54821__ = new_new_n54817__ & new_new_n54820__;
  assign new_new_n54822__ = ys__n24819 & new_new_n52316__;
  assign new_new_n54823__ = ys__n24816 & new_new_n52318__;
  assign new_new_n54824__ = ~new_new_n54822__ & ~new_new_n54823__;
  assign new_new_n54825__ = ys__n24813 & new_new_n52322__;
  assign new_new_n54826__ = ys__n39768 & new_new_n52324__;
  assign new_new_n54827__ = ~new_new_n54825__ & ~new_new_n54826__;
  assign new_new_n54828__ = new_new_n54824__ & new_new_n54827__;
  assign new_new_n54829__ = new_new_n54821__ & new_new_n54828__;
  assign new_new_n54830__ = ~new_new_n54814__ & ~new_new_n54829__;
  assign new_new_n54831__ = ys__n39754 & new_new_n52449__;
  assign new_new_n54832__ = ys__n39752 & new_new_n52448__;
  assign new_new_n54833__ = ~new_new_n54831__ & ~new_new_n54832__;
  assign new_new_n54834__ = ys__n33719 & new_new_n52462__;
  assign new_new_n54835__ = ~ys__n33719 & new_new_n52465__;
  assign new_new_n54836__ = ~new_new_n54834__ & ~new_new_n54835__;
  assign new_new_n54837__ = new_new_n54833__ & new_new_n54836__;
  assign new_new_n54838__ = ys__n24801 & new_new_n52454__;
  assign new_new_n54839__ = ys__n24798 & new_new_n52457__;
  assign new_new_n54840__ = ~new_new_n54838__ & ~new_new_n54839__;
  assign new_new_n54841__ = ys__n24795 & new_new_n52456__;
  assign new_new_n54842__ = ys__n39756 & new_new_n52446__;
  assign new_new_n54843__ = ~new_new_n54841__ & ~new_new_n54842__;
  assign new_new_n54844__ = new_new_n54840__ & new_new_n54843__;
  assign new_new_n54845__ = new_new_n54837__ & new_new_n54844__;
  assign new_new_n54846__ = ~new_new_n54814__ & ~new_new_n54845__;
  assign new_new_n54847__ = ~new_new_n54829__ & ~new_new_n54845__;
  assign new_new_n54848__ = ~new_new_n54846__ & ~new_new_n54847__;
  assign new_new_n54849__ = ~new_new_n54830__ & new_new_n54848__;
  assign new_new_n54850__ = ~new_new_n54799__ & ~new_new_n54849__;
  assign new_new_n54851__ = ys__n39742 & new_new_n52359__;
  assign new_new_n54852__ = ys__n39740 & new_new_n52358__;
  assign new_new_n54853__ = ~new_new_n54851__ & ~new_new_n54852__;
  assign new_new_n54854__ = ys__n33707 & new_new_n52372__;
  assign new_new_n54855__ = ~ys__n33707 & new_new_n52375__;
  assign new_new_n54856__ = ~new_new_n54854__ & ~new_new_n54855__;
  assign new_new_n54857__ = new_new_n54853__ & new_new_n54856__;
  assign new_new_n54858__ = ys__n24783 & new_new_n52364__;
  assign new_new_n54859__ = ys__n24780 & new_new_n52367__;
  assign new_new_n54860__ = ~new_new_n54858__ & ~new_new_n54859__;
  assign new_new_n54861__ = ys__n24777 & new_new_n52366__;
  assign new_new_n54862__ = ys__n39744 & new_new_n52356__;
  assign new_new_n54863__ = ~new_new_n54861__ & ~new_new_n54862__;
  assign new_new_n54864__ = new_new_n54860__ & new_new_n54863__;
  assign new_new_n54865__ = new_new_n54857__ & new_new_n54864__;
  assign new_new_n54866__ = ys__n39748 & new_new_n52334__;
  assign new_new_n54867__ = ys__n39746 & new_new_n52333__;
  assign new_new_n54868__ = ~new_new_n54866__ & ~new_new_n54867__;
  assign new_new_n54869__ = ys__n33713 & new_new_n52347__;
  assign new_new_n54870__ = ~ys__n33713 & new_new_n52350__;
  assign new_new_n54871__ = ~new_new_n54869__ & ~new_new_n54870__;
  assign new_new_n54872__ = new_new_n54868__ & new_new_n54871__;
  assign new_new_n54873__ = ys__n24792 & new_new_n52339__;
  assign new_new_n54874__ = ys__n24789 & new_new_n52342__;
  assign new_new_n54875__ = ~new_new_n54873__ & ~new_new_n54874__;
  assign new_new_n54876__ = ys__n24786 & new_new_n52341__;
  assign new_new_n54877__ = ys__n39750 & new_new_n52331__;
  assign new_new_n54878__ = ~new_new_n54876__ & ~new_new_n54877__;
  assign new_new_n54879__ = new_new_n54875__ & new_new_n54878__;
  assign new_new_n54880__ = new_new_n54872__ & new_new_n54879__;
  assign new_new_n54881__ = ~new_new_n54865__ & ~new_new_n54880__;
  assign new_new_n54882__ = ys__n24774 & new_new_n52383__;
  assign new_new_n54883__ = ys__n24771 & new_new_n52384__;
  assign new_new_n54884__ = ~new_new_n54882__ & ~new_new_n54883__;
  assign new_new_n54885__ = ys__n39738 & new_new_n52391__;
  assign new_new_n54886__ = ys__n39736 & new_new_n52392__;
  assign new_new_n54887__ = ~new_new_n54885__ & ~new_new_n54886__;
  assign new_new_n54888__ = new_new_n54884__ & new_new_n54887__;
  assign new_new_n54889__ = ~new_new_n54865__ & ~new_new_n54888__;
  assign new_new_n54890__ = ~new_new_n54880__ & ~new_new_n54888__;
  assign new_new_n54891__ = ~new_new_n54889__ & ~new_new_n54890__;
  assign new_new_n54892__ = ~new_new_n54881__ & new_new_n54891__;
  assign new_new_n54893__ = ~new_new_n54799__ & ~new_new_n54892__;
  assign new_new_n54894__ = ~new_new_n54849__ & ~new_new_n54892__;
  assign new_new_n54895__ = ~new_new_n54893__ & ~new_new_n54894__;
  assign new_new_n54896__ = ~new_new_n54850__ & new_new_n54895__;
  assign new_new_n54897__ = ~new_new_n54778__ & ~new_new_n54896__;
  assign new_new_n54898__ = ~new_new_n54788__ & ~new_new_n54896__;
  assign new_new_n54899__ = ~new_new_n54897__ & ~new_new_n54898__;
  assign ys__n43187 = new_new_n54789__ | ~new_new_n54899__;
  assign new_new_n54901__ = ~new_new_n54788__ & new_new_n54897__;
  assign new_new_n54902__ = new_new_n54788__ & ~new_new_n54896__;
  assign new_new_n54903__ = new_new_n54778__ & new_new_n54902__;
  assign new_new_n54904__ = ~new_new_n54788__ & new_new_n54896__;
  assign new_new_n54905__ = new_new_n54778__ & new_new_n54904__;
  assign new_new_n54906__ = new_new_n54788__ & new_new_n54896__;
  assign new_new_n54907__ = ~new_new_n54778__ & new_new_n54906__;
  assign new_new_n54908__ = ~new_new_n54905__ & ~new_new_n54907__;
  assign new_new_n54909__ = ~new_new_n54903__ & new_new_n54908__;
  assign ys__n43192 = new_new_n54901__ | ~new_new_n54909__;
  assign new_new_n54911__ = ~new_new_n54849__ & new_new_n54893__;
  assign new_new_n54912__ = new_new_n54849__ & ~new_new_n54892__;
  assign new_new_n54913__ = new_new_n54799__ & new_new_n54912__;
  assign new_new_n54914__ = ~new_new_n54849__ & new_new_n54892__;
  assign new_new_n54915__ = new_new_n54799__ & new_new_n54914__;
  assign new_new_n54916__ = new_new_n54849__ & new_new_n54892__;
  assign new_new_n54917__ = ~new_new_n54799__ & new_new_n54916__;
  assign new_new_n54918__ = ~new_new_n54915__ & ~new_new_n54917__;
  assign new_new_n54919__ = ~new_new_n54913__ & new_new_n54918__;
  assign new_new_n54920__ = ~new_new_n54911__ & new_new_n54919__;
  assign new_new_n54921__ = ~new_new_n54687__ & new_new_n54704__;
  assign new_new_n54922__ = new_new_n54672__ & new_new_n54703__;
  assign new_new_n54923__ = ~new_new_n54687__ & new_new_n54922__;
  assign new_new_n54924__ = ~new_new_n54921__ & ~new_new_n54923__;
  assign new_new_n54925__ = ~new_new_n54672__ & new_new_n54703__;
  assign new_new_n54926__ = new_new_n54687__ & new_new_n54925__;
  assign new_new_n54927__ = new_new_n54672__ & ~new_new_n54703__;
  assign new_new_n54928__ = new_new_n54687__ & new_new_n54927__;
  assign new_new_n54929__ = ~new_new_n54926__ & ~new_new_n54928__;
  assign new_new_n54930__ = new_new_n54924__ & new_new_n54929__;
  assign new_new_n54931__ = ~new_new_n54920__ & ~new_new_n54930__;
  assign new_new_n54932__ = ~new_new_n54880__ & new_new_n54889__;
  assign new_new_n54933__ = new_new_n54865__ & new_new_n54888__;
  assign new_new_n54934__ = ~new_new_n54880__ & new_new_n54933__;
  assign new_new_n54935__ = ~new_new_n54932__ & ~new_new_n54934__;
  assign new_new_n54936__ = ~new_new_n54865__ & new_new_n54888__;
  assign new_new_n54937__ = new_new_n54880__ & new_new_n54936__;
  assign new_new_n54938__ = new_new_n54865__ & ~new_new_n54888__;
  assign new_new_n54939__ = new_new_n54880__ & new_new_n54938__;
  assign new_new_n54940__ = ~new_new_n54937__ & ~new_new_n54939__;
  assign new_new_n54941__ = new_new_n54935__ & new_new_n54940__;
  assign new_new_n54942__ = ys__n39758 & new_new_n52412__;
  assign new_new_n54943__ = ys__n39756 & new_new_n52411__;
  assign new_new_n54944__ = ~new_new_n54942__ & ~new_new_n54943__;
  assign new_new_n54945__ = ys__n33723 & new_new_n52425__;
  assign new_new_n54946__ = ~ys__n33723 & new_new_n52428__;
  assign new_new_n54947__ = ~new_new_n54945__ & ~new_new_n54946__;
  assign new_new_n54948__ = new_new_n54944__ & new_new_n54947__;
  assign new_new_n54949__ = ys__n24807 & new_new_n52417__;
  assign new_new_n54950__ = ys__n24804 & new_new_n52420__;
  assign new_new_n54951__ = ~new_new_n54949__ & ~new_new_n54950__;
  assign new_new_n54952__ = ys__n24801 & new_new_n52419__;
  assign new_new_n54953__ = ys__n39760 & new_new_n52409__;
  assign new_new_n54954__ = ~new_new_n54952__ & ~new_new_n54953__;
  assign new_new_n54955__ = new_new_n54951__ & new_new_n54954__;
  assign new_new_n54956__ = new_new_n54948__ & new_new_n54955__;
  assign new_new_n54957__ = ys__n39764 & new_new_n52301__;
  assign new_new_n54958__ = ys__n39762 & new_new_n52304__;
  assign new_new_n54959__ = ~new_new_n54957__ & ~new_new_n54958__;
  assign new_new_n54960__ = ys__n33729 & new_new_n52308__;
  assign new_new_n54961__ = ~ys__n33729 & new_new_n52311__;
  assign new_new_n54962__ = ~new_new_n54960__ & ~new_new_n54961__;
  assign new_new_n54963__ = new_new_n54959__ & new_new_n54962__;
  assign new_new_n54964__ = ys__n24816 & new_new_n52316__;
  assign new_new_n54965__ = ys__n24813 & new_new_n52318__;
  assign new_new_n54966__ = ~new_new_n54964__ & ~new_new_n54965__;
  assign new_new_n54967__ = ys__n24810 & new_new_n52322__;
  assign new_new_n54968__ = ys__n39766 & new_new_n52324__;
  assign new_new_n54969__ = ~new_new_n54967__ & ~new_new_n54968__;
  assign new_new_n54970__ = new_new_n54966__ & new_new_n54969__;
  assign new_new_n54971__ = new_new_n54963__ & new_new_n54970__;
  assign new_new_n54972__ = ~new_new_n54956__ & ~new_new_n54971__;
  assign new_new_n54973__ = ys__n39752 & new_new_n52449__;
  assign new_new_n54974__ = ys__n39750 & new_new_n52448__;
  assign new_new_n54975__ = ~new_new_n54973__ & ~new_new_n54974__;
  assign new_new_n54976__ = ys__n33717 & new_new_n52462__;
  assign new_new_n54977__ = ~ys__n33717 & new_new_n52465__;
  assign new_new_n54978__ = ~new_new_n54976__ & ~new_new_n54977__;
  assign new_new_n54979__ = new_new_n54975__ & new_new_n54978__;
  assign new_new_n54980__ = ys__n24798 & new_new_n52454__;
  assign new_new_n54981__ = ys__n24795 & new_new_n52457__;
  assign new_new_n54982__ = ~new_new_n54980__ & ~new_new_n54981__;
  assign new_new_n54983__ = ys__n24792 & new_new_n52456__;
  assign new_new_n54984__ = ys__n39754 & new_new_n52446__;
  assign new_new_n54985__ = ~new_new_n54983__ & ~new_new_n54984__;
  assign new_new_n54986__ = new_new_n54982__ & new_new_n54985__;
  assign new_new_n54987__ = new_new_n54979__ & new_new_n54986__;
  assign new_new_n54988__ = ~new_new_n54956__ & ~new_new_n54987__;
  assign new_new_n54989__ = ~new_new_n54971__ & ~new_new_n54987__;
  assign new_new_n54990__ = ~new_new_n54988__ & ~new_new_n54989__;
  assign new_new_n54991__ = ~new_new_n54972__ & new_new_n54990__;
  assign new_new_n54992__ = ~new_new_n54941__ & ~new_new_n54991__;
  assign new_new_n54993__ = ys__n39740 & new_new_n52359__;
  assign new_new_n54994__ = ys__n39738 & new_new_n52358__;
  assign new_new_n54995__ = ~new_new_n54993__ & ~new_new_n54994__;
  assign new_new_n54996__ = ys__n33705 & new_new_n52372__;
  assign new_new_n54997__ = ~ys__n33705 & new_new_n52375__;
  assign new_new_n54998__ = ~new_new_n54996__ & ~new_new_n54997__;
  assign new_new_n54999__ = new_new_n54995__ & new_new_n54998__;
  assign new_new_n55000__ = ys__n24780 & new_new_n52364__;
  assign new_new_n55001__ = ys__n24777 & new_new_n52367__;
  assign new_new_n55002__ = ~new_new_n55000__ & ~new_new_n55001__;
  assign new_new_n55003__ = ys__n24774 & new_new_n52366__;
  assign new_new_n55004__ = ys__n39742 & new_new_n52356__;
  assign new_new_n55005__ = ~new_new_n55003__ & ~new_new_n55004__;
  assign new_new_n55006__ = new_new_n55002__ & new_new_n55005__;
  assign new_new_n55007__ = new_new_n54999__ & new_new_n55006__;
  assign new_new_n55008__ = ys__n39746 & new_new_n52334__;
  assign new_new_n55009__ = ys__n39744 & new_new_n52333__;
  assign new_new_n55010__ = ~new_new_n55008__ & ~new_new_n55009__;
  assign new_new_n55011__ = ys__n33711 & new_new_n52347__;
  assign new_new_n55012__ = ~ys__n33711 & new_new_n52350__;
  assign new_new_n55013__ = ~new_new_n55011__ & ~new_new_n55012__;
  assign new_new_n55014__ = new_new_n55010__ & new_new_n55013__;
  assign new_new_n55015__ = ys__n24789 & new_new_n52339__;
  assign new_new_n55016__ = ys__n24786 & new_new_n52342__;
  assign new_new_n55017__ = ~new_new_n55015__ & ~new_new_n55016__;
  assign new_new_n55018__ = ys__n24783 & new_new_n52341__;
  assign new_new_n55019__ = ys__n39748 & new_new_n52331__;
  assign new_new_n55020__ = ~new_new_n55018__ & ~new_new_n55019__;
  assign new_new_n55021__ = new_new_n55017__ & new_new_n55020__;
  assign new_new_n55022__ = new_new_n55014__ & new_new_n55021__;
  assign new_new_n55023__ = ~new_new_n55007__ & ~new_new_n55022__;
  assign new_new_n55024__ = ys__n24771 & new_new_n52383__;
  assign new_new_n55025__ = ys__n24768 & new_new_n52384__;
  assign new_new_n55026__ = ~new_new_n55024__ & ~new_new_n55025__;
  assign new_new_n55027__ = ys__n39736 & new_new_n52391__;
  assign new_new_n55028__ = ys__n39734 & new_new_n52392__;
  assign new_new_n55029__ = ~new_new_n55027__ & ~new_new_n55028__;
  assign new_new_n55030__ = new_new_n55026__ & new_new_n55029__;
  assign new_new_n55031__ = ~new_new_n55007__ & ~new_new_n55030__;
  assign new_new_n55032__ = ~new_new_n55022__ & ~new_new_n55030__;
  assign new_new_n55033__ = ~new_new_n55031__ & ~new_new_n55032__;
  assign new_new_n55034__ = ~new_new_n55023__ & new_new_n55033__;
  assign new_new_n55035__ = ~new_new_n54941__ & ~new_new_n55034__;
  assign new_new_n55036__ = ~new_new_n54991__ & ~new_new_n55034__;
  assign new_new_n55037__ = ~new_new_n55035__ & ~new_new_n55036__;
  assign new_new_n55038__ = ~new_new_n54992__ & new_new_n55037__;
  assign new_new_n55039__ = ~new_new_n54920__ & ~new_new_n55038__;
  assign new_new_n55040__ = ~new_new_n54930__ & ~new_new_n55038__;
  assign new_new_n55041__ = ~new_new_n55039__ & ~new_new_n55040__;
  assign ys__n43241 = new_new_n54931__ | ~new_new_n55041__;
  assign new_new_n55043__ = ~new_new_n54930__ & new_new_n55039__;
  assign new_new_n55044__ = new_new_n54930__ & ~new_new_n55038__;
  assign new_new_n55045__ = new_new_n54920__ & new_new_n55044__;
  assign new_new_n55046__ = ~new_new_n54930__ & new_new_n55038__;
  assign new_new_n55047__ = new_new_n54920__ & new_new_n55046__;
  assign new_new_n55048__ = new_new_n54930__ & new_new_n55038__;
  assign new_new_n55049__ = ~new_new_n54920__ & new_new_n55048__;
  assign new_new_n55050__ = ~new_new_n55047__ & ~new_new_n55049__;
  assign new_new_n55051__ = ~new_new_n55045__ & new_new_n55050__;
  assign ys__n43246 = new_new_n55043__ | ~new_new_n55051__;
  assign new_new_n55053__ = ~new_new_n54991__ & new_new_n55035__;
  assign new_new_n55054__ = new_new_n54991__ & ~new_new_n55034__;
  assign new_new_n55055__ = new_new_n54941__ & new_new_n55054__;
  assign new_new_n55056__ = ~new_new_n54991__ & new_new_n55034__;
  assign new_new_n55057__ = new_new_n54941__ & new_new_n55056__;
  assign new_new_n55058__ = new_new_n54991__ & new_new_n55034__;
  assign new_new_n55059__ = ~new_new_n54941__ & new_new_n55058__;
  assign new_new_n55060__ = ~new_new_n55057__ & ~new_new_n55059__;
  assign new_new_n55061__ = ~new_new_n55055__ & new_new_n55060__;
  assign new_new_n55062__ = ~new_new_n55053__ & new_new_n55061__;
  assign new_new_n55063__ = ~new_new_n54829__ & new_new_n54846__;
  assign new_new_n55064__ = new_new_n54814__ & new_new_n54845__;
  assign new_new_n55065__ = ~new_new_n54829__ & new_new_n55064__;
  assign new_new_n55066__ = ~new_new_n55063__ & ~new_new_n55065__;
  assign new_new_n55067__ = ~new_new_n54814__ & new_new_n54845__;
  assign new_new_n55068__ = new_new_n54829__ & new_new_n55067__;
  assign new_new_n55069__ = new_new_n54814__ & ~new_new_n54845__;
  assign new_new_n55070__ = new_new_n54829__ & new_new_n55069__;
  assign new_new_n55071__ = ~new_new_n55068__ & ~new_new_n55070__;
  assign new_new_n55072__ = new_new_n55066__ & new_new_n55071__;
  assign new_new_n55073__ = ~new_new_n55062__ & ~new_new_n55072__;
  assign new_new_n55074__ = ~new_new_n55022__ & new_new_n55031__;
  assign new_new_n55075__ = new_new_n55007__ & new_new_n55030__;
  assign new_new_n55076__ = ~new_new_n55022__ & new_new_n55075__;
  assign new_new_n55077__ = ~new_new_n55074__ & ~new_new_n55076__;
  assign new_new_n55078__ = ~new_new_n55007__ & new_new_n55030__;
  assign new_new_n55079__ = new_new_n55022__ & new_new_n55078__;
  assign new_new_n55080__ = new_new_n55007__ & ~new_new_n55030__;
  assign new_new_n55081__ = new_new_n55022__ & new_new_n55080__;
  assign new_new_n55082__ = ~new_new_n55079__ & ~new_new_n55081__;
  assign new_new_n55083__ = new_new_n55077__ & new_new_n55082__;
  assign new_new_n55084__ = ys__n39756 & new_new_n52412__;
  assign new_new_n55085__ = ys__n39754 & new_new_n52411__;
  assign new_new_n55086__ = ~new_new_n55084__ & ~new_new_n55085__;
  assign new_new_n55087__ = ys__n33721 & new_new_n52425__;
  assign new_new_n55088__ = ~ys__n33721 & new_new_n52428__;
  assign new_new_n55089__ = ~new_new_n55087__ & ~new_new_n55088__;
  assign new_new_n55090__ = new_new_n55086__ & new_new_n55089__;
  assign new_new_n55091__ = ys__n24804 & new_new_n52417__;
  assign new_new_n55092__ = ys__n24801 & new_new_n52420__;
  assign new_new_n55093__ = ~new_new_n55091__ & ~new_new_n55092__;
  assign new_new_n55094__ = ys__n24798 & new_new_n52419__;
  assign new_new_n55095__ = ys__n39758 & new_new_n52409__;
  assign new_new_n55096__ = ~new_new_n55094__ & ~new_new_n55095__;
  assign new_new_n55097__ = new_new_n55093__ & new_new_n55096__;
  assign new_new_n55098__ = new_new_n55090__ & new_new_n55097__;
  assign new_new_n55099__ = ys__n39762 & new_new_n52301__;
  assign new_new_n55100__ = ys__n39760 & new_new_n52304__;
  assign new_new_n55101__ = ~new_new_n55099__ & ~new_new_n55100__;
  assign new_new_n55102__ = ys__n33727 & new_new_n52308__;
  assign new_new_n55103__ = ~ys__n33727 & new_new_n52311__;
  assign new_new_n55104__ = ~new_new_n55102__ & ~new_new_n55103__;
  assign new_new_n55105__ = new_new_n55101__ & new_new_n55104__;
  assign new_new_n55106__ = ys__n24813 & new_new_n52316__;
  assign new_new_n55107__ = ys__n24810 & new_new_n52318__;
  assign new_new_n55108__ = ~new_new_n55106__ & ~new_new_n55107__;
  assign new_new_n55109__ = ys__n24807 & new_new_n52322__;
  assign new_new_n55110__ = ys__n39764 & new_new_n52324__;
  assign new_new_n55111__ = ~new_new_n55109__ & ~new_new_n55110__;
  assign new_new_n55112__ = new_new_n55108__ & new_new_n55111__;
  assign new_new_n55113__ = new_new_n55105__ & new_new_n55112__;
  assign new_new_n55114__ = ~new_new_n55098__ & ~new_new_n55113__;
  assign new_new_n55115__ = ys__n39750 & new_new_n52449__;
  assign new_new_n55116__ = ys__n39748 & new_new_n52448__;
  assign new_new_n55117__ = ~new_new_n55115__ & ~new_new_n55116__;
  assign new_new_n55118__ = ys__n33715 & new_new_n52462__;
  assign new_new_n55119__ = ~ys__n33715 & new_new_n52465__;
  assign new_new_n55120__ = ~new_new_n55118__ & ~new_new_n55119__;
  assign new_new_n55121__ = new_new_n55117__ & new_new_n55120__;
  assign new_new_n55122__ = ys__n24795 & new_new_n52454__;
  assign new_new_n55123__ = ys__n24792 & new_new_n52457__;
  assign new_new_n55124__ = ~new_new_n55122__ & ~new_new_n55123__;
  assign new_new_n55125__ = ys__n24789 & new_new_n52456__;
  assign new_new_n55126__ = ys__n39752 & new_new_n52446__;
  assign new_new_n55127__ = ~new_new_n55125__ & ~new_new_n55126__;
  assign new_new_n55128__ = new_new_n55124__ & new_new_n55127__;
  assign new_new_n55129__ = new_new_n55121__ & new_new_n55128__;
  assign new_new_n55130__ = ~new_new_n55098__ & ~new_new_n55129__;
  assign new_new_n55131__ = ~new_new_n55113__ & ~new_new_n55129__;
  assign new_new_n55132__ = ~new_new_n55130__ & ~new_new_n55131__;
  assign new_new_n55133__ = ~new_new_n55114__ & new_new_n55132__;
  assign new_new_n55134__ = ~new_new_n55083__ & ~new_new_n55133__;
  assign new_new_n55135__ = ys__n39738 & new_new_n52359__;
  assign new_new_n55136__ = ys__n39736 & new_new_n52358__;
  assign new_new_n55137__ = ~new_new_n55135__ & ~new_new_n55136__;
  assign new_new_n55138__ = ys__n33703 & new_new_n52372__;
  assign new_new_n55139__ = ~ys__n33703 & new_new_n52375__;
  assign new_new_n55140__ = ~new_new_n55138__ & ~new_new_n55139__;
  assign new_new_n55141__ = new_new_n55137__ & new_new_n55140__;
  assign new_new_n55142__ = ys__n24777 & new_new_n52364__;
  assign new_new_n55143__ = ys__n24774 & new_new_n52367__;
  assign new_new_n55144__ = ~new_new_n55142__ & ~new_new_n55143__;
  assign new_new_n55145__ = ys__n24771 & new_new_n52366__;
  assign new_new_n55146__ = ys__n39740 & new_new_n52356__;
  assign new_new_n55147__ = ~new_new_n55145__ & ~new_new_n55146__;
  assign new_new_n55148__ = new_new_n55144__ & new_new_n55147__;
  assign new_new_n55149__ = new_new_n55141__ & new_new_n55148__;
  assign new_new_n55150__ = ys__n39744 & new_new_n52334__;
  assign new_new_n55151__ = ys__n39742 & new_new_n52333__;
  assign new_new_n55152__ = ~new_new_n55150__ & ~new_new_n55151__;
  assign new_new_n55153__ = ys__n33709 & new_new_n52347__;
  assign new_new_n55154__ = ~ys__n33709 & new_new_n52350__;
  assign new_new_n55155__ = ~new_new_n55153__ & ~new_new_n55154__;
  assign new_new_n55156__ = new_new_n55152__ & new_new_n55155__;
  assign new_new_n55157__ = ys__n24786 & new_new_n52339__;
  assign new_new_n55158__ = ys__n24783 & new_new_n52342__;
  assign new_new_n55159__ = ~new_new_n55157__ & ~new_new_n55158__;
  assign new_new_n55160__ = ys__n24780 & new_new_n52341__;
  assign new_new_n55161__ = ys__n39746 & new_new_n52331__;
  assign new_new_n55162__ = ~new_new_n55160__ & ~new_new_n55161__;
  assign new_new_n55163__ = new_new_n55159__ & new_new_n55162__;
  assign new_new_n55164__ = new_new_n55156__ & new_new_n55163__;
  assign new_new_n55165__ = ~new_new_n55149__ & ~new_new_n55164__;
  assign new_new_n55166__ = ys__n24768 & new_new_n52383__;
  assign new_new_n55167__ = ys__n24765 & new_new_n52384__;
  assign new_new_n55168__ = ~new_new_n55166__ & ~new_new_n55167__;
  assign new_new_n55169__ = ys__n39734 & new_new_n52391__;
  assign new_new_n55170__ = ys__n39732 & new_new_n52392__;
  assign new_new_n55171__ = ~new_new_n55169__ & ~new_new_n55170__;
  assign new_new_n55172__ = new_new_n55168__ & new_new_n55171__;
  assign new_new_n55173__ = ~new_new_n55149__ & ~new_new_n55172__;
  assign new_new_n55174__ = ~new_new_n55164__ & ~new_new_n55172__;
  assign new_new_n55175__ = ~new_new_n55173__ & ~new_new_n55174__;
  assign new_new_n55176__ = ~new_new_n55165__ & new_new_n55175__;
  assign new_new_n55177__ = ~new_new_n55083__ & ~new_new_n55176__;
  assign new_new_n55178__ = ~new_new_n55133__ & ~new_new_n55176__;
  assign new_new_n55179__ = ~new_new_n55177__ & ~new_new_n55178__;
  assign new_new_n55180__ = ~new_new_n55134__ & new_new_n55179__;
  assign new_new_n55181__ = ~new_new_n55062__ & ~new_new_n55180__;
  assign new_new_n55182__ = ~new_new_n55072__ & ~new_new_n55180__;
  assign new_new_n55183__ = ~new_new_n55181__ & ~new_new_n55182__;
  assign ys__n43295 = new_new_n55073__ | ~new_new_n55183__;
  assign new_new_n55185__ = ~new_new_n55072__ & new_new_n55181__;
  assign new_new_n55186__ = new_new_n55072__ & ~new_new_n55180__;
  assign new_new_n55187__ = new_new_n55062__ & new_new_n55186__;
  assign new_new_n55188__ = ~new_new_n55072__ & new_new_n55180__;
  assign new_new_n55189__ = new_new_n55062__ & new_new_n55188__;
  assign new_new_n55190__ = new_new_n55072__ & new_new_n55180__;
  assign new_new_n55191__ = ~new_new_n55062__ & new_new_n55190__;
  assign new_new_n55192__ = ~new_new_n55189__ & ~new_new_n55191__;
  assign new_new_n55193__ = ~new_new_n55187__ & new_new_n55192__;
  assign ys__n43300 = new_new_n55185__ | ~new_new_n55193__;
  assign new_new_n55195__ = ~new_new_n55133__ & new_new_n55177__;
  assign new_new_n55196__ = new_new_n55133__ & ~new_new_n55176__;
  assign new_new_n55197__ = new_new_n55083__ & new_new_n55196__;
  assign new_new_n55198__ = ~new_new_n55133__ & new_new_n55176__;
  assign new_new_n55199__ = new_new_n55083__ & new_new_n55198__;
  assign new_new_n55200__ = new_new_n55133__ & new_new_n55176__;
  assign new_new_n55201__ = ~new_new_n55083__ & new_new_n55200__;
  assign new_new_n55202__ = ~new_new_n55199__ & ~new_new_n55201__;
  assign new_new_n55203__ = ~new_new_n55197__ & new_new_n55202__;
  assign new_new_n55204__ = ~new_new_n55195__ & new_new_n55203__;
  assign new_new_n55205__ = ~new_new_n54971__ & new_new_n54988__;
  assign new_new_n55206__ = new_new_n54956__ & new_new_n54987__;
  assign new_new_n55207__ = ~new_new_n54971__ & new_new_n55206__;
  assign new_new_n55208__ = ~new_new_n55205__ & ~new_new_n55207__;
  assign new_new_n55209__ = ~new_new_n54956__ & new_new_n54987__;
  assign new_new_n55210__ = new_new_n54971__ & new_new_n55209__;
  assign new_new_n55211__ = new_new_n54956__ & ~new_new_n54987__;
  assign new_new_n55212__ = new_new_n54971__ & new_new_n55211__;
  assign new_new_n55213__ = ~new_new_n55210__ & ~new_new_n55212__;
  assign new_new_n55214__ = new_new_n55208__ & new_new_n55213__;
  assign new_new_n55215__ = ~new_new_n55204__ & ~new_new_n55214__;
  assign new_new_n55216__ = ~new_new_n55164__ & new_new_n55173__;
  assign new_new_n55217__ = new_new_n55149__ & new_new_n55172__;
  assign new_new_n55218__ = ~new_new_n55164__ & new_new_n55217__;
  assign new_new_n55219__ = ~new_new_n55216__ & ~new_new_n55218__;
  assign new_new_n55220__ = ~new_new_n55149__ & new_new_n55172__;
  assign new_new_n55221__ = new_new_n55164__ & new_new_n55220__;
  assign new_new_n55222__ = new_new_n55149__ & ~new_new_n55172__;
  assign new_new_n55223__ = new_new_n55164__ & new_new_n55222__;
  assign new_new_n55224__ = ~new_new_n55221__ & ~new_new_n55223__;
  assign new_new_n55225__ = new_new_n55219__ & new_new_n55224__;
  assign new_new_n55226__ = ys__n39754 & new_new_n52412__;
  assign new_new_n55227__ = ys__n39752 & new_new_n52411__;
  assign new_new_n55228__ = ~new_new_n55226__ & ~new_new_n55227__;
  assign new_new_n55229__ = ys__n33719 & new_new_n52425__;
  assign new_new_n55230__ = ~ys__n33719 & new_new_n52428__;
  assign new_new_n55231__ = ~new_new_n55229__ & ~new_new_n55230__;
  assign new_new_n55232__ = new_new_n55228__ & new_new_n55231__;
  assign new_new_n55233__ = ys__n24801 & new_new_n52417__;
  assign new_new_n55234__ = ys__n24798 & new_new_n52420__;
  assign new_new_n55235__ = ~new_new_n55233__ & ~new_new_n55234__;
  assign new_new_n55236__ = ys__n24795 & new_new_n52419__;
  assign new_new_n55237__ = ys__n39756 & new_new_n52409__;
  assign new_new_n55238__ = ~new_new_n55236__ & ~new_new_n55237__;
  assign new_new_n55239__ = new_new_n55235__ & new_new_n55238__;
  assign new_new_n55240__ = new_new_n55232__ & new_new_n55239__;
  assign new_new_n55241__ = ys__n39760 & new_new_n52301__;
  assign new_new_n55242__ = ys__n39758 & new_new_n52304__;
  assign new_new_n55243__ = ~new_new_n55241__ & ~new_new_n55242__;
  assign new_new_n55244__ = ys__n33725 & new_new_n52308__;
  assign new_new_n55245__ = ~ys__n33725 & new_new_n52311__;
  assign new_new_n55246__ = ~new_new_n55244__ & ~new_new_n55245__;
  assign new_new_n55247__ = new_new_n55243__ & new_new_n55246__;
  assign new_new_n55248__ = ys__n24810 & new_new_n52316__;
  assign new_new_n55249__ = ys__n24807 & new_new_n52318__;
  assign new_new_n55250__ = ~new_new_n55248__ & ~new_new_n55249__;
  assign new_new_n55251__ = ys__n24804 & new_new_n52322__;
  assign new_new_n55252__ = ys__n39762 & new_new_n52324__;
  assign new_new_n55253__ = ~new_new_n55251__ & ~new_new_n55252__;
  assign new_new_n55254__ = new_new_n55250__ & new_new_n55253__;
  assign new_new_n55255__ = new_new_n55247__ & new_new_n55254__;
  assign new_new_n55256__ = ~new_new_n55240__ & ~new_new_n55255__;
  assign new_new_n55257__ = ys__n39748 & new_new_n52449__;
  assign new_new_n55258__ = ys__n39746 & new_new_n52448__;
  assign new_new_n55259__ = ~new_new_n55257__ & ~new_new_n55258__;
  assign new_new_n55260__ = ys__n33713 & new_new_n52462__;
  assign new_new_n55261__ = ~ys__n33713 & new_new_n52465__;
  assign new_new_n55262__ = ~new_new_n55260__ & ~new_new_n55261__;
  assign new_new_n55263__ = new_new_n55259__ & new_new_n55262__;
  assign new_new_n55264__ = ys__n24792 & new_new_n52454__;
  assign new_new_n55265__ = ys__n24789 & new_new_n52457__;
  assign new_new_n55266__ = ~new_new_n55264__ & ~new_new_n55265__;
  assign new_new_n55267__ = ys__n24786 & new_new_n52456__;
  assign new_new_n55268__ = ys__n39750 & new_new_n52446__;
  assign new_new_n55269__ = ~new_new_n55267__ & ~new_new_n55268__;
  assign new_new_n55270__ = new_new_n55266__ & new_new_n55269__;
  assign new_new_n55271__ = new_new_n55263__ & new_new_n55270__;
  assign new_new_n55272__ = ~new_new_n55240__ & ~new_new_n55271__;
  assign new_new_n55273__ = ~new_new_n55255__ & ~new_new_n55271__;
  assign new_new_n55274__ = ~new_new_n55272__ & ~new_new_n55273__;
  assign new_new_n55275__ = ~new_new_n55256__ & new_new_n55274__;
  assign new_new_n55276__ = ~new_new_n55225__ & ~new_new_n55275__;
  assign new_new_n55277__ = ys__n39736 & new_new_n52359__;
  assign new_new_n55278__ = ys__n39734 & new_new_n52358__;
  assign new_new_n55279__ = ~new_new_n55277__ & ~new_new_n55278__;
  assign new_new_n55280__ = ys__n33701 & new_new_n52372__;
  assign new_new_n55281__ = ~ys__n33701 & new_new_n52375__;
  assign new_new_n55282__ = ~new_new_n55280__ & ~new_new_n55281__;
  assign new_new_n55283__ = new_new_n55279__ & new_new_n55282__;
  assign new_new_n55284__ = ys__n24774 & new_new_n52364__;
  assign new_new_n55285__ = ys__n24771 & new_new_n52367__;
  assign new_new_n55286__ = ~new_new_n55284__ & ~new_new_n55285__;
  assign new_new_n55287__ = ys__n24768 & new_new_n52366__;
  assign new_new_n55288__ = ys__n39738 & new_new_n52356__;
  assign new_new_n55289__ = ~new_new_n55287__ & ~new_new_n55288__;
  assign new_new_n55290__ = new_new_n55286__ & new_new_n55289__;
  assign new_new_n55291__ = new_new_n55283__ & new_new_n55290__;
  assign new_new_n55292__ = ys__n39742 & new_new_n52334__;
  assign new_new_n55293__ = ys__n39740 & new_new_n52333__;
  assign new_new_n55294__ = ~new_new_n55292__ & ~new_new_n55293__;
  assign new_new_n55295__ = ys__n33707 & new_new_n52347__;
  assign new_new_n55296__ = ~ys__n33707 & new_new_n52350__;
  assign new_new_n55297__ = ~new_new_n55295__ & ~new_new_n55296__;
  assign new_new_n55298__ = new_new_n55294__ & new_new_n55297__;
  assign new_new_n55299__ = ys__n24783 & new_new_n52339__;
  assign new_new_n55300__ = ys__n24780 & new_new_n52342__;
  assign new_new_n55301__ = ~new_new_n55299__ & ~new_new_n55300__;
  assign new_new_n55302__ = ys__n24777 & new_new_n52341__;
  assign new_new_n55303__ = ys__n39744 & new_new_n52331__;
  assign new_new_n55304__ = ~new_new_n55302__ & ~new_new_n55303__;
  assign new_new_n55305__ = new_new_n55301__ & new_new_n55304__;
  assign new_new_n55306__ = new_new_n55298__ & new_new_n55305__;
  assign new_new_n55307__ = ~new_new_n55291__ & ~new_new_n55306__;
  assign new_new_n55308__ = ys__n24765 & new_new_n52383__;
  assign new_new_n55309__ = ys__n24762 & new_new_n52384__;
  assign new_new_n55310__ = ~new_new_n55308__ & ~new_new_n55309__;
  assign new_new_n55311__ = ys__n39732 & new_new_n52391__;
  assign new_new_n55312__ = ys__n39730 & new_new_n52392__;
  assign new_new_n55313__ = ~new_new_n55311__ & ~new_new_n55312__;
  assign new_new_n55314__ = new_new_n55310__ & new_new_n55313__;
  assign new_new_n55315__ = ~new_new_n55291__ & ~new_new_n55314__;
  assign new_new_n55316__ = ~new_new_n55306__ & ~new_new_n55314__;
  assign new_new_n55317__ = ~new_new_n55315__ & ~new_new_n55316__;
  assign new_new_n55318__ = ~new_new_n55307__ & new_new_n55317__;
  assign new_new_n55319__ = ~new_new_n55225__ & ~new_new_n55318__;
  assign new_new_n55320__ = ~new_new_n55275__ & ~new_new_n55318__;
  assign new_new_n55321__ = ~new_new_n55319__ & ~new_new_n55320__;
  assign new_new_n55322__ = ~new_new_n55276__ & new_new_n55321__;
  assign new_new_n55323__ = ~new_new_n55204__ & ~new_new_n55322__;
  assign new_new_n55324__ = ~new_new_n55214__ & ~new_new_n55322__;
  assign new_new_n55325__ = ~new_new_n55323__ & ~new_new_n55324__;
  assign ys__n43349 = new_new_n55215__ | ~new_new_n55325__;
  assign new_new_n55327__ = ~new_new_n55214__ & new_new_n55323__;
  assign new_new_n55328__ = new_new_n55214__ & ~new_new_n55322__;
  assign new_new_n55329__ = new_new_n55204__ & new_new_n55328__;
  assign new_new_n55330__ = ~new_new_n55214__ & new_new_n55322__;
  assign new_new_n55331__ = new_new_n55204__ & new_new_n55330__;
  assign new_new_n55332__ = new_new_n55214__ & new_new_n55322__;
  assign new_new_n55333__ = ~new_new_n55204__ & new_new_n55332__;
  assign new_new_n55334__ = ~new_new_n55331__ & ~new_new_n55333__;
  assign new_new_n55335__ = ~new_new_n55329__ & new_new_n55334__;
  assign ys__n43354 = new_new_n55327__ | ~new_new_n55335__;
  assign new_new_n55337__ = ~new_new_n55275__ & new_new_n55319__;
  assign new_new_n55338__ = new_new_n55275__ & ~new_new_n55318__;
  assign new_new_n55339__ = new_new_n55225__ & new_new_n55338__;
  assign new_new_n55340__ = ~new_new_n55275__ & new_new_n55318__;
  assign new_new_n55341__ = new_new_n55225__ & new_new_n55340__;
  assign new_new_n55342__ = new_new_n55275__ & new_new_n55318__;
  assign new_new_n55343__ = ~new_new_n55225__ & new_new_n55342__;
  assign new_new_n55344__ = ~new_new_n55341__ & ~new_new_n55343__;
  assign new_new_n55345__ = ~new_new_n55339__ & new_new_n55344__;
  assign new_new_n55346__ = ~new_new_n55337__ & new_new_n55345__;
  assign new_new_n55347__ = ~new_new_n55113__ & new_new_n55130__;
  assign new_new_n55348__ = new_new_n55098__ & new_new_n55129__;
  assign new_new_n55349__ = ~new_new_n55113__ & new_new_n55348__;
  assign new_new_n55350__ = ~new_new_n55347__ & ~new_new_n55349__;
  assign new_new_n55351__ = ~new_new_n55098__ & new_new_n55129__;
  assign new_new_n55352__ = new_new_n55113__ & new_new_n55351__;
  assign new_new_n55353__ = new_new_n55098__ & ~new_new_n55129__;
  assign new_new_n55354__ = new_new_n55113__ & new_new_n55353__;
  assign new_new_n55355__ = ~new_new_n55352__ & ~new_new_n55354__;
  assign new_new_n55356__ = new_new_n55350__ & new_new_n55355__;
  assign new_new_n55357__ = ~new_new_n55346__ & ~new_new_n55356__;
  assign new_new_n55358__ = ~new_new_n55306__ & new_new_n55315__;
  assign new_new_n55359__ = new_new_n55291__ & new_new_n55314__;
  assign new_new_n55360__ = ~new_new_n55306__ & new_new_n55359__;
  assign new_new_n55361__ = ~new_new_n55358__ & ~new_new_n55360__;
  assign new_new_n55362__ = ~new_new_n55291__ & new_new_n55314__;
  assign new_new_n55363__ = new_new_n55306__ & new_new_n55362__;
  assign new_new_n55364__ = new_new_n55291__ & ~new_new_n55314__;
  assign new_new_n55365__ = new_new_n55306__ & new_new_n55364__;
  assign new_new_n55366__ = ~new_new_n55363__ & ~new_new_n55365__;
  assign new_new_n55367__ = new_new_n55361__ & new_new_n55366__;
  assign new_new_n55368__ = ys__n39752 & new_new_n52412__;
  assign new_new_n55369__ = ys__n39750 & new_new_n52411__;
  assign new_new_n55370__ = ~new_new_n55368__ & ~new_new_n55369__;
  assign new_new_n55371__ = ys__n33717 & new_new_n52425__;
  assign new_new_n55372__ = ~ys__n33717 & new_new_n52428__;
  assign new_new_n55373__ = ~new_new_n55371__ & ~new_new_n55372__;
  assign new_new_n55374__ = new_new_n55370__ & new_new_n55373__;
  assign new_new_n55375__ = ys__n24798 & new_new_n52417__;
  assign new_new_n55376__ = ys__n24795 & new_new_n52420__;
  assign new_new_n55377__ = ~new_new_n55375__ & ~new_new_n55376__;
  assign new_new_n55378__ = ys__n24792 & new_new_n52419__;
  assign new_new_n55379__ = ys__n39754 & new_new_n52409__;
  assign new_new_n55380__ = ~new_new_n55378__ & ~new_new_n55379__;
  assign new_new_n55381__ = new_new_n55377__ & new_new_n55380__;
  assign new_new_n55382__ = new_new_n55374__ & new_new_n55381__;
  assign new_new_n55383__ = ys__n39758 & new_new_n52301__;
  assign new_new_n55384__ = ys__n39756 & new_new_n52304__;
  assign new_new_n55385__ = ~new_new_n55383__ & ~new_new_n55384__;
  assign new_new_n55386__ = ys__n33723 & new_new_n52308__;
  assign new_new_n55387__ = ~ys__n33723 & new_new_n52311__;
  assign new_new_n55388__ = ~new_new_n55386__ & ~new_new_n55387__;
  assign new_new_n55389__ = new_new_n55385__ & new_new_n55388__;
  assign new_new_n55390__ = ys__n24807 & new_new_n52316__;
  assign new_new_n55391__ = ys__n24804 & new_new_n52318__;
  assign new_new_n55392__ = ~new_new_n55390__ & ~new_new_n55391__;
  assign new_new_n55393__ = ys__n24801 & new_new_n52322__;
  assign new_new_n55394__ = ys__n39760 & new_new_n52324__;
  assign new_new_n55395__ = ~new_new_n55393__ & ~new_new_n55394__;
  assign new_new_n55396__ = new_new_n55392__ & new_new_n55395__;
  assign new_new_n55397__ = new_new_n55389__ & new_new_n55396__;
  assign new_new_n55398__ = ~new_new_n55382__ & ~new_new_n55397__;
  assign new_new_n55399__ = ys__n39746 & new_new_n52449__;
  assign new_new_n55400__ = ys__n39744 & new_new_n52448__;
  assign new_new_n55401__ = ~new_new_n55399__ & ~new_new_n55400__;
  assign new_new_n55402__ = ys__n33711 & new_new_n52462__;
  assign new_new_n55403__ = ~ys__n33711 & new_new_n52465__;
  assign new_new_n55404__ = ~new_new_n55402__ & ~new_new_n55403__;
  assign new_new_n55405__ = new_new_n55401__ & new_new_n55404__;
  assign new_new_n55406__ = ys__n24789 & new_new_n52454__;
  assign new_new_n55407__ = ys__n24786 & new_new_n52457__;
  assign new_new_n55408__ = ~new_new_n55406__ & ~new_new_n55407__;
  assign new_new_n55409__ = ys__n24783 & new_new_n52456__;
  assign new_new_n55410__ = ys__n39748 & new_new_n52446__;
  assign new_new_n55411__ = ~new_new_n55409__ & ~new_new_n55410__;
  assign new_new_n55412__ = new_new_n55408__ & new_new_n55411__;
  assign new_new_n55413__ = new_new_n55405__ & new_new_n55412__;
  assign new_new_n55414__ = ~new_new_n55382__ & ~new_new_n55413__;
  assign new_new_n55415__ = ~new_new_n55397__ & ~new_new_n55413__;
  assign new_new_n55416__ = ~new_new_n55414__ & ~new_new_n55415__;
  assign new_new_n55417__ = ~new_new_n55398__ & new_new_n55416__;
  assign new_new_n55418__ = ~new_new_n55367__ & ~new_new_n55417__;
  assign new_new_n55419__ = ys__n39734 & new_new_n52359__;
  assign new_new_n55420__ = ys__n39732 & new_new_n52358__;
  assign new_new_n55421__ = ~new_new_n55419__ & ~new_new_n55420__;
  assign new_new_n55422__ = ys__n33699 & new_new_n52372__;
  assign new_new_n55423__ = ~ys__n33699 & new_new_n52375__;
  assign new_new_n55424__ = ~new_new_n55422__ & ~new_new_n55423__;
  assign new_new_n55425__ = new_new_n55421__ & new_new_n55424__;
  assign new_new_n55426__ = ys__n24771 & new_new_n52364__;
  assign new_new_n55427__ = ys__n24768 & new_new_n52367__;
  assign new_new_n55428__ = ~new_new_n55426__ & ~new_new_n55427__;
  assign new_new_n55429__ = ys__n24765 & new_new_n52366__;
  assign new_new_n55430__ = ys__n39736 & new_new_n52356__;
  assign new_new_n55431__ = ~new_new_n55429__ & ~new_new_n55430__;
  assign new_new_n55432__ = new_new_n55428__ & new_new_n55431__;
  assign new_new_n55433__ = new_new_n55425__ & new_new_n55432__;
  assign new_new_n55434__ = ys__n39740 & new_new_n52334__;
  assign new_new_n55435__ = ys__n39738 & new_new_n52333__;
  assign new_new_n55436__ = ~new_new_n55434__ & ~new_new_n55435__;
  assign new_new_n55437__ = ys__n33705 & new_new_n52347__;
  assign new_new_n55438__ = ~ys__n33705 & new_new_n52350__;
  assign new_new_n55439__ = ~new_new_n55437__ & ~new_new_n55438__;
  assign new_new_n55440__ = new_new_n55436__ & new_new_n55439__;
  assign new_new_n55441__ = ys__n24780 & new_new_n52339__;
  assign new_new_n55442__ = ys__n24777 & new_new_n52342__;
  assign new_new_n55443__ = ~new_new_n55441__ & ~new_new_n55442__;
  assign new_new_n55444__ = ys__n24774 & new_new_n52341__;
  assign new_new_n55445__ = ys__n39742 & new_new_n52331__;
  assign new_new_n55446__ = ~new_new_n55444__ & ~new_new_n55445__;
  assign new_new_n55447__ = new_new_n55443__ & new_new_n55446__;
  assign new_new_n55448__ = new_new_n55440__ & new_new_n55447__;
  assign new_new_n55449__ = ~new_new_n55433__ & ~new_new_n55448__;
  assign new_new_n55450__ = ys__n24762 & new_new_n52383__;
  assign new_new_n55451__ = ys__n24759 & new_new_n52384__;
  assign new_new_n55452__ = ~new_new_n55450__ & ~new_new_n55451__;
  assign new_new_n55453__ = ys__n39730 & new_new_n52391__;
  assign new_new_n55454__ = ys__n39728 & new_new_n52392__;
  assign new_new_n55455__ = ~new_new_n55453__ & ~new_new_n55454__;
  assign new_new_n55456__ = new_new_n55452__ & new_new_n55455__;
  assign new_new_n55457__ = ~new_new_n55433__ & ~new_new_n55456__;
  assign new_new_n55458__ = ~new_new_n55448__ & ~new_new_n55456__;
  assign new_new_n55459__ = ~new_new_n55457__ & ~new_new_n55458__;
  assign new_new_n55460__ = ~new_new_n55449__ & new_new_n55459__;
  assign new_new_n55461__ = ~new_new_n55367__ & ~new_new_n55460__;
  assign new_new_n55462__ = ~new_new_n55417__ & ~new_new_n55460__;
  assign new_new_n55463__ = ~new_new_n55461__ & ~new_new_n55462__;
  assign new_new_n55464__ = ~new_new_n55418__ & new_new_n55463__;
  assign new_new_n55465__ = ~new_new_n55346__ & ~new_new_n55464__;
  assign new_new_n55466__ = ~new_new_n55356__ & ~new_new_n55464__;
  assign new_new_n55467__ = ~new_new_n55465__ & ~new_new_n55466__;
  assign ys__n43403 = new_new_n55357__ | ~new_new_n55467__;
  assign new_new_n55469__ = ~new_new_n55356__ & new_new_n55465__;
  assign new_new_n55470__ = new_new_n55356__ & ~new_new_n55464__;
  assign new_new_n55471__ = new_new_n55346__ & new_new_n55470__;
  assign new_new_n55472__ = ~new_new_n55356__ & new_new_n55464__;
  assign new_new_n55473__ = new_new_n55346__ & new_new_n55472__;
  assign new_new_n55474__ = new_new_n55356__ & new_new_n55464__;
  assign new_new_n55475__ = ~new_new_n55346__ & new_new_n55474__;
  assign new_new_n55476__ = ~new_new_n55473__ & ~new_new_n55475__;
  assign new_new_n55477__ = ~new_new_n55471__ & new_new_n55476__;
  assign ys__n43408 = new_new_n55469__ | ~new_new_n55477__;
  assign new_new_n55479__ = ~new_new_n55417__ & new_new_n55461__;
  assign new_new_n55480__ = new_new_n55417__ & ~new_new_n55460__;
  assign new_new_n55481__ = new_new_n55367__ & new_new_n55480__;
  assign new_new_n55482__ = ~new_new_n55417__ & new_new_n55460__;
  assign new_new_n55483__ = new_new_n55367__ & new_new_n55482__;
  assign new_new_n55484__ = new_new_n55417__ & new_new_n55460__;
  assign new_new_n55485__ = ~new_new_n55367__ & new_new_n55484__;
  assign new_new_n55486__ = ~new_new_n55483__ & ~new_new_n55485__;
  assign new_new_n55487__ = ~new_new_n55481__ & new_new_n55486__;
  assign new_new_n55488__ = ~new_new_n55479__ & new_new_n55487__;
  assign new_new_n55489__ = ~new_new_n55255__ & new_new_n55272__;
  assign new_new_n55490__ = new_new_n55240__ & new_new_n55271__;
  assign new_new_n55491__ = ~new_new_n55255__ & new_new_n55490__;
  assign new_new_n55492__ = ~new_new_n55489__ & ~new_new_n55491__;
  assign new_new_n55493__ = ~new_new_n55240__ & new_new_n55271__;
  assign new_new_n55494__ = new_new_n55255__ & new_new_n55493__;
  assign new_new_n55495__ = new_new_n55240__ & ~new_new_n55271__;
  assign new_new_n55496__ = new_new_n55255__ & new_new_n55495__;
  assign new_new_n55497__ = ~new_new_n55494__ & ~new_new_n55496__;
  assign new_new_n55498__ = new_new_n55492__ & new_new_n55497__;
  assign new_new_n55499__ = ~new_new_n55488__ & ~new_new_n55498__;
  assign new_new_n55500__ = ~new_new_n55448__ & new_new_n55457__;
  assign new_new_n55501__ = new_new_n55433__ & new_new_n55456__;
  assign new_new_n55502__ = ~new_new_n55448__ & new_new_n55501__;
  assign new_new_n55503__ = ~new_new_n55500__ & ~new_new_n55502__;
  assign new_new_n55504__ = ~new_new_n55433__ & new_new_n55456__;
  assign new_new_n55505__ = new_new_n55448__ & new_new_n55504__;
  assign new_new_n55506__ = new_new_n55433__ & ~new_new_n55456__;
  assign new_new_n55507__ = new_new_n55448__ & new_new_n55506__;
  assign new_new_n55508__ = ~new_new_n55505__ & ~new_new_n55507__;
  assign new_new_n55509__ = new_new_n55503__ & new_new_n55508__;
  assign new_new_n55510__ = ys__n39750 & new_new_n52412__;
  assign new_new_n55511__ = ys__n39748 & new_new_n52411__;
  assign new_new_n55512__ = ~new_new_n55510__ & ~new_new_n55511__;
  assign new_new_n55513__ = ys__n33715 & new_new_n52425__;
  assign new_new_n55514__ = ~ys__n33715 & new_new_n52428__;
  assign new_new_n55515__ = ~new_new_n55513__ & ~new_new_n55514__;
  assign new_new_n55516__ = new_new_n55512__ & new_new_n55515__;
  assign new_new_n55517__ = ys__n24795 & new_new_n52417__;
  assign new_new_n55518__ = ys__n24792 & new_new_n52420__;
  assign new_new_n55519__ = ~new_new_n55517__ & ~new_new_n55518__;
  assign new_new_n55520__ = ys__n24789 & new_new_n52419__;
  assign new_new_n55521__ = ys__n39752 & new_new_n52409__;
  assign new_new_n55522__ = ~new_new_n55520__ & ~new_new_n55521__;
  assign new_new_n55523__ = new_new_n55519__ & new_new_n55522__;
  assign new_new_n55524__ = new_new_n55516__ & new_new_n55523__;
  assign new_new_n55525__ = ys__n39756 & new_new_n52301__;
  assign new_new_n55526__ = ys__n39754 & new_new_n52304__;
  assign new_new_n55527__ = ~new_new_n55525__ & ~new_new_n55526__;
  assign new_new_n55528__ = ys__n33721 & new_new_n52308__;
  assign new_new_n55529__ = ~ys__n33721 & new_new_n52311__;
  assign new_new_n55530__ = ~new_new_n55528__ & ~new_new_n55529__;
  assign new_new_n55531__ = new_new_n55527__ & new_new_n55530__;
  assign new_new_n55532__ = ys__n24804 & new_new_n52316__;
  assign new_new_n55533__ = ys__n24801 & new_new_n52318__;
  assign new_new_n55534__ = ~new_new_n55532__ & ~new_new_n55533__;
  assign new_new_n55535__ = ys__n24798 & new_new_n52322__;
  assign new_new_n55536__ = ys__n39758 & new_new_n52324__;
  assign new_new_n55537__ = ~new_new_n55535__ & ~new_new_n55536__;
  assign new_new_n55538__ = new_new_n55534__ & new_new_n55537__;
  assign new_new_n55539__ = new_new_n55531__ & new_new_n55538__;
  assign new_new_n55540__ = ~new_new_n55524__ & ~new_new_n55539__;
  assign new_new_n55541__ = ys__n39744 & new_new_n52449__;
  assign new_new_n55542__ = ys__n39742 & new_new_n52448__;
  assign new_new_n55543__ = ~new_new_n55541__ & ~new_new_n55542__;
  assign new_new_n55544__ = ys__n33709 & new_new_n52462__;
  assign new_new_n55545__ = ~ys__n33709 & new_new_n52465__;
  assign new_new_n55546__ = ~new_new_n55544__ & ~new_new_n55545__;
  assign new_new_n55547__ = new_new_n55543__ & new_new_n55546__;
  assign new_new_n55548__ = ys__n24786 & new_new_n52454__;
  assign new_new_n55549__ = ys__n24783 & new_new_n52457__;
  assign new_new_n55550__ = ~new_new_n55548__ & ~new_new_n55549__;
  assign new_new_n55551__ = ys__n24780 & new_new_n52456__;
  assign new_new_n55552__ = ys__n39746 & new_new_n52446__;
  assign new_new_n55553__ = ~new_new_n55551__ & ~new_new_n55552__;
  assign new_new_n55554__ = new_new_n55550__ & new_new_n55553__;
  assign new_new_n55555__ = new_new_n55547__ & new_new_n55554__;
  assign new_new_n55556__ = ~new_new_n55524__ & ~new_new_n55555__;
  assign new_new_n55557__ = ~new_new_n55539__ & ~new_new_n55555__;
  assign new_new_n55558__ = ~new_new_n55556__ & ~new_new_n55557__;
  assign new_new_n55559__ = ~new_new_n55540__ & new_new_n55558__;
  assign new_new_n55560__ = ~new_new_n55509__ & ~new_new_n55559__;
  assign new_new_n55561__ = ys__n39732 & new_new_n52359__;
  assign new_new_n55562__ = ys__n39730 & new_new_n52358__;
  assign new_new_n55563__ = ~new_new_n55561__ & ~new_new_n55562__;
  assign new_new_n55564__ = ys__n33697 & new_new_n52372__;
  assign new_new_n55565__ = ~ys__n33697 & new_new_n52375__;
  assign new_new_n55566__ = ~new_new_n55564__ & ~new_new_n55565__;
  assign new_new_n55567__ = new_new_n55563__ & new_new_n55566__;
  assign new_new_n55568__ = ys__n24768 & new_new_n52364__;
  assign new_new_n55569__ = ys__n24765 & new_new_n52367__;
  assign new_new_n55570__ = ~new_new_n55568__ & ~new_new_n55569__;
  assign new_new_n55571__ = ys__n24762 & new_new_n52366__;
  assign new_new_n55572__ = ys__n39734 & new_new_n52356__;
  assign new_new_n55573__ = ~new_new_n55571__ & ~new_new_n55572__;
  assign new_new_n55574__ = new_new_n55570__ & new_new_n55573__;
  assign new_new_n55575__ = new_new_n55567__ & new_new_n55574__;
  assign new_new_n55576__ = ys__n39738 & new_new_n52334__;
  assign new_new_n55577__ = ys__n39736 & new_new_n52333__;
  assign new_new_n55578__ = ~new_new_n55576__ & ~new_new_n55577__;
  assign new_new_n55579__ = ys__n33703 & new_new_n52347__;
  assign new_new_n55580__ = ~ys__n33703 & new_new_n52350__;
  assign new_new_n55581__ = ~new_new_n55579__ & ~new_new_n55580__;
  assign new_new_n55582__ = new_new_n55578__ & new_new_n55581__;
  assign new_new_n55583__ = ys__n24777 & new_new_n52339__;
  assign new_new_n55584__ = ys__n24774 & new_new_n52342__;
  assign new_new_n55585__ = ~new_new_n55583__ & ~new_new_n55584__;
  assign new_new_n55586__ = ys__n24771 & new_new_n52341__;
  assign new_new_n55587__ = ys__n39740 & new_new_n52331__;
  assign new_new_n55588__ = ~new_new_n55586__ & ~new_new_n55587__;
  assign new_new_n55589__ = new_new_n55585__ & new_new_n55588__;
  assign new_new_n55590__ = new_new_n55582__ & new_new_n55589__;
  assign new_new_n55591__ = ~new_new_n55575__ & ~new_new_n55590__;
  assign new_new_n55592__ = ys__n24759 & new_new_n52383__;
  assign new_new_n55593__ = ys__n24756 & new_new_n52384__;
  assign new_new_n55594__ = ~new_new_n55592__ & ~new_new_n55593__;
  assign new_new_n55595__ = ys__n39728 & new_new_n52391__;
  assign new_new_n55596__ = ys__n39726 & new_new_n52392__;
  assign new_new_n55597__ = ~new_new_n55595__ & ~new_new_n55596__;
  assign new_new_n55598__ = new_new_n55594__ & new_new_n55597__;
  assign new_new_n55599__ = ~new_new_n55575__ & ~new_new_n55598__;
  assign new_new_n55600__ = ~new_new_n55590__ & ~new_new_n55598__;
  assign new_new_n55601__ = ~new_new_n55599__ & ~new_new_n55600__;
  assign new_new_n55602__ = ~new_new_n55591__ & new_new_n55601__;
  assign new_new_n55603__ = ~new_new_n55509__ & ~new_new_n55602__;
  assign new_new_n55604__ = ~new_new_n55559__ & ~new_new_n55602__;
  assign new_new_n55605__ = ~new_new_n55603__ & ~new_new_n55604__;
  assign new_new_n55606__ = ~new_new_n55560__ & new_new_n55605__;
  assign new_new_n55607__ = ~new_new_n55488__ & ~new_new_n55606__;
  assign new_new_n55608__ = ~new_new_n55498__ & ~new_new_n55606__;
  assign new_new_n55609__ = ~new_new_n55607__ & ~new_new_n55608__;
  assign ys__n43457 = new_new_n55499__ | ~new_new_n55609__;
  assign new_new_n55611__ = ~new_new_n55498__ & new_new_n55607__;
  assign new_new_n55612__ = new_new_n55498__ & ~new_new_n55606__;
  assign new_new_n55613__ = new_new_n55488__ & new_new_n55612__;
  assign new_new_n55614__ = ~new_new_n55498__ & new_new_n55606__;
  assign new_new_n55615__ = new_new_n55488__ & new_new_n55614__;
  assign new_new_n55616__ = new_new_n55498__ & new_new_n55606__;
  assign new_new_n55617__ = ~new_new_n55488__ & new_new_n55616__;
  assign new_new_n55618__ = ~new_new_n55615__ & ~new_new_n55617__;
  assign new_new_n55619__ = ~new_new_n55613__ & new_new_n55618__;
  assign ys__n43462 = new_new_n55611__ | ~new_new_n55619__;
  assign new_new_n55621__ = ~new_new_n55559__ & new_new_n55603__;
  assign new_new_n55622__ = new_new_n55559__ & ~new_new_n55602__;
  assign new_new_n55623__ = new_new_n55509__ & new_new_n55622__;
  assign new_new_n55624__ = ~new_new_n55559__ & new_new_n55602__;
  assign new_new_n55625__ = new_new_n55509__ & new_new_n55624__;
  assign new_new_n55626__ = new_new_n55559__ & new_new_n55602__;
  assign new_new_n55627__ = ~new_new_n55509__ & new_new_n55626__;
  assign new_new_n55628__ = ~new_new_n55625__ & ~new_new_n55627__;
  assign new_new_n55629__ = ~new_new_n55623__ & new_new_n55628__;
  assign new_new_n55630__ = ~new_new_n55621__ & new_new_n55629__;
  assign new_new_n55631__ = ~new_new_n55397__ & new_new_n55414__;
  assign new_new_n55632__ = new_new_n55382__ & new_new_n55413__;
  assign new_new_n55633__ = ~new_new_n55397__ & new_new_n55632__;
  assign new_new_n55634__ = ~new_new_n55631__ & ~new_new_n55633__;
  assign new_new_n55635__ = ~new_new_n55382__ & new_new_n55413__;
  assign new_new_n55636__ = new_new_n55397__ & new_new_n55635__;
  assign new_new_n55637__ = new_new_n55382__ & ~new_new_n55413__;
  assign new_new_n55638__ = new_new_n55397__ & new_new_n55637__;
  assign new_new_n55639__ = ~new_new_n55636__ & ~new_new_n55638__;
  assign new_new_n55640__ = new_new_n55634__ & new_new_n55639__;
  assign new_new_n55641__ = ~new_new_n55630__ & ~new_new_n55640__;
  assign new_new_n55642__ = ~new_new_n55590__ & new_new_n55599__;
  assign new_new_n55643__ = new_new_n55575__ & new_new_n55598__;
  assign new_new_n55644__ = ~new_new_n55590__ & new_new_n55643__;
  assign new_new_n55645__ = ~new_new_n55642__ & ~new_new_n55644__;
  assign new_new_n55646__ = ~new_new_n55575__ & new_new_n55598__;
  assign new_new_n55647__ = new_new_n55590__ & new_new_n55646__;
  assign new_new_n55648__ = new_new_n55575__ & ~new_new_n55598__;
  assign new_new_n55649__ = new_new_n55590__ & new_new_n55648__;
  assign new_new_n55650__ = ~new_new_n55647__ & ~new_new_n55649__;
  assign new_new_n55651__ = new_new_n55645__ & new_new_n55650__;
  assign new_new_n55652__ = ys__n39748 & new_new_n52412__;
  assign new_new_n55653__ = ys__n39746 & new_new_n52411__;
  assign new_new_n55654__ = ~new_new_n55652__ & ~new_new_n55653__;
  assign new_new_n55655__ = ys__n33713 & new_new_n52425__;
  assign new_new_n55656__ = ~ys__n33713 & new_new_n52428__;
  assign new_new_n55657__ = ~new_new_n55655__ & ~new_new_n55656__;
  assign new_new_n55658__ = new_new_n55654__ & new_new_n55657__;
  assign new_new_n55659__ = ys__n24792 & new_new_n52417__;
  assign new_new_n55660__ = ys__n24789 & new_new_n52420__;
  assign new_new_n55661__ = ~new_new_n55659__ & ~new_new_n55660__;
  assign new_new_n55662__ = ys__n24786 & new_new_n52419__;
  assign new_new_n55663__ = ys__n39750 & new_new_n52409__;
  assign new_new_n55664__ = ~new_new_n55662__ & ~new_new_n55663__;
  assign new_new_n55665__ = new_new_n55661__ & new_new_n55664__;
  assign new_new_n55666__ = new_new_n55658__ & new_new_n55665__;
  assign new_new_n55667__ = ys__n39754 & new_new_n52301__;
  assign new_new_n55668__ = ys__n39752 & new_new_n52304__;
  assign new_new_n55669__ = ~new_new_n55667__ & ~new_new_n55668__;
  assign new_new_n55670__ = ys__n33719 & new_new_n52308__;
  assign new_new_n55671__ = ~ys__n33719 & new_new_n52311__;
  assign new_new_n55672__ = ~new_new_n55670__ & ~new_new_n55671__;
  assign new_new_n55673__ = new_new_n55669__ & new_new_n55672__;
  assign new_new_n55674__ = ys__n24801 & new_new_n52316__;
  assign new_new_n55675__ = ys__n24798 & new_new_n52318__;
  assign new_new_n55676__ = ~new_new_n55674__ & ~new_new_n55675__;
  assign new_new_n55677__ = ys__n24795 & new_new_n52322__;
  assign new_new_n55678__ = ys__n39756 & new_new_n52324__;
  assign new_new_n55679__ = ~new_new_n55677__ & ~new_new_n55678__;
  assign new_new_n55680__ = new_new_n55676__ & new_new_n55679__;
  assign new_new_n55681__ = new_new_n55673__ & new_new_n55680__;
  assign new_new_n55682__ = ~new_new_n55666__ & ~new_new_n55681__;
  assign new_new_n55683__ = ys__n39742 & new_new_n52449__;
  assign new_new_n55684__ = ys__n39740 & new_new_n52448__;
  assign new_new_n55685__ = ~new_new_n55683__ & ~new_new_n55684__;
  assign new_new_n55686__ = ys__n33707 & new_new_n52462__;
  assign new_new_n55687__ = ~ys__n33707 & new_new_n52465__;
  assign new_new_n55688__ = ~new_new_n55686__ & ~new_new_n55687__;
  assign new_new_n55689__ = new_new_n55685__ & new_new_n55688__;
  assign new_new_n55690__ = ys__n24783 & new_new_n52454__;
  assign new_new_n55691__ = ys__n24780 & new_new_n52457__;
  assign new_new_n55692__ = ~new_new_n55690__ & ~new_new_n55691__;
  assign new_new_n55693__ = ys__n24777 & new_new_n52456__;
  assign new_new_n55694__ = ys__n39744 & new_new_n52446__;
  assign new_new_n55695__ = ~new_new_n55693__ & ~new_new_n55694__;
  assign new_new_n55696__ = new_new_n55692__ & new_new_n55695__;
  assign new_new_n55697__ = new_new_n55689__ & new_new_n55696__;
  assign new_new_n55698__ = ~new_new_n55666__ & ~new_new_n55697__;
  assign new_new_n55699__ = ~new_new_n55681__ & ~new_new_n55697__;
  assign new_new_n55700__ = ~new_new_n55698__ & ~new_new_n55699__;
  assign new_new_n55701__ = ~new_new_n55682__ & new_new_n55700__;
  assign new_new_n55702__ = ~new_new_n55651__ & ~new_new_n55701__;
  assign new_new_n55703__ = ys__n39730 & new_new_n52359__;
  assign new_new_n55704__ = ys__n39728 & new_new_n52358__;
  assign new_new_n55705__ = ~new_new_n55703__ & ~new_new_n55704__;
  assign new_new_n55706__ = ys__n33695 & new_new_n52372__;
  assign new_new_n55707__ = ~ys__n33695 & new_new_n52375__;
  assign new_new_n55708__ = ~new_new_n55706__ & ~new_new_n55707__;
  assign new_new_n55709__ = new_new_n55705__ & new_new_n55708__;
  assign new_new_n55710__ = ys__n24765 & new_new_n52364__;
  assign new_new_n55711__ = ys__n24762 & new_new_n52367__;
  assign new_new_n55712__ = ~new_new_n55710__ & ~new_new_n55711__;
  assign new_new_n55713__ = ys__n24759 & new_new_n52366__;
  assign new_new_n55714__ = ys__n39732 & new_new_n52356__;
  assign new_new_n55715__ = ~new_new_n55713__ & ~new_new_n55714__;
  assign new_new_n55716__ = new_new_n55712__ & new_new_n55715__;
  assign new_new_n55717__ = new_new_n55709__ & new_new_n55716__;
  assign new_new_n55718__ = ys__n39736 & new_new_n52334__;
  assign new_new_n55719__ = ys__n39734 & new_new_n52333__;
  assign new_new_n55720__ = ~new_new_n55718__ & ~new_new_n55719__;
  assign new_new_n55721__ = ys__n33701 & new_new_n52347__;
  assign new_new_n55722__ = ~ys__n33701 & new_new_n52350__;
  assign new_new_n55723__ = ~new_new_n55721__ & ~new_new_n55722__;
  assign new_new_n55724__ = new_new_n55720__ & new_new_n55723__;
  assign new_new_n55725__ = ys__n24774 & new_new_n52339__;
  assign new_new_n55726__ = ys__n24771 & new_new_n52342__;
  assign new_new_n55727__ = ~new_new_n55725__ & ~new_new_n55726__;
  assign new_new_n55728__ = ys__n24768 & new_new_n52341__;
  assign new_new_n55729__ = ys__n39738 & new_new_n52331__;
  assign new_new_n55730__ = ~new_new_n55728__ & ~new_new_n55729__;
  assign new_new_n55731__ = new_new_n55727__ & new_new_n55730__;
  assign new_new_n55732__ = new_new_n55724__ & new_new_n55731__;
  assign new_new_n55733__ = ~new_new_n55717__ & ~new_new_n55732__;
  assign new_new_n55734__ = ys__n24756 & new_new_n52383__;
  assign new_new_n55735__ = ys__n24753 & new_new_n52384__;
  assign new_new_n55736__ = ~new_new_n55734__ & ~new_new_n55735__;
  assign new_new_n55737__ = ys__n39726 & new_new_n52391__;
  assign new_new_n55738__ = ys__n39724 & new_new_n52392__;
  assign new_new_n55739__ = ~new_new_n55737__ & ~new_new_n55738__;
  assign new_new_n55740__ = new_new_n55736__ & new_new_n55739__;
  assign new_new_n55741__ = ~new_new_n55717__ & ~new_new_n55740__;
  assign new_new_n55742__ = ~new_new_n55732__ & ~new_new_n55740__;
  assign new_new_n55743__ = ~new_new_n55741__ & ~new_new_n55742__;
  assign new_new_n55744__ = ~new_new_n55733__ & new_new_n55743__;
  assign new_new_n55745__ = ~new_new_n55651__ & ~new_new_n55744__;
  assign new_new_n55746__ = ~new_new_n55701__ & ~new_new_n55744__;
  assign new_new_n55747__ = ~new_new_n55745__ & ~new_new_n55746__;
  assign new_new_n55748__ = ~new_new_n55702__ & new_new_n55747__;
  assign new_new_n55749__ = ~new_new_n55630__ & ~new_new_n55748__;
  assign new_new_n55750__ = ~new_new_n55640__ & ~new_new_n55748__;
  assign new_new_n55751__ = ~new_new_n55749__ & ~new_new_n55750__;
  assign ys__n43511 = new_new_n55641__ | ~new_new_n55751__;
  assign new_new_n55753__ = ~new_new_n55640__ & new_new_n55749__;
  assign new_new_n55754__ = new_new_n55640__ & ~new_new_n55748__;
  assign new_new_n55755__ = new_new_n55630__ & new_new_n55754__;
  assign new_new_n55756__ = ~new_new_n55640__ & new_new_n55748__;
  assign new_new_n55757__ = new_new_n55630__ & new_new_n55756__;
  assign new_new_n55758__ = new_new_n55640__ & new_new_n55748__;
  assign new_new_n55759__ = ~new_new_n55630__ & new_new_n55758__;
  assign new_new_n55760__ = ~new_new_n55757__ & ~new_new_n55759__;
  assign new_new_n55761__ = ~new_new_n55755__ & new_new_n55760__;
  assign ys__n43516 = new_new_n55753__ | ~new_new_n55761__;
  assign new_new_n55763__ = ~new_new_n55701__ & new_new_n55745__;
  assign new_new_n55764__ = new_new_n55701__ & ~new_new_n55744__;
  assign new_new_n55765__ = new_new_n55651__ & new_new_n55764__;
  assign new_new_n55766__ = ~new_new_n55701__ & new_new_n55744__;
  assign new_new_n55767__ = new_new_n55651__ & new_new_n55766__;
  assign new_new_n55768__ = new_new_n55701__ & new_new_n55744__;
  assign new_new_n55769__ = ~new_new_n55651__ & new_new_n55768__;
  assign new_new_n55770__ = ~new_new_n55767__ & ~new_new_n55769__;
  assign new_new_n55771__ = ~new_new_n55765__ & new_new_n55770__;
  assign new_new_n55772__ = ~new_new_n55763__ & new_new_n55771__;
  assign new_new_n55773__ = ~new_new_n55539__ & new_new_n55556__;
  assign new_new_n55774__ = new_new_n55524__ & new_new_n55555__;
  assign new_new_n55775__ = ~new_new_n55539__ & new_new_n55774__;
  assign new_new_n55776__ = ~new_new_n55773__ & ~new_new_n55775__;
  assign new_new_n55777__ = ~new_new_n55524__ & new_new_n55555__;
  assign new_new_n55778__ = new_new_n55539__ & new_new_n55777__;
  assign new_new_n55779__ = new_new_n55524__ & ~new_new_n55555__;
  assign new_new_n55780__ = new_new_n55539__ & new_new_n55779__;
  assign new_new_n55781__ = ~new_new_n55778__ & ~new_new_n55780__;
  assign new_new_n55782__ = new_new_n55776__ & new_new_n55781__;
  assign new_new_n55783__ = ~new_new_n55772__ & ~new_new_n55782__;
  assign new_new_n55784__ = ~new_new_n55732__ & new_new_n55741__;
  assign new_new_n55785__ = new_new_n55717__ & new_new_n55740__;
  assign new_new_n55786__ = ~new_new_n55732__ & new_new_n55785__;
  assign new_new_n55787__ = ~new_new_n55784__ & ~new_new_n55786__;
  assign new_new_n55788__ = ~new_new_n55717__ & new_new_n55740__;
  assign new_new_n55789__ = new_new_n55732__ & new_new_n55788__;
  assign new_new_n55790__ = new_new_n55717__ & ~new_new_n55740__;
  assign new_new_n55791__ = new_new_n55732__ & new_new_n55790__;
  assign new_new_n55792__ = ~new_new_n55789__ & ~new_new_n55791__;
  assign new_new_n55793__ = new_new_n55787__ & new_new_n55792__;
  assign new_new_n55794__ = ys__n39746 & new_new_n52412__;
  assign new_new_n55795__ = ys__n39744 & new_new_n52411__;
  assign new_new_n55796__ = ~new_new_n55794__ & ~new_new_n55795__;
  assign new_new_n55797__ = ys__n33711 & new_new_n52425__;
  assign new_new_n55798__ = ~ys__n33711 & new_new_n52428__;
  assign new_new_n55799__ = ~new_new_n55797__ & ~new_new_n55798__;
  assign new_new_n55800__ = new_new_n55796__ & new_new_n55799__;
  assign new_new_n55801__ = ys__n24789 & new_new_n52417__;
  assign new_new_n55802__ = ys__n24786 & new_new_n52420__;
  assign new_new_n55803__ = ~new_new_n55801__ & ~new_new_n55802__;
  assign new_new_n55804__ = ys__n24783 & new_new_n52419__;
  assign new_new_n55805__ = ys__n39748 & new_new_n52409__;
  assign new_new_n55806__ = ~new_new_n55804__ & ~new_new_n55805__;
  assign new_new_n55807__ = new_new_n55803__ & new_new_n55806__;
  assign new_new_n55808__ = new_new_n55800__ & new_new_n55807__;
  assign new_new_n55809__ = ys__n39752 & new_new_n52301__;
  assign new_new_n55810__ = ys__n39750 & new_new_n52304__;
  assign new_new_n55811__ = ~new_new_n55809__ & ~new_new_n55810__;
  assign new_new_n55812__ = ys__n33717 & new_new_n52308__;
  assign new_new_n55813__ = ~ys__n33717 & new_new_n52311__;
  assign new_new_n55814__ = ~new_new_n55812__ & ~new_new_n55813__;
  assign new_new_n55815__ = new_new_n55811__ & new_new_n55814__;
  assign new_new_n55816__ = ys__n24798 & new_new_n52316__;
  assign new_new_n55817__ = ys__n24795 & new_new_n52318__;
  assign new_new_n55818__ = ~new_new_n55816__ & ~new_new_n55817__;
  assign new_new_n55819__ = ys__n24792 & new_new_n52322__;
  assign new_new_n55820__ = ys__n39754 & new_new_n52324__;
  assign new_new_n55821__ = ~new_new_n55819__ & ~new_new_n55820__;
  assign new_new_n55822__ = new_new_n55818__ & new_new_n55821__;
  assign new_new_n55823__ = new_new_n55815__ & new_new_n55822__;
  assign new_new_n55824__ = ~new_new_n55808__ & ~new_new_n55823__;
  assign new_new_n55825__ = ys__n39740 & new_new_n52449__;
  assign new_new_n55826__ = ys__n39738 & new_new_n52448__;
  assign new_new_n55827__ = ~new_new_n55825__ & ~new_new_n55826__;
  assign new_new_n55828__ = ys__n33705 & new_new_n52462__;
  assign new_new_n55829__ = ~ys__n33705 & new_new_n52465__;
  assign new_new_n55830__ = ~new_new_n55828__ & ~new_new_n55829__;
  assign new_new_n55831__ = new_new_n55827__ & new_new_n55830__;
  assign new_new_n55832__ = ys__n24780 & new_new_n52454__;
  assign new_new_n55833__ = ys__n24777 & new_new_n52457__;
  assign new_new_n55834__ = ~new_new_n55832__ & ~new_new_n55833__;
  assign new_new_n55835__ = ys__n24774 & new_new_n52456__;
  assign new_new_n55836__ = ys__n39742 & new_new_n52446__;
  assign new_new_n55837__ = ~new_new_n55835__ & ~new_new_n55836__;
  assign new_new_n55838__ = new_new_n55834__ & new_new_n55837__;
  assign new_new_n55839__ = new_new_n55831__ & new_new_n55838__;
  assign new_new_n55840__ = ~new_new_n55808__ & ~new_new_n55839__;
  assign new_new_n55841__ = ~new_new_n55823__ & ~new_new_n55839__;
  assign new_new_n55842__ = ~new_new_n55840__ & ~new_new_n55841__;
  assign new_new_n55843__ = ~new_new_n55824__ & new_new_n55842__;
  assign new_new_n55844__ = ~new_new_n55793__ & ~new_new_n55843__;
  assign new_new_n55845__ = ys__n39728 & new_new_n52359__;
  assign new_new_n55846__ = ys__n39726 & new_new_n52358__;
  assign new_new_n55847__ = ~new_new_n55845__ & ~new_new_n55846__;
  assign new_new_n55848__ = ys__n33693 & new_new_n52372__;
  assign new_new_n55849__ = ~ys__n33693 & new_new_n52375__;
  assign new_new_n55850__ = ~new_new_n55848__ & ~new_new_n55849__;
  assign new_new_n55851__ = new_new_n55847__ & new_new_n55850__;
  assign new_new_n55852__ = ys__n24762 & new_new_n52364__;
  assign new_new_n55853__ = ys__n24759 & new_new_n52367__;
  assign new_new_n55854__ = ~new_new_n55852__ & ~new_new_n55853__;
  assign new_new_n55855__ = ys__n24756 & new_new_n52366__;
  assign new_new_n55856__ = ys__n39730 & new_new_n52356__;
  assign new_new_n55857__ = ~new_new_n55855__ & ~new_new_n55856__;
  assign new_new_n55858__ = new_new_n55854__ & new_new_n55857__;
  assign new_new_n55859__ = new_new_n55851__ & new_new_n55858__;
  assign new_new_n55860__ = ys__n39734 & new_new_n52334__;
  assign new_new_n55861__ = ys__n39732 & new_new_n52333__;
  assign new_new_n55862__ = ~new_new_n55860__ & ~new_new_n55861__;
  assign new_new_n55863__ = ys__n33699 & new_new_n52347__;
  assign new_new_n55864__ = ~ys__n33699 & new_new_n52350__;
  assign new_new_n55865__ = ~new_new_n55863__ & ~new_new_n55864__;
  assign new_new_n55866__ = new_new_n55862__ & new_new_n55865__;
  assign new_new_n55867__ = ys__n24771 & new_new_n52339__;
  assign new_new_n55868__ = ys__n24768 & new_new_n52342__;
  assign new_new_n55869__ = ~new_new_n55867__ & ~new_new_n55868__;
  assign new_new_n55870__ = ys__n24765 & new_new_n52341__;
  assign new_new_n55871__ = ys__n39736 & new_new_n52331__;
  assign new_new_n55872__ = ~new_new_n55870__ & ~new_new_n55871__;
  assign new_new_n55873__ = new_new_n55869__ & new_new_n55872__;
  assign new_new_n55874__ = new_new_n55866__ & new_new_n55873__;
  assign new_new_n55875__ = ~new_new_n55859__ & ~new_new_n55874__;
  assign new_new_n55876__ = ys__n24753 & new_new_n52383__;
  assign new_new_n55877__ = ys__n24750 & new_new_n52384__;
  assign new_new_n55878__ = ~new_new_n55876__ & ~new_new_n55877__;
  assign new_new_n55879__ = ys__n39724 & new_new_n52391__;
  assign new_new_n55880__ = ys__n39722 & new_new_n52392__;
  assign new_new_n55881__ = ~new_new_n55879__ & ~new_new_n55880__;
  assign new_new_n55882__ = new_new_n55878__ & new_new_n55881__;
  assign new_new_n55883__ = ~new_new_n55859__ & ~new_new_n55882__;
  assign new_new_n55884__ = ~new_new_n55874__ & ~new_new_n55882__;
  assign new_new_n55885__ = ~new_new_n55883__ & ~new_new_n55884__;
  assign new_new_n55886__ = ~new_new_n55875__ & new_new_n55885__;
  assign new_new_n55887__ = ~new_new_n55793__ & ~new_new_n55886__;
  assign new_new_n55888__ = ~new_new_n55843__ & ~new_new_n55886__;
  assign new_new_n55889__ = ~new_new_n55887__ & ~new_new_n55888__;
  assign new_new_n55890__ = ~new_new_n55844__ & new_new_n55889__;
  assign new_new_n55891__ = ~new_new_n55772__ & ~new_new_n55890__;
  assign new_new_n55892__ = ~new_new_n55782__ & ~new_new_n55890__;
  assign new_new_n55893__ = ~new_new_n55891__ & ~new_new_n55892__;
  assign ys__n43565 = new_new_n55783__ | ~new_new_n55893__;
  assign new_new_n55895__ = ~new_new_n55782__ & new_new_n55891__;
  assign new_new_n55896__ = new_new_n55782__ & ~new_new_n55890__;
  assign new_new_n55897__ = new_new_n55772__ & new_new_n55896__;
  assign new_new_n55898__ = ~new_new_n55782__ & new_new_n55890__;
  assign new_new_n55899__ = new_new_n55772__ & new_new_n55898__;
  assign new_new_n55900__ = new_new_n55782__ & new_new_n55890__;
  assign new_new_n55901__ = ~new_new_n55772__ & new_new_n55900__;
  assign new_new_n55902__ = ~new_new_n55899__ & ~new_new_n55901__;
  assign new_new_n55903__ = ~new_new_n55897__ & new_new_n55902__;
  assign ys__n43570 = new_new_n55895__ | ~new_new_n55903__;
  assign new_new_n55905__ = ~new_new_n55843__ & new_new_n55887__;
  assign new_new_n55906__ = new_new_n55843__ & ~new_new_n55886__;
  assign new_new_n55907__ = new_new_n55793__ & new_new_n55906__;
  assign new_new_n55908__ = ~new_new_n55843__ & new_new_n55886__;
  assign new_new_n55909__ = new_new_n55793__ & new_new_n55908__;
  assign new_new_n55910__ = new_new_n55843__ & new_new_n55886__;
  assign new_new_n55911__ = ~new_new_n55793__ & new_new_n55910__;
  assign new_new_n55912__ = ~new_new_n55909__ & ~new_new_n55911__;
  assign new_new_n55913__ = ~new_new_n55907__ & new_new_n55912__;
  assign new_new_n55914__ = ~new_new_n55905__ & new_new_n55913__;
  assign new_new_n55915__ = ~new_new_n55681__ & new_new_n55698__;
  assign new_new_n55916__ = new_new_n55666__ & new_new_n55697__;
  assign new_new_n55917__ = ~new_new_n55681__ & new_new_n55916__;
  assign new_new_n55918__ = ~new_new_n55915__ & ~new_new_n55917__;
  assign new_new_n55919__ = ~new_new_n55666__ & new_new_n55697__;
  assign new_new_n55920__ = new_new_n55681__ & new_new_n55919__;
  assign new_new_n55921__ = new_new_n55666__ & ~new_new_n55697__;
  assign new_new_n55922__ = new_new_n55681__ & new_new_n55921__;
  assign new_new_n55923__ = ~new_new_n55920__ & ~new_new_n55922__;
  assign new_new_n55924__ = new_new_n55918__ & new_new_n55923__;
  assign new_new_n55925__ = ~new_new_n55914__ & ~new_new_n55924__;
  assign new_new_n55926__ = ~new_new_n55874__ & new_new_n55883__;
  assign new_new_n55927__ = new_new_n55859__ & new_new_n55882__;
  assign new_new_n55928__ = ~new_new_n55874__ & new_new_n55927__;
  assign new_new_n55929__ = ~new_new_n55926__ & ~new_new_n55928__;
  assign new_new_n55930__ = ~new_new_n55859__ & new_new_n55882__;
  assign new_new_n55931__ = new_new_n55874__ & new_new_n55930__;
  assign new_new_n55932__ = new_new_n55859__ & ~new_new_n55882__;
  assign new_new_n55933__ = new_new_n55874__ & new_new_n55932__;
  assign new_new_n55934__ = ~new_new_n55931__ & ~new_new_n55933__;
  assign new_new_n55935__ = new_new_n55929__ & new_new_n55934__;
  assign new_new_n55936__ = ys__n39744 & new_new_n52412__;
  assign new_new_n55937__ = ys__n39742 & new_new_n52411__;
  assign new_new_n55938__ = ~new_new_n55936__ & ~new_new_n55937__;
  assign new_new_n55939__ = ys__n33709 & new_new_n52425__;
  assign new_new_n55940__ = ~ys__n33709 & new_new_n52428__;
  assign new_new_n55941__ = ~new_new_n55939__ & ~new_new_n55940__;
  assign new_new_n55942__ = new_new_n55938__ & new_new_n55941__;
  assign new_new_n55943__ = ys__n24786 & new_new_n52417__;
  assign new_new_n55944__ = ys__n24783 & new_new_n52420__;
  assign new_new_n55945__ = ~new_new_n55943__ & ~new_new_n55944__;
  assign new_new_n55946__ = ys__n24780 & new_new_n52419__;
  assign new_new_n55947__ = ys__n39746 & new_new_n52409__;
  assign new_new_n55948__ = ~new_new_n55946__ & ~new_new_n55947__;
  assign new_new_n55949__ = new_new_n55945__ & new_new_n55948__;
  assign new_new_n55950__ = new_new_n55942__ & new_new_n55949__;
  assign new_new_n55951__ = ys__n39750 & new_new_n52301__;
  assign new_new_n55952__ = ys__n39748 & new_new_n52304__;
  assign new_new_n55953__ = ~new_new_n55951__ & ~new_new_n55952__;
  assign new_new_n55954__ = ys__n33715 & new_new_n52308__;
  assign new_new_n55955__ = ~ys__n33715 & new_new_n52311__;
  assign new_new_n55956__ = ~new_new_n55954__ & ~new_new_n55955__;
  assign new_new_n55957__ = new_new_n55953__ & new_new_n55956__;
  assign new_new_n55958__ = ys__n24795 & new_new_n52316__;
  assign new_new_n55959__ = ys__n24792 & new_new_n52318__;
  assign new_new_n55960__ = ~new_new_n55958__ & ~new_new_n55959__;
  assign new_new_n55961__ = ys__n24789 & new_new_n52322__;
  assign new_new_n55962__ = ys__n39752 & new_new_n52324__;
  assign new_new_n55963__ = ~new_new_n55961__ & ~new_new_n55962__;
  assign new_new_n55964__ = new_new_n55960__ & new_new_n55963__;
  assign new_new_n55965__ = new_new_n55957__ & new_new_n55964__;
  assign new_new_n55966__ = ~new_new_n55950__ & ~new_new_n55965__;
  assign new_new_n55967__ = ys__n39738 & new_new_n52449__;
  assign new_new_n55968__ = ys__n39736 & new_new_n52448__;
  assign new_new_n55969__ = ~new_new_n55967__ & ~new_new_n55968__;
  assign new_new_n55970__ = ys__n33703 & new_new_n52462__;
  assign new_new_n55971__ = ~ys__n33703 & new_new_n52465__;
  assign new_new_n55972__ = ~new_new_n55970__ & ~new_new_n55971__;
  assign new_new_n55973__ = new_new_n55969__ & new_new_n55972__;
  assign new_new_n55974__ = ys__n24777 & new_new_n52454__;
  assign new_new_n55975__ = ys__n24774 & new_new_n52457__;
  assign new_new_n55976__ = ~new_new_n55974__ & ~new_new_n55975__;
  assign new_new_n55977__ = ys__n24771 & new_new_n52456__;
  assign new_new_n55978__ = ys__n39740 & new_new_n52446__;
  assign new_new_n55979__ = ~new_new_n55977__ & ~new_new_n55978__;
  assign new_new_n55980__ = new_new_n55976__ & new_new_n55979__;
  assign new_new_n55981__ = new_new_n55973__ & new_new_n55980__;
  assign new_new_n55982__ = ~new_new_n55950__ & ~new_new_n55981__;
  assign new_new_n55983__ = ~new_new_n55965__ & ~new_new_n55981__;
  assign new_new_n55984__ = ~new_new_n55982__ & ~new_new_n55983__;
  assign new_new_n55985__ = ~new_new_n55966__ & new_new_n55984__;
  assign new_new_n55986__ = ~new_new_n55935__ & ~new_new_n55985__;
  assign new_new_n55987__ = ys__n39726 & new_new_n52359__;
  assign new_new_n55988__ = ys__n39724 & new_new_n52358__;
  assign new_new_n55989__ = ~new_new_n55987__ & ~new_new_n55988__;
  assign new_new_n55990__ = ys__n33691 & new_new_n52372__;
  assign new_new_n55991__ = ~ys__n33691 & new_new_n52375__;
  assign new_new_n55992__ = ~new_new_n55990__ & ~new_new_n55991__;
  assign new_new_n55993__ = new_new_n55989__ & new_new_n55992__;
  assign new_new_n55994__ = ys__n24759 & new_new_n52364__;
  assign new_new_n55995__ = ys__n24756 & new_new_n52367__;
  assign new_new_n55996__ = ~new_new_n55994__ & ~new_new_n55995__;
  assign new_new_n55997__ = ys__n24753 & new_new_n52366__;
  assign new_new_n55998__ = ys__n39728 & new_new_n52356__;
  assign new_new_n55999__ = ~new_new_n55997__ & ~new_new_n55998__;
  assign new_new_n56000__ = new_new_n55996__ & new_new_n55999__;
  assign new_new_n56001__ = new_new_n55993__ & new_new_n56000__;
  assign new_new_n56002__ = ys__n39732 & new_new_n52334__;
  assign new_new_n56003__ = ys__n39730 & new_new_n52333__;
  assign new_new_n56004__ = ~new_new_n56002__ & ~new_new_n56003__;
  assign new_new_n56005__ = ys__n33697 & new_new_n52347__;
  assign new_new_n56006__ = ~ys__n33697 & new_new_n52350__;
  assign new_new_n56007__ = ~new_new_n56005__ & ~new_new_n56006__;
  assign new_new_n56008__ = new_new_n56004__ & new_new_n56007__;
  assign new_new_n56009__ = ys__n24768 & new_new_n52339__;
  assign new_new_n56010__ = ys__n24765 & new_new_n52342__;
  assign new_new_n56011__ = ~new_new_n56009__ & ~new_new_n56010__;
  assign new_new_n56012__ = ys__n24762 & new_new_n52341__;
  assign new_new_n56013__ = ys__n39734 & new_new_n52331__;
  assign new_new_n56014__ = ~new_new_n56012__ & ~new_new_n56013__;
  assign new_new_n56015__ = new_new_n56011__ & new_new_n56014__;
  assign new_new_n56016__ = new_new_n56008__ & new_new_n56015__;
  assign new_new_n56017__ = ~new_new_n56001__ & ~new_new_n56016__;
  assign new_new_n56018__ = ys__n24750 & new_new_n52383__;
  assign new_new_n56019__ = ys__n24747 & new_new_n52384__;
  assign new_new_n56020__ = ~new_new_n56018__ & ~new_new_n56019__;
  assign new_new_n56021__ = ys__n39722 & new_new_n52391__;
  assign new_new_n56022__ = ys__n39720 & new_new_n52392__;
  assign new_new_n56023__ = ~new_new_n56021__ & ~new_new_n56022__;
  assign new_new_n56024__ = new_new_n56020__ & new_new_n56023__;
  assign new_new_n56025__ = ~new_new_n56001__ & ~new_new_n56024__;
  assign new_new_n56026__ = ~new_new_n56016__ & ~new_new_n56024__;
  assign new_new_n56027__ = ~new_new_n56025__ & ~new_new_n56026__;
  assign new_new_n56028__ = ~new_new_n56017__ & new_new_n56027__;
  assign new_new_n56029__ = ~new_new_n55935__ & ~new_new_n56028__;
  assign new_new_n56030__ = ~new_new_n55985__ & ~new_new_n56028__;
  assign new_new_n56031__ = ~new_new_n56029__ & ~new_new_n56030__;
  assign new_new_n56032__ = ~new_new_n55986__ & new_new_n56031__;
  assign new_new_n56033__ = ~new_new_n55914__ & ~new_new_n56032__;
  assign new_new_n56034__ = ~new_new_n55924__ & ~new_new_n56032__;
  assign new_new_n56035__ = ~new_new_n56033__ & ~new_new_n56034__;
  assign ys__n43619 = new_new_n55925__ | ~new_new_n56035__;
  assign new_new_n56037__ = ~new_new_n55924__ & new_new_n56033__;
  assign new_new_n56038__ = new_new_n55924__ & ~new_new_n56032__;
  assign new_new_n56039__ = new_new_n55914__ & new_new_n56038__;
  assign new_new_n56040__ = ~new_new_n55924__ & new_new_n56032__;
  assign new_new_n56041__ = new_new_n55914__ & new_new_n56040__;
  assign new_new_n56042__ = new_new_n55924__ & new_new_n56032__;
  assign new_new_n56043__ = ~new_new_n55914__ & new_new_n56042__;
  assign new_new_n56044__ = ~new_new_n56041__ & ~new_new_n56043__;
  assign new_new_n56045__ = ~new_new_n56039__ & new_new_n56044__;
  assign ys__n43624 = new_new_n56037__ | ~new_new_n56045__;
  assign new_new_n56047__ = ~new_new_n55985__ & new_new_n56029__;
  assign new_new_n56048__ = new_new_n55985__ & ~new_new_n56028__;
  assign new_new_n56049__ = new_new_n55935__ & new_new_n56048__;
  assign new_new_n56050__ = ~new_new_n55985__ & new_new_n56028__;
  assign new_new_n56051__ = new_new_n55935__ & new_new_n56050__;
  assign new_new_n56052__ = new_new_n55985__ & new_new_n56028__;
  assign new_new_n56053__ = ~new_new_n55935__ & new_new_n56052__;
  assign new_new_n56054__ = ~new_new_n56051__ & ~new_new_n56053__;
  assign new_new_n56055__ = ~new_new_n56049__ & new_new_n56054__;
  assign new_new_n56056__ = ~new_new_n56047__ & new_new_n56055__;
  assign new_new_n56057__ = ~new_new_n55823__ & new_new_n55840__;
  assign new_new_n56058__ = new_new_n55808__ & new_new_n55839__;
  assign new_new_n56059__ = ~new_new_n55823__ & new_new_n56058__;
  assign new_new_n56060__ = ~new_new_n56057__ & ~new_new_n56059__;
  assign new_new_n56061__ = ~new_new_n55808__ & new_new_n55839__;
  assign new_new_n56062__ = new_new_n55823__ & new_new_n56061__;
  assign new_new_n56063__ = new_new_n55808__ & ~new_new_n55839__;
  assign new_new_n56064__ = new_new_n55823__ & new_new_n56063__;
  assign new_new_n56065__ = ~new_new_n56062__ & ~new_new_n56064__;
  assign new_new_n56066__ = new_new_n56060__ & new_new_n56065__;
  assign new_new_n56067__ = ~new_new_n56056__ & ~new_new_n56066__;
  assign new_new_n56068__ = ~new_new_n56016__ & new_new_n56025__;
  assign new_new_n56069__ = new_new_n56001__ & new_new_n56024__;
  assign new_new_n56070__ = ~new_new_n56016__ & new_new_n56069__;
  assign new_new_n56071__ = ~new_new_n56068__ & ~new_new_n56070__;
  assign new_new_n56072__ = ~new_new_n56001__ & new_new_n56024__;
  assign new_new_n56073__ = new_new_n56016__ & new_new_n56072__;
  assign new_new_n56074__ = new_new_n56001__ & ~new_new_n56024__;
  assign new_new_n56075__ = new_new_n56016__ & new_new_n56074__;
  assign new_new_n56076__ = ~new_new_n56073__ & ~new_new_n56075__;
  assign new_new_n56077__ = new_new_n56071__ & new_new_n56076__;
  assign new_new_n56078__ = ys__n39742 & new_new_n52412__;
  assign new_new_n56079__ = ys__n39740 & new_new_n52411__;
  assign new_new_n56080__ = ~new_new_n56078__ & ~new_new_n56079__;
  assign new_new_n56081__ = ys__n33707 & new_new_n52425__;
  assign new_new_n56082__ = ~ys__n33707 & new_new_n52428__;
  assign new_new_n56083__ = ~new_new_n56081__ & ~new_new_n56082__;
  assign new_new_n56084__ = new_new_n56080__ & new_new_n56083__;
  assign new_new_n56085__ = ys__n24783 & new_new_n52417__;
  assign new_new_n56086__ = ys__n24780 & new_new_n52420__;
  assign new_new_n56087__ = ~new_new_n56085__ & ~new_new_n56086__;
  assign new_new_n56088__ = ys__n24777 & new_new_n52419__;
  assign new_new_n56089__ = ys__n39744 & new_new_n52409__;
  assign new_new_n56090__ = ~new_new_n56088__ & ~new_new_n56089__;
  assign new_new_n56091__ = new_new_n56087__ & new_new_n56090__;
  assign new_new_n56092__ = new_new_n56084__ & new_new_n56091__;
  assign new_new_n56093__ = ys__n39748 & new_new_n52301__;
  assign new_new_n56094__ = ys__n39746 & new_new_n52304__;
  assign new_new_n56095__ = ~new_new_n56093__ & ~new_new_n56094__;
  assign new_new_n56096__ = ys__n33713 & new_new_n52308__;
  assign new_new_n56097__ = ~ys__n33713 & new_new_n52311__;
  assign new_new_n56098__ = ~new_new_n56096__ & ~new_new_n56097__;
  assign new_new_n56099__ = new_new_n56095__ & new_new_n56098__;
  assign new_new_n56100__ = ys__n24792 & new_new_n52316__;
  assign new_new_n56101__ = ys__n24789 & new_new_n52318__;
  assign new_new_n56102__ = ~new_new_n56100__ & ~new_new_n56101__;
  assign new_new_n56103__ = ys__n24786 & new_new_n52322__;
  assign new_new_n56104__ = ys__n39750 & new_new_n52324__;
  assign new_new_n56105__ = ~new_new_n56103__ & ~new_new_n56104__;
  assign new_new_n56106__ = new_new_n56102__ & new_new_n56105__;
  assign new_new_n56107__ = new_new_n56099__ & new_new_n56106__;
  assign new_new_n56108__ = ~new_new_n56092__ & ~new_new_n56107__;
  assign new_new_n56109__ = ys__n39736 & new_new_n52449__;
  assign new_new_n56110__ = ys__n39734 & new_new_n52448__;
  assign new_new_n56111__ = ~new_new_n56109__ & ~new_new_n56110__;
  assign new_new_n56112__ = ys__n33701 & new_new_n52462__;
  assign new_new_n56113__ = ~ys__n33701 & new_new_n52465__;
  assign new_new_n56114__ = ~new_new_n56112__ & ~new_new_n56113__;
  assign new_new_n56115__ = new_new_n56111__ & new_new_n56114__;
  assign new_new_n56116__ = ys__n24774 & new_new_n52454__;
  assign new_new_n56117__ = ys__n24771 & new_new_n52457__;
  assign new_new_n56118__ = ~new_new_n56116__ & ~new_new_n56117__;
  assign new_new_n56119__ = ys__n24768 & new_new_n52456__;
  assign new_new_n56120__ = ys__n39738 & new_new_n52446__;
  assign new_new_n56121__ = ~new_new_n56119__ & ~new_new_n56120__;
  assign new_new_n56122__ = new_new_n56118__ & new_new_n56121__;
  assign new_new_n56123__ = new_new_n56115__ & new_new_n56122__;
  assign new_new_n56124__ = ~new_new_n56092__ & ~new_new_n56123__;
  assign new_new_n56125__ = ~new_new_n56107__ & ~new_new_n56123__;
  assign new_new_n56126__ = ~new_new_n56124__ & ~new_new_n56125__;
  assign new_new_n56127__ = ~new_new_n56108__ & new_new_n56126__;
  assign new_new_n56128__ = ~new_new_n56077__ & ~new_new_n56127__;
  assign new_new_n56129__ = ys__n39724 & new_new_n52359__;
  assign new_new_n56130__ = ys__n39722 & new_new_n52358__;
  assign new_new_n56131__ = ~new_new_n56129__ & ~new_new_n56130__;
  assign new_new_n56132__ = ys__n33689 & new_new_n52372__;
  assign new_new_n56133__ = ~ys__n33689 & new_new_n52375__;
  assign new_new_n56134__ = ~new_new_n56132__ & ~new_new_n56133__;
  assign new_new_n56135__ = new_new_n56131__ & new_new_n56134__;
  assign new_new_n56136__ = ys__n24756 & new_new_n52364__;
  assign new_new_n56137__ = ys__n24753 & new_new_n52367__;
  assign new_new_n56138__ = ~new_new_n56136__ & ~new_new_n56137__;
  assign new_new_n56139__ = ys__n24750 & new_new_n52366__;
  assign new_new_n56140__ = ys__n39726 & new_new_n52356__;
  assign new_new_n56141__ = ~new_new_n56139__ & ~new_new_n56140__;
  assign new_new_n56142__ = new_new_n56138__ & new_new_n56141__;
  assign new_new_n56143__ = new_new_n56135__ & new_new_n56142__;
  assign new_new_n56144__ = ys__n39730 & new_new_n52334__;
  assign new_new_n56145__ = ys__n39728 & new_new_n52333__;
  assign new_new_n56146__ = ~new_new_n56144__ & ~new_new_n56145__;
  assign new_new_n56147__ = ys__n33695 & new_new_n52347__;
  assign new_new_n56148__ = ~ys__n33695 & new_new_n52350__;
  assign new_new_n56149__ = ~new_new_n56147__ & ~new_new_n56148__;
  assign new_new_n56150__ = new_new_n56146__ & new_new_n56149__;
  assign new_new_n56151__ = ys__n24765 & new_new_n52339__;
  assign new_new_n56152__ = ys__n24762 & new_new_n52342__;
  assign new_new_n56153__ = ~new_new_n56151__ & ~new_new_n56152__;
  assign new_new_n56154__ = ys__n24759 & new_new_n52341__;
  assign new_new_n56155__ = ys__n39732 & new_new_n52331__;
  assign new_new_n56156__ = ~new_new_n56154__ & ~new_new_n56155__;
  assign new_new_n56157__ = new_new_n56153__ & new_new_n56156__;
  assign new_new_n56158__ = new_new_n56150__ & new_new_n56157__;
  assign new_new_n56159__ = ~new_new_n56143__ & ~new_new_n56158__;
  assign new_new_n56160__ = ys__n24747 & new_new_n52383__;
  assign new_new_n56161__ = ys__n24744 & new_new_n52384__;
  assign new_new_n56162__ = ~new_new_n56160__ & ~new_new_n56161__;
  assign new_new_n56163__ = ys__n39720 & new_new_n52391__;
  assign new_new_n56164__ = ys__n39718 & new_new_n52392__;
  assign new_new_n56165__ = ~new_new_n56163__ & ~new_new_n56164__;
  assign new_new_n56166__ = new_new_n56162__ & new_new_n56165__;
  assign new_new_n56167__ = ~new_new_n56143__ & ~new_new_n56166__;
  assign new_new_n56168__ = ~new_new_n56158__ & ~new_new_n56166__;
  assign new_new_n56169__ = ~new_new_n56167__ & ~new_new_n56168__;
  assign new_new_n56170__ = ~new_new_n56159__ & new_new_n56169__;
  assign new_new_n56171__ = ~new_new_n56077__ & ~new_new_n56170__;
  assign new_new_n56172__ = ~new_new_n56127__ & ~new_new_n56170__;
  assign new_new_n56173__ = ~new_new_n56171__ & ~new_new_n56172__;
  assign new_new_n56174__ = ~new_new_n56128__ & new_new_n56173__;
  assign new_new_n56175__ = ~new_new_n56056__ & ~new_new_n56174__;
  assign new_new_n56176__ = ~new_new_n56066__ & ~new_new_n56174__;
  assign new_new_n56177__ = ~new_new_n56175__ & ~new_new_n56176__;
  assign ys__n43673 = new_new_n56067__ | ~new_new_n56177__;
  assign new_new_n56179__ = ~new_new_n56066__ & new_new_n56175__;
  assign new_new_n56180__ = new_new_n56066__ & ~new_new_n56174__;
  assign new_new_n56181__ = new_new_n56056__ & new_new_n56180__;
  assign new_new_n56182__ = ~new_new_n56066__ & new_new_n56174__;
  assign new_new_n56183__ = new_new_n56056__ & new_new_n56182__;
  assign new_new_n56184__ = new_new_n56066__ & new_new_n56174__;
  assign new_new_n56185__ = ~new_new_n56056__ & new_new_n56184__;
  assign new_new_n56186__ = ~new_new_n56183__ & ~new_new_n56185__;
  assign new_new_n56187__ = ~new_new_n56181__ & new_new_n56186__;
  assign ys__n43678 = new_new_n56179__ | ~new_new_n56187__;
  assign new_new_n56189__ = ~new_new_n56127__ & new_new_n56171__;
  assign new_new_n56190__ = new_new_n56127__ & ~new_new_n56170__;
  assign new_new_n56191__ = new_new_n56077__ & new_new_n56190__;
  assign new_new_n56192__ = ~new_new_n56127__ & new_new_n56170__;
  assign new_new_n56193__ = new_new_n56077__ & new_new_n56192__;
  assign new_new_n56194__ = new_new_n56127__ & new_new_n56170__;
  assign new_new_n56195__ = ~new_new_n56077__ & new_new_n56194__;
  assign new_new_n56196__ = ~new_new_n56193__ & ~new_new_n56195__;
  assign new_new_n56197__ = ~new_new_n56191__ & new_new_n56196__;
  assign new_new_n56198__ = ~new_new_n56189__ & new_new_n56197__;
  assign new_new_n56199__ = ~new_new_n55965__ & new_new_n55982__;
  assign new_new_n56200__ = new_new_n55950__ & new_new_n55981__;
  assign new_new_n56201__ = ~new_new_n55965__ & new_new_n56200__;
  assign new_new_n56202__ = ~new_new_n56199__ & ~new_new_n56201__;
  assign new_new_n56203__ = ~new_new_n55950__ & new_new_n55981__;
  assign new_new_n56204__ = new_new_n55965__ & new_new_n56203__;
  assign new_new_n56205__ = new_new_n55950__ & ~new_new_n55981__;
  assign new_new_n56206__ = new_new_n55965__ & new_new_n56205__;
  assign new_new_n56207__ = ~new_new_n56204__ & ~new_new_n56206__;
  assign new_new_n56208__ = new_new_n56202__ & new_new_n56207__;
  assign new_new_n56209__ = ~new_new_n56198__ & ~new_new_n56208__;
  assign new_new_n56210__ = ~new_new_n56158__ & new_new_n56167__;
  assign new_new_n56211__ = new_new_n56143__ & new_new_n56166__;
  assign new_new_n56212__ = ~new_new_n56158__ & new_new_n56211__;
  assign new_new_n56213__ = ~new_new_n56210__ & ~new_new_n56212__;
  assign new_new_n56214__ = ~new_new_n56143__ & new_new_n56166__;
  assign new_new_n56215__ = new_new_n56158__ & new_new_n56214__;
  assign new_new_n56216__ = new_new_n56143__ & ~new_new_n56166__;
  assign new_new_n56217__ = new_new_n56158__ & new_new_n56216__;
  assign new_new_n56218__ = ~new_new_n56215__ & ~new_new_n56217__;
  assign new_new_n56219__ = new_new_n56213__ & new_new_n56218__;
  assign new_new_n56220__ = ys__n39740 & new_new_n52412__;
  assign new_new_n56221__ = ys__n39738 & new_new_n52411__;
  assign new_new_n56222__ = ~new_new_n56220__ & ~new_new_n56221__;
  assign new_new_n56223__ = ys__n33705 & new_new_n52425__;
  assign new_new_n56224__ = ~ys__n33705 & new_new_n52428__;
  assign new_new_n56225__ = ~new_new_n56223__ & ~new_new_n56224__;
  assign new_new_n56226__ = new_new_n56222__ & new_new_n56225__;
  assign new_new_n56227__ = ys__n24780 & new_new_n52417__;
  assign new_new_n56228__ = ys__n24777 & new_new_n52420__;
  assign new_new_n56229__ = ~new_new_n56227__ & ~new_new_n56228__;
  assign new_new_n56230__ = ys__n24774 & new_new_n52419__;
  assign new_new_n56231__ = ys__n39742 & new_new_n52409__;
  assign new_new_n56232__ = ~new_new_n56230__ & ~new_new_n56231__;
  assign new_new_n56233__ = new_new_n56229__ & new_new_n56232__;
  assign new_new_n56234__ = new_new_n56226__ & new_new_n56233__;
  assign new_new_n56235__ = ys__n39746 & new_new_n52301__;
  assign new_new_n56236__ = ys__n39744 & new_new_n52304__;
  assign new_new_n56237__ = ~new_new_n56235__ & ~new_new_n56236__;
  assign new_new_n56238__ = ys__n33711 & new_new_n52308__;
  assign new_new_n56239__ = ~ys__n33711 & new_new_n52311__;
  assign new_new_n56240__ = ~new_new_n56238__ & ~new_new_n56239__;
  assign new_new_n56241__ = new_new_n56237__ & new_new_n56240__;
  assign new_new_n56242__ = ys__n24789 & new_new_n52316__;
  assign new_new_n56243__ = ys__n24786 & new_new_n52318__;
  assign new_new_n56244__ = ~new_new_n56242__ & ~new_new_n56243__;
  assign new_new_n56245__ = ys__n24783 & new_new_n52322__;
  assign new_new_n56246__ = ys__n39748 & new_new_n52324__;
  assign new_new_n56247__ = ~new_new_n56245__ & ~new_new_n56246__;
  assign new_new_n56248__ = new_new_n56244__ & new_new_n56247__;
  assign new_new_n56249__ = new_new_n56241__ & new_new_n56248__;
  assign new_new_n56250__ = ~new_new_n56234__ & ~new_new_n56249__;
  assign new_new_n56251__ = ys__n39734 & new_new_n52449__;
  assign new_new_n56252__ = ys__n39732 & new_new_n52448__;
  assign new_new_n56253__ = ~new_new_n56251__ & ~new_new_n56252__;
  assign new_new_n56254__ = ys__n33699 & new_new_n52462__;
  assign new_new_n56255__ = ~ys__n33699 & new_new_n52465__;
  assign new_new_n56256__ = ~new_new_n56254__ & ~new_new_n56255__;
  assign new_new_n56257__ = new_new_n56253__ & new_new_n56256__;
  assign new_new_n56258__ = ys__n24771 & new_new_n52454__;
  assign new_new_n56259__ = ys__n24768 & new_new_n52457__;
  assign new_new_n56260__ = ~new_new_n56258__ & ~new_new_n56259__;
  assign new_new_n56261__ = ys__n24765 & new_new_n52456__;
  assign new_new_n56262__ = ys__n39736 & new_new_n52446__;
  assign new_new_n56263__ = ~new_new_n56261__ & ~new_new_n56262__;
  assign new_new_n56264__ = new_new_n56260__ & new_new_n56263__;
  assign new_new_n56265__ = new_new_n56257__ & new_new_n56264__;
  assign new_new_n56266__ = ~new_new_n56234__ & ~new_new_n56265__;
  assign new_new_n56267__ = ~new_new_n56249__ & ~new_new_n56265__;
  assign new_new_n56268__ = ~new_new_n56266__ & ~new_new_n56267__;
  assign new_new_n56269__ = ~new_new_n56250__ & new_new_n56268__;
  assign new_new_n56270__ = ~new_new_n56219__ & ~new_new_n56269__;
  assign new_new_n56271__ = ys__n39722 & new_new_n52359__;
  assign new_new_n56272__ = ys__n39720 & new_new_n52358__;
  assign new_new_n56273__ = ~new_new_n56271__ & ~new_new_n56272__;
  assign new_new_n56274__ = ys__n33687 & new_new_n52372__;
  assign new_new_n56275__ = ~ys__n33687 & new_new_n52375__;
  assign new_new_n56276__ = ~new_new_n56274__ & ~new_new_n56275__;
  assign new_new_n56277__ = new_new_n56273__ & new_new_n56276__;
  assign new_new_n56278__ = ys__n24753 & new_new_n52364__;
  assign new_new_n56279__ = ys__n24750 & new_new_n52367__;
  assign new_new_n56280__ = ~new_new_n56278__ & ~new_new_n56279__;
  assign new_new_n56281__ = ys__n24747 & new_new_n52366__;
  assign new_new_n56282__ = ys__n39724 & new_new_n52356__;
  assign new_new_n56283__ = ~new_new_n56281__ & ~new_new_n56282__;
  assign new_new_n56284__ = new_new_n56280__ & new_new_n56283__;
  assign new_new_n56285__ = new_new_n56277__ & new_new_n56284__;
  assign new_new_n56286__ = ys__n39728 & new_new_n52334__;
  assign new_new_n56287__ = ys__n39726 & new_new_n52333__;
  assign new_new_n56288__ = ~new_new_n56286__ & ~new_new_n56287__;
  assign new_new_n56289__ = ys__n33693 & new_new_n52347__;
  assign new_new_n56290__ = ~ys__n33693 & new_new_n52350__;
  assign new_new_n56291__ = ~new_new_n56289__ & ~new_new_n56290__;
  assign new_new_n56292__ = new_new_n56288__ & new_new_n56291__;
  assign new_new_n56293__ = ys__n24762 & new_new_n52339__;
  assign new_new_n56294__ = ys__n24759 & new_new_n52342__;
  assign new_new_n56295__ = ~new_new_n56293__ & ~new_new_n56294__;
  assign new_new_n56296__ = ys__n24756 & new_new_n52341__;
  assign new_new_n56297__ = ys__n39730 & new_new_n52331__;
  assign new_new_n56298__ = ~new_new_n56296__ & ~new_new_n56297__;
  assign new_new_n56299__ = new_new_n56295__ & new_new_n56298__;
  assign new_new_n56300__ = new_new_n56292__ & new_new_n56299__;
  assign new_new_n56301__ = ~new_new_n56285__ & ~new_new_n56300__;
  assign new_new_n56302__ = ys__n24744 & new_new_n52383__;
  assign new_new_n56303__ = ys__n24741 & new_new_n52384__;
  assign new_new_n56304__ = ~new_new_n56302__ & ~new_new_n56303__;
  assign new_new_n56305__ = ys__n39718 & new_new_n52391__;
  assign new_new_n56306__ = ys__n24741 & new_new_n52392__;
  assign new_new_n56307__ = ~new_new_n56305__ & ~new_new_n56306__;
  assign new_new_n56308__ = new_new_n56304__ & new_new_n56307__;
  assign new_new_n56309__ = ~new_new_n56285__ & ~new_new_n56308__;
  assign new_new_n56310__ = ~new_new_n56300__ & ~new_new_n56308__;
  assign new_new_n56311__ = ~new_new_n56309__ & ~new_new_n56310__;
  assign new_new_n56312__ = ~new_new_n56301__ & new_new_n56311__;
  assign new_new_n56313__ = ~new_new_n56219__ & ~new_new_n56312__;
  assign new_new_n56314__ = ~new_new_n56269__ & ~new_new_n56312__;
  assign new_new_n56315__ = ~new_new_n56313__ & ~new_new_n56314__;
  assign new_new_n56316__ = ~new_new_n56270__ & new_new_n56315__;
  assign new_new_n56317__ = ~new_new_n56198__ & ~new_new_n56316__;
  assign new_new_n56318__ = ~new_new_n56208__ & ~new_new_n56316__;
  assign new_new_n56319__ = ~new_new_n56317__ & ~new_new_n56318__;
  assign ys__n43727 = new_new_n56209__ | ~new_new_n56319__;
  assign new_new_n56321__ = ~new_new_n56208__ & new_new_n56317__;
  assign new_new_n56322__ = new_new_n56208__ & ~new_new_n56316__;
  assign new_new_n56323__ = new_new_n56198__ & new_new_n56322__;
  assign new_new_n56324__ = ~new_new_n56208__ & new_new_n56316__;
  assign new_new_n56325__ = new_new_n56198__ & new_new_n56324__;
  assign new_new_n56326__ = new_new_n56208__ & new_new_n56316__;
  assign new_new_n56327__ = ~new_new_n56198__ & new_new_n56326__;
  assign new_new_n56328__ = ~new_new_n56325__ & ~new_new_n56327__;
  assign new_new_n56329__ = ~new_new_n56323__ & new_new_n56328__;
  assign ys__n43732 = new_new_n56321__ | ~new_new_n56329__;
  assign new_new_n56331__ = ~new_new_n56269__ & new_new_n56313__;
  assign new_new_n56332__ = new_new_n56269__ & ~new_new_n56312__;
  assign new_new_n56333__ = new_new_n56219__ & new_new_n56332__;
  assign new_new_n56334__ = ~new_new_n56269__ & new_new_n56312__;
  assign new_new_n56335__ = new_new_n56219__ & new_new_n56334__;
  assign new_new_n56336__ = new_new_n56269__ & new_new_n56312__;
  assign new_new_n56337__ = ~new_new_n56219__ & new_new_n56336__;
  assign new_new_n56338__ = ~new_new_n56335__ & ~new_new_n56337__;
  assign new_new_n56339__ = ~new_new_n56333__ & new_new_n56338__;
  assign new_new_n56340__ = ~new_new_n56331__ & new_new_n56339__;
  assign new_new_n56341__ = ~new_new_n56107__ & new_new_n56124__;
  assign new_new_n56342__ = new_new_n56092__ & new_new_n56123__;
  assign new_new_n56343__ = ~new_new_n56107__ & new_new_n56342__;
  assign new_new_n56344__ = ~new_new_n56341__ & ~new_new_n56343__;
  assign new_new_n56345__ = ~new_new_n56092__ & new_new_n56123__;
  assign new_new_n56346__ = new_new_n56107__ & new_new_n56345__;
  assign new_new_n56347__ = new_new_n56092__ & ~new_new_n56123__;
  assign new_new_n56348__ = new_new_n56107__ & new_new_n56347__;
  assign new_new_n56349__ = ~new_new_n56346__ & ~new_new_n56348__;
  assign new_new_n56350__ = new_new_n56344__ & new_new_n56349__;
  assign new_new_n56351__ = ~new_new_n56340__ & ~new_new_n56350__;
  assign new_new_n56352__ = ~new_new_n56300__ & new_new_n56309__;
  assign new_new_n56353__ = new_new_n56285__ & new_new_n56308__;
  assign new_new_n56354__ = ~new_new_n56300__ & new_new_n56353__;
  assign new_new_n56355__ = ~new_new_n56352__ & ~new_new_n56354__;
  assign new_new_n56356__ = ~new_new_n56285__ & new_new_n56308__;
  assign new_new_n56357__ = new_new_n56300__ & new_new_n56356__;
  assign new_new_n56358__ = new_new_n56285__ & ~new_new_n56308__;
  assign new_new_n56359__ = new_new_n56300__ & new_new_n56358__;
  assign new_new_n56360__ = ~new_new_n56357__ & ~new_new_n56359__;
  assign new_new_n56361__ = new_new_n56355__ & new_new_n56360__;
  assign new_new_n56362__ = ys__n39738 & new_new_n52412__;
  assign new_new_n56363__ = ys__n39736 & new_new_n52411__;
  assign new_new_n56364__ = ~new_new_n56362__ & ~new_new_n56363__;
  assign new_new_n56365__ = ys__n33703 & new_new_n52425__;
  assign new_new_n56366__ = ~ys__n33703 & new_new_n52428__;
  assign new_new_n56367__ = ~new_new_n56365__ & ~new_new_n56366__;
  assign new_new_n56368__ = new_new_n56364__ & new_new_n56367__;
  assign new_new_n56369__ = ys__n24777 & new_new_n52417__;
  assign new_new_n56370__ = ys__n24774 & new_new_n52420__;
  assign new_new_n56371__ = ~new_new_n56369__ & ~new_new_n56370__;
  assign new_new_n56372__ = ys__n24771 & new_new_n52419__;
  assign new_new_n56373__ = ys__n39740 & new_new_n52409__;
  assign new_new_n56374__ = ~new_new_n56372__ & ~new_new_n56373__;
  assign new_new_n56375__ = new_new_n56371__ & new_new_n56374__;
  assign new_new_n56376__ = new_new_n56368__ & new_new_n56375__;
  assign new_new_n56377__ = ys__n39744 & new_new_n52301__;
  assign new_new_n56378__ = ys__n39742 & new_new_n52304__;
  assign new_new_n56379__ = ~new_new_n56377__ & ~new_new_n56378__;
  assign new_new_n56380__ = ys__n33709 & new_new_n52308__;
  assign new_new_n56381__ = ~ys__n33709 & new_new_n52311__;
  assign new_new_n56382__ = ~new_new_n56380__ & ~new_new_n56381__;
  assign new_new_n56383__ = new_new_n56379__ & new_new_n56382__;
  assign new_new_n56384__ = ys__n24786 & new_new_n52316__;
  assign new_new_n56385__ = ys__n24783 & new_new_n52318__;
  assign new_new_n56386__ = ~new_new_n56384__ & ~new_new_n56385__;
  assign new_new_n56387__ = ys__n24780 & new_new_n52322__;
  assign new_new_n56388__ = ys__n39746 & new_new_n52324__;
  assign new_new_n56389__ = ~new_new_n56387__ & ~new_new_n56388__;
  assign new_new_n56390__ = new_new_n56386__ & new_new_n56389__;
  assign new_new_n56391__ = new_new_n56383__ & new_new_n56390__;
  assign new_new_n56392__ = ~new_new_n56376__ & ~new_new_n56391__;
  assign new_new_n56393__ = ys__n39732 & new_new_n52449__;
  assign new_new_n56394__ = ys__n39730 & new_new_n52448__;
  assign new_new_n56395__ = ~new_new_n56393__ & ~new_new_n56394__;
  assign new_new_n56396__ = ys__n33697 & new_new_n52462__;
  assign new_new_n56397__ = ~ys__n33697 & new_new_n52465__;
  assign new_new_n56398__ = ~new_new_n56396__ & ~new_new_n56397__;
  assign new_new_n56399__ = new_new_n56395__ & new_new_n56398__;
  assign new_new_n56400__ = ys__n24768 & new_new_n52454__;
  assign new_new_n56401__ = ys__n24765 & new_new_n52457__;
  assign new_new_n56402__ = ~new_new_n56400__ & ~new_new_n56401__;
  assign new_new_n56403__ = ys__n24762 & new_new_n52456__;
  assign new_new_n56404__ = ys__n39734 & new_new_n52446__;
  assign new_new_n56405__ = ~new_new_n56403__ & ~new_new_n56404__;
  assign new_new_n56406__ = new_new_n56402__ & new_new_n56405__;
  assign new_new_n56407__ = new_new_n56399__ & new_new_n56406__;
  assign new_new_n56408__ = ~new_new_n56376__ & ~new_new_n56407__;
  assign new_new_n56409__ = ~new_new_n56391__ & ~new_new_n56407__;
  assign new_new_n56410__ = ~new_new_n56408__ & ~new_new_n56409__;
  assign new_new_n56411__ = ~new_new_n56392__ & new_new_n56410__;
  assign new_new_n56412__ = ~new_new_n56361__ & ~new_new_n56411__;
  assign new_new_n56413__ = ys__n39720 & new_new_n52359__;
  assign new_new_n56414__ = ys__n39718 & new_new_n52358__;
  assign new_new_n56415__ = ~new_new_n56413__ & ~new_new_n56414__;
  assign new_new_n56416__ = ys__n33685 & new_new_n52372__;
  assign new_new_n56417__ = ~ys__n33685 & new_new_n52375__;
  assign new_new_n56418__ = ~new_new_n56416__ & ~new_new_n56417__;
  assign new_new_n56419__ = new_new_n56415__ & new_new_n56418__;
  assign new_new_n56420__ = ys__n24750 & new_new_n52364__;
  assign new_new_n56421__ = ys__n24747 & new_new_n52367__;
  assign new_new_n56422__ = ~new_new_n56420__ & ~new_new_n56421__;
  assign new_new_n56423__ = ys__n24744 & new_new_n52366__;
  assign new_new_n56424__ = ys__n39722 & new_new_n52356__;
  assign new_new_n56425__ = ~new_new_n56423__ & ~new_new_n56424__;
  assign new_new_n56426__ = new_new_n56422__ & new_new_n56425__;
  assign new_new_n56427__ = new_new_n56419__ & new_new_n56426__;
  assign new_new_n56428__ = ys__n39726 & new_new_n52334__;
  assign new_new_n56429__ = ys__n39724 & new_new_n52333__;
  assign new_new_n56430__ = ~new_new_n56428__ & ~new_new_n56429__;
  assign new_new_n56431__ = ys__n33691 & new_new_n52347__;
  assign new_new_n56432__ = ~ys__n33691 & new_new_n52350__;
  assign new_new_n56433__ = ~new_new_n56431__ & ~new_new_n56432__;
  assign new_new_n56434__ = new_new_n56430__ & new_new_n56433__;
  assign new_new_n56435__ = ys__n24759 & new_new_n52339__;
  assign new_new_n56436__ = ys__n24756 & new_new_n52342__;
  assign new_new_n56437__ = ~new_new_n56435__ & ~new_new_n56436__;
  assign new_new_n56438__ = ys__n24753 & new_new_n52341__;
  assign new_new_n56439__ = ys__n39728 & new_new_n52331__;
  assign new_new_n56440__ = ~new_new_n56438__ & ~new_new_n56439__;
  assign new_new_n56441__ = new_new_n56437__ & new_new_n56440__;
  assign new_new_n56442__ = new_new_n56434__ & new_new_n56441__;
  assign new_new_n56443__ = ~new_new_n56427__ & ~new_new_n56442__;
  assign new_new_n56444__ = ys__n24741 & new_new_n52383__;
  assign new_new_n56445__ = ys__n24741 & new_new_n52391__;
  assign new_new_n56446__ = ~new_new_n56444__ & ~new_new_n56445__;
  assign new_new_n56447__ = ~new_new_n56427__ & ~new_new_n56446__;
  assign new_new_n56448__ = ~new_new_n56442__ & ~new_new_n56446__;
  assign new_new_n56449__ = ~new_new_n56447__ & ~new_new_n56448__;
  assign new_new_n56450__ = ~new_new_n56443__ & new_new_n56449__;
  assign new_new_n56451__ = ~new_new_n56361__ & ~new_new_n56450__;
  assign new_new_n56452__ = ~new_new_n56411__ & ~new_new_n56450__;
  assign new_new_n56453__ = ~new_new_n56451__ & ~new_new_n56452__;
  assign new_new_n56454__ = ~new_new_n56412__ & new_new_n56453__;
  assign new_new_n56455__ = ~new_new_n56340__ & ~new_new_n56454__;
  assign new_new_n56456__ = ~new_new_n56350__ & ~new_new_n56454__;
  assign new_new_n56457__ = ~new_new_n56455__ & ~new_new_n56456__;
  assign ys__n43781 = new_new_n56351__ | ~new_new_n56457__;
  assign new_new_n56459__ = ~new_new_n56350__ & new_new_n56455__;
  assign new_new_n56460__ = new_new_n56350__ & ~new_new_n56454__;
  assign new_new_n56461__ = new_new_n56340__ & new_new_n56460__;
  assign new_new_n56462__ = ~new_new_n56350__ & new_new_n56454__;
  assign new_new_n56463__ = new_new_n56340__ & new_new_n56462__;
  assign new_new_n56464__ = new_new_n56350__ & new_new_n56454__;
  assign new_new_n56465__ = ~new_new_n56340__ & new_new_n56464__;
  assign new_new_n56466__ = ~new_new_n56463__ & ~new_new_n56465__;
  assign new_new_n56467__ = ~new_new_n56461__ & new_new_n56466__;
  assign ys__n43786 = new_new_n56459__ | ~new_new_n56467__;
  assign new_new_n56469__ = ~new_new_n56411__ & new_new_n56451__;
  assign new_new_n56470__ = new_new_n56411__ & ~new_new_n56450__;
  assign new_new_n56471__ = new_new_n56361__ & new_new_n56470__;
  assign new_new_n56472__ = ~new_new_n56411__ & new_new_n56450__;
  assign new_new_n56473__ = new_new_n56361__ & new_new_n56472__;
  assign new_new_n56474__ = new_new_n56411__ & new_new_n56450__;
  assign new_new_n56475__ = ~new_new_n56361__ & new_new_n56474__;
  assign new_new_n56476__ = ~new_new_n56473__ & ~new_new_n56475__;
  assign new_new_n56477__ = ~new_new_n56471__ & new_new_n56476__;
  assign new_new_n56478__ = ~new_new_n56469__ & new_new_n56477__;
  assign new_new_n56479__ = ~new_new_n56249__ & new_new_n56266__;
  assign new_new_n56480__ = new_new_n56234__ & new_new_n56265__;
  assign new_new_n56481__ = ~new_new_n56249__ & new_new_n56480__;
  assign new_new_n56482__ = ~new_new_n56479__ & ~new_new_n56481__;
  assign new_new_n56483__ = ~new_new_n56234__ & new_new_n56265__;
  assign new_new_n56484__ = new_new_n56249__ & new_new_n56483__;
  assign new_new_n56485__ = new_new_n56234__ & ~new_new_n56265__;
  assign new_new_n56486__ = new_new_n56249__ & new_new_n56485__;
  assign new_new_n56487__ = ~new_new_n56484__ & ~new_new_n56486__;
  assign new_new_n56488__ = new_new_n56482__ & new_new_n56487__;
  assign new_new_n56489__ = ~new_new_n56478__ & ~new_new_n56488__;
  assign new_new_n56490__ = ~new_new_n56442__ & new_new_n56447__;
  assign new_new_n56491__ = new_new_n56427__ & new_new_n56446__;
  assign new_new_n56492__ = ~new_new_n56442__ & new_new_n56491__;
  assign new_new_n56493__ = ~new_new_n56490__ & ~new_new_n56492__;
  assign new_new_n56494__ = ~new_new_n56427__ & new_new_n56446__;
  assign new_new_n56495__ = new_new_n56442__ & new_new_n56494__;
  assign new_new_n56496__ = new_new_n56427__ & ~new_new_n56446__;
  assign new_new_n56497__ = new_new_n56442__ & new_new_n56496__;
  assign new_new_n56498__ = ~new_new_n56495__ & ~new_new_n56497__;
  assign new_new_n56499__ = new_new_n56493__ & new_new_n56498__;
  assign new_new_n56500__ = ys__n39736 & new_new_n52412__;
  assign new_new_n56501__ = ys__n39734 & new_new_n52411__;
  assign new_new_n56502__ = ~new_new_n56500__ & ~new_new_n56501__;
  assign new_new_n56503__ = ys__n33701 & new_new_n52425__;
  assign new_new_n56504__ = ~ys__n33701 & new_new_n52428__;
  assign new_new_n56505__ = ~new_new_n56503__ & ~new_new_n56504__;
  assign new_new_n56506__ = new_new_n56502__ & new_new_n56505__;
  assign new_new_n56507__ = ys__n24774 & new_new_n52417__;
  assign new_new_n56508__ = ys__n24771 & new_new_n52420__;
  assign new_new_n56509__ = ~new_new_n56507__ & ~new_new_n56508__;
  assign new_new_n56510__ = ys__n24768 & new_new_n52419__;
  assign new_new_n56511__ = ys__n39738 & new_new_n52409__;
  assign new_new_n56512__ = ~new_new_n56510__ & ~new_new_n56511__;
  assign new_new_n56513__ = new_new_n56509__ & new_new_n56512__;
  assign new_new_n56514__ = new_new_n56506__ & new_new_n56513__;
  assign new_new_n56515__ = ys__n39742 & new_new_n52301__;
  assign new_new_n56516__ = ys__n39740 & new_new_n52304__;
  assign new_new_n56517__ = ~new_new_n56515__ & ~new_new_n56516__;
  assign new_new_n56518__ = ys__n33707 & new_new_n52308__;
  assign new_new_n56519__ = ~ys__n33707 & new_new_n52311__;
  assign new_new_n56520__ = ~new_new_n56518__ & ~new_new_n56519__;
  assign new_new_n56521__ = new_new_n56517__ & new_new_n56520__;
  assign new_new_n56522__ = ys__n24783 & new_new_n52316__;
  assign new_new_n56523__ = ys__n24780 & new_new_n52318__;
  assign new_new_n56524__ = ~new_new_n56522__ & ~new_new_n56523__;
  assign new_new_n56525__ = ys__n24777 & new_new_n52322__;
  assign new_new_n56526__ = ys__n39744 & new_new_n52324__;
  assign new_new_n56527__ = ~new_new_n56525__ & ~new_new_n56526__;
  assign new_new_n56528__ = new_new_n56524__ & new_new_n56527__;
  assign new_new_n56529__ = new_new_n56521__ & new_new_n56528__;
  assign new_new_n56530__ = ~new_new_n56514__ & ~new_new_n56529__;
  assign new_new_n56531__ = ys__n39730 & new_new_n52449__;
  assign new_new_n56532__ = ys__n39728 & new_new_n52448__;
  assign new_new_n56533__ = ~new_new_n56531__ & ~new_new_n56532__;
  assign new_new_n56534__ = ys__n33695 & new_new_n52462__;
  assign new_new_n56535__ = ~ys__n33695 & new_new_n52465__;
  assign new_new_n56536__ = ~new_new_n56534__ & ~new_new_n56535__;
  assign new_new_n56537__ = new_new_n56533__ & new_new_n56536__;
  assign new_new_n56538__ = ys__n24765 & new_new_n52454__;
  assign new_new_n56539__ = ys__n24762 & new_new_n52457__;
  assign new_new_n56540__ = ~new_new_n56538__ & ~new_new_n56539__;
  assign new_new_n56541__ = ys__n24759 & new_new_n52456__;
  assign new_new_n56542__ = ys__n39732 & new_new_n52446__;
  assign new_new_n56543__ = ~new_new_n56541__ & ~new_new_n56542__;
  assign new_new_n56544__ = new_new_n56540__ & new_new_n56543__;
  assign new_new_n56545__ = new_new_n56537__ & new_new_n56544__;
  assign new_new_n56546__ = ~new_new_n56514__ & ~new_new_n56545__;
  assign new_new_n56547__ = ~new_new_n56529__ & ~new_new_n56545__;
  assign new_new_n56548__ = ~new_new_n56546__ & ~new_new_n56547__;
  assign new_new_n56549__ = ~new_new_n56530__ & new_new_n56548__;
  assign new_new_n56550__ = ~new_new_n56499__ & ~new_new_n56549__;
  assign new_new_n56551__ = ys__n39718 & new_new_n52359__;
  assign new_new_n56552__ = ys__n24741 & new_new_n52358__;
  assign new_new_n56553__ = ~new_new_n56551__ & ~new_new_n56552__;
  assign new_new_n56554__ = ys__n33683 & new_new_n52372__;
  assign new_new_n56555__ = ~ys__n33683 & new_new_n52375__;
  assign new_new_n56556__ = ~new_new_n56554__ & ~new_new_n56555__;
  assign new_new_n56557__ = new_new_n56553__ & new_new_n56556__;
  assign new_new_n56558__ = ys__n24747 & new_new_n52364__;
  assign new_new_n56559__ = ys__n24744 & new_new_n52367__;
  assign new_new_n56560__ = ~new_new_n56558__ & ~new_new_n56559__;
  assign new_new_n56561__ = ys__n24741 & new_new_n52366__;
  assign new_new_n56562__ = ys__n39720 & new_new_n52356__;
  assign new_new_n56563__ = ~new_new_n56561__ & ~new_new_n56562__;
  assign new_new_n56564__ = new_new_n56560__ & new_new_n56563__;
  assign new_new_n56565__ = new_new_n56557__ & new_new_n56564__;
  assign new_new_n56566__ = ys__n39724 & new_new_n52334__;
  assign new_new_n56567__ = ys__n39722 & new_new_n52333__;
  assign new_new_n56568__ = ~new_new_n56566__ & ~new_new_n56567__;
  assign new_new_n56569__ = ys__n33689 & new_new_n52347__;
  assign new_new_n56570__ = ~ys__n33689 & new_new_n52350__;
  assign new_new_n56571__ = ~new_new_n56569__ & ~new_new_n56570__;
  assign new_new_n56572__ = new_new_n56568__ & new_new_n56571__;
  assign new_new_n56573__ = ys__n24756 & new_new_n52339__;
  assign new_new_n56574__ = ys__n24753 & new_new_n52342__;
  assign new_new_n56575__ = ~new_new_n56573__ & ~new_new_n56574__;
  assign new_new_n56576__ = ys__n24750 & new_new_n52341__;
  assign new_new_n56577__ = ys__n39726 & new_new_n52331__;
  assign new_new_n56578__ = ~new_new_n56576__ & ~new_new_n56577__;
  assign new_new_n56579__ = new_new_n56575__ & new_new_n56578__;
  assign new_new_n56580__ = new_new_n56572__ & new_new_n56579__;
  assign new_new_n56581__ = ~new_new_n56565__ & ~new_new_n56580__;
  assign new_new_n56582__ = ~new_new_n56499__ & new_new_n56581__;
  assign new_new_n56583__ = ~new_new_n56549__ & new_new_n56581__;
  assign new_new_n56584__ = ~new_new_n56582__ & ~new_new_n56583__;
  assign new_new_n56585__ = ~new_new_n56550__ & new_new_n56584__;
  assign new_new_n56586__ = ~new_new_n56478__ & ~new_new_n56585__;
  assign new_new_n56587__ = ~new_new_n56488__ & ~new_new_n56585__;
  assign new_new_n56588__ = ~new_new_n56586__ & ~new_new_n56587__;
  assign ys__n43835 = new_new_n56489__ | ~new_new_n56588__;
  assign new_new_n56590__ = ~new_new_n56488__ & new_new_n56586__;
  assign new_new_n56591__ = new_new_n56488__ & ~new_new_n56585__;
  assign new_new_n56592__ = new_new_n56478__ & new_new_n56591__;
  assign new_new_n56593__ = ~new_new_n56488__ & new_new_n56585__;
  assign new_new_n56594__ = new_new_n56478__ & new_new_n56593__;
  assign new_new_n56595__ = new_new_n56488__ & new_new_n56585__;
  assign new_new_n56596__ = ~new_new_n56478__ & new_new_n56595__;
  assign new_new_n56597__ = ~new_new_n56594__ & ~new_new_n56596__;
  assign new_new_n56598__ = ~new_new_n56592__ & new_new_n56597__;
  assign ys__n43840 = new_new_n56590__ | ~new_new_n56598__;
  assign new_new_n56600__ = ~new_new_n56549__ & new_new_n56582__;
  assign new_new_n56601__ = new_new_n56549__ & new_new_n56581__;
  assign new_new_n56602__ = new_new_n56499__ & new_new_n56601__;
  assign new_new_n56603__ = ~new_new_n56549__ & ~new_new_n56581__;
  assign new_new_n56604__ = new_new_n56499__ & new_new_n56603__;
  assign new_new_n56605__ = new_new_n56549__ & ~new_new_n56581__;
  assign new_new_n56606__ = ~new_new_n56499__ & new_new_n56605__;
  assign new_new_n56607__ = ~new_new_n56604__ & ~new_new_n56606__;
  assign new_new_n56608__ = ~new_new_n56602__ & new_new_n56607__;
  assign new_new_n56609__ = ~new_new_n56600__ & new_new_n56608__;
  assign new_new_n56610__ = ~new_new_n56391__ & new_new_n56408__;
  assign new_new_n56611__ = new_new_n56376__ & new_new_n56407__;
  assign new_new_n56612__ = ~new_new_n56391__ & new_new_n56611__;
  assign new_new_n56613__ = ~new_new_n56610__ & ~new_new_n56612__;
  assign new_new_n56614__ = ~new_new_n56376__ & new_new_n56407__;
  assign new_new_n56615__ = new_new_n56391__ & new_new_n56614__;
  assign new_new_n56616__ = new_new_n56376__ & ~new_new_n56407__;
  assign new_new_n56617__ = new_new_n56391__ & new_new_n56616__;
  assign new_new_n56618__ = ~new_new_n56615__ & ~new_new_n56617__;
  assign new_new_n56619__ = new_new_n56613__ & new_new_n56618__;
  assign new_new_n56620__ = ~new_new_n56609__ & ~new_new_n56619__;
  assign new_new_n56621__ = new_new_n56565__ & ~new_new_n56580__;
  assign new_new_n56622__ = ~new_new_n56565__ & new_new_n56580__;
  assign new_new_n56623__ = ~new_new_n56621__ & ~new_new_n56622__;
  assign new_new_n56624__ = ys__n39734 & new_new_n52412__;
  assign new_new_n56625__ = ys__n39732 & new_new_n52411__;
  assign new_new_n56626__ = ~new_new_n56624__ & ~new_new_n56625__;
  assign new_new_n56627__ = ys__n33699 & new_new_n52425__;
  assign new_new_n56628__ = ~ys__n33699 & new_new_n52428__;
  assign new_new_n56629__ = ~new_new_n56627__ & ~new_new_n56628__;
  assign new_new_n56630__ = new_new_n56626__ & new_new_n56629__;
  assign new_new_n56631__ = ys__n24771 & new_new_n52417__;
  assign new_new_n56632__ = ys__n24768 & new_new_n52420__;
  assign new_new_n56633__ = ~new_new_n56631__ & ~new_new_n56632__;
  assign new_new_n56634__ = ys__n24765 & new_new_n52419__;
  assign new_new_n56635__ = ys__n39736 & new_new_n52409__;
  assign new_new_n56636__ = ~new_new_n56634__ & ~new_new_n56635__;
  assign new_new_n56637__ = new_new_n56633__ & new_new_n56636__;
  assign new_new_n56638__ = new_new_n56630__ & new_new_n56637__;
  assign new_new_n56639__ = ys__n39740 & new_new_n52301__;
  assign new_new_n56640__ = ys__n39738 & new_new_n52304__;
  assign new_new_n56641__ = ~new_new_n56639__ & ~new_new_n56640__;
  assign new_new_n56642__ = ys__n33705 & new_new_n52308__;
  assign new_new_n56643__ = ~ys__n33705 & new_new_n52311__;
  assign new_new_n56644__ = ~new_new_n56642__ & ~new_new_n56643__;
  assign new_new_n56645__ = new_new_n56641__ & new_new_n56644__;
  assign new_new_n56646__ = ys__n24780 & new_new_n52316__;
  assign new_new_n56647__ = ys__n24777 & new_new_n52318__;
  assign new_new_n56648__ = ~new_new_n56646__ & ~new_new_n56647__;
  assign new_new_n56649__ = ys__n24774 & new_new_n52322__;
  assign new_new_n56650__ = ys__n39742 & new_new_n52324__;
  assign new_new_n56651__ = ~new_new_n56649__ & ~new_new_n56650__;
  assign new_new_n56652__ = new_new_n56648__ & new_new_n56651__;
  assign new_new_n56653__ = new_new_n56645__ & new_new_n56652__;
  assign new_new_n56654__ = ~new_new_n56638__ & ~new_new_n56653__;
  assign new_new_n56655__ = ys__n39728 & new_new_n52449__;
  assign new_new_n56656__ = ys__n39726 & new_new_n52448__;
  assign new_new_n56657__ = ~new_new_n56655__ & ~new_new_n56656__;
  assign new_new_n56658__ = ys__n33693 & new_new_n52462__;
  assign new_new_n56659__ = ~ys__n33693 & new_new_n52465__;
  assign new_new_n56660__ = ~new_new_n56658__ & ~new_new_n56659__;
  assign new_new_n56661__ = new_new_n56657__ & new_new_n56660__;
  assign new_new_n56662__ = ys__n24762 & new_new_n52454__;
  assign new_new_n56663__ = ys__n24759 & new_new_n52457__;
  assign new_new_n56664__ = ~new_new_n56662__ & ~new_new_n56663__;
  assign new_new_n56665__ = ys__n24756 & new_new_n52456__;
  assign new_new_n56666__ = ys__n39730 & new_new_n52446__;
  assign new_new_n56667__ = ~new_new_n56665__ & ~new_new_n56666__;
  assign new_new_n56668__ = new_new_n56664__ & new_new_n56667__;
  assign new_new_n56669__ = new_new_n56661__ & new_new_n56668__;
  assign new_new_n56670__ = ~new_new_n56638__ & ~new_new_n56669__;
  assign new_new_n56671__ = ~new_new_n56653__ & ~new_new_n56669__;
  assign new_new_n56672__ = ~new_new_n56670__ & ~new_new_n56671__;
  assign new_new_n56673__ = ~new_new_n56654__ & new_new_n56672__;
  assign new_new_n56674__ = ~new_new_n56623__ & ~new_new_n56673__;
  assign new_new_n56675__ = ys__n24744 & new_new_n52364__;
  assign new_new_n56676__ = ys__n24741 & new_new_n52367__;
  assign new_new_n56677__ = ~new_new_n56675__ & ~new_new_n56676__;
  assign new_new_n56678__ = ys__n39718 & new_new_n52356__;
  assign new_new_n56679__ = ys__n24741 & new_new_n52359__;
  assign new_new_n56680__ = ~new_new_n56678__ & ~new_new_n56679__;
  assign new_new_n56681__ = ys__n33681 & new_new_n52372__;
  assign new_new_n56682__ = ~ys__n33681 & new_new_n52375__;
  assign new_new_n56683__ = ~new_new_n56681__ & ~new_new_n56682__;
  assign new_new_n56684__ = new_new_n56680__ & new_new_n56683__;
  assign new_new_n56685__ = new_new_n56677__ & new_new_n56684__;
  assign new_new_n56686__ = ys__n39722 & new_new_n52334__;
  assign new_new_n56687__ = ys__n39720 & new_new_n52333__;
  assign new_new_n56688__ = ~new_new_n56686__ & ~new_new_n56687__;
  assign new_new_n56689__ = ys__n33687 & new_new_n52347__;
  assign new_new_n56690__ = ~ys__n33687 & new_new_n52350__;
  assign new_new_n56691__ = ~new_new_n56689__ & ~new_new_n56690__;
  assign new_new_n56692__ = new_new_n56688__ & new_new_n56691__;
  assign new_new_n56693__ = ys__n24753 & new_new_n52339__;
  assign new_new_n56694__ = ys__n24750 & new_new_n52342__;
  assign new_new_n56695__ = ~new_new_n56693__ & ~new_new_n56694__;
  assign new_new_n56696__ = ys__n24747 & new_new_n52341__;
  assign new_new_n56697__ = ys__n39724 & new_new_n52331__;
  assign new_new_n56698__ = ~new_new_n56696__ & ~new_new_n56697__;
  assign new_new_n56699__ = new_new_n56695__ & new_new_n56698__;
  assign new_new_n56700__ = new_new_n56692__ & new_new_n56699__;
  assign new_new_n56701__ = ~new_new_n56685__ & ~new_new_n56700__;
  assign new_new_n56702__ = ~new_new_n56623__ & new_new_n56701__;
  assign new_new_n56703__ = ~new_new_n56673__ & new_new_n56701__;
  assign new_new_n56704__ = ~new_new_n56702__ & ~new_new_n56703__;
  assign new_new_n56705__ = ~new_new_n56674__ & new_new_n56704__;
  assign new_new_n56706__ = ~new_new_n56609__ & ~new_new_n56705__;
  assign new_new_n56707__ = ~new_new_n56619__ & ~new_new_n56705__;
  assign new_new_n56708__ = ~new_new_n56706__ & ~new_new_n56707__;
  assign ys__n43889 = new_new_n56620__ | ~new_new_n56708__;
  assign new_new_n56710__ = ~new_new_n56619__ & new_new_n56706__;
  assign new_new_n56711__ = new_new_n56619__ & ~new_new_n56705__;
  assign new_new_n56712__ = new_new_n56609__ & new_new_n56711__;
  assign new_new_n56713__ = ~new_new_n56619__ & new_new_n56705__;
  assign new_new_n56714__ = new_new_n56609__ & new_new_n56713__;
  assign new_new_n56715__ = new_new_n56619__ & new_new_n56705__;
  assign new_new_n56716__ = ~new_new_n56609__ & new_new_n56715__;
  assign new_new_n56717__ = ~new_new_n56714__ & ~new_new_n56716__;
  assign new_new_n56718__ = ~new_new_n56712__ & new_new_n56717__;
  assign ys__n43894 = new_new_n56710__ | ~new_new_n56718__;
  assign new_new_n56720__ = ~new_new_n56673__ & new_new_n56702__;
  assign new_new_n56721__ = new_new_n56623__ & ~new_new_n56701__;
  assign new_new_n56722__ = ~new_new_n56673__ & new_new_n56721__;
  assign new_new_n56723__ = ~new_new_n56720__ & ~new_new_n56722__;
  assign new_new_n56724__ = ~new_new_n56623__ & ~new_new_n56701__;
  assign new_new_n56725__ = new_new_n56673__ & new_new_n56724__;
  assign new_new_n56726__ = new_new_n56623__ & new_new_n56701__;
  assign new_new_n56727__ = new_new_n56673__ & new_new_n56726__;
  assign new_new_n56728__ = ~new_new_n56725__ & ~new_new_n56727__;
  assign new_new_n56729__ = new_new_n56723__ & new_new_n56728__;
  assign new_new_n56730__ = ~new_new_n56529__ & new_new_n56546__;
  assign new_new_n56731__ = new_new_n56514__ & new_new_n56545__;
  assign new_new_n56732__ = ~new_new_n56529__ & new_new_n56731__;
  assign new_new_n56733__ = ~new_new_n56730__ & ~new_new_n56732__;
  assign new_new_n56734__ = ~new_new_n56514__ & new_new_n56545__;
  assign new_new_n56735__ = new_new_n56529__ & new_new_n56734__;
  assign new_new_n56736__ = new_new_n56514__ & ~new_new_n56545__;
  assign new_new_n56737__ = new_new_n56529__ & new_new_n56736__;
  assign new_new_n56738__ = ~new_new_n56735__ & ~new_new_n56737__;
  assign new_new_n56739__ = new_new_n56733__ & new_new_n56738__;
  assign new_new_n56740__ = ~new_new_n56729__ & ~new_new_n56739__;
  assign new_new_n56741__ = new_new_n56685__ & ~new_new_n56700__;
  assign new_new_n56742__ = ~new_new_n56685__ & new_new_n56700__;
  assign new_new_n56743__ = ~new_new_n56741__ & ~new_new_n56742__;
  assign new_new_n56744__ = ys__n39732 & new_new_n52412__;
  assign new_new_n56745__ = ys__n39730 & new_new_n52411__;
  assign new_new_n56746__ = ~new_new_n56744__ & ~new_new_n56745__;
  assign new_new_n56747__ = ys__n33697 & new_new_n52425__;
  assign new_new_n56748__ = ~ys__n33697 & new_new_n52428__;
  assign new_new_n56749__ = ~new_new_n56747__ & ~new_new_n56748__;
  assign new_new_n56750__ = new_new_n56746__ & new_new_n56749__;
  assign new_new_n56751__ = ys__n24768 & new_new_n52417__;
  assign new_new_n56752__ = ys__n24765 & new_new_n52420__;
  assign new_new_n56753__ = ~new_new_n56751__ & ~new_new_n56752__;
  assign new_new_n56754__ = ys__n24762 & new_new_n52419__;
  assign new_new_n56755__ = ys__n39734 & new_new_n52409__;
  assign new_new_n56756__ = ~new_new_n56754__ & ~new_new_n56755__;
  assign new_new_n56757__ = new_new_n56753__ & new_new_n56756__;
  assign new_new_n56758__ = new_new_n56750__ & new_new_n56757__;
  assign new_new_n56759__ = ys__n39738 & new_new_n52301__;
  assign new_new_n56760__ = ys__n39736 & new_new_n52304__;
  assign new_new_n56761__ = ~new_new_n56759__ & ~new_new_n56760__;
  assign new_new_n56762__ = ys__n33703 & new_new_n52308__;
  assign new_new_n56763__ = ~ys__n33703 & new_new_n52311__;
  assign new_new_n56764__ = ~new_new_n56762__ & ~new_new_n56763__;
  assign new_new_n56765__ = new_new_n56761__ & new_new_n56764__;
  assign new_new_n56766__ = ys__n24777 & new_new_n52316__;
  assign new_new_n56767__ = ys__n24774 & new_new_n52318__;
  assign new_new_n56768__ = ~new_new_n56766__ & ~new_new_n56767__;
  assign new_new_n56769__ = ys__n24771 & new_new_n52322__;
  assign new_new_n56770__ = ys__n39740 & new_new_n52324__;
  assign new_new_n56771__ = ~new_new_n56769__ & ~new_new_n56770__;
  assign new_new_n56772__ = new_new_n56768__ & new_new_n56771__;
  assign new_new_n56773__ = new_new_n56765__ & new_new_n56772__;
  assign new_new_n56774__ = ~new_new_n56758__ & ~new_new_n56773__;
  assign new_new_n56775__ = ys__n39726 & new_new_n52449__;
  assign new_new_n56776__ = ys__n39724 & new_new_n52448__;
  assign new_new_n56777__ = ~new_new_n56775__ & ~new_new_n56776__;
  assign new_new_n56778__ = ys__n33691 & new_new_n52462__;
  assign new_new_n56779__ = ~ys__n33691 & new_new_n52465__;
  assign new_new_n56780__ = ~new_new_n56778__ & ~new_new_n56779__;
  assign new_new_n56781__ = new_new_n56777__ & new_new_n56780__;
  assign new_new_n56782__ = ys__n24759 & new_new_n52454__;
  assign new_new_n56783__ = ys__n24756 & new_new_n52457__;
  assign new_new_n56784__ = ~new_new_n56782__ & ~new_new_n56783__;
  assign new_new_n56785__ = ys__n24753 & new_new_n52456__;
  assign new_new_n56786__ = ys__n39728 & new_new_n52446__;
  assign new_new_n56787__ = ~new_new_n56785__ & ~new_new_n56786__;
  assign new_new_n56788__ = new_new_n56784__ & new_new_n56787__;
  assign new_new_n56789__ = new_new_n56781__ & new_new_n56788__;
  assign new_new_n56790__ = ~new_new_n56758__ & ~new_new_n56789__;
  assign new_new_n56791__ = ~new_new_n56773__ & ~new_new_n56789__;
  assign new_new_n56792__ = ~new_new_n56790__ & ~new_new_n56791__;
  assign new_new_n56793__ = ~new_new_n56774__ & new_new_n56792__;
  assign new_new_n56794__ = ~new_new_n56743__ & ~new_new_n56793__;
  assign new_new_n56795__ = ys__n24741 & new_new_n52364__;
  assign new_new_n56796__ = ys__n24741 & new_new_n52356__;
  assign new_new_n56797__ = ~new_new_n56795__ & ~new_new_n56796__;
  assign new_new_n56798__ = ys__n24741 & new_new_n52372__;
  assign new_new_n56799__ = ~ys__n24741 & new_new_n52375__;
  assign new_new_n56800__ = ~new_new_n56798__ & ~new_new_n56799__;
  assign new_new_n56801__ = new_new_n56797__ & new_new_n56800__;
  assign new_new_n56802__ = ys__n39720 & new_new_n52334__;
  assign new_new_n56803__ = ys__n39718 & new_new_n52333__;
  assign new_new_n56804__ = ~new_new_n56802__ & ~new_new_n56803__;
  assign new_new_n56805__ = ys__n33685 & new_new_n52347__;
  assign new_new_n56806__ = ~ys__n33685 & new_new_n52350__;
  assign new_new_n56807__ = ~new_new_n56805__ & ~new_new_n56806__;
  assign new_new_n56808__ = new_new_n56804__ & new_new_n56807__;
  assign new_new_n56809__ = ys__n24750 & new_new_n52339__;
  assign new_new_n56810__ = ys__n24747 & new_new_n52342__;
  assign new_new_n56811__ = ~new_new_n56809__ & ~new_new_n56810__;
  assign new_new_n56812__ = ys__n24744 & new_new_n52341__;
  assign new_new_n56813__ = ys__n39722 & new_new_n52331__;
  assign new_new_n56814__ = ~new_new_n56812__ & ~new_new_n56813__;
  assign new_new_n56815__ = new_new_n56811__ & new_new_n56814__;
  assign new_new_n56816__ = new_new_n56808__ & new_new_n56815__;
  assign new_new_n56817__ = ~new_new_n56801__ & ~new_new_n56816__;
  assign new_new_n56818__ = new_new_n52375__ & ~new_new_n56801__;
  assign new_new_n56819__ = new_new_n52375__ & ~new_new_n56816__;
  assign new_new_n56820__ = ~new_new_n56818__ & ~new_new_n56819__;
  assign new_new_n56821__ = ~new_new_n56817__ & new_new_n56820__;
  assign new_new_n56822__ = ~new_new_n56743__ & ~new_new_n56821__;
  assign new_new_n56823__ = ~new_new_n56793__ & ~new_new_n56821__;
  assign new_new_n56824__ = ~new_new_n56822__ & ~new_new_n56823__;
  assign new_new_n56825__ = ~new_new_n56794__ & new_new_n56824__;
  assign new_new_n56826__ = ~new_new_n56729__ & ~new_new_n56825__;
  assign new_new_n56827__ = ~new_new_n56739__ & ~new_new_n56825__;
  assign new_new_n56828__ = ~new_new_n56826__ & ~new_new_n56827__;
  assign ys__n43932 = new_new_n56740__ | ~new_new_n56828__;
  assign new_new_n56830__ = ~new_new_n56739__ & new_new_n56826__;
  assign new_new_n56831__ = ~new_new_n56739__ & new_new_n56825__;
  assign new_new_n56832__ = new_new_n56729__ & new_new_n56831__;
  assign new_new_n56833__ = ~new_new_n56830__ & ~new_new_n56832__;
  assign new_new_n56834__ = new_new_n56739__ & new_new_n56825__;
  assign new_new_n56835__ = ~new_new_n56729__ & new_new_n56834__;
  assign new_new_n56836__ = new_new_n56739__ & ~new_new_n56825__;
  assign new_new_n56837__ = new_new_n56729__ & new_new_n56836__;
  assign new_new_n56838__ = ~new_new_n56835__ & ~new_new_n56837__;
  assign ys__n43937 = ~new_new_n56833__ | ~new_new_n56838__;
  assign new_new_n56840__ = ~new_new_n56793__ & new_new_n56822__;
  assign new_new_n56841__ = new_new_n56743__ & new_new_n56821__;
  assign new_new_n56842__ = ~new_new_n56793__ & new_new_n56841__;
  assign new_new_n56843__ = ~new_new_n56840__ & ~new_new_n56842__;
  assign new_new_n56844__ = ~new_new_n56743__ & new_new_n56821__;
  assign new_new_n56845__ = new_new_n56793__ & new_new_n56844__;
  assign new_new_n56846__ = new_new_n56743__ & ~new_new_n56821__;
  assign new_new_n56847__ = new_new_n56793__ & new_new_n56846__;
  assign new_new_n56848__ = ~new_new_n56845__ & ~new_new_n56847__;
  assign new_new_n56849__ = new_new_n56843__ & new_new_n56848__;
  assign new_new_n56850__ = ~new_new_n56653__ & new_new_n56670__;
  assign new_new_n56851__ = new_new_n56638__ & new_new_n56669__;
  assign new_new_n56852__ = ~new_new_n56653__ & new_new_n56851__;
  assign new_new_n56853__ = ~new_new_n56850__ & ~new_new_n56852__;
  assign new_new_n56854__ = ~new_new_n56638__ & new_new_n56669__;
  assign new_new_n56855__ = new_new_n56653__ & new_new_n56854__;
  assign new_new_n56856__ = new_new_n56638__ & ~new_new_n56669__;
  assign new_new_n56857__ = new_new_n56653__ & new_new_n56856__;
  assign new_new_n56858__ = ~new_new_n56855__ & ~new_new_n56857__;
  assign new_new_n56859__ = new_new_n56853__ & new_new_n56858__;
  assign new_new_n56860__ = ~new_new_n56849__ & ~new_new_n56859__;
  assign new_new_n56861__ = ~new_new_n56816__ & new_new_n56818__;
  assign new_new_n56862__ = ~new_new_n52375__ & new_new_n56801__;
  assign new_new_n56863__ = ~new_new_n56816__ & new_new_n56862__;
  assign new_new_n56864__ = ~new_new_n56861__ & ~new_new_n56863__;
  assign new_new_n56865__ = ~new_new_n52375__ & ~new_new_n56801__;
  assign new_new_n56866__ = new_new_n56816__ & new_new_n56865__;
  assign new_new_n56867__ = new_new_n52375__ & new_new_n56801__;
  assign new_new_n56868__ = new_new_n56816__ & new_new_n56867__;
  assign new_new_n56869__ = ~new_new_n56866__ & ~new_new_n56868__;
  assign new_new_n56870__ = new_new_n56864__ & new_new_n56869__;
  assign new_new_n56871__ = ys__n39730 & new_new_n52412__;
  assign new_new_n56872__ = ys__n39728 & new_new_n52411__;
  assign new_new_n56873__ = ~new_new_n56871__ & ~new_new_n56872__;
  assign new_new_n56874__ = ys__n33695 & new_new_n52425__;
  assign new_new_n56875__ = ~ys__n33695 & new_new_n52428__;
  assign new_new_n56876__ = ~new_new_n56874__ & ~new_new_n56875__;
  assign new_new_n56877__ = new_new_n56873__ & new_new_n56876__;
  assign new_new_n56878__ = ys__n24765 & new_new_n52417__;
  assign new_new_n56879__ = ys__n24762 & new_new_n52420__;
  assign new_new_n56880__ = ~new_new_n56878__ & ~new_new_n56879__;
  assign new_new_n56881__ = ys__n24759 & new_new_n52419__;
  assign new_new_n56882__ = ys__n39732 & new_new_n52409__;
  assign new_new_n56883__ = ~new_new_n56881__ & ~new_new_n56882__;
  assign new_new_n56884__ = new_new_n56880__ & new_new_n56883__;
  assign new_new_n56885__ = new_new_n56877__ & new_new_n56884__;
  assign new_new_n56886__ = ys__n39736 & new_new_n52301__;
  assign new_new_n56887__ = ys__n39734 & new_new_n52304__;
  assign new_new_n56888__ = ~new_new_n56886__ & ~new_new_n56887__;
  assign new_new_n56889__ = ys__n33701 & new_new_n52308__;
  assign new_new_n56890__ = ~ys__n33701 & new_new_n52311__;
  assign new_new_n56891__ = ~new_new_n56889__ & ~new_new_n56890__;
  assign new_new_n56892__ = new_new_n56888__ & new_new_n56891__;
  assign new_new_n56893__ = ys__n24774 & new_new_n52316__;
  assign new_new_n56894__ = ys__n24771 & new_new_n52318__;
  assign new_new_n56895__ = ~new_new_n56893__ & ~new_new_n56894__;
  assign new_new_n56896__ = ys__n24768 & new_new_n52322__;
  assign new_new_n56897__ = ys__n39738 & new_new_n52324__;
  assign new_new_n56898__ = ~new_new_n56896__ & ~new_new_n56897__;
  assign new_new_n56899__ = new_new_n56895__ & new_new_n56898__;
  assign new_new_n56900__ = new_new_n56892__ & new_new_n56899__;
  assign new_new_n56901__ = ~new_new_n56885__ & ~new_new_n56900__;
  assign new_new_n56902__ = ys__n39724 & new_new_n52449__;
  assign new_new_n56903__ = ys__n39722 & new_new_n52448__;
  assign new_new_n56904__ = ~new_new_n56902__ & ~new_new_n56903__;
  assign new_new_n56905__ = ys__n33689 & new_new_n52462__;
  assign new_new_n56906__ = ~ys__n33689 & new_new_n52465__;
  assign new_new_n56907__ = ~new_new_n56905__ & ~new_new_n56906__;
  assign new_new_n56908__ = new_new_n56904__ & new_new_n56907__;
  assign new_new_n56909__ = ys__n24756 & new_new_n52454__;
  assign new_new_n56910__ = ys__n24753 & new_new_n52457__;
  assign new_new_n56911__ = ~new_new_n56909__ & ~new_new_n56910__;
  assign new_new_n56912__ = ys__n24750 & new_new_n52456__;
  assign new_new_n56913__ = ys__n39726 & new_new_n52446__;
  assign new_new_n56914__ = ~new_new_n56912__ & ~new_new_n56913__;
  assign new_new_n56915__ = new_new_n56911__ & new_new_n56914__;
  assign new_new_n56916__ = new_new_n56908__ & new_new_n56915__;
  assign new_new_n56917__ = ~new_new_n56885__ & ~new_new_n56916__;
  assign new_new_n56918__ = ~new_new_n56900__ & ~new_new_n56916__;
  assign new_new_n56919__ = ~new_new_n56917__ & ~new_new_n56918__;
  assign new_new_n56920__ = ~new_new_n56901__ & new_new_n56919__;
  assign new_new_n56921__ = ~new_new_n56870__ & ~new_new_n56920__;
  assign new_new_n56922__ = ~new_new_n56849__ & new_new_n56921__;
  assign new_new_n56923__ = ~new_new_n56859__ & new_new_n56921__;
  assign new_new_n56924__ = ~new_new_n56922__ & ~new_new_n56923__;
  assign ys__n43975 = new_new_n56860__ | ~new_new_n56924__;
  assign new_new_n56926__ = ~new_new_n56859__ & new_new_n56922__;
  assign new_new_n56927__ = new_new_n56859__ & new_new_n56921__;
  assign new_new_n56928__ = new_new_n56849__ & new_new_n56927__;
  assign new_new_n56929__ = ~new_new_n56859__ & ~new_new_n56921__;
  assign new_new_n56930__ = new_new_n56849__ & new_new_n56929__;
  assign new_new_n56931__ = new_new_n56859__ & ~new_new_n56921__;
  assign new_new_n56932__ = ~new_new_n56849__ & new_new_n56931__;
  assign new_new_n56933__ = ~new_new_n56930__ & ~new_new_n56932__;
  assign new_new_n56934__ = ~new_new_n56928__ & new_new_n56933__;
  assign ys__n43980 = new_new_n56926__ | ~new_new_n56934__;
  assign new_new_n56936__ = new_new_n56870__ & ~new_new_n56920__;
  assign new_new_n56937__ = ~new_new_n56870__ & new_new_n56920__;
  assign new_new_n56938__ = ~new_new_n56936__ & ~new_new_n56937__;
  assign new_new_n56939__ = ~new_new_n56773__ & new_new_n56790__;
  assign new_new_n56940__ = new_new_n56758__ & new_new_n56789__;
  assign new_new_n56941__ = ~new_new_n56773__ & new_new_n56940__;
  assign new_new_n56942__ = ~new_new_n56939__ & ~new_new_n56941__;
  assign new_new_n56943__ = ~new_new_n56758__ & new_new_n56789__;
  assign new_new_n56944__ = new_new_n56773__ & new_new_n56943__;
  assign new_new_n56945__ = new_new_n56758__ & ~new_new_n56789__;
  assign new_new_n56946__ = new_new_n56773__ & new_new_n56945__;
  assign new_new_n56947__ = ~new_new_n56944__ & ~new_new_n56946__;
  assign new_new_n56948__ = new_new_n56942__ & new_new_n56947__;
  assign new_new_n56949__ = ~new_new_n56938__ & ~new_new_n56948__;
  assign new_new_n56950__ = ys__n39718 & new_new_n52334__;
  assign new_new_n56951__ = ys__n24741 & new_new_n52333__;
  assign new_new_n56952__ = ~new_new_n56950__ & ~new_new_n56951__;
  assign new_new_n56953__ = ys__n33683 & new_new_n52347__;
  assign new_new_n56954__ = ~ys__n33683 & new_new_n52350__;
  assign new_new_n56955__ = ~new_new_n56953__ & ~new_new_n56954__;
  assign new_new_n56956__ = new_new_n56952__ & new_new_n56955__;
  assign new_new_n56957__ = ys__n24747 & new_new_n52339__;
  assign new_new_n56958__ = ys__n24744 & new_new_n52342__;
  assign new_new_n56959__ = ~new_new_n56957__ & ~new_new_n56958__;
  assign new_new_n56960__ = ys__n24741 & new_new_n52341__;
  assign new_new_n56961__ = ys__n39720 & new_new_n52331__;
  assign new_new_n56962__ = ~new_new_n56960__ & ~new_new_n56961__;
  assign new_new_n56963__ = new_new_n56959__ & new_new_n56962__;
  assign new_new_n56964__ = new_new_n56956__ & new_new_n56963__;
  assign new_new_n56965__ = ys__n39728 & new_new_n52412__;
  assign new_new_n56966__ = ys__n39726 & new_new_n52411__;
  assign new_new_n56967__ = ~new_new_n56965__ & ~new_new_n56966__;
  assign new_new_n56968__ = ys__n33693 & new_new_n52425__;
  assign new_new_n56969__ = ~ys__n33693 & new_new_n52428__;
  assign new_new_n56970__ = ~new_new_n56968__ & ~new_new_n56969__;
  assign new_new_n56971__ = new_new_n56967__ & new_new_n56970__;
  assign new_new_n56972__ = ys__n24762 & new_new_n52417__;
  assign new_new_n56973__ = ys__n24759 & new_new_n52420__;
  assign new_new_n56974__ = ~new_new_n56972__ & ~new_new_n56973__;
  assign new_new_n56975__ = ys__n24756 & new_new_n52419__;
  assign new_new_n56976__ = ys__n39730 & new_new_n52409__;
  assign new_new_n56977__ = ~new_new_n56975__ & ~new_new_n56976__;
  assign new_new_n56978__ = new_new_n56974__ & new_new_n56977__;
  assign new_new_n56979__ = new_new_n56971__ & new_new_n56978__;
  assign new_new_n56980__ = ys__n39734 & new_new_n52301__;
  assign new_new_n56981__ = ys__n39732 & new_new_n52304__;
  assign new_new_n56982__ = ~new_new_n56980__ & ~new_new_n56981__;
  assign new_new_n56983__ = ys__n33699 & new_new_n52308__;
  assign new_new_n56984__ = ~ys__n33699 & new_new_n52311__;
  assign new_new_n56985__ = ~new_new_n56983__ & ~new_new_n56984__;
  assign new_new_n56986__ = new_new_n56982__ & new_new_n56985__;
  assign new_new_n56987__ = ys__n24771 & new_new_n52316__;
  assign new_new_n56988__ = ys__n24768 & new_new_n52318__;
  assign new_new_n56989__ = ~new_new_n56987__ & ~new_new_n56988__;
  assign new_new_n56990__ = ys__n24765 & new_new_n52322__;
  assign new_new_n56991__ = ys__n39736 & new_new_n52324__;
  assign new_new_n56992__ = ~new_new_n56990__ & ~new_new_n56991__;
  assign new_new_n56993__ = new_new_n56989__ & new_new_n56992__;
  assign new_new_n56994__ = new_new_n56986__ & new_new_n56993__;
  assign new_new_n56995__ = ~new_new_n56979__ & ~new_new_n56994__;
  assign new_new_n56996__ = ys__n39722 & new_new_n52449__;
  assign new_new_n56997__ = ys__n39720 & new_new_n52448__;
  assign new_new_n56998__ = ~new_new_n56996__ & ~new_new_n56997__;
  assign new_new_n56999__ = ys__n33687 & new_new_n52462__;
  assign new_new_n57000__ = ~ys__n33687 & new_new_n52465__;
  assign new_new_n57001__ = ~new_new_n56999__ & ~new_new_n57000__;
  assign new_new_n57002__ = new_new_n56998__ & new_new_n57001__;
  assign new_new_n57003__ = ys__n24753 & new_new_n52454__;
  assign new_new_n57004__ = ys__n24750 & new_new_n52457__;
  assign new_new_n57005__ = ~new_new_n57003__ & ~new_new_n57004__;
  assign new_new_n57006__ = ys__n24747 & new_new_n52456__;
  assign new_new_n57007__ = ys__n39724 & new_new_n52446__;
  assign new_new_n57008__ = ~new_new_n57006__ & ~new_new_n57007__;
  assign new_new_n57009__ = new_new_n57005__ & new_new_n57008__;
  assign new_new_n57010__ = new_new_n57002__ & new_new_n57009__;
  assign new_new_n57011__ = ~new_new_n56979__ & ~new_new_n57010__;
  assign new_new_n57012__ = ~new_new_n56994__ & ~new_new_n57010__;
  assign new_new_n57013__ = ~new_new_n57011__ & ~new_new_n57012__;
  assign new_new_n57014__ = ~new_new_n56995__ & new_new_n57013__;
  assign new_new_n57015__ = ~new_new_n56964__ & ~new_new_n57014__;
  assign new_new_n57016__ = ~new_new_n56938__ & new_new_n57015__;
  assign new_new_n57017__ = ~new_new_n56948__ & new_new_n57015__;
  assign new_new_n57018__ = ~new_new_n57016__ & ~new_new_n57017__;
  assign ys__n44018 = new_new_n56949__ | ~new_new_n57018__;
  assign new_new_n57020__ = ~new_new_n56948__ & new_new_n57016__;
  assign new_new_n57021__ = new_new_n56948__ & new_new_n57015__;
  assign new_new_n57022__ = new_new_n56938__ & new_new_n57021__;
  assign new_new_n57023__ = ~new_new_n56948__ & ~new_new_n57015__;
  assign new_new_n57024__ = new_new_n56938__ & new_new_n57023__;
  assign new_new_n57025__ = new_new_n56948__ & ~new_new_n57015__;
  assign new_new_n57026__ = ~new_new_n56938__ & new_new_n57025__;
  assign new_new_n57027__ = ~new_new_n57024__ & ~new_new_n57026__;
  assign new_new_n57028__ = ~new_new_n57022__ & new_new_n57027__;
  assign ys__n44023 = new_new_n57020__ | ~new_new_n57028__;
  assign new_new_n57030__ = ys__n24744 & new_new_n52339__;
  assign new_new_n57031__ = ys__n24741 & new_new_n52342__;
  assign new_new_n57032__ = ~new_new_n57030__ & ~new_new_n57031__;
  assign new_new_n57033__ = ys__n39718 & new_new_n52331__;
  assign new_new_n57034__ = ys__n24741 & new_new_n52334__;
  assign new_new_n57035__ = ~new_new_n57033__ & ~new_new_n57034__;
  assign new_new_n57036__ = ys__n33681 & new_new_n52347__;
  assign new_new_n57037__ = ~ys__n33681 & new_new_n52350__;
  assign new_new_n57038__ = ~new_new_n57036__ & ~new_new_n57037__;
  assign new_new_n57039__ = new_new_n57035__ & new_new_n57038__;
  assign new_new_n57040__ = new_new_n57032__ & new_new_n57039__;
  assign new_new_n57041__ = ys__n39726 & new_new_n52412__;
  assign new_new_n57042__ = ys__n39724 & new_new_n52411__;
  assign new_new_n57043__ = ~new_new_n57041__ & ~new_new_n57042__;
  assign new_new_n57044__ = ys__n33691 & new_new_n52425__;
  assign new_new_n57045__ = ~ys__n33691 & new_new_n52428__;
  assign new_new_n57046__ = ~new_new_n57044__ & ~new_new_n57045__;
  assign new_new_n57047__ = new_new_n57043__ & new_new_n57046__;
  assign new_new_n57048__ = ys__n24759 & new_new_n52417__;
  assign new_new_n57049__ = ys__n24756 & new_new_n52420__;
  assign new_new_n57050__ = ~new_new_n57048__ & ~new_new_n57049__;
  assign new_new_n57051__ = ys__n24753 & new_new_n52419__;
  assign new_new_n57052__ = ys__n39728 & new_new_n52409__;
  assign new_new_n57053__ = ~new_new_n57051__ & ~new_new_n57052__;
  assign new_new_n57054__ = new_new_n57050__ & new_new_n57053__;
  assign new_new_n57055__ = new_new_n57047__ & new_new_n57054__;
  assign new_new_n57056__ = ys__n39732 & new_new_n52301__;
  assign new_new_n57057__ = ys__n39730 & new_new_n52304__;
  assign new_new_n57058__ = ~new_new_n57056__ & ~new_new_n57057__;
  assign new_new_n57059__ = ys__n33697 & new_new_n52308__;
  assign new_new_n57060__ = ~ys__n33697 & new_new_n52311__;
  assign new_new_n57061__ = ~new_new_n57059__ & ~new_new_n57060__;
  assign new_new_n57062__ = new_new_n57058__ & new_new_n57061__;
  assign new_new_n57063__ = ys__n24768 & new_new_n52316__;
  assign new_new_n57064__ = ys__n24765 & new_new_n52318__;
  assign new_new_n57065__ = ~new_new_n57063__ & ~new_new_n57064__;
  assign new_new_n57066__ = ys__n24762 & new_new_n52322__;
  assign new_new_n57067__ = ys__n39734 & new_new_n52324__;
  assign new_new_n57068__ = ~new_new_n57066__ & ~new_new_n57067__;
  assign new_new_n57069__ = new_new_n57065__ & new_new_n57068__;
  assign new_new_n57070__ = new_new_n57062__ & new_new_n57069__;
  assign new_new_n57071__ = ~new_new_n57055__ & ~new_new_n57070__;
  assign new_new_n57072__ = ys__n39720 & new_new_n52449__;
  assign new_new_n57073__ = ys__n39718 & new_new_n52448__;
  assign new_new_n57074__ = ~new_new_n57072__ & ~new_new_n57073__;
  assign new_new_n57075__ = ys__n33685 & new_new_n52462__;
  assign new_new_n57076__ = ~ys__n33685 & new_new_n52465__;
  assign new_new_n57077__ = ~new_new_n57075__ & ~new_new_n57076__;
  assign new_new_n57078__ = new_new_n57074__ & new_new_n57077__;
  assign new_new_n57079__ = ys__n24750 & new_new_n52454__;
  assign new_new_n57080__ = ys__n24747 & new_new_n52457__;
  assign new_new_n57081__ = ~new_new_n57079__ & ~new_new_n57080__;
  assign new_new_n57082__ = ys__n24744 & new_new_n52456__;
  assign new_new_n57083__ = ys__n39722 & new_new_n52446__;
  assign new_new_n57084__ = ~new_new_n57082__ & ~new_new_n57083__;
  assign new_new_n57085__ = new_new_n57081__ & new_new_n57084__;
  assign new_new_n57086__ = new_new_n57078__ & new_new_n57085__;
  assign new_new_n57087__ = ~new_new_n57055__ & ~new_new_n57086__;
  assign new_new_n57088__ = ~new_new_n57070__ & ~new_new_n57086__;
  assign new_new_n57089__ = ~new_new_n57087__ & ~new_new_n57088__;
  assign new_new_n57090__ = ~new_new_n57071__ & new_new_n57089__;
  assign new_new_n57091__ = ~new_new_n57040__ & ~new_new_n57090__;
  assign new_new_n57092__ = ys__n24741 & new_new_n52339__;
  assign new_new_n57093__ = ys__n24741 & new_new_n52331__;
  assign new_new_n57094__ = ~new_new_n57092__ & ~new_new_n57093__;
  assign new_new_n57095__ = ys__n24741 & new_new_n52347__;
  assign new_new_n57096__ = ~ys__n24741 & new_new_n52350__;
  assign new_new_n57097__ = ~new_new_n57095__ & ~new_new_n57096__;
  assign new_new_n57098__ = new_new_n57094__ & new_new_n57097__;
  assign new_new_n57099__ = new_new_n52350__ & ~new_new_n57098__;
  assign new_new_n57100__ = ~new_new_n57040__ & new_new_n57099__;
  assign new_new_n57101__ = ~new_new_n57090__ & new_new_n57099__;
  assign new_new_n57102__ = ~new_new_n57100__ & ~new_new_n57101__;
  assign new_new_n57103__ = ~new_new_n57091__ & new_new_n57102__;
  assign new_new_n57104__ = ~new_new_n56900__ & new_new_n56917__;
  assign new_new_n57105__ = new_new_n56885__ & new_new_n56916__;
  assign new_new_n57106__ = ~new_new_n56900__ & new_new_n57105__;
  assign new_new_n57107__ = ~new_new_n57104__ & ~new_new_n57106__;
  assign new_new_n57108__ = ~new_new_n56885__ & new_new_n56916__;
  assign new_new_n57109__ = new_new_n56900__ & new_new_n57108__;
  assign new_new_n57110__ = new_new_n56885__ & ~new_new_n56916__;
  assign new_new_n57111__ = new_new_n56900__ & new_new_n57110__;
  assign new_new_n57112__ = ~new_new_n57109__ & ~new_new_n57111__;
  assign new_new_n57113__ = new_new_n57107__ & new_new_n57112__;
  assign new_new_n57114__ = ~new_new_n57103__ & ~new_new_n57113__;
  assign new_new_n57115__ = new_new_n56964__ & ~new_new_n57014__;
  assign new_new_n57116__ = ~new_new_n56964__ & new_new_n57014__;
  assign new_new_n57117__ = ~new_new_n57115__ & ~new_new_n57116__;
  assign new_new_n57118__ = ~new_new_n57103__ & ~new_new_n57117__;
  assign new_new_n57119__ = ~new_new_n57113__ & ~new_new_n57117__;
  assign new_new_n57120__ = ~new_new_n57118__ & ~new_new_n57119__;
  assign ys__n44048 = new_new_n57114__ | ~new_new_n57120__;
  assign new_new_n57122__ = ~new_new_n57113__ & new_new_n57118__;
  assign new_new_n57123__ = new_new_n57113__ & new_new_n57117__;
  assign new_new_n57124__ = ~new_new_n57103__ & new_new_n57123__;
  assign new_new_n57125__ = ~new_new_n57113__ & new_new_n57117__;
  assign new_new_n57126__ = new_new_n57103__ & new_new_n57125__;
  assign new_new_n57127__ = new_new_n57113__ & ~new_new_n57117__;
  assign new_new_n57128__ = new_new_n57103__ & new_new_n57127__;
  assign new_new_n57129__ = ~new_new_n57126__ & ~new_new_n57128__;
  assign new_new_n57130__ = ~new_new_n57124__ & new_new_n57129__;
  assign ys__n44053 = new_new_n57122__ | ~new_new_n57130__;
  assign new_new_n57132__ = ~new_new_n57090__ & new_new_n57100__;
  assign new_new_n57133__ = new_new_n57040__ & ~new_new_n57099__;
  assign new_new_n57134__ = ~new_new_n57090__ & new_new_n57133__;
  assign new_new_n57135__ = ~new_new_n57132__ & ~new_new_n57134__;
  assign new_new_n57136__ = ~new_new_n57040__ & ~new_new_n57099__;
  assign new_new_n57137__ = new_new_n57090__ & new_new_n57136__;
  assign new_new_n57138__ = new_new_n57040__ & new_new_n57099__;
  assign new_new_n57139__ = new_new_n57090__ & new_new_n57138__;
  assign new_new_n57140__ = ~new_new_n57137__ & ~new_new_n57139__;
  assign new_new_n57141__ = new_new_n57135__ & new_new_n57140__;
  assign new_new_n57142__ = ~new_new_n56994__ & new_new_n57011__;
  assign new_new_n57143__ = new_new_n56979__ & new_new_n57010__;
  assign new_new_n57144__ = ~new_new_n56994__ & new_new_n57143__;
  assign new_new_n57145__ = ~new_new_n57142__ & ~new_new_n57144__;
  assign new_new_n57146__ = ~new_new_n56979__ & new_new_n57010__;
  assign new_new_n57147__ = new_new_n56994__ & new_new_n57146__;
  assign new_new_n57148__ = new_new_n56979__ & ~new_new_n57010__;
  assign new_new_n57149__ = new_new_n56994__ & new_new_n57148__;
  assign new_new_n57150__ = ~new_new_n57147__ & ~new_new_n57149__;
  assign new_new_n57151__ = new_new_n57145__ & new_new_n57150__;
  assign new_new_n57152__ = ~new_new_n57141__ & ~new_new_n57151__;
  assign new_new_n57153__ = ~new_new_n52350__ & ~new_new_n57098__;
  assign new_new_n57154__ = new_new_n52350__ & new_new_n57098__;
  assign new_new_n57155__ = ~new_new_n57153__ & ~new_new_n57154__;
  assign new_new_n57156__ = ys__n39724 & new_new_n52412__;
  assign new_new_n57157__ = ys__n39722 & new_new_n52411__;
  assign new_new_n57158__ = ~new_new_n57156__ & ~new_new_n57157__;
  assign new_new_n57159__ = ys__n33689 & new_new_n52425__;
  assign new_new_n57160__ = ~ys__n33689 & new_new_n52428__;
  assign new_new_n57161__ = ~new_new_n57159__ & ~new_new_n57160__;
  assign new_new_n57162__ = new_new_n57158__ & new_new_n57161__;
  assign new_new_n57163__ = ys__n24756 & new_new_n52417__;
  assign new_new_n57164__ = ys__n24753 & new_new_n52420__;
  assign new_new_n57165__ = ~new_new_n57163__ & ~new_new_n57164__;
  assign new_new_n57166__ = ys__n24750 & new_new_n52419__;
  assign new_new_n57167__ = ys__n39726 & new_new_n52409__;
  assign new_new_n57168__ = ~new_new_n57166__ & ~new_new_n57167__;
  assign new_new_n57169__ = new_new_n57165__ & new_new_n57168__;
  assign new_new_n57170__ = new_new_n57162__ & new_new_n57169__;
  assign new_new_n57171__ = ys__n39730 & new_new_n52301__;
  assign new_new_n57172__ = ys__n39728 & new_new_n52304__;
  assign new_new_n57173__ = ~new_new_n57171__ & ~new_new_n57172__;
  assign new_new_n57174__ = ys__n33695 & new_new_n52308__;
  assign new_new_n57175__ = ~ys__n33695 & new_new_n52311__;
  assign new_new_n57176__ = ~new_new_n57174__ & ~new_new_n57175__;
  assign new_new_n57177__ = new_new_n57173__ & new_new_n57176__;
  assign new_new_n57178__ = ys__n24765 & new_new_n52316__;
  assign new_new_n57179__ = ys__n24762 & new_new_n52318__;
  assign new_new_n57180__ = ~new_new_n57178__ & ~new_new_n57179__;
  assign new_new_n57181__ = ys__n24759 & new_new_n52322__;
  assign new_new_n57182__ = ys__n39732 & new_new_n52324__;
  assign new_new_n57183__ = ~new_new_n57181__ & ~new_new_n57182__;
  assign new_new_n57184__ = new_new_n57180__ & new_new_n57183__;
  assign new_new_n57185__ = new_new_n57177__ & new_new_n57184__;
  assign new_new_n57186__ = ~new_new_n57170__ & ~new_new_n57185__;
  assign new_new_n57187__ = ys__n39718 & new_new_n52449__;
  assign new_new_n57188__ = ys__n24741 & new_new_n52448__;
  assign new_new_n57189__ = ~new_new_n57187__ & ~new_new_n57188__;
  assign new_new_n57190__ = ys__n33683 & new_new_n52462__;
  assign new_new_n57191__ = ~ys__n33683 & new_new_n52465__;
  assign new_new_n57192__ = ~new_new_n57190__ & ~new_new_n57191__;
  assign new_new_n57193__ = new_new_n57189__ & new_new_n57192__;
  assign new_new_n57194__ = ys__n24747 & new_new_n52454__;
  assign new_new_n57195__ = ys__n24744 & new_new_n52457__;
  assign new_new_n57196__ = ~new_new_n57194__ & ~new_new_n57195__;
  assign new_new_n57197__ = ys__n24741 & new_new_n52456__;
  assign new_new_n57198__ = ys__n39720 & new_new_n52446__;
  assign new_new_n57199__ = ~new_new_n57197__ & ~new_new_n57198__;
  assign new_new_n57200__ = new_new_n57196__ & new_new_n57199__;
  assign new_new_n57201__ = new_new_n57193__ & new_new_n57200__;
  assign new_new_n57202__ = ~new_new_n57170__ & ~new_new_n57201__;
  assign new_new_n57203__ = ~new_new_n57185__ & ~new_new_n57201__;
  assign new_new_n57204__ = ~new_new_n57202__ & ~new_new_n57203__;
  assign new_new_n57205__ = ~new_new_n57186__ & new_new_n57204__;
  assign new_new_n57206__ = ~new_new_n57155__ & ~new_new_n57205__;
  assign new_new_n57207__ = ~new_new_n57141__ & new_new_n57206__;
  assign new_new_n57208__ = ~new_new_n57151__ & new_new_n57206__;
  assign new_new_n57209__ = ~new_new_n57207__ & ~new_new_n57208__;
  assign ys__n44089 = new_new_n57152__ | ~new_new_n57209__;
  assign new_new_n57211__ = ~new_new_n57151__ & new_new_n57207__;
  assign new_new_n57212__ = new_new_n57151__ & new_new_n57206__;
  assign new_new_n57213__ = new_new_n57141__ & new_new_n57212__;
  assign new_new_n57214__ = ~new_new_n57151__ & ~new_new_n57206__;
  assign new_new_n57215__ = new_new_n57141__ & new_new_n57214__;
  assign new_new_n57216__ = new_new_n57151__ & ~new_new_n57206__;
  assign new_new_n57217__ = ~new_new_n57141__ & new_new_n57216__;
  assign new_new_n57218__ = ~new_new_n57215__ & ~new_new_n57217__;
  assign new_new_n57219__ = ~new_new_n57213__ & new_new_n57218__;
  assign ys__n44094 = new_new_n57211__ | ~new_new_n57219__;
  assign new_new_n57221__ = new_new_n57155__ & ~new_new_n57205__;
  assign new_new_n57222__ = ~new_new_n57155__ & new_new_n57205__;
  assign new_new_n57223__ = ~new_new_n57221__ & ~new_new_n57222__;
  assign new_new_n57224__ = ~new_new_n57070__ & new_new_n57087__;
  assign new_new_n57225__ = new_new_n57055__ & new_new_n57086__;
  assign new_new_n57226__ = ~new_new_n57070__ & new_new_n57225__;
  assign new_new_n57227__ = ~new_new_n57224__ & ~new_new_n57226__;
  assign new_new_n57228__ = ~new_new_n57055__ & new_new_n57086__;
  assign new_new_n57229__ = new_new_n57070__ & new_new_n57228__;
  assign new_new_n57230__ = new_new_n57055__ & ~new_new_n57086__;
  assign new_new_n57231__ = new_new_n57070__ & new_new_n57230__;
  assign new_new_n57232__ = ~new_new_n57229__ & ~new_new_n57231__;
  assign new_new_n57233__ = new_new_n57227__ & new_new_n57232__;
  assign ys__n44119 = ~new_new_n57223__ & ~new_new_n57233__;
  assign new_new_n57235__ = new_new_n57223__ & ~new_new_n57233__;
  assign new_new_n57236__ = ~new_new_n57223__ & new_new_n57233__;
  assign ys__n44122 = new_new_n57235__ | new_new_n57236__;
  assign new_new_n57238__ = ys__n39722 & new_new_n52412__;
  assign new_new_n57239__ = ys__n39720 & new_new_n52411__;
  assign new_new_n57240__ = ~new_new_n57238__ & ~new_new_n57239__;
  assign new_new_n57241__ = ys__n33687 & new_new_n52425__;
  assign new_new_n57242__ = ~ys__n33687 & new_new_n52428__;
  assign new_new_n57243__ = ~new_new_n57241__ & ~new_new_n57242__;
  assign new_new_n57244__ = new_new_n57240__ & new_new_n57243__;
  assign new_new_n57245__ = ys__n24753 & new_new_n52417__;
  assign new_new_n57246__ = ys__n24750 & new_new_n52420__;
  assign new_new_n57247__ = ~new_new_n57245__ & ~new_new_n57246__;
  assign new_new_n57248__ = ys__n24747 & new_new_n52419__;
  assign new_new_n57249__ = ys__n39724 & new_new_n52409__;
  assign new_new_n57250__ = ~new_new_n57248__ & ~new_new_n57249__;
  assign new_new_n57251__ = new_new_n57247__ & new_new_n57250__;
  assign new_new_n57252__ = new_new_n57244__ & new_new_n57251__;
  assign new_new_n57253__ = ys__n39728 & new_new_n52301__;
  assign new_new_n57254__ = ys__n39726 & new_new_n52304__;
  assign new_new_n57255__ = ~new_new_n57253__ & ~new_new_n57254__;
  assign new_new_n57256__ = ys__n33693 & new_new_n52308__;
  assign new_new_n57257__ = ~ys__n33693 & new_new_n52311__;
  assign new_new_n57258__ = ~new_new_n57256__ & ~new_new_n57257__;
  assign new_new_n57259__ = new_new_n57255__ & new_new_n57258__;
  assign new_new_n57260__ = ys__n24762 & new_new_n52316__;
  assign new_new_n57261__ = ys__n24759 & new_new_n52318__;
  assign new_new_n57262__ = ~new_new_n57260__ & ~new_new_n57261__;
  assign new_new_n57263__ = ys__n24756 & new_new_n52322__;
  assign new_new_n57264__ = ys__n39730 & new_new_n52324__;
  assign new_new_n57265__ = ~new_new_n57263__ & ~new_new_n57264__;
  assign new_new_n57266__ = new_new_n57262__ & new_new_n57265__;
  assign new_new_n57267__ = new_new_n57259__ & new_new_n57266__;
  assign new_new_n57268__ = ~new_new_n57252__ & ~new_new_n57267__;
  assign new_new_n57269__ = ys__n24744 & new_new_n52454__;
  assign new_new_n57270__ = ys__n24741 & new_new_n52457__;
  assign new_new_n57271__ = ~new_new_n57269__ & ~new_new_n57270__;
  assign new_new_n57272__ = ys__n39718 & new_new_n52446__;
  assign new_new_n57273__ = ys__n24741 & new_new_n52449__;
  assign new_new_n57274__ = ~new_new_n57272__ & ~new_new_n57273__;
  assign new_new_n57275__ = ys__n33681 & new_new_n52462__;
  assign new_new_n57276__ = ~ys__n33681 & new_new_n52465__;
  assign new_new_n57277__ = ~new_new_n57275__ & ~new_new_n57276__;
  assign new_new_n57278__ = new_new_n57274__ & new_new_n57277__;
  assign new_new_n57279__ = new_new_n57271__ & new_new_n57278__;
  assign new_new_n57280__ = ~new_new_n57252__ & ~new_new_n57279__;
  assign new_new_n57281__ = ~new_new_n57267__ & ~new_new_n57279__;
  assign new_new_n57282__ = ~new_new_n57280__ & ~new_new_n57281__;
  assign new_new_n57283__ = ~new_new_n57268__ & new_new_n57282__;
  assign new_new_n57284__ = ~new_new_n57185__ & new_new_n57202__;
  assign new_new_n57285__ = new_new_n57170__ & new_new_n57201__;
  assign new_new_n57286__ = ~new_new_n57185__ & new_new_n57285__;
  assign new_new_n57287__ = ~new_new_n57284__ & ~new_new_n57286__;
  assign new_new_n57288__ = ~new_new_n57170__ & new_new_n57201__;
  assign new_new_n57289__ = new_new_n57185__ & new_new_n57288__;
  assign new_new_n57290__ = new_new_n57170__ & ~new_new_n57201__;
  assign new_new_n57291__ = new_new_n57185__ & new_new_n57290__;
  assign new_new_n57292__ = ~new_new_n57289__ & ~new_new_n57291__;
  assign new_new_n57293__ = new_new_n57287__ & new_new_n57292__;
  assign ys__n44136 = ~new_new_n57283__ & ~new_new_n57293__;
  assign new_new_n57295__ = new_new_n57283__ & ~new_new_n57293__;
  assign new_new_n57296__ = ~new_new_n57283__ & new_new_n57293__;
  assign ys__n44139 = new_new_n57295__ | new_new_n57296__;
  assign new_new_n57298__ = ys__n39720 & new_new_n52412__;
  assign new_new_n57299__ = ys__n39718 & new_new_n52411__;
  assign new_new_n57300__ = ~new_new_n57298__ & ~new_new_n57299__;
  assign new_new_n57301__ = ys__n33685 & new_new_n52425__;
  assign new_new_n57302__ = ~ys__n33685 & new_new_n52428__;
  assign new_new_n57303__ = ~new_new_n57301__ & ~new_new_n57302__;
  assign new_new_n57304__ = new_new_n57300__ & new_new_n57303__;
  assign new_new_n57305__ = ys__n24750 & new_new_n52417__;
  assign new_new_n57306__ = ys__n24747 & new_new_n52420__;
  assign new_new_n57307__ = ~new_new_n57305__ & ~new_new_n57306__;
  assign new_new_n57308__ = ys__n24744 & new_new_n52419__;
  assign new_new_n57309__ = ys__n39722 & new_new_n52409__;
  assign new_new_n57310__ = ~new_new_n57308__ & ~new_new_n57309__;
  assign new_new_n57311__ = new_new_n57307__ & new_new_n57310__;
  assign new_new_n57312__ = new_new_n57304__ & new_new_n57311__;
  assign new_new_n57313__ = ys__n39726 & new_new_n52301__;
  assign new_new_n57314__ = ys__n39724 & new_new_n52304__;
  assign new_new_n57315__ = ~new_new_n57313__ & ~new_new_n57314__;
  assign new_new_n57316__ = ys__n33691 & new_new_n52308__;
  assign new_new_n57317__ = ~ys__n33691 & new_new_n52311__;
  assign new_new_n57318__ = ~new_new_n57316__ & ~new_new_n57317__;
  assign new_new_n57319__ = new_new_n57315__ & new_new_n57318__;
  assign new_new_n57320__ = ys__n24759 & new_new_n52316__;
  assign new_new_n57321__ = ys__n24756 & new_new_n52318__;
  assign new_new_n57322__ = ~new_new_n57320__ & ~new_new_n57321__;
  assign new_new_n57323__ = ys__n24753 & new_new_n52322__;
  assign new_new_n57324__ = ys__n39728 & new_new_n52324__;
  assign new_new_n57325__ = ~new_new_n57323__ & ~new_new_n57324__;
  assign new_new_n57326__ = new_new_n57322__ & new_new_n57325__;
  assign new_new_n57327__ = new_new_n57319__ & new_new_n57326__;
  assign new_new_n57328__ = ~new_new_n57312__ & ~new_new_n57327__;
  assign new_new_n57329__ = ys__n24741 & new_new_n52454__;
  assign new_new_n57330__ = ys__n24741 & new_new_n52446__;
  assign new_new_n57331__ = ~new_new_n57329__ & ~new_new_n57330__;
  assign new_new_n57332__ = ys__n24741 & new_new_n52462__;
  assign new_new_n57333__ = ~ys__n24741 & new_new_n52465__;
  assign new_new_n57334__ = ~new_new_n57332__ & ~new_new_n57333__;
  assign new_new_n57335__ = new_new_n57331__ & new_new_n57334__;
  assign new_new_n57336__ = ~new_new_n57312__ & ~new_new_n57335__;
  assign new_new_n57337__ = ~new_new_n57327__ & ~new_new_n57335__;
  assign new_new_n57338__ = ~new_new_n57336__ & ~new_new_n57337__;
  assign new_new_n57339__ = ~new_new_n57328__ & new_new_n57338__;
  assign new_new_n57340__ = ~new_new_n57267__ & new_new_n57280__;
  assign new_new_n57341__ = new_new_n57252__ & new_new_n57279__;
  assign new_new_n57342__ = ~new_new_n57267__ & new_new_n57341__;
  assign new_new_n57343__ = ~new_new_n57340__ & ~new_new_n57342__;
  assign new_new_n57344__ = ~new_new_n57252__ & new_new_n57279__;
  assign new_new_n57345__ = new_new_n57267__ & new_new_n57344__;
  assign new_new_n57346__ = new_new_n57252__ & ~new_new_n57279__;
  assign new_new_n57347__ = new_new_n57267__ & new_new_n57346__;
  assign new_new_n57348__ = ~new_new_n57345__ & ~new_new_n57347__;
  assign new_new_n57349__ = new_new_n57343__ & new_new_n57348__;
  assign new_new_n57350__ = ~new_new_n57339__ & ~new_new_n57349__;
  assign new_new_n57351__ = ys__n39718 & new_new_n52412__;
  assign new_new_n57352__ = ys__n24741 & new_new_n52411__;
  assign new_new_n57353__ = ~new_new_n57351__ & ~new_new_n57352__;
  assign new_new_n57354__ = ys__n33683 & new_new_n52425__;
  assign new_new_n57355__ = ~ys__n33683 & new_new_n52428__;
  assign new_new_n57356__ = ~new_new_n57354__ & ~new_new_n57355__;
  assign new_new_n57357__ = new_new_n57353__ & new_new_n57356__;
  assign new_new_n57358__ = ys__n24747 & new_new_n52417__;
  assign new_new_n57359__ = ys__n24744 & new_new_n52420__;
  assign new_new_n57360__ = ~new_new_n57358__ & ~new_new_n57359__;
  assign new_new_n57361__ = ys__n24741 & new_new_n52419__;
  assign new_new_n57362__ = ys__n39720 & new_new_n52409__;
  assign new_new_n57363__ = ~new_new_n57361__ & ~new_new_n57362__;
  assign new_new_n57364__ = new_new_n57360__ & new_new_n57363__;
  assign new_new_n57365__ = new_new_n57357__ & new_new_n57364__;
  assign new_new_n57366__ = ys__n39724 & new_new_n52301__;
  assign new_new_n57367__ = ys__n39722 & new_new_n52304__;
  assign new_new_n57368__ = ~new_new_n57366__ & ~new_new_n57367__;
  assign new_new_n57369__ = ys__n33689 & new_new_n52308__;
  assign new_new_n57370__ = ~ys__n33689 & new_new_n52311__;
  assign new_new_n57371__ = ~new_new_n57369__ & ~new_new_n57370__;
  assign new_new_n57372__ = new_new_n57368__ & new_new_n57371__;
  assign new_new_n57373__ = ys__n24756 & new_new_n52316__;
  assign new_new_n57374__ = ys__n24753 & new_new_n52318__;
  assign new_new_n57375__ = ~new_new_n57373__ & ~new_new_n57374__;
  assign new_new_n57376__ = ys__n24750 & new_new_n52322__;
  assign new_new_n57377__ = ys__n39726 & new_new_n52324__;
  assign new_new_n57378__ = ~new_new_n57376__ & ~new_new_n57377__;
  assign new_new_n57379__ = new_new_n57375__ & new_new_n57378__;
  assign new_new_n57380__ = new_new_n57372__ & new_new_n57379__;
  assign new_new_n57381__ = ~new_new_n57365__ & ~new_new_n57380__;
  assign new_new_n57382__ = new_new_n52465__ & new_new_n57381__;
  assign new_new_n57383__ = ~new_new_n57339__ & new_new_n57382__;
  assign new_new_n57384__ = ~new_new_n57349__ & new_new_n57382__;
  assign new_new_n57385__ = ~new_new_n57383__ & ~new_new_n57384__;
  assign ys__n44155 = new_new_n57350__ | ~new_new_n57385__;
  assign new_new_n57387__ = ~new_new_n57349__ & new_new_n57383__;
  assign new_new_n57388__ = new_new_n57339__ & ~new_new_n57382__;
  assign new_new_n57389__ = ~new_new_n57349__ & new_new_n57388__;
  assign new_new_n57390__ = ~new_new_n57387__ & ~new_new_n57389__;
  assign new_new_n57391__ = ~new_new_n57339__ & ~new_new_n57382__;
  assign new_new_n57392__ = new_new_n57349__ & new_new_n57391__;
  assign new_new_n57393__ = new_new_n57339__ & new_new_n57382__;
  assign new_new_n57394__ = new_new_n57349__ & new_new_n57393__;
  assign new_new_n57395__ = ~new_new_n57392__ & ~new_new_n57394__;
  assign ys__n44160 = ~new_new_n57390__ | ~new_new_n57395__;
  assign new_new_n57397__ = ~new_new_n52465__ & new_new_n57381__;
  assign new_new_n57398__ = new_new_n52465__ & ~new_new_n57381__;
  assign new_new_n57399__ = ~new_new_n57397__ & ~new_new_n57398__;
  assign new_new_n57400__ = ~new_new_n57327__ & new_new_n57336__;
  assign new_new_n57401__ = new_new_n57312__ & new_new_n57335__;
  assign new_new_n57402__ = ~new_new_n57327__ & new_new_n57401__;
  assign new_new_n57403__ = ~new_new_n57400__ & ~new_new_n57402__;
  assign new_new_n57404__ = ~new_new_n57312__ & new_new_n57335__;
  assign new_new_n57405__ = new_new_n57327__ & new_new_n57404__;
  assign new_new_n57406__ = new_new_n57312__ & ~new_new_n57335__;
  assign new_new_n57407__ = new_new_n57327__ & new_new_n57406__;
  assign new_new_n57408__ = ~new_new_n57405__ & ~new_new_n57407__;
  assign new_new_n57409__ = new_new_n57403__ & new_new_n57408__;
  assign ys__n44183 = ~new_new_n57399__ & ~new_new_n57409__;
  assign new_new_n57411__ = new_new_n57399__ & ~new_new_n57409__;
  assign new_new_n57412__ = ~new_new_n57399__ & new_new_n57409__;
  assign ys__n44186 = new_new_n57411__ | new_new_n57412__;
  assign new_new_n57414__ = ys__n24744 & new_new_n52417__;
  assign new_new_n57415__ = ys__n24741 & new_new_n52420__;
  assign new_new_n57416__ = ~new_new_n57414__ & ~new_new_n57415__;
  assign new_new_n57417__ = ys__n39718 & new_new_n52409__;
  assign new_new_n57418__ = ys__n24741 & new_new_n52412__;
  assign new_new_n57419__ = ~new_new_n57417__ & ~new_new_n57418__;
  assign new_new_n57420__ = ys__n33681 & new_new_n52425__;
  assign new_new_n57421__ = ~ys__n33681 & new_new_n52428__;
  assign new_new_n57422__ = ~new_new_n57420__ & ~new_new_n57421__;
  assign new_new_n57423__ = new_new_n57419__ & new_new_n57422__;
  assign new_new_n57424__ = new_new_n57416__ & new_new_n57423__;
  assign new_new_n57425__ = ys__n39722 & new_new_n52301__;
  assign new_new_n57426__ = ys__n39720 & new_new_n52304__;
  assign new_new_n57427__ = ~new_new_n57425__ & ~new_new_n57426__;
  assign new_new_n57428__ = ys__n33687 & new_new_n52308__;
  assign new_new_n57429__ = ~ys__n33687 & new_new_n52311__;
  assign new_new_n57430__ = ~new_new_n57428__ & ~new_new_n57429__;
  assign new_new_n57431__ = new_new_n57427__ & new_new_n57430__;
  assign new_new_n57432__ = ys__n24753 & new_new_n52316__;
  assign new_new_n57433__ = ys__n24750 & new_new_n52318__;
  assign new_new_n57434__ = ~new_new_n57432__ & ~new_new_n57433__;
  assign new_new_n57435__ = ys__n24747 & new_new_n52322__;
  assign new_new_n57436__ = ys__n39724 & new_new_n52324__;
  assign new_new_n57437__ = ~new_new_n57435__ & ~new_new_n57436__;
  assign new_new_n57438__ = new_new_n57434__ & new_new_n57437__;
  assign new_new_n57439__ = new_new_n57431__ & new_new_n57438__;
  assign new_new_n57440__ = ~new_new_n57424__ & ~new_new_n57439__;
  assign new_new_n57441__ = new_new_n57365__ & ~new_new_n57380__;
  assign new_new_n57442__ = ~new_new_n57365__ & new_new_n57380__;
  assign new_new_n57443__ = ~new_new_n57441__ & ~new_new_n57442__;
  assign ys__n44189 = new_new_n57440__ & ~new_new_n57443__;
  assign new_new_n57445__ = ~new_new_n57440__ & ~new_new_n57443__;
  assign new_new_n57446__ = new_new_n57440__ & new_new_n57443__;
  assign ys__n44192 = new_new_n57445__ | new_new_n57446__;
  assign new_new_n57448__ = ys__n24741 & new_new_n52417__;
  assign new_new_n57449__ = ys__n24741 & new_new_n52409__;
  assign new_new_n57450__ = ~new_new_n57448__ & ~new_new_n57449__;
  assign new_new_n57451__ = ys__n24741 & new_new_n52425__;
  assign new_new_n57452__ = ~ys__n24741 & new_new_n52428__;
  assign new_new_n57453__ = ~new_new_n57451__ & ~new_new_n57452__;
  assign new_new_n57454__ = new_new_n57450__ & new_new_n57453__;
  assign new_new_n57455__ = ys__n39720 & new_new_n52301__;
  assign new_new_n57456__ = ys__n39718 & new_new_n52304__;
  assign new_new_n57457__ = ~new_new_n57455__ & ~new_new_n57456__;
  assign new_new_n57458__ = ys__n33685 & new_new_n52308__;
  assign new_new_n57459__ = ~ys__n33685 & new_new_n52311__;
  assign new_new_n57460__ = ~new_new_n57458__ & ~new_new_n57459__;
  assign new_new_n57461__ = new_new_n57457__ & new_new_n57460__;
  assign new_new_n57462__ = ys__n24750 & new_new_n52316__;
  assign new_new_n57463__ = ys__n24747 & new_new_n52318__;
  assign new_new_n57464__ = ~new_new_n57462__ & ~new_new_n57463__;
  assign new_new_n57465__ = ys__n24744 & new_new_n52322__;
  assign new_new_n57466__ = ys__n39722 & new_new_n52324__;
  assign new_new_n57467__ = ~new_new_n57465__ & ~new_new_n57466__;
  assign new_new_n57468__ = new_new_n57464__ & new_new_n57467__;
  assign new_new_n57469__ = new_new_n57461__ & new_new_n57468__;
  assign new_new_n57470__ = ~new_new_n57454__ & ~new_new_n57469__;
  assign new_new_n57471__ = new_new_n52428__ & ~new_new_n57454__;
  assign new_new_n57472__ = new_new_n52428__ & ~new_new_n57469__;
  assign new_new_n57473__ = ~new_new_n57471__ & ~new_new_n57472__;
  assign new_new_n57474__ = ~new_new_n57470__ & new_new_n57473__;
  assign new_new_n57475__ = new_new_n57424__ & ~new_new_n57439__;
  assign new_new_n57476__ = ~new_new_n57424__ & new_new_n57439__;
  assign new_new_n57477__ = ~new_new_n57475__ & ~new_new_n57476__;
  assign ys__n44195 = ~new_new_n57474__ & ~new_new_n57477__;
  assign new_new_n57479__ = new_new_n57474__ & ~new_new_n57477__;
  assign new_new_n57480__ = ~new_new_n57474__ & new_new_n57477__;
  assign ys__n44198 = new_new_n57479__ | new_new_n57480__;
  assign new_new_n57482__ = ~new_new_n57469__ & new_new_n57471__;
  assign new_new_n57483__ = ~new_new_n52428__ & new_new_n57454__;
  assign new_new_n57484__ = ~new_new_n57469__ & new_new_n57483__;
  assign new_new_n57485__ = ~new_new_n57482__ & ~new_new_n57484__;
  assign new_new_n57486__ = ~new_new_n52428__ & ~new_new_n57454__;
  assign new_new_n57487__ = new_new_n57469__ & new_new_n57486__;
  assign new_new_n57488__ = new_new_n52428__ & new_new_n57454__;
  assign new_new_n57489__ = new_new_n57469__ & new_new_n57488__;
  assign new_new_n57490__ = ~new_new_n57487__ & ~new_new_n57489__;
  assign ys__n44205 = ~new_new_n57485__ | ~new_new_n57490__;
  assign new_new_n57492__ = ys__n24741 & new_new_n52316__;
  assign new_new_n57493__ = ys__n24741 & new_new_n52324__;
  assign new_new_n57494__ = ~new_new_n57492__ & ~new_new_n57493__;
  assign new_new_n57495__ = ys__n24741 & new_new_n52308__;
  assign new_new_n57496__ = ~ys__n24741 & new_new_n52311__;
  assign new_new_n57497__ = ~new_new_n57495__ & ~new_new_n57496__;
  assign new_new_n57498__ = new_new_n57494__ & new_new_n57497__;
  assign new_new_n57499__ = new_new_n52311__ & ~new_new_n57498__;
  assign new_new_n57500__ = ys__n24744 & new_new_n52316__;
  assign new_new_n57501__ = ys__n24741 & new_new_n52318__;
  assign new_new_n57502__ = ~new_new_n57500__ & ~new_new_n57501__;
  assign new_new_n57503__ = ys__n39718 & new_new_n52324__;
  assign new_new_n57504__ = ys__n24741 & new_new_n52301__;
  assign new_new_n57505__ = ~new_new_n57503__ & ~new_new_n57504__;
  assign new_new_n57506__ = ys__n33681 & new_new_n52308__;
  assign new_new_n57507__ = ~ys__n33681 & new_new_n52311__;
  assign new_new_n57508__ = ~new_new_n57506__ & ~new_new_n57507__;
  assign new_new_n57509__ = new_new_n57505__ & new_new_n57508__;
  assign new_new_n57510__ = new_new_n57502__ & new_new_n57509__;
  assign ys__n44213 = new_new_n57499__ & ~new_new_n57510__;
  assign new_new_n57512__ = ~new_new_n57499__ & ~new_new_n57510__;
  assign new_new_n57513__ = new_new_n57499__ & new_new_n57510__;
  assign ys__n44216 = new_new_n57512__ | new_new_n57513__;
  assign new_new_n57515__ = ~new_new_n52311__ & ~new_new_n57498__;
  assign new_new_n57516__ = new_new_n52311__ & new_new_n57498__;
  assign ys__n44219 = new_new_n57515__ | new_new_n57516__;
  assign new_new_n57518__ = new_new_n12338__ & new_new_n12607__;
  assign new_new_n57519__ = ys__n948 & new_new_n57518__;
  assign ys__n44838 = ys__n44836 | new_new_n57519__;
  assign ys__n44841 = ys__n44840 & ~ys__n4566;
  assign ys__n44843 = ys__n44842 & ~ys__n4566;
  assign new_new_n57523__ = ys__n160 & ys__n344;
  assign new_new_n57524__ = ys__n352 & new_new_n57523__;
  assign new_new_n57525__ = new_new_n12600__ & new_new_n57524__;
  assign new_new_n57526__ = new_new_n12349__ & new_new_n57525__;
  assign new_new_n57527__ = new_new_n41396__ & ~new_new_n57526__;
  assign ys__n44844 = ys__n948 & ~new_new_n57527__;
  assign ys__n44845 = ys__n948 & ~new_new_n51829__;
  assign new_new_n57530__ = new_new_n12592__ & new_new_n51817__;
  assign new_new_n57531__ = new_new_n51819__ & new_new_n57530__;
  assign new_new_n57532__ = new_new_n51821__ & new_new_n57530__;
  assign new_new_n57533__ = ~new_new_n57531__ & ~new_new_n57532__;
  assign new_new_n57534__ = new_new_n12598__ & new_new_n57530__;
  assign new_new_n57535__ = ys__n352 & new_new_n51825__;
  assign new_new_n57536__ = new_new_n57530__ & new_new_n57535__;
  assign new_new_n57537__ = ~new_new_n57534__ & ~new_new_n57536__;
  assign new_new_n57538__ = new_new_n57533__ & new_new_n57537__;
  assign ys__n44846 = ys__n948 & ~new_new_n57538__;
  assign ys__n44848 = ys__n44847 & ~ys__n4566;
  assign ys__n44850 = ys__n44849 & ~ys__n4566;
  assign new_new_n57542__ = new_new_n12604__ & new_new_n51830__;
  assign new_new_n57543__ = ~new_new_n41395__ & ~new_new_n51822__;
  assign new_new_n57544__ = ~new_new_n51827__ & ~new_new_n57532__;
  assign new_new_n57545__ = ~new_new_n57536__ & new_new_n57544__;
  assign new_new_n57546__ = new_new_n57543__ & new_new_n57545__;
  assign new_new_n57547__ = new_new_n57542__ & new_new_n57546__;
  assign new_new_n57548__ = ~new_new_n41394__ & ~new_new_n51820__;
  assign new_new_n57549__ = ~new_new_n51824__ & ~new_new_n57531__;
  assign new_new_n57550__ = ~new_new_n57534__ & new_new_n57549__;
  assign new_new_n57551__ = new_new_n57548__ & new_new_n57550__;
  assign new_new_n57552__ = new_new_n57547__ & new_new_n57551__;
  assign new_new_n57553__ = ~new_new_n57547__ & ~new_new_n57552__;
  assign ys__n44851 = ys__n948 & new_new_n57553__;
  assign new_new_n57555__ = new_new_n57542__ & new_new_n57551__;
  assign new_new_n57556__ = ~new_new_n57552__ & ~new_new_n57555__;
  assign ys__n44852 = ys__n948 & new_new_n57556__;
  assign ys__n44853 = ys__n948 & ~new_new_n41390__;
  assign new_new_n57559__ = ~new_new_n51822__ & ~new_new_n57532__;
  assign new_new_n57560__ = ~new_new_n51820__ & ~new_new_n57531__;
  assign new_new_n57561__ = new_new_n41390__ & new_new_n57560__;
  assign new_new_n57562__ = new_new_n57559__ & new_new_n57561__;
  assign new_new_n57563__ = ys__n948 & ~new_new_n57559__;
  assign ys__n44854 = ~new_new_n57562__ & new_new_n57563__;
  assign new_new_n57565__ = ys__n948 & ~new_new_n57561__;
  assign ys__n44855 = ~new_new_n57562__ & new_new_n57565__;
  assign new_new_n57567__ = ys__n152 & ~ys__n158;
  assign new_new_n57568__ = ys__n148 & new_new_n41374__;
  assign new_new_n57569__ = new_new_n57567__ & new_new_n57568__;
  assign new_new_n57570__ = new_new_n41370__ & new_new_n57568__;
  assign new_new_n57571__ = ~new_new_n57569__ & ~new_new_n57570__;
  assign new_new_n57572__ = new_new_n41380__ & new_new_n57571__;
  assign new_new_n57573__ = new_new_n41373__ & new_new_n57572__;
  assign new_new_n57574__ = ~new_new_n41369__ & new_new_n57572__;
  assign new_new_n57575__ = ~ys__n30837 & ~new_new_n57574__;
  assign new_new_n57576__ = ~new_new_n57573__ & new_new_n57575__;
  assign new_new_n57577__ = ~new_new_n41372__ & new_new_n57572__;
  assign new_new_n57578__ = ~ys__n30837 & ~new_new_n57573__;
  assign new_new_n57579__ = ~new_new_n57577__ & new_new_n57578__;
  assign new_new_n57580__ = ~new_new_n57576__ & ~new_new_n57579__;
  assign new_new_n57581__ = ~ys__n4839 & ~ys__n4840;
  assign new_new_n57582__ = ~ys__n402 & ~new_new_n16247__;
  assign new_new_n57583__ = new_new_n16268__ & new_new_n57582__;
  assign new_new_n57584__ = new_new_n57581__ & ~new_new_n57583__;
  assign new_new_n57585__ = ~new_new_n57580__ & new_new_n57584__;
  assign new_new_n57586__ = new_new_n57556__ & new_new_n57576__;
  assign new_new_n57587__ = new_new_n57553__ & new_new_n57579__;
  assign new_new_n57588__ = ~new_new_n57586__ & ~new_new_n57587__;
  assign new_new_n57589__ = new_new_n51832__ & ~new_new_n57518__;
  assign new_new_n57590__ = ~new_new_n57588__ & ~new_new_n57589__;
  assign new_new_n57591__ = ~new_new_n57585__ & ~new_new_n57590__;
  assign new_new_n57592__ = ys__n948 & ~new_new_n57591__;
  assign new_new_n57593__ = new_new_n41367__ & new_new_n41375__;
  assign new_new_n57594__ = ys__n148 & new_new_n57593__;
  assign new_new_n57595__ = new_new_n41367__ & new_new_n57567__;
  assign new_new_n57596__ = ys__n148 & new_new_n57595__;
  assign new_new_n57597__ = ~new_new_n57594__ & ~new_new_n57596__;
  assign new_new_n57598__ = ~ys__n30837 & new_new_n57596__;
  assign new_new_n57599__ = ~new_new_n57597__ & new_new_n57598__;
  assign new_new_n57600__ = new_new_n57553__ & new_new_n57599__;
  assign new_new_n57601__ = ~ys__n30837 & new_new_n57594__;
  assign new_new_n57602__ = ~new_new_n57597__ & new_new_n57601__;
  assign new_new_n57603__ = new_new_n57556__ & new_new_n57602__;
  assign new_new_n57604__ = ~new_new_n57599__ & ~new_new_n57602__;
  assign new_new_n57605__ = ~new_new_n57583__ & ~new_new_n57604__;
  assign new_new_n57606__ = new_new_n57581__ & new_new_n57605__;
  assign new_new_n57607__ = ys__n30820 & new_new_n57602__;
  assign new_new_n57608__ = ys__n30819 & new_new_n57599__;
  assign new_new_n57609__ = ~new_new_n57607__ & ~new_new_n57608__;
  assign new_new_n57610__ = ys__n2779 & ~new_new_n57609__;
  assign new_new_n57611__ = ys__n44849 & new_new_n57602__;
  assign new_new_n57612__ = ys__n44847 & new_new_n57599__;
  assign new_new_n57613__ = ~new_new_n57611__ & ~new_new_n57612__;
  assign new_new_n57614__ = ~new_new_n57610__ & new_new_n57613__;
  assign new_new_n57615__ = ~new_new_n57606__ & new_new_n57614__;
  assign new_new_n57616__ = ~new_new_n57603__ & new_new_n57615__;
  assign new_new_n57617__ = ~new_new_n57600__ & new_new_n57616__;
  assign new_new_n57618__ = ys__n948 & ~new_new_n57617__;
  assign new_new_n57619__ = new_new_n16267__ & new_new_n41402__;
  assign new_new_n57620__ = new_new_n41390__ & new_new_n57619__;
  assign new_new_n57621__ = new_new_n57551__ & new_new_n57620__;
  assign new_new_n57622__ = new_new_n57546__ & new_new_n57551__;
  assign new_new_n57623__ = new_new_n57620__ & new_new_n57622__;
  assign new_new_n57624__ = ~new_new_n57621__ & ~new_new_n57623__;
  assign new_new_n57625__ = new_new_n57546__ & new_new_n57620__;
  assign new_new_n57626__ = ~new_new_n57623__ & ~new_new_n57625__;
  assign new_new_n57627__ = ~new_new_n57624__ & ~new_new_n57626__;
  assign new_new_n57628__ = ~ys__n4836 & ~ys__n4837;
  assign new_new_n57629__ = ~new_new_n57582__ & new_new_n57628__;
  assign new_new_n57630__ = ~ys__n4566 & ys__n30832;
  assign new_new_n57631__ = new_new_n57629__ & new_new_n57630__;
  assign new_new_n57632__ = ~new_new_n57627__ & new_new_n57631__;
  assign new_new_n57633__ = new_new_n12342__ & new_new_n41391__;
  assign new_new_n57634__ = new_new_n12342__ & new_new_n41384__;
  assign new_new_n57635__ = ~new_new_n57633__ & ~new_new_n57634__;
  assign new_new_n57636__ = new_new_n57633__ & ~new_new_n57635__;
  assign new_new_n57637__ = ys__n30819 & new_new_n57636__;
  assign new_new_n57638__ = new_new_n57634__ & ~new_new_n57635__;
  assign new_new_n57639__ = ys__n30820 & new_new_n57638__;
  assign new_new_n57640__ = ~new_new_n57637__ & ~new_new_n57639__;
  assign new_new_n57641__ = ys__n2779 & ~new_new_n57640__;
  assign new_new_n57642__ = ~new_new_n57636__ & ~new_new_n57638__;
  assign new_new_n57643__ = new_new_n57629__ & ~new_new_n57642__;
  assign new_new_n57644__ = ys__n44847 & new_new_n57636__;
  assign new_new_n57645__ = ys__n44849 & new_new_n57638__;
  assign new_new_n57646__ = ~new_new_n57644__ & ~new_new_n57645__;
  assign new_new_n57647__ = ~new_new_n57643__ & new_new_n57646__;
  assign new_new_n57648__ = ~new_new_n57641__ & new_new_n57647__;
  assign new_new_n57649__ = new_new_n57630__ & ~new_new_n57648__;
  assign new_new_n57650__ = ~new_new_n57582__ & new_new_n57630__;
  assign new_new_n57651__ = ~new_new_n16268__ & new_new_n57650__;
  assign new_new_n57652__ = ~ys__n30837 & ~new_new_n57571__;
  assign new_new_n57653__ = ~ys__n4566 & new_new_n57652__;
  assign new_new_n57654__ = ~ys__n30832 & new_new_n57653__;
  assign new_new_n57655__ = ~new_new_n57583__ & new_new_n57654__;
  assign new_new_n57656__ = new_new_n41383__ & ~new_new_n51832__;
  assign new_new_n57657__ = ~new_new_n57655__ & ~new_new_n57656__;
  assign new_new_n57658__ = ~new_new_n57651__ & new_new_n57657__;
  assign new_new_n57659__ = ~new_new_n57649__ & new_new_n57658__;
  assign new_new_n57660__ = ~new_new_n57632__ & new_new_n57659__;
  assign new_new_n57661__ = ~new_new_n57618__ & new_new_n57660__;
  assign ys__n44858 = new_new_n57592__ | ~new_new_n57661__;
  assign ys__n44948 = ~ys__n4566 & new_new_n57599__;
  assign ys__n44949 = ~ys__n4566 & new_new_n57602__;
  assign new_new_n57665__ = new_new_n41373__ & new_new_n57597__;
  assign new_new_n57666__ = new_new_n57572__ & new_new_n57665__;
  assign new_new_n57667__ = ~ys__n30837 & ~ys__n30832;
  assign new_new_n57668__ = ~new_new_n57666__ & new_new_n57667__;
  assign new_new_n57669__ = ys__n352 & ys__n30832;
  assign new_new_n57670__ = ~new_new_n57668__ & ~new_new_n57669__;
  assign ys__n44950 = ~ys__n4566 & ~new_new_n57670__;
  assign new_new_n57672__ = ~ys__n22792 & ys__n38927;
  assign ys__n44985 = ys__n46954 & new_new_n57672__;
  assign new_new_n57674__ = ~ys__n38236 & ~ys__n38237;
  assign new_new_n57675__ = ~ys__n33364 & ~new_new_n57674__;
  assign ys__n44987 = new_new_n13884__ & new_new_n57675__;
  assign new_new_n57677__ = ~new_new_n51119__ & new_new_n51127__;
  assign ys__n46131 = ys__n46130 | new_new_n57677__;
  assign new_new_n57679__ = ~new_new_n51119__ & new_new_n51126__;
  assign ys__n46133 = ys__n46132 | new_new_n57679__;
  assign new_new_n57681__ = ~new_new_n51119__ & new_new_n51124__;
  assign ys__n46135 = ys__n46134 | new_new_n57681__;
  assign new_new_n57683__ = ~new_new_n51119__ & new_new_n51123__;
  assign ys__n46137 = ys__n46136 | new_new_n57683__;
  assign new_new_n57685__ = ~ys__n35028 & ys__n26573;
  assign new_new_n57686__ = ~ys__n30863 & ~new_new_n57685__;
  assign new_new_n57687__ = ~ys__n46141 & ys__n46142;
  assign new_new_n57688__ = ys__n46141 & ~ys__n46142;
  assign new_new_n57689__ = ~new_new_n57687__ & ~new_new_n57688__;
  assign ys__n46143 = ~new_new_n57686__ & new_new_n57689__;
  assign new_new_n57691__ = ~ys__n34988 & ys__n26555;
  assign new_new_n57692__ = ~ys__n34966 & new_new_n57691__;
  assign new_new_n57693__ = ys__n34966 & ~new_new_n57691__;
  assign ys__n46146 = new_new_n57692__ | new_new_n57693__;
  assign new_new_n57695__ = ys__n18317 & ~new_new_n32347__;
  assign ys__n46159 = ~ys__n34962 & new_new_n57695__;
  assign new_new_n57697__ = ~ys__n35033 & ys__n46159;
  assign new_new_n57698__ = ~ys__n35047 & ~new_new_n57697__;
  assign new_new_n57699__ = ~ys__n46152 & ys__n46153;
  assign new_new_n57700__ = ys__n46152 & ~ys__n46153;
  assign new_new_n57701__ = ~new_new_n57699__ & ~new_new_n57700__;
  assign ys__n46154 = ~new_new_n57698__ & new_new_n57701__;
  assign new_new_n57703__ = ys__n46150 & ~ys__n46151;
  assign new_new_n57704__ = ~ys__n46150 & ys__n46151;
  assign new_new_n57705__ = ~ys__n26565 & ~new_new_n57704__;
  assign new_new_n57706__ = ~new_new_n57703__ & new_new_n57705__;
  assign new_new_n57707__ = ~ys__n30941 & ~ys__n35031;
  assign ys__n46163 = ~ys__n26291 & new_new_n57707__;
  assign new_new_n57709__ = ~ys__n34976 & ys__n46163;
  assign ys__n46155 = ~new_new_n57706__ & ~new_new_n57709__;
  assign new_new_n57711__ = ~ys__n34972 & new_new_n57697__;
  assign new_new_n57712__ = ys__n34972 & ~new_new_n57697__;
  assign ys__n46158 = new_new_n57711__ | new_new_n57712__;
  assign new_new_n57714__ = ~ys__n34978 & new_new_n57709__;
  assign new_new_n57715__ = ys__n34978 & ~new_new_n57709__;
  assign ys__n46162 = new_new_n57714__ | new_new_n57715__;
  assign new_new_n57717__ = ~ys__n35035 & ys__n26288;
  assign new_new_n57718__ = ~ys__n26561 & ~new_new_n57717__;
  assign new_new_n57719__ = ~ys__n46170 & ys__n46171;
  assign new_new_n57720__ = ys__n46170 & ~ys__n46171;
  assign new_new_n57721__ = ~new_new_n57719__ & ~new_new_n57720__;
  assign ys__n46172 = ~new_new_n57718__ & new_new_n57721__;
  assign new_new_n57723__ = ys__n46168 & ~ys__n46169;
  assign new_new_n57724__ = ~ys__n46168 & ys__n46169;
  assign new_new_n57725__ = ~ys__n46166 & ~new_new_n57724__;
  assign new_new_n57726__ = ~new_new_n57723__ & new_new_n57725__;
  assign ys__n46173 = ~new_new_n57691__ & ~new_new_n57726__;
  assign new_new_n57728__ = ~ys__n34984 & new_new_n57717__;
  assign new_new_n57729__ = ys__n34984 & ~new_new_n57717__;
  assign ys__n46176 = new_new_n57728__ | new_new_n57729__;
  assign new_new_n57731__ = ~ys__n34990 & new_new_n57691__;
  assign new_new_n57732__ = ys__n34990 & ~new_new_n57691__;
  assign ys__n46179 = new_new_n57731__ | new_new_n57732__;
  assign new_new_n57734__ = ~ys__n35037 & ys__n26294;
  assign new_new_n57735__ = ~ys__n46180 & ~new_new_n57734__;
  assign new_new_n57736__ = ~ys__n46186 & ys__n46187;
  assign new_new_n57737__ = ys__n46186 & ~ys__n46187;
  assign new_new_n57738__ = ~new_new_n57736__ & ~new_new_n57737__;
  assign ys__n46188 = ~new_new_n57735__ & new_new_n57738__;
  assign new_new_n57740__ = ys__n46184 & ~ys__n46185;
  assign new_new_n57741__ = ~ys__n46184 & ys__n46185;
  assign new_new_n57742__ = ~ys__n26553 & ~new_new_n57741__;
  assign new_new_n57743__ = ~new_new_n57740__ & new_new_n57742__;
  assign new_new_n57744__ = ~ys__n35000 & ys__n26282;
  assign ys__n46189 = ~new_new_n57743__ & ~new_new_n57744__;
  assign new_new_n57746__ = ~ys__n34996 & new_new_n57734__;
  assign new_new_n57747__ = ys__n34996 & ~new_new_n57734__;
  assign ys__n46192 = new_new_n57746__ | new_new_n57747__;
  assign new_new_n57749__ = ~ys__n35002 & new_new_n57744__;
  assign new_new_n57750__ = ys__n35002 & ~new_new_n57744__;
  assign ys__n46195 = new_new_n57749__ | new_new_n57750__;
  assign new_new_n57752__ = ~ys__n35039 & ys__n26284;
  assign new_new_n57753__ = ~ys__n26554 & ~new_new_n57752__;
  assign new_new_n57754__ = ~ys__n46202 & ys__n46203;
  assign new_new_n57755__ = ys__n46202 & ~ys__n46203;
  assign new_new_n57756__ = ~new_new_n57754__ & ~new_new_n57755__;
  assign ys__n46204 = ~new_new_n57753__ & new_new_n57756__;
  assign new_new_n57758__ = ys__n46200 & ~ys__n46201;
  assign new_new_n57759__ = ~ys__n46200 & ys__n46201;
  assign new_new_n57760__ = ~ys__n46198 & ~new_new_n57759__;
  assign new_new_n57761__ = ~new_new_n57758__ & new_new_n57760__;
  assign new_new_n57762__ = ~ys__n35012 & ys__n26293;
  assign ys__n46205 = ~new_new_n57761__ & ~new_new_n57762__;
  assign new_new_n57764__ = ~ys__n35008 & new_new_n57752__;
  assign new_new_n57765__ = ys__n35008 & ~new_new_n57752__;
  assign ys__n46208 = new_new_n57764__ | new_new_n57765__;
  assign new_new_n57767__ = ~ys__n35014 & new_new_n57762__;
  assign new_new_n57768__ = ys__n35014 & ~new_new_n57762__;
  assign ys__n46211 = new_new_n57767__ | new_new_n57768__;
  assign new_new_n57770__ = ~ys__n35041 & ys__n26286;
  assign new_new_n57771__ = ~ys__n26560 & ~new_new_n57770__;
  assign new_new_n57772__ = ~ys__n46218 & ys__n46219;
  assign new_new_n57773__ = ys__n46218 & ~ys__n46219;
  assign new_new_n57774__ = ~new_new_n57772__ & ~new_new_n57773__;
  assign ys__n46220 = ~new_new_n57771__ & new_new_n57774__;
  assign new_new_n57776__ = ys__n46216 & ~ys__n46217;
  assign new_new_n57777__ = ~ys__n46216 & ys__n46217;
  assign new_new_n57778__ = ~ys__n46214 & ~new_new_n57777__;
  assign new_new_n57779__ = ~new_new_n57776__ & new_new_n57778__;
  assign new_new_n57780__ = ~ys__n35024 & ys__n37738;
  assign ys__n46221 = ~new_new_n57779__ & ~new_new_n57780__;
  assign new_new_n57782__ = ~ys__n35020 & new_new_n57770__;
  assign new_new_n57783__ = ys__n35020 & ~new_new_n57770__;
  assign ys__n46224 = new_new_n57782__ | new_new_n57783__;
  assign new_new_n57785__ = ~ys__n35026 & new_new_n57780__;
  assign new_new_n57786__ = ys__n35026 & ~new_new_n57780__;
  assign ys__n46227 = new_new_n57785__ | new_new_n57786__;
  assign ys__n46233 = ~ys__n26562 & ys__n26563;
  assign new_new_n57789__ = ~ys__n25470 & ys__n30863;
  assign ys__n46234 = ys__n46166 | new_new_n57789__;
  assign new_new_n57791__ = ys__n312 & ~ys__n622;
  assign new_new_n57792__ = ~ys__n312 & ys__n622;
  assign ys__n48339 = new_new_n57791__ | new_new_n57792__;
  assign new_new_n57794__ = ~ys__n620 & new_new_n16490__;
  assign new_new_n57795__ = ys__n620 & ~new_new_n16490__;
  assign ys__n48340 = new_new_n57794__ | new_new_n57795__;
  assign new_new_n57797__ = ys__n620 & new_new_n16490__;
  assign new_new_n57798__ = ~ys__n618 & new_new_n57797__;
  assign new_new_n57799__ = ys__n618 & ~new_new_n57797__;
  assign ys__n48341 = new_new_n57798__ | new_new_n57799__;
  assign new_new_n57801__ = ~ys__n614 & new_new_n16492__;
  assign new_new_n57802__ = ys__n614 & ~new_new_n16492__;
  assign ys__n48342 = new_new_n57801__ | new_new_n57802__;
  assign new_new_n57804__ = ys__n614 & new_new_n16492__;
  assign new_new_n57805__ = ~ys__n612 & new_new_n57804__;
  assign new_new_n57806__ = ys__n612 & ~new_new_n57804__;
  assign ys__n48343 = new_new_n57805__ | new_new_n57806__;
  assign new_new_n57808__ = new_new_n16492__ & new_new_n16493__;
  assign new_new_n57809__ = ~ys__n616 & new_new_n57808__;
  assign new_new_n57810__ = ys__n616 & ~new_new_n57808__;
  assign ys__n48344 = new_new_n57809__ | new_new_n57810__;
  assign new_new_n57812__ = new_new_n40673__ & new_new_n40689__;
  assign new_new_n57813__ = ~new_new_n40673__ & ~new_new_n40689__;
  assign ys__n48349 = new_new_n57812__ | new_new_n57813__;
  assign new_new_n57815__ = ~new_new_n40673__ & new_new_n40689__;
  assign new_new_n57816__ = ~new_new_n40693__ & ~new_new_n57815__;
  assign new_new_n57817__ = new_new_n40682__ & ~new_new_n57816__;
  assign new_new_n57818__ = ~new_new_n40682__ & new_new_n57816__;
  assign ys__n48350 = new_new_n57817__ | new_new_n57818__;
  assign new_new_n57820__ = ~new_new_n40696__ & new_new_n40733__;
  assign new_new_n57821__ = new_new_n40696__ & ~new_new_n40733__;
  assign ys__n48351 = new_new_n57820__ | new_new_n57821__;
  assign new_new_n57823__ = ~new_new_n40696__ & ~new_new_n40733__;
  assign new_new_n57824__ = ~new_new_n40738__ & ~new_new_n57823__;
  assign new_new_n57825__ = new_new_n40730__ & ~new_new_n57824__;
  assign new_new_n57826__ = ~new_new_n40730__ & new_new_n57824__;
  assign ys__n48352 = new_new_n57825__ | new_new_n57826__;
  assign new_new_n57828__ = ~new_new_n40696__ & new_new_n40734__;
  assign new_new_n57829__ = new_new_n40740__ & ~new_new_n57828__;
  assign new_new_n57830__ = new_new_n40720__ & ~new_new_n57829__;
  assign new_new_n57831__ = ~new_new_n40720__ & new_new_n57829__;
  assign ys__n48353 = new_new_n57830__ | new_new_n57831__;
  assign new_new_n57833__ = ~new_new_n40720__ & ~new_new_n57829__;
  assign new_new_n57834__ = ~new_new_n40743__ & ~new_new_n57833__;
  assign new_new_n57835__ = new_new_n40711__ & ~new_new_n57834__;
  assign new_new_n57836__ = ~new_new_n40711__ & new_new_n57834__;
  assign ys__n48354 = new_new_n57835__ | new_new_n57836__;
  assign new_new_n57838__ = ~new_new_n40747__ & new_new_n40817__;
  assign new_new_n57839__ = new_new_n40747__ & ~new_new_n40817__;
  assign ys__n48355 = new_new_n57838__ | new_new_n57839__;
  assign new_new_n57841__ = ~new_new_n40747__ & ~new_new_n40817__;
  assign new_new_n57842__ = ~new_new_n40823__ & ~new_new_n57841__;
  assign new_new_n57843__ = new_new_n40814__ & ~new_new_n57842__;
  assign new_new_n57844__ = ~new_new_n40814__ & new_new_n57842__;
  assign ys__n48356 = new_new_n57843__ | new_new_n57844__;
  assign new_new_n57846__ = ~new_new_n40747__ & new_new_n40818__;
  assign new_new_n57847__ = new_new_n40825__ & ~new_new_n57846__;
  assign new_new_n57848__ = new_new_n40804__ & ~new_new_n57847__;
  assign new_new_n57849__ = ~new_new_n40804__ & new_new_n57847__;
  assign ys__n48357 = new_new_n57848__ | new_new_n57849__;
  assign new_new_n57851__ = ~new_new_n40804__ & ~new_new_n57847__;
  assign new_new_n57852__ = ~new_new_n40828__ & ~new_new_n57851__;
  assign new_new_n57853__ = new_new_n40795__ & ~new_new_n57852__;
  assign new_new_n57854__ = ~new_new_n40795__ & new_new_n57852__;
  assign ys__n48358 = new_new_n57853__ | new_new_n57854__;
  assign new_new_n57856__ = ~new_new_n40747__ & new_new_n40819__;
  assign new_new_n57857__ = new_new_n40831__ & ~new_new_n57856__;
  assign new_new_n57858__ = new_new_n40784__ & ~new_new_n57857__;
  assign new_new_n57859__ = ~new_new_n40784__ & new_new_n57857__;
  assign ys__n48359 = new_new_n57858__ | new_new_n57859__;
  assign new_new_n57861__ = ~new_new_n40784__ & ~new_new_n57857__;
  assign new_new_n57862__ = ~new_new_n40834__ & ~new_new_n57861__;
  assign new_new_n57863__ = new_new_n40775__ & ~new_new_n57862__;
  assign new_new_n57864__ = ~new_new_n40775__ & new_new_n57862__;
  assign ys__n48360 = new_new_n57863__ | new_new_n57864__;
  assign new_new_n57866__ = new_new_n40785__ & ~new_new_n57857__;
  assign new_new_n57867__ = new_new_n40836__ & ~new_new_n57866__;
  assign new_new_n57868__ = new_new_n40765__ & ~new_new_n57867__;
  assign new_new_n57869__ = ~new_new_n40765__ & new_new_n57867__;
  assign ys__n48361 = new_new_n57868__ | new_new_n57869__;
  assign new_new_n57871__ = ~new_new_n40765__ & ~new_new_n57867__;
  assign new_new_n57872__ = ~new_new_n40839__ & ~new_new_n57871__;
  assign new_new_n57873__ = new_new_n40756__ & ~new_new_n57872__;
  assign new_new_n57874__ = ~new_new_n40756__ & new_new_n57872__;
  assign ys__n48362 = new_new_n57873__ | new_new_n57874__;
  assign ys__n280 = ~ys__n20273;
  assign ys__n313 = ~ys__n312;
  assign ys__n319 = ~ys__n318;
  assign ys__n415 = ~ys__n414;
  assign ys__n417 = ~ys__n416;
  assign ys__n455 = ~ys__n454;
  assign ys__n457 = ~ys__n456;
  assign ys__n565 = ~ys__n564;
  assign ys__n890 = ~ys__n874;
  assign ys__n18131 = ~ys__n33515;
  assign ys__n18386 = ~ys__n33324;
  assign ys__n18391 = ~ys__n33317;
  assign ys__n23340 = ~ys__n28243;
  assign ys__n33420 = ~ys__n18121;
  assign ys__n33437 = ~ys__n33438;
  assign ys__n33439 = ~ys__n24177;
  assign ys__n33453 = ~ys__n33454;
  assign ys__n33456 = ~ys__n33455;
  assign ys__n33513 = ~ys__n33514;
  assign ys__n33535 = ~ys__n24590;
  assign ys__n4175 = ys__n738;
  assign ys__n28269 = ys__n23340;
  assign ys__n28334 = ys__n28276;
  assign ys__n38338 = ys__n38334;
  assign ys__n48348 = ys__n35144;
  assign ys__n33333 = ~ys__n33332;
  assign new_new_n98_9_ = ys__n29707 & ~ys__n29709;
  assign new_new_n99_9_ = ys__n29708 & ys__n29709;
  assign ys__n29710 = new_new_n98_9_ | new_new_n99_9_;
  assign new_new_n101_9_ = ~ys__n29709 & ys__n29711;
  assign new_new_n102_9_ = ys__n29709 & ys__n29712;
  assign ys__n29713 = new_new_n101_9_ | new_new_n102_9_;
  assign new_new_n104_9_ = ~ys__n29709 & ys__n29714;
  assign new_new_n105_9_ = ys__n29709 & ys__n29715;
  assign ys__n29716 = new_new_n104_9_ | new_new_n105_9_;
  assign new_new_n107_9_ = ~ys__n29709 & ys__n29717;
  assign new_new_n108_9_ = ys__n29709 & ys__n29718;
  assign ys__n29719 = new_new_n107_9_ | new_new_n108_9_;
  assign new_new_n110_9_ = ~ys__n29709 & ys__n29720;
  assign new_new_n111_9_ = ys__n29709 & ys__n29721;
  assign ys__n29722 = new_new_n110_9_ | new_new_n111_9_;
  assign new_new_n113_9_ = ~ys__n29709 & ys__n29723;
  assign new_new_n114_9_ = ys__n29709 & ys__n29724;
  assign ys__n29725 = new_new_n113_9_ | new_new_n114_9_;
  assign new_new_n116_9_ = ~ys__n29709 & ys__n29726;
  assign new_new_n117_9_ = ys__n29709 & ys__n29727;
  assign ys__n29728 = new_new_n116_9_ | new_new_n117_9_;
  assign new_new_n119_9_ = ~ys__n29709 & ys__n29729;
  assign new_new_n120_9_ = ys__n29709 & ys__n29730;
  assign ys__n29731 = new_new_n119_9_ | new_new_n120_9_;
  assign new_new_n122_9_ = ~ys__n29709 & ys__n29732;
  assign new_new_n123_9_ = ys__n29709 & ys__n29733;
  assign ys__n29734 = new_new_n122_9_ | new_new_n123_9_;
  assign new_new_n125_9_ = ~ys__n29709 & ys__n29735;
  assign new_new_n126_9_ = ys__n29709 & ys__n29736;
  assign ys__n29737 = new_new_n125_9_ | new_new_n126_9_;
  assign new_new_n128_9_ = ~ys__n29709 & ys__n29738;
  assign new_new_n129_9_ = ys__n29709 & ys__n29739;
  assign ys__n29740 = new_new_n128_9_ | new_new_n129_9_;
  assign new_new_n131_9_ = ~ys__n29709 & ys__n29741;
  assign new_new_n132_9_ = ys__n29709 & ys__n29742;
  assign ys__n29743 = new_new_n131_9_ | new_new_n132_9_;
  assign new_new_n134_9_ = ~ys__n29709 & ys__n29744;
  assign new_new_n135_9_ = ys__n29709 & ys__n29745;
  assign ys__n29746 = new_new_n134_9_ | new_new_n135_9_;
  assign new_new_n137_9_ = ~ys__n29709 & ys__n29747;
  assign new_new_n138_9_ = ys__n29709 & ys__n29748;
  assign ys__n29749 = new_new_n137_9_ | new_new_n138_9_;
  assign new_new_n140_9_ = ~ys__n29709 & ys__n29750;
  assign new_new_n141_9_ = ys__n29709 & ys__n29751;
  assign ys__n29752 = new_new_n140_9_ | new_new_n141_9_;
  assign new_new_n143_9_ = ~ys__n29709 & ys__n29753;
  assign new_new_n144_9_ = ys__n29709 & ys__n29754;
  assign ys__n29755 = new_new_n143_9_ | new_new_n144_9_;
  assign new_new_n146_9_ = ~ys__n29709 & ys__n29756;
  assign new_new_n147_9_ = ys__n29709 & ys__n29757;
  assign ys__n29758 = new_new_n146_9_ | new_new_n147_9_;
  assign new_new_n149_9_ = ~ys__n29709 & ys__n29759;
  assign new_new_n150_9_ = ys__n29709 & ys__n29760;
  assign ys__n29761 = new_new_n149_9_ | new_new_n150_9_;
  assign new_new_n152_9_ = ~ys__n29709 & ys__n29762;
  assign new_new_n153_9_ = ys__n29709 & ys__n29763;
  assign ys__n29764 = new_new_n152_9_ | new_new_n153_9_;
  assign new_new_n155_9_ = ~ys__n29709 & ys__n29765;
  assign new_new_n156_9_ = ys__n29709 & ys__n29766;
  assign ys__n29767 = new_new_n155_9_ | new_new_n156_9_;
  assign new_new_n158_9_ = ~ys__n29709 & ys__n29768;
  assign new_new_n159_9_ = ys__n29709 & ys__n29769;
  assign ys__n29770 = new_new_n158_9_ | new_new_n159_9_;
  assign new_new_n161_9_ = ~ys__n29709 & ys__n29771;
  assign new_new_n162_9_ = ys__n29709 & ys__n29772;
  assign ys__n29773 = new_new_n161_9_ | new_new_n162_9_;
  assign new_new_n164_9_ = ~ys__n29709 & ys__n29774;
  assign new_new_n165_9_ = ys__n29709 & ys__n29775;
  assign ys__n29776 = new_new_n164_9_ | new_new_n165_9_;
  assign new_new_n167_9_ = ~ys__n29709 & ys__n29777;
  assign new_new_n168_9_ = ys__n29709 & ys__n29778;
  assign ys__n29779 = new_new_n167_9_ | new_new_n168_9_;
  assign new_new_n170_9_ = ~ys__n29709 & ys__n29780;
  assign new_new_n171_9_ = ys__n29709 & ys__n29781;
  assign ys__n29782 = new_new_n170_9_ | new_new_n171_9_;
  assign new_new_n173_9_ = ~ys__n29709 & ys__n29783;
  assign new_new_n174_9_ = ys__n29709 & ys__n29784;
  assign ys__n29785 = new_new_n173_9_ | new_new_n174_9_;
  assign new_new_n176_9_ = ~ys__n29709 & ys__n29786;
  assign new_new_n177_9_ = ys__n29709 & ys__n29787;
  assign ys__n29788 = new_new_n176_9_ | new_new_n177_9_;
  assign new_new_n179_9_ = ~ys__n29709 & ys__n29789;
  assign new_new_n180_9_ = ys__n29709 & ys__n29790;
  assign ys__n29791 = new_new_n179_9_ | new_new_n180_9_;
  assign new_new_n182_9_ = ~ys__n29709 & ys__n29792;
  assign new_new_n183_9_ = ys__n29709 & ys__n29793;
  assign ys__n29794 = new_new_n182_9_ | new_new_n183_9_;
  assign new_new_n185_9_ = ~ys__n29709 & ys__n29795;
  assign new_new_n186_9_ = ys__n29709 & ys__n29796;
  assign ys__n29797 = new_new_n185_9_ | new_new_n186_9_;
  assign new_new_n188_9_ = ~ys__n29709 & ys__n29798;
  assign new_new_n189_9_ = ys__n29709 & ys__n29799;
  assign ys__n29800 = new_new_n188_9_ | new_new_n189_9_;
  assign new_new_n191_9_ = ~ys__n29709 & ys__n29801;
  assign new_new_n192_9_ = ys__n29709 & ys__n29802;
  assign ys__n29803 = new_new_n191_9_ | new_new_n192_9_;
  assign ys__n33339 = ~ys__n33338;
  assign ys__n264 = 1'b0;
  assign ys__n28247 = 1'b0;
  assign ys__n28249 = 1'b1;
  assign ys__n28250 = 1'b0;
  assign ys__n28251 = 1'b0;
  assign ys__n28252 = 1'b0;
  assign ys__n28254 = 1'b0;
  assign ys__n28256 = 1'b1;
  assign ys__n28259 = 1'b0;
  assign ys__n28261 = 1'b0;
  assign ys__n28263 = 1'b0;
  assign ys__n28265 = 1'b0;
  assign ys__n28266 = 1'b0;
  assign ys__n28268 = 1'b0;
  assign ys__n28270 = 1'b0;
  assign ys__n28271 = 1'b0;
  assign ys__n28272 = 1'b0;
  assign ys__n28274 = 1'b0;
  assign ys__n28858 = 1'b0;
  assign ys__n30836 = 1'b0;
  assign ys__n30856 = 1'b0;
  assign ys__n30858 = 1'b0;
  assign ys__n30860 = 1'b0;
  assign ys__n38185 = 1'b0;
  assign ys__n38186 = 1'b0;
  assign ys__n38188 = 1'b0;
  assign ys__n38191 = 1'b0;
endmodule


