// Benchmark "merged" written by ABC on Wed Sep  6 14:54:47 2023

module merged ( 
    ys__n14, ys__n16, ys__n22, ys__n24, ys__n26, ys__n28, ys__n30, ys__n32,
    ys__n34, ys__n36, ys__n38, ys__n40, ys__n42, ys__n44, ys__n46, ys__n48,
    ys__n50, ys__n52, ys__n54, ys__n56, ys__n58, ys__n60, ys__n62, ys__n66,
    ys__n70, ys__n72, ys__n74, ys__n76, ys__n78, ys__n80, ys__n82, ys__n84,
    ys__n86, ys__n88, ys__n90, ys__n96, ys__n98, ys__n100, ys__n108,
    ys__n110, ys__n112, ys__n114, ys__n116, ys__n118, ys__n120, ys__n122,
    ys__n124, ys__n126, ys__n128, ys__n130, ys__n132, ys__n134, ys__n136,
    ys__n138, ys__n140, ys__n142, ys__n148, ys__n150, ys__n152, ys__n156,
    ys__n158, ys__n160, ys__n162, ys__n164, ys__n166, ys__n168, ys__n170,
    ys__n172, ys__n174, ys__n176, ys__n178, ys__n182, ys__n184, ys__n186,
    ys__n190, ys__n192, ys__n194, ys__n196, ys__n198, ys__n202, ys__n204,
    ys__n206, ys__n208, ys__n210, ys__n212, ys__n214, ys__n216, ys__n218,
    ys__n220, ys__n222, ys__n226, ys__n232, ys__n238, ys__n240, ys__n242,
    ys__n244, ys__n248, ys__n256, ys__n258, ys__n262, ys__n290, ys__n294,
    ys__n296, ys__n298, ys__n300, ys__n302, ys__n304, ys__n306, ys__n308,
    ys__n310, ys__n312, ys__n314, ys__n316, ys__n318, ys__n326, ys__n328,
    ys__n330, ys__n332, ys__n336, ys__n338, ys__n340, ys__n342, ys__n344,
    ys__n346, ys__n348, ys__n350, ys__n352, ys__n354, ys__n356, ys__n358,
    ys__n360, ys__n362, ys__n364, ys__n366, ys__n368, ys__n370, ys__n372,
    ys__n374, ys__n376, ys__n378, ys__n380, ys__n382, ys__n384, ys__n386,
    ys__n392, ys__n394, ys__n396, ys__n398, ys__n402, ys__n408, ys__n414,
    ys__n416, ys__n418, ys__n420, ys__n422, ys__n424, ys__n426, ys__n428,
    ys__n430, ys__n432, ys__n434, ys__n436, ys__n438, ys__n440, ys__n442,
    ys__n444, ys__n446, ys__n448, ys__n450, ys__n452, ys__n454, ys__n456,
    ys__n464, ys__n488, ys__n490, ys__n500, ys__n504, ys__n512, ys__n514,
    ys__n516, ys__n518, ys__n520, ys__n522, ys__n524, ys__n526, ys__n528,
    ys__n530, ys__n532, ys__n536, ys__n538, ys__n544, ys__n546, ys__n548,
    ys__n550, ys__n556, ys__n558, ys__n562, ys__n564, ys__n566, ys__n568,
    ys__n570, ys__n572, ys__n580, ys__n582, ys__n584, ys__n586, ys__n588,
    ys__n598, ys__n600, ys__n602, ys__n604, ys__n606, ys__n608, ys__n610,
    ys__n612, ys__n614, ys__n616, ys__n618, ys__n620, ys__n622, ys__n624,
    ys__n626, ys__n632, ys__n634, ys__n636, ys__n638, ys__n640, ys__n642,
    ys__n644, ys__n646, ys__n648, ys__n650, ys__n652, ys__n654, ys__n656,
    ys__n658, ys__n660, ys__n662, ys__n664, ys__n666, ys__n668, ys__n670,
    ys__n672, ys__n674, ys__n676, ys__n678, ys__n680, ys__n682, ys__n684,
    ys__n686, ys__n688, ys__n690, ys__n692, ys__n694, ys__n696, ys__n698,
    ys__n700, ys__n702, ys__n704, ys__n706, ys__n708, ys__n710, ys__n712,
    ys__n718, ys__n720, ys__n722, ys__n724, ys__n726, ys__n728, ys__n736,
    ys__n742, ys__n744, ys__n746, ys__n748, ys__n750, ys__n752, ys__n758,
    ys__n760, ys__n762, ys__n764, ys__n766, ys__n768, ys__n770, ys__n772,
    ys__n774, ys__n776, ys__n778, ys__n780, ys__n782, ys__n784, ys__n816,
    ys__n818, ys__n820, ys__n822, ys__n824, ys__n826, ys__n828, ys__n830,
    ys__n832, ys__n834, ys__n836, ys__n838, ys__n840, ys__n842, ys__n844,
    ys__n846, ys__n848, ys__n850, ys__n852, ys__n854, ys__n856, ys__n858,
    ys__n860, ys__n874, ys__n889, ys__n935, ys__n1029, ys__n1036,
    ys__n1038, ys__n1048, ys__n1072, ys__n1076, ys__n1078, ys__n1084,
    ys__n1094, ys__n1098, ys__n1099, ys__n1106, ys__n1107, ys__n1109,
    ys__n1110, ys__n1116, ys__n1117, ys__n1119, ys__n1120, ys__n1129,
    ys__n1147, ys__n1151, ys__n1153, ys__n1154, ys__n1156, ys__n1157,
    ys__n1301, ys__n1309, ys__n1489, ys__n1490, ys__n1492, ys__n1493,
    ys__n1495, ys__n1496, ys__n1498, ys__n1499, ys__n1502, ys__n1503,
    ys__n1505, ys__n1506, ys__n1508, ys__n1509, ys__n1511, ys__n1535,
    ys__n2024, ys__n2233, ys__n2239, ys__n2245, ys__n2247, ys__n2251,
    ys__n2276, ys__n2282, ys__n2306, ys__n2308, ys__n2312, ys__n2427,
    ys__n2429, ys__n2433, ys__n2644, ys__n2652, ys__n2693, ys__n2716,
    ys__n2779, ys__n2830, ys__n2924, ys__n3214, ys__n4168, ys__n4176,
    ys__n4177, ys__n4184, ys__n4185, ys__n4190, ys__n4291, ys__n4292,
    ys__n4294, ys__n4296, ys__n4297, ys__n4299, ys__n4300, ys__n4305,
    ys__n4340, ys__n4448, ys__n4449, ys__n4451, ys__n4452, ys__n4454,
    ys__n4455, ys__n4457, ys__n4458, ys__n4460, ys__n4461, ys__n4465,
    ys__n4478, ys__n4480, ys__n4488, ys__n4494, ys__n4496, ys__n4613,
    ys__n4625, ys__n4627, ys__n4688, ys__n4698, ys__n4736, ys__n4744,
    ys__n4746, ys__n4750, ys__n4751, ys__n4753, ys__n4754, ys__n4756,
    ys__n4757, ys__n4759, ys__n4761, ys__n4783, ys__n4784, ys__n4810,
    ys__n4826, ys__n4832, ys__n4833, ys__n4836, ys__n4837, ys__n6112,
    ys__n6113, ys__n6115, ys__n6118, ys__n6119, ys__n6120, ys__n6121,
    ys__n6123, ys__n6124, ys__n6126, ys__n6127, ys__n6129, ys__n6130,
    ys__n6133, ys__n6134, ys__n17803, ys__n17804, ys__n17806, ys__n17807,
    ys__n17809, ys__n17810, ys__n17812, ys__n17813, ys__n17815, ys__n17816,
    ys__n17818, ys__n17819, ys__n17821, ys__n17822, ys__n17824, ys__n17825,
    ys__n17827, ys__n17828, ys__n17830, ys__n17831, ys__n17833, ys__n17834,
    ys__n17836, ys__n17837, ys__n17839, ys__n17840, ys__n17842, ys__n17843,
    ys__n17845, ys__n17846, ys__n17848, ys__n17849, ys__n17866, ys__n17867,
    ys__n17869, ys__n17870, ys__n17872, ys__n17873, ys__n17875, ys__n17876,
    ys__n17878, ys__n17879, ys__n17881, ys__n17882, ys__n17884, ys__n17885,
    ys__n17887, ys__n17888, ys__n17890, ys__n17891, ys__n17893, ys__n17894,
    ys__n17896, ys__n17897, ys__n17899, ys__n17900, ys__n17902, ys__n17903,
    ys__n17905, ys__n17906, ys__n17908, ys__n17909, ys__n17911, ys__n17912,
    ys__n17941, ys__n17943, ys__n18041, ys__n18043, ys__n18045, ys__n18047,
    ys__n18049, ys__n18051, ys__n18053, ys__n18055, ys__n18057, ys__n18059,
    ys__n18061, ys__n18063, ys__n18065, ys__n18067, ys__n18070, ys__n18071,
    ys__n18090, ys__n18101, ys__n18105, ys__n18106, ys__n18109, ys__n18111,
    ys__n18112, ys__n18114, ys__n18116, ys__n18118, ys__n18121, ys__n18122,
    ys__n18124, ys__n18143, ys__n18149, ys__n18150, ys__n18156, ys__n18173,
    ys__n18208, ys__n18226, ys__n18229, ys__n18231, ys__n18240, ys__n18242,
    ys__n18243, ys__n18270, ys__n18271, ys__n18277, ys__n18280, ys__n18283,
    ys__n18286, ys__n18317, ys__n18378, ys__n18381, ys__n18384, ys__n18389,
    ys__n18393, ys__n18448, ys__n18451, ys__n18454, ys__n18457, ys__n18460,
    ys__n18463, ys__n18466, ys__n18469, ys__n18472, ys__n18475, ys__n18478,
    ys__n18481, ys__n18484, ys__n18487, ys__n18490, ys__n18493, ys__n18496,
    ys__n18499, ys__n18502, ys__n18505, ys__n18508, ys__n18511, ys__n18514,
    ys__n18517, ys__n18520, ys__n18523, ys__n18526, ys__n18529, ys__n18532,
    ys__n18535, ys__n18538, ys__n18541, ys__n18544, ys__n18546, ys__n18556,
    ys__n18558, ys__n18560, ys__n18562, ys__n18565, ys__n18568, ys__n18569,
    ys__n18571, ys__n18572, ys__n18574, ys__n18575, ys__n18577, ys__n18578,
    ys__n18580, ys__n18581, ys__n18583, ys__n18584, ys__n18586, ys__n18587,
    ys__n18589, ys__n18590, ys__n18592, ys__n18593, ys__n18595, ys__n18596,
    ys__n18598, ys__n18599, ys__n18601, ys__n18602, ys__n18604, ys__n18605,
    ys__n18607, ys__n18608, ys__n18610, ys__n18611, ys__n18613, ys__n18614,
    ys__n18616, ys__n18617, ys__n18619, ys__n18620, ys__n18622, ys__n18623,
    ys__n18625, ys__n18626, ys__n18628, ys__n18630, ys__n18632, ys__n18634,
    ys__n18636, ys__n18638, ys__n18639, ys__n18641, ys__n18642, ys__n18644,
    ys__n18645, ys__n18647, ys__n18650, ys__n18651, ys__n18749, ys__n18752,
    ys__n18755, ys__n18758, ys__n18761, ys__n18762, ys__n18765, ys__n18767,
    ys__n18769, ys__n18771, ys__n18773, ys__n18775, ys__n18777, ys__n18779,
    ys__n18781, ys__n18783, ys__n18785, ys__n18787, ys__n18789, ys__n18791,
    ys__n18793, ys__n18795, ys__n18797, ys__n18799, ys__n18801, ys__n18803,
    ys__n18805, ys__n18807, ys__n18809, ys__n18811, ys__n18813, ys__n18815,
    ys__n18817, ys__n18819, ys__n18821, ys__n18823, ys__n18825, ys__n18827,
    ys__n18829, ys__n18831, ys__n18833, ys__n18835, ys__n18837, ys__n18839,
    ys__n18841, ys__n18843, ys__n18845, ys__n18847, ys__n18849, ys__n18851,
    ys__n18853, ys__n18855, ys__n18857, ys__n18859, ys__n18861, ys__n18863,
    ys__n18865, ys__n18867, ys__n18869, ys__n18871, ys__n18873, ys__n18875,
    ys__n18877, ys__n18879, ys__n18881, ys__n18883, ys__n18885, ys__n18887,
    ys__n18889, ys__n18891, ys__n18956, ys__n18957, ys__n18958, ys__n18959,
    ys__n18960, ys__n18961, ys__n18962, ys__n18963, ys__n18964, ys__n18965,
    ys__n18966, ys__n18967, ys__n18968, ys__n18969, ys__n18970, ys__n18971,
    ys__n18972, ys__n18973, ys__n18974, ys__n18975, ys__n18976, ys__n18977,
    ys__n18978, ys__n18979, ys__n18980, ys__n18981, ys__n18982, ys__n18983,
    ys__n18984, ys__n18985, ys__n18986, ys__n18987, ys__n18989, ys__n18991,
    ys__n18993, ys__n18995, ys__n18997, ys__n18999, ys__n19001, ys__n19003,
    ys__n19005, ys__n19007, ys__n19009, ys__n19011, ys__n19013, ys__n19015,
    ys__n19017, ys__n19019, ys__n19021, ys__n19023, ys__n19025, ys__n19027,
    ys__n19029, ys__n19031, ys__n19033, ys__n19035, ys__n19037, ys__n19039,
    ys__n19041, ys__n19043, ys__n19045, ys__n19047, ys__n19049, ys__n19051,
    ys__n19116, ys__n19117, ys__n19118, ys__n19119, ys__n19120, ys__n19121,
    ys__n19122, ys__n19123, ys__n19124, ys__n19125, ys__n19126, ys__n19127,
    ys__n19128, ys__n19129, ys__n19130, ys__n19131, ys__n19132, ys__n19133,
    ys__n19134, ys__n19135, ys__n19136, ys__n19137, ys__n19138, ys__n19139,
    ys__n19140, ys__n19141, ys__n19142, ys__n19143, ys__n19144, ys__n19145,
    ys__n19146, ys__n19147, ys__n19156, ys__n19157, ys__n19166, ys__n19171,
    ys__n19203, ys__n19215, ys__n19245, ys__n19251, ys__n19253, ys__n19259,
    ys__n19261, ys__n19263, ys__n19843, ys__n19844, ys__n19845, ys__n19846,
    ys__n19847, ys__n19848, ys__n19849, ys__n19850, ys__n19851, ys__n19852,
    ys__n19853, ys__n19854, ys__n19855, ys__n19856, ys__n19857, ys__n19858,
    ys__n19859, ys__n19860, ys__n19861, ys__n19862, ys__n19863, ys__n19864,
    ys__n19865, ys__n19866, ys__n19867, ys__n19868, ys__n19869, ys__n19870,
    ys__n19871, ys__n19872, ys__n19873, ys__n19874, ys__n19875, ys__n19972,
    ys__n19973, ys__n19974, ys__n19975, ys__n19976, ys__n19977, ys__n19978,
    ys__n19979, ys__n19980, ys__n19981, ys__n19982, ys__n19983, ys__n19984,
    ys__n19985, ys__n19986, ys__n19987, ys__n19988, ys__n19989, ys__n19990,
    ys__n19991, ys__n19992, ys__n19993, ys__n19994, ys__n19995, ys__n19996,
    ys__n19997, ys__n19998, ys__n19999, ys__n20000, ys__n20001, ys__n20002,
    ys__n20003, ys__n20004, ys__n20035, ys__n20058, ys__n20061, ys__n20064,
    ys__n20067, ys__n20070, ys__n20073, ys__n20076, ys__n20079, ys__n20138,
    ys__n20140, ys__n20142, ys__n20144, ys__n20146, ys__n20148, ys__n20150,
    ys__n20152, ys__n20186, ys__n20188, ys__n20190, ys__n20192, ys__n20194,
    ys__n20196, ys__n20198, ys__n20200, ys__n20202, ys__n20204, ys__n20206,
    ys__n20208, ys__n20210, ys__n20212, ys__n20214, ys__n20216, ys__n20273,
    ys__n20279, ys__n20280, ys__n20540, ys__n20542, ys__n20544, ys__n20546,
    ys__n20548, ys__n20550, ys__n20552, ys__n20554, ys__n20556, ys__n20558,
    ys__n20560, ys__n20562, ys__n20564, ys__n20566, ys__n20568, ys__n20570,
    ys__n20572, ys__n20574, ys__n20576, ys__n20578, ys__n20580, ys__n20582,
    ys__n20584, ys__n20586, ys__n20588, ys__n20590, ys__n20592, ys__n20594,
    ys__n20596, ys__n20598, ys__n20600, ys__n20602, ys__n20604, ys__n20606,
    ys__n20608, ys__n20610, ys__n20612, ys__n20614, ys__n20616, ys__n20618,
    ys__n20620, ys__n20622, ys__n20624, ys__n20626, ys__n20628, ys__n20630,
    ys__n20632, ys__n20634, ys__n20636, ys__n20638, ys__n20640, ys__n20642,
    ys__n20644, ys__n20646, ys__n20648, ys__n20650, ys__n20652, ys__n20654,
    ys__n20656, ys__n20658, ys__n20660, ys__n20662, ys__n20664, ys__n20666,
    ys__n20668, ys__n20670, ys__n20672, ys__n20674, ys__n20676, ys__n20678,
    ys__n20680, ys__n20682, ys__n20684, ys__n20686, ys__n20688, ys__n20690,
    ys__n20692, ys__n20694, ys__n20696, ys__n20698, ys__n20700, ys__n20702,
    ys__n20704, ys__n20706, ys__n20708, ys__n20710, ys__n20712, ys__n20714,
    ys__n20716, ys__n20718, ys__n20720, ys__n20722, ys__n20724, ys__n20726,
    ys__n20728, ys__n20730, ys__n20732, ys__n20734, ys__n20736, ys__n20738,
    ys__n20740, ys__n20742, ys__n20744, ys__n20746, ys__n20748, ys__n20750,
    ys__n20752, ys__n20754, ys__n20756, ys__n20758, ys__n20760, ys__n20762,
    ys__n20764, ys__n20766, ys__n20768, ys__n20770, ys__n20772, ys__n20774,
    ys__n20776, ys__n20778, ys__n20780, ys__n20782, ys__n20784, ys__n20786,
    ys__n20788, ys__n20790, ys__n20792, ys__n20794, ys__n20796, ys__n20798,
    ys__n20800, ys__n20802, ys__n20804, ys__n20806, ys__n20808, ys__n20810,
    ys__n20812, ys__n20814, ys__n20816, ys__n20818, ys__n20820, ys__n20822,
    ys__n20824, ys__n20826, ys__n20828, ys__n20830, ys__n20832, ys__n20834,
    ys__n20836, ys__n20838, ys__n20840, ys__n20842, ys__n20844, ys__n20846,
    ys__n20848, ys__n20850, ys__n20852, ys__n20854, ys__n20856, ys__n20858,
    ys__n20860, ys__n20862, ys__n20864, ys__n20866, ys__n20868, ys__n20870,
    ys__n20872, ys__n20874, ys__n20876, ys__n20878, ys__n20880, ys__n20882,
    ys__n20884, ys__n20886, ys__n20888, ys__n20890, ys__n20892, ys__n20894,
    ys__n20896, ys__n20898, ys__n20900, ys__n20902, ys__n20904, ys__n20906,
    ys__n20908, ys__n20910, ys__n20912, ys__n20914, ys__n20916, ys__n20918,
    ys__n20920, ys__n20922, ys__n20924, ys__n20925, ys__n20926, ys__n20927,
    ys__n20928, ys__n20929, ys__n20930, ys__n20931, ys__n20932, ys__n20933,
    ys__n20934, ys__n20935, ys__n20936, ys__n20937, ys__n20938, ys__n20939,
    ys__n20940, ys__n20941, ys__n20942, ys__n20943, ys__n20944, ys__n20945,
    ys__n20946, ys__n20947, ys__n20948, ys__n20949, ys__n20950, ys__n20951,
    ys__n20952, ys__n20953, ys__n20954, ys__n20955, ys__n20956, ys__n20958,
    ys__n20960, ys__n20962, ys__n20964, ys__n20966, ys__n20968, ys__n20970,
    ys__n20972, ys__n20974, ys__n20976, ys__n20978, ys__n20980, ys__n20982,
    ys__n20984, ys__n20986, ys__n20988, ys__n20990, ys__n20992, ys__n20994,
    ys__n20996, ys__n20998, ys__n21000, ys__n21002, ys__n21004, ys__n21006,
    ys__n21008, ys__n21010, ys__n21012, ys__n21014, ys__n21016, ys__n21018,
    ys__n21020, ys__n21022, ys__n21024, ys__n21026, ys__n21028, ys__n21030,
    ys__n21032, ys__n21034, ys__n21036, ys__n21038, ys__n21040, ys__n21042,
    ys__n21044, ys__n21046, ys__n21048, ys__n21050, ys__n21052, ys__n21054,
    ys__n21056, ys__n21058, ys__n21060, ys__n21062, ys__n21064, ys__n21066,
    ys__n21068, ys__n21070, ys__n21072, ys__n21074, ys__n21076, ys__n21078,
    ys__n21080, ys__n21082, ys__n21084, ys__n21086, ys__n21088, ys__n21090,
    ys__n21092, ys__n21094, ys__n21096, ys__n21098, ys__n21100, ys__n21102,
    ys__n21104, ys__n21106, ys__n21108, ys__n21110, ys__n21112, ys__n21114,
    ys__n21116, ys__n21118, ys__n21120, ys__n21122, ys__n21124, ys__n21126,
    ys__n21128, ys__n21130, ys__n21132, ys__n21134, ys__n21136, ys__n21138,
    ys__n21140, ys__n21142, ys__n21144, ys__n21146, ys__n21148, ys__n21150,
    ys__n21152, ys__n21154, ys__n21156, ys__n21158, ys__n21160, ys__n21162,
    ys__n21164, ys__n21166, ys__n21168, ys__n21170, ys__n21172, ys__n21174,
    ys__n21176, ys__n21178, ys__n21180, ys__n21182, ys__n21184, ys__n21186,
    ys__n21188, ys__n21190, ys__n21192, ys__n21194, ys__n21196, ys__n21198,
    ys__n21200, ys__n21202, ys__n21204, ys__n21206, ys__n21208, ys__n21210,
    ys__n21212, ys__n21214, ys__n21216, ys__n21218, ys__n21220, ys__n21222,
    ys__n21224, ys__n21226, ys__n21228, ys__n21230, ys__n21232, ys__n21234,
    ys__n21236, ys__n21238, ys__n21240, ys__n21242, ys__n21244, ys__n21246,
    ys__n21248, ys__n21250, ys__n21252, ys__n21254, ys__n21256, ys__n21258,
    ys__n21260, ys__n21262, ys__n21264, ys__n21266, ys__n21268, ys__n21270,
    ys__n21272, ys__n21274, ys__n21276, ys__n21278, ys__n21280, ys__n21282,
    ys__n21284, ys__n21286, ys__n21288, ys__n21290, ys__n21292, ys__n21294,
    ys__n21296, ys__n21298, ys__n21300, ys__n21302, ys__n21304, ys__n21306,
    ys__n21308, ys__n21310, ys__n21312, ys__n21314, ys__n21316, ys__n21318,
    ys__n21320, ys__n21322, ys__n21324, ys__n21326, ys__n21328, ys__n21330,
    ys__n21332, ys__n21334, ys__n21336, ys__n21338, ys__n21340, ys__n21342,
    ys__n21344, ys__n21346, ys__n21348, ys__n21350, ys__n21352, ys__n21354,
    ys__n21356, ys__n21358, ys__n21360, ys__n21362, ys__n21364, ys__n21366,
    ys__n21368, ys__n21370, ys__n21372, ys__n21374, ys__n21376, ys__n21378,
    ys__n21380, ys__n21382, ys__n21384, ys__n21386, ys__n21388, ys__n21390,
    ys__n21392, ys__n21394, ys__n21396, ys__n21398, ys__n21400, ys__n21402,
    ys__n21404, ys__n21405, ys__n21406, ys__n21407, ys__n21408, ys__n21409,
    ys__n21410, ys__n21411, ys__n21412, ys__n21413, ys__n21414, ys__n21415,
    ys__n21416, ys__n21417, ys__n21418, ys__n21419, ys__n21420, ys__n21421,
    ys__n21422, ys__n21423, ys__n21424, ys__n21425, ys__n21426, ys__n21427,
    ys__n21428, ys__n21429, ys__n21430, ys__n21431, ys__n21432, ys__n21433,
    ys__n21434, ys__n21435, ys__n21500, ys__n21502, ys__n21504, ys__n21506,
    ys__n21508, ys__n21510, ys__n21512, ys__n21514, ys__n21516, ys__n21518,
    ys__n21520, ys__n21522, ys__n21524, ys__n21526, ys__n21528, ys__n21530,
    ys__n21532, ys__n21534, ys__n21536, ys__n21538, ys__n21540, ys__n21542,
    ys__n21544, ys__n21546, ys__n21548, ys__n21550, ys__n21552, ys__n21554,
    ys__n21556, ys__n21558, ys__n21560, ys__n21562, ys__n21564, ys__n21566,
    ys__n21568, ys__n21570, ys__n21572, ys__n21574, ys__n21576, ys__n21578,
    ys__n21580, ys__n21582, ys__n21584, ys__n21586, ys__n21588, ys__n21590,
    ys__n21592, ys__n21594, ys__n21596, ys__n21598, ys__n21600, ys__n21602,
    ys__n21604, ys__n21606, ys__n21608, ys__n21610, ys__n21612, ys__n21614,
    ys__n21616, ys__n21618, ys__n21620, ys__n21622, ys__n21624, ys__n21626,
    ys__n21628, ys__n21630, ys__n21632, ys__n21634, ys__n21636, ys__n21638,
    ys__n21640, ys__n21642, ys__n21644, ys__n21646, ys__n21648, ys__n21650,
    ys__n21652, ys__n21654, ys__n21656, ys__n21658, ys__n21660, ys__n21662,
    ys__n21664, ys__n21666, ys__n21668, ys__n21670, ys__n21672, ys__n21674,
    ys__n21676, ys__n21678, ys__n21680, ys__n21682, ys__n21684, ys__n21686,
    ys__n21688, ys__n21690, ys__n21692, ys__n21694, ys__n21696, ys__n21698,
    ys__n21700, ys__n21702, ys__n21704, ys__n21706, ys__n21708, ys__n21710,
    ys__n21712, ys__n21714, ys__n21716, ys__n21718, ys__n21720, ys__n21722,
    ys__n21724, ys__n21726, ys__n21728, ys__n21730, ys__n21732, ys__n21734,
    ys__n21736, ys__n21738, ys__n21740, ys__n21742, ys__n21744, ys__n21746,
    ys__n21748, ys__n21750, ys__n21752, ys__n21754, ys__n21756, ys__n21758,
    ys__n21760, ys__n21762, ys__n21764, ys__n21766, ys__n21768, ys__n21770,
    ys__n21772, ys__n21774, ys__n21776, ys__n21778, ys__n21780, ys__n21782,
    ys__n21784, ys__n21786, ys__n21788, ys__n21790, ys__n21792, ys__n21794,
    ys__n21796, ys__n21798, ys__n21800, ys__n21802, ys__n21804, ys__n21806,
    ys__n21808, ys__n21810, ys__n21812, ys__n21814, ys__n21816, ys__n21818,
    ys__n21820, ys__n21822, ys__n21824, ys__n21826, ys__n21828, ys__n21830,
    ys__n21832, ys__n21834, ys__n21836, ys__n21838, ys__n21840, ys__n21842,
    ys__n21844, ys__n21846, ys__n21848, ys__n21850, ys__n21852, ys__n21854,
    ys__n21856, ys__n21858, ys__n21860, ys__n21862, ys__n21864, ys__n21866,
    ys__n21868, ys__n21870, ys__n21872, ys__n21874, ys__n21876, ys__n21878,
    ys__n21880, ys__n21882, ys__n21884, ys__n21886, ys__n21888, ys__n21890,
    ys__n21892, ys__n21894, ys__n21896, ys__n21898, ys__n21900, ys__n21902,
    ys__n21904, ys__n21906, ys__n21908, ys__n21910, ys__n21912, ys__n21914,
    ys__n21916, ys__n21918, ys__n21920, ys__n21922, ys__n21924, ys__n21926,
    ys__n21928, ys__n21930, ys__n21932, ys__n21934, ys__n21936, ys__n21938,
    ys__n21940, ys__n21942, ys__n21944, ys__n21946, ys__n21948, ys__n21949,
    ys__n21950, ys__n21951, ys__n21952, ys__n21953, ys__n21954, ys__n21955,
    ys__n21956, ys__n21957, ys__n21958, ys__n21959, ys__n21960, ys__n21961,
    ys__n21962, ys__n21963, ys__n21964, ys__n21965, ys__n21966, ys__n21967,
    ys__n21968, ys__n21969, ys__n21970, ys__n21971, ys__n21972, ys__n21973,
    ys__n21974, ys__n21975, ys__n21976, ys__n21977, ys__n21978, ys__n21979,
    ys__n21980, ys__n21982, ys__n21984, ys__n21986, ys__n21988, ys__n21990,
    ys__n21992, ys__n21994, ys__n21996, ys__n21998, ys__n22000, ys__n22002,
    ys__n22004, ys__n22006, ys__n22008, ys__n22010, ys__n22012, ys__n22014,
    ys__n22016, ys__n22018, ys__n22020, ys__n22022, ys__n22024, ys__n22026,
    ys__n22028, ys__n22030, ys__n22032, ys__n22034, ys__n22036, ys__n22038,
    ys__n22040, ys__n22042, ys__n22044, ys__n22046, ys__n22048, ys__n22050,
    ys__n22052, ys__n22054, ys__n22056, ys__n22058, ys__n22060, ys__n22062,
    ys__n22064, ys__n22066, ys__n22068, ys__n22070, ys__n22072, ys__n22074,
    ys__n22076, ys__n22078, ys__n22080, ys__n22082, ys__n22084, ys__n22086,
    ys__n22088, ys__n22090, ys__n22092, ys__n22094, ys__n22096, ys__n22098,
    ys__n22100, ys__n22102, ys__n22104, ys__n22106, ys__n22108, ys__n22110,
    ys__n22112, ys__n22114, ys__n22116, ys__n22118, ys__n22120, ys__n22122,
    ys__n22124, ys__n22126, ys__n22128, ys__n22130, ys__n22132, ys__n22134,
    ys__n22136, ys__n22138, ys__n22140, ys__n22142, ys__n22144, ys__n22146,
    ys__n22148, ys__n22150, ys__n22152, ys__n22154, ys__n22156, ys__n22158,
    ys__n22160, ys__n22162, ys__n22164, ys__n22166, ys__n22168, ys__n22170,
    ys__n22172, ys__n22174, ys__n22176, ys__n22178, ys__n22180, ys__n22182,
    ys__n22184, ys__n22186, ys__n22188, ys__n22190, ys__n22192, ys__n22194,
    ys__n22196, ys__n22198, ys__n22200, ys__n22202, ys__n22204, ys__n22206,
    ys__n22208, ys__n22210, ys__n22212, ys__n22214, ys__n22216, ys__n22218,
    ys__n22220, ys__n22222, ys__n22224, ys__n22226, ys__n22228, ys__n22230,
    ys__n22232, ys__n22234, ys__n22236, ys__n22238, ys__n22240, ys__n22242,
    ys__n22244, ys__n22246, ys__n22248, ys__n22250, ys__n22252, ys__n22254,
    ys__n22256, ys__n22258, ys__n22260, ys__n22262, ys__n22264, ys__n22266,
    ys__n22268, ys__n22270, ys__n22272, ys__n22274, ys__n22276, ys__n22278,
    ys__n22280, ys__n22282, ys__n22284, ys__n22286, ys__n22288, ys__n22290,
    ys__n22292, ys__n22294, ys__n22296, ys__n22298, ys__n22300, ys__n22302,
    ys__n22304, ys__n22306, ys__n22308, ys__n22310, ys__n22312, ys__n22314,
    ys__n22316, ys__n22318, ys__n22320, ys__n22322, ys__n22324, ys__n22326,
    ys__n22328, ys__n22330, ys__n22332, ys__n22334, ys__n22336, ys__n22338,
    ys__n22340, ys__n22342, ys__n22344, ys__n22346, ys__n22348, ys__n22350,
    ys__n22352, ys__n22354, ys__n22356, ys__n22358, ys__n22360, ys__n22362,
    ys__n22364, ys__n22366, ys__n22368, ys__n22370, ys__n22372, ys__n22374,
    ys__n22376, ys__n22378, ys__n22380, ys__n22382, ys__n22384, ys__n22386,
    ys__n22388, ys__n22390, ys__n22392, ys__n22394, ys__n22396, ys__n22398,
    ys__n22400, ys__n22402, ys__n22404, ys__n22406, ys__n22408, ys__n22410,
    ys__n22412, ys__n22414, ys__n22416, ys__n22418, ys__n22420, ys__n22422,
    ys__n22424, ys__n22426, ys__n22428, ys__n22429, ys__n22430, ys__n22431,
    ys__n22432, ys__n22433, ys__n22434, ys__n22435, ys__n22436, ys__n22437,
    ys__n22438, ys__n22439, ys__n22440, ys__n22441, ys__n22442, ys__n22443,
    ys__n22444, ys__n22445, ys__n22446, ys__n22447, ys__n22448, ys__n22449,
    ys__n22450, ys__n22451, ys__n22452, ys__n22453, ys__n22454, ys__n22455,
    ys__n22456, ys__n22457, ys__n22458, ys__n22459, ys__n22464, ys__n22465,
    ys__n22564, ys__n22566, ys__n22568, ys__n22570, ys__n22572, ys__n22574,
    ys__n22576, ys__n22578, ys__n22580, ys__n22582, ys__n22584, ys__n22586,
    ys__n22588, ys__n22590, ys__n22592, ys__n22594, ys__n22596, ys__n22598,
    ys__n22600, ys__n22602, ys__n22604, ys__n22606, ys__n22608, ys__n22610,
    ys__n22612, ys__n22614, ys__n22616, ys__n22618, ys__n22620, ys__n22622,
    ys__n22624, ys__n22626, ys__n22630, ys__n22632, ys__n22634, ys__n22636,
    ys__n22640, ys__n22642, ys__n22644, ys__n22646, ys__n22648, ys__n22650,
    ys__n22652, ys__n22654, ys__n22668, ys__n22670, ys__n22673, ys__n22675,
    ys__n22677, ys__n22679, ys__n22681, ys__n22683, ys__n22685, ys__n22687,
    ys__n22689, ys__n22715, ys__n22717, ys__n22719, ys__n22721, ys__n22723,
    ys__n22725, ys__n22727, ys__n22729, ys__n22731, ys__n22733, ys__n22735,
    ys__n22737, ys__n22739, ys__n22741, ys__n22743, ys__n22745, ys__n22747,
    ys__n22749, ys__n22751, ys__n22753, ys__n22755, ys__n22757, ys__n22759,
    ys__n22761, ys__n22763, ys__n22765, ys__n22767, ys__n22769, ys__n22771,
    ys__n22773, ys__n22775, ys__n22777, ys__n22779, ys__n22781, ys__n22783,
    ys__n22785, ys__n22787, ys__n22789, ys__n22792, ys__n22794, ys__n22799,
    ys__n22818, ys__n22820, ys__n22822, ys__n22824, ys__n22826, ys__n22828,
    ys__n22830, ys__n22832, ys__n22834, ys__n22836, ys__n22838, ys__n22840,
    ys__n22842, ys__n22844, ys__n22846, ys__n22848, ys__n22850, ys__n22852,
    ys__n22854, ys__n22856, ys__n22858, ys__n22860, ys__n22862, ys__n22864,
    ys__n22866, ys__n22868, ys__n22870, ys__n22872, ys__n22874, ys__n22876,
    ys__n22878, ys__n22880, ys__n22882, ys__n22884, ys__n22885, ys__n22886,
    ys__n22887, ys__n22888, ys__n22889, ys__n22890, ys__n22891, ys__n22892,
    ys__n22893, ys__n22894, ys__n22895, ys__n22896, ys__n22897, ys__n22898,
    ys__n22899, ys__n22900, ys__n22901, ys__n22902, ys__n22903, ys__n22904,
    ys__n22905, ys__n22906, ys__n22907, ys__n22908, ys__n22909, ys__n22910,
    ys__n22911, ys__n22912, ys__n22913, ys__n22914, ys__n22915, ys__n22916,
    ys__n22918, ys__n22921, ys__n22924, ys__n22927, ys__n22930, ys__n22933,
    ys__n22936, ys__n22939, ys__n22942, ys__n22945, ys__n22948, ys__n22951,
    ys__n22954, ys__n22957, ys__n22960, ys__n22963, ys__n22966, ys__n22969,
    ys__n22972, ys__n22975, ys__n22978, ys__n22981, ys__n22984, ys__n22987,
    ys__n22990, ys__n22993, ys__n22996, ys__n22999, ys__n23002, ys__n23005,
    ys__n23008, ys__n23011, ys__n23014, ys__n23016, ys__n23018, ys__n23020,
    ys__n23022, ys__n23024, ys__n23026, ys__n23028, ys__n23030, ys__n23032,
    ys__n23034, ys__n23036, ys__n23038, ys__n23040, ys__n23042, ys__n23044,
    ys__n23046, ys__n23048, ys__n23050, ys__n23052, ys__n23054, ys__n23056,
    ys__n23058, ys__n23060, ys__n23062, ys__n23064, ys__n23066, ys__n23068,
    ys__n23070, ys__n23072, ys__n23074, ys__n23076, ys__n23077, ys__n23078,
    ys__n23079, ys__n23080, ys__n23081, ys__n23082, ys__n23083, ys__n23084,
    ys__n23085, ys__n23086, ys__n23087, ys__n23088, ys__n23089, ys__n23090,
    ys__n23091, ys__n23092, ys__n23093, ys__n23094, ys__n23095, ys__n23096,
    ys__n23097, ys__n23098, ys__n23099, ys__n23100, ys__n23101, ys__n23102,
    ys__n23103, ys__n23104, ys__n23105, ys__n23106, ys__n23107, ys__n23108,
    ys__n23111, ys__n23114, ys__n23117, ys__n23120, ys__n23123, ys__n23126,
    ys__n23129, ys__n23132, ys__n23135, ys__n23138, ys__n23141, ys__n23144,
    ys__n23147, ys__n23150, ys__n23153, ys__n23156, ys__n23159, ys__n23162,
    ys__n23165, ys__n23168, ys__n23171, ys__n23174, ys__n23177, ys__n23180,
    ys__n23183, ys__n23186, ys__n23189, ys__n23192, ys__n23195, ys__n23198,
    ys__n23203, ys__n23205, ys__n23207, ys__n23209, ys__n23211, ys__n23213,
    ys__n23215, ys__n23217, ys__n23219, ys__n23221, ys__n23223, ys__n23225,
    ys__n23227, ys__n23229, ys__n23231, ys__n23233, ys__n23235, ys__n23237,
    ys__n23239, ys__n23241, ys__n23243, ys__n23245, ys__n23247, ys__n23249,
    ys__n23251, ys__n23253, ys__n23255, ys__n23257, ys__n23259, ys__n23261,
    ys__n23269, ys__n23271, ys__n23272, ys__n23274, ys__n23276, ys__n23278,
    ys__n23280, ys__n23282, ys__n23284, ys__n23286, ys__n23288, ys__n23290,
    ys__n23292, ys__n23294, ys__n23296, ys__n23298, ys__n23300, ys__n23302,
    ys__n23304, ys__n23306, ys__n23308, ys__n23310, ys__n23312, ys__n23314,
    ys__n23316, ys__n23318, ys__n23320, ys__n23322, ys__n23324, ys__n23326,
    ys__n23328, ys__n23330, ys__n23332, ys__n23335, ys__n23339, ys__n23480,
    ys__n23548, ys__n23550, ys__n23552, ys__n23554, ys__n23556, ys__n23558,
    ys__n23560, ys__n23562, ys__n23564, ys__n23566, ys__n23568, ys__n23570,
    ys__n23572, ys__n23574, ys__n23627, ys__n23629, ys__n23641, ys__n23644,
    ys__n23645, ys__n23647, ys__n23650, ys__n23652, ys__n23655, ys__n23658,
    ys__n23661, ys__n23663, ys__n23705, ys__n23706, ys__n23707, ys__n23708,
    ys__n23709, ys__n23710, ys__n23711, ys__n23712, ys__n23713, ys__n23714,
    ys__n23715, ys__n23717, ys__n23729, ys__n23730, ys__n23763, ys__n23818,
    ys__n23819, ys__n23820, ys__n23821, ys__n23822, ys__n23834, ys__n23836,
    ys__n23838, ys__n23840, ys__n23842, ys__n23850, ys__n23888, ys__n23889,
    ys__n23890, ys__n23891, ys__n23892, ys__n23904, ys__n23906, ys__n23908,
    ys__n23910, ys__n23912, ys__n23956, ys__n23957, ys__n23958, ys__n23959,
    ys__n23960, ys__n23977, ys__n23979, ys__n23981, ys__n23983, ys__n23985,
    ys__n24106, ys__n24107, ys__n24108, ys__n24112, ys__n24123, ys__n24124,
    ys__n24131, ys__n24143, ys__n24158, ys__n24167, ys__n24168, ys__n24177,
    ys__n24197, ys__n24199, ys__n24201, ys__n24203, ys__n24205, ys__n24207,
    ys__n24209, ys__n24211, ys__n24213, ys__n24215, ys__n24217, ys__n24219,
    ys__n24228, ys__n24233, ys__n24235, ys__n24243, ys__n24248, ys__n24279,
    ys__n24280, ys__n24303, ys__n24306, ys__n24308, ys__n24310, ys__n24312,
    ys__n24314, ys__n24316, ys__n24318, ys__n24337, ys__n24340, ys__n24342,
    ys__n24344, ys__n24346, ys__n24348, ys__n24350, ys__n24352, ys__n24371,
    ys__n24374, ys__n24376, ys__n24378, ys__n24380, ys__n24382, ys__n24384,
    ys__n24386, ys__n24389, ys__n24406, ys__n24409, ys__n24411, ys__n24413,
    ys__n24415, ys__n24417, ys__n24419, ys__n24421, ys__n24427, ys__n24433,
    ys__n24434, ys__n24461, ys__n24463, ys__n24464, ys__n24483, ys__n24485,
    ys__n24506, ys__n24519, ys__n24567, ys__n24575, ys__n24578, ys__n24590,
    ys__n24591, ys__n24615, ys__n24616, ys__n24617, ys__n24618, ys__n24619,
    ys__n24620, ys__n24621, ys__n24622, ys__n24623, ys__n24624, ys__n24625,
    ys__n24626, ys__n24627, ys__n24628, ys__n24629, ys__n24630, ys__n24631,
    ys__n24632, ys__n24633, ys__n24634, ys__n24635, ys__n24636, ys__n24637,
    ys__n24638, ys__n24639, ys__n24640, ys__n24641, ys__n24642, ys__n24643,
    ys__n24644, ys__n24645, ys__n24646, ys__n24647, ys__n24648, ys__n24649,
    ys__n24650, ys__n24651, ys__n24652, ys__n24653, ys__n24654, ys__n24655,
    ys__n24656, ys__n24657, ys__n24658, ys__n24659, ys__n24660, ys__n24661,
    ys__n24662, ys__n24663, ys__n24664, ys__n24665, ys__n24666, ys__n24667,
    ys__n24668, ys__n24669, ys__n24670, ys__n24671, ys__n24672, ys__n24673,
    ys__n24674, ys__n24675, ys__n24677, ys__n24679, ys__n24681, ys__n24683,
    ys__n24684, ys__n24685, ys__n24686, ys__n24687, ys__n24688, ys__n24689,
    ys__n24690, ys__n24691, ys__n24692, ys__n24693, ys__n24694, ys__n24695,
    ys__n24696, ys__n24697, ys__n24698, ys__n24699, ys__n24700, ys__n24701,
    ys__n24702, ys__n24703, ys__n24704, ys__n24705, ys__n24706, ys__n24707,
    ys__n24708, ys__n24709, ys__n24710, ys__n24711, ys__n24712, ys__n24741,
    ys__n24744, ys__n24747, ys__n24750, ys__n24753, ys__n24756, ys__n24759,
    ys__n24762, ys__n24765, ys__n24768, ys__n24771, ys__n24774, ys__n24777,
    ys__n24780, ys__n24783, ys__n24786, ys__n24789, ys__n24792, ys__n24795,
    ys__n24798, ys__n24801, ys__n24804, ys__n24807, ys__n24810, ys__n24813,
    ys__n24816, ys__n24819, ys__n24822, ys__n24825, ys__n24828, ys__n24831,
    ys__n24834, ys__n25292, ys__n25300, ys__n25381, ys__n25382, ys__n25383,
    ys__n25384, ys__n25470, ys__n25564, ys__n25567, ys__n25570, ys__n25573,
    ys__n25576, ys__n25579, ys__n25582, ys__n25585, ys__n25588, ys__n25591,
    ys__n25594, ys__n25597, ys__n25600, ys__n25603, ys__n25606, ys__n25609,
    ys__n25612, ys__n25615, ys__n25618, ys__n25621, ys__n25624, ys__n25627,
    ys__n25630, ys__n25633, ys__n25636, ys__n25639, ys__n25642, ys__n25645,
    ys__n25648, ys__n25651, ys__n25654, ys__n25657, ys__n25727, ys__n25730,
    ys__n25733, ys__n25736, ys__n25853, ys__n25856, ys__n25859, ys__n25862,
    ys__n25980, ys__n25984, ys__n25987, ys__n25990, ys__n25993, ys__n25996,
    ys__n25999, ys__n26002, ys__n26005, ys__n26008, ys__n26011, ys__n26014,
    ys__n26017, ys__n26020, ys__n26023, ys__n26026, ys__n26029, ys__n26032,
    ys__n26035, ys__n26038, ys__n26041, ys__n26044, ys__n26047, ys__n26050,
    ys__n26053, ys__n26056, ys__n26059, ys__n26062, ys__n26065, ys__n26068,
    ys__n26071, ys__n26074, ys__n26143, ys__n26145, ys__n26147, ys__n26149,
    ys__n26151, ys__n26153, ys__n26155, ys__n26157, ys__n26159, ys__n26161,
    ys__n26162, ys__n26164, ys__n26166, ys__n26168, ys__n26170, ys__n26172,
    ys__n26174, ys__n26176, ys__n26178, ys__n26180, ys__n26182, ys__n26184,
    ys__n26186, ys__n26188, ys__n26190, ys__n26192, ys__n26194, ys__n26196,
    ys__n26198, ys__n26200, ys__n26202, ys__n26204, ys__n26206, ys__n26208,
    ys__n26210, ys__n26212, ys__n26214, ys__n26216, ys__n26218, ys__n26279,
    ys__n26285, ys__n26359, ys__n26362, ys__n26425, ys__n26428, ys__n26431,
    ys__n26434, ys__n26437, ys__n26440, ys__n26443, ys__n26446, ys__n26449,
    ys__n26452, ys__n26455, ys__n26460, ys__n26463, ys__n26466, ys__n26469,
    ys__n26472, ys__n26475, ys__n26478, ys__n26481, ys__n26484, ys__n26487,
    ys__n26490, ys__n26493, ys__n26496, ys__n26499, ys__n26502, ys__n26505,
    ys__n26508, ys__n26511, ys__n26514, ys__n26517, ys__n26552, ys__n26553,
    ys__n26554, ys__n26556, ys__n26557, ys__n26558, ys__n26559, ys__n26560,
    ys__n26561, ys__n26562, ys__n26563, ys__n26564, ys__n26565, ys__n26567,
    ys__n26568, ys__n26569, ys__n26570, ys__n26571, ys__n26572, ys__n26766,
    ys__n26768, ys__n26770, ys__n26772, ys__n27479, ys__n27481, ys__n27485,
    ys__n27488, ys__n27496, ys__n27498, ys__n27499, ys__n27507, ys__n27509,
    ys__n27510, ys__n27518, ys__n27520, ys__n27607, ys__n27608, ys__n27611,
    ys__n27612, ys__n27614, ys__n27615, ys__n27617, ys__n27618, ys__n27620,
    ys__n27621, ys__n27623, ys__n27624, ys__n27626, ys__n27627, ys__n27629,
    ys__n27630, ys__n27632, ys__n27633, ys__n27635, ys__n27636, ys__n27638,
    ys__n27639, ys__n27641, ys__n27642, ys__n27644, ys__n27645, ys__n27647,
    ys__n27648, ys__n27650, ys__n27651, ys__n27653, ys__n27654, ys__n27656,
    ys__n27657, ys__n27659, ys__n27660, ys__n27662, ys__n27663, ys__n27665,
    ys__n27666, ys__n27668, ys__n27669, ys__n27671, ys__n27672, ys__n27674,
    ys__n27675, ys__n27677, ys__n27678, ys__n27680, ys__n27681, ys__n27683,
    ys__n27684, ys__n27686, ys__n27687, ys__n27689, ys__n27690, ys__n27692,
    ys__n27693, ys__n27695, ys__n27696, ys__n27698, ys__n27699, ys__n27701,
    ys__n27702, ys__n27737, ys__n27738, ys__n27740, ys__n27743, ys__n27747,
    ys__n27750, ys__n27753, ys__n27756, ys__n27759, ys__n27762, ys__n27765,
    ys__n27768, ys__n27771, ys__n27774, ys__n27777, ys__n27780, ys__n27783,
    ys__n27786, ys__n27789, ys__n27792, ys__n27795, ys__n27798, ys__n27801,
    ys__n27804, ys__n27807, ys__n27810, ys__n27813, ys__n27816, ys__n27819,
    ys__n27822, ys__n27825, ys__n27828, ys__n27831, ys__n27834, ys__n27837,
    ys__n27855, ys__n27857, ys__n27859, ys__n27861, ys__n27863, ys__n27865,
    ys__n27867, ys__n27869, ys__n27871, ys__n27873, ys__n27875, ys__n27877,
    ys__n27879, ys__n27881, ys__n27883, ys__n27885, ys__n28015, ys__n28016,
    ys__n28017, ys__n28018, ys__n28019, ys__n28020, ys__n28021, ys__n28022,
    ys__n28023, ys__n28024, ys__n28025, ys__n28026, ys__n28027, ys__n28028,
    ys__n28029, ys__n28030, ys__n28243, ys__n28287, ys__n28288, ys__n28290,
    ys__n28292, ys__n28294, ys__n28296, ys__n28424, ys__n28426, ys__n28428,
    ys__n28430, ys__n28432, ys__n28434, ys__n28436, ys__n28438, ys__n28446,
    ys__n28453, ys__n28455, ys__n28457, ys__n28459, ys__n28462, ys__n28464,
    ys__n28466, ys__n28468, ys__n28470, ys__n28472, ys__n28632, ys__n28633,
    ys__n28634, ys__n28635, ys__n28636, ys__n28637, ys__n28638, ys__n28639,
    ys__n28640, ys__n28641, ys__n28718, ys__n28719, ys__n28720, ys__n28859,
    ys__n28863, ys__n28866, ys__n28869, ys__n28872, ys__n28875, ys__n28878,
    ys__n28881, ys__n28884, ys__n28887, ys__n28890, ys__n28893, ys__n28896,
    ys__n28899, ys__n28902, ys__n28905, ys__n28908, ys__n28911, ys__n28914,
    ys__n28917, ys__n28920, ys__n28923, ys__n28926, ys__n28929, ys__n28932,
    ys__n28935, ys__n28938, ys__n28941, ys__n28944, ys__n28947, ys__n28950,
    ys__n28953, ys__n29117, ys__n29119, ys__n29120, ys__n29121, ys__n29123,
    ys__n29124, ys__n29126, ys__n29127, ys__n29129, ys__n29130, ys__n29132,
    ys__n29133, ys__n29135, ys__n29136, ys__n29138, ys__n29139, ys__n29141,
    ys__n29142, ys__n29144, ys__n29145, ys__n29147, ys__n29148, ys__n29150,
    ys__n29151, ys__n29153, ys__n29154, ys__n29156, ys__n29157, ys__n29159,
    ys__n29160, ys__n29162, ys__n29163, ys__n29165, ys__n29166, ys__n29168,
    ys__n29169, ys__n29171, ys__n29172, ys__n29174, ys__n29175, ys__n29177,
    ys__n29178, ys__n29180, ys__n29181, ys__n29183, ys__n29184, ys__n29186,
    ys__n29187, ys__n29189, ys__n29190, ys__n29192, ys__n29193, ys__n29195,
    ys__n29196, ys__n29198, ys__n29199, ys__n29201, ys__n29202, ys__n29204,
    ys__n29205, ys__n29207, ys__n29208, ys__n29210, ys__n29211, ys__n29213,
    ys__n29214, ys__n29218, ys__n29220, ys__n29224, ys__n29237, ys__n29240,
    ys__n29242, ys__n29244, ys__n29246, ys__n29248, ys__n29250, ys__n29252,
    ys__n29254, ys__n29256, ys__n29258, ys__n29260, ys__n29262, ys__n29264,
    ys__n29266, ys__n29268, ys__n29270, ys__n29272, ys__n29274, ys__n29276,
    ys__n29278, ys__n29280, ys__n29282, ys__n29284, ys__n29286, ys__n29288,
    ys__n29290, ys__n29292, ys__n29294, ys__n29296, ys__n29298, ys__n29300,
    ys__n29432, ys__n29433, ys__n29434, ys__n29436, ys__n29437, ys__n29439,
    ys__n29440, ys__n29442, ys__n29443, ys__n29445, ys__n29446, ys__n29448,
    ys__n29449, ys__n29451, ys__n29452, ys__n29454, ys__n29455, ys__n29457,
    ys__n29458, ys__n29460, ys__n29461, ys__n29463, ys__n29464, ys__n29466,
    ys__n29467, ys__n29469, ys__n29470, ys__n29472, ys__n29473, ys__n29475,
    ys__n29476, ys__n29478, ys__n29479, ys__n29481, ys__n29482, ys__n29484,
    ys__n29485, ys__n29487, ys__n29488, ys__n29490, ys__n29491, ys__n29493,
    ys__n29494, ys__n29496, ys__n29497, ys__n29499, ys__n29500, ys__n29502,
    ys__n29503, ys__n29505, ys__n29506, ys__n29508, ys__n29509, ys__n29511,
    ys__n29512, ys__n29514, ys__n29515, ys__n29517, ys__n29518, ys__n29520,
    ys__n29521, ys__n29523, ys__n29524, ys__n29526, ys__n29527, ys__n29531,
    ys__n29533, ys__n29537, ys__n29550, ys__n29552, ys__n29553, ys__n29554,
    ys__n29555, ys__n29556, ys__n29557, ys__n29558, ys__n29559, ys__n29560,
    ys__n29561, ys__n29562, ys__n29563, ys__n29564, ys__n29565, ys__n29566,
    ys__n29567, ys__n29568, ys__n29569, ys__n29570, ys__n29571, ys__n29572,
    ys__n29573, ys__n29574, ys__n29575, ys__n29576, ys__n29577, ys__n29578,
    ys__n29579, ys__n29580, ys__n29581, ys__n29582, ys__n29583, ys__n29584,
    ys__n29585, ys__n29586, ys__n29587, ys__n29588, ys__n29589, ys__n29590,
    ys__n29591, ys__n29592, ys__n29593, ys__n29594, ys__n29595, ys__n29596,
    ys__n29597, ys__n29598, ys__n29599, ys__n29600, ys__n29601, ys__n29602,
    ys__n29603, ys__n29604, ys__n29605, ys__n29606, ys__n29607, ys__n29608,
    ys__n29707, ys__n29708, ys__n29709, ys__n29711, ys__n29712, ys__n29714,
    ys__n29715, ys__n29717, ys__n29718, ys__n29720, ys__n29721, ys__n29723,
    ys__n29724, ys__n29726, ys__n29727, ys__n29729, ys__n29730, ys__n29732,
    ys__n29733, ys__n29735, ys__n29736, ys__n29738, ys__n29739, ys__n29741,
    ys__n29742, ys__n29744, ys__n29745, ys__n29747, ys__n29748, ys__n29750,
    ys__n29751, ys__n29753, ys__n29754, ys__n29756, ys__n29757, ys__n29759,
    ys__n29760, ys__n29762, ys__n29763, ys__n29765, ys__n29766, ys__n29768,
    ys__n29769, ys__n29771, ys__n29772, ys__n29774, ys__n29775, ys__n29777,
    ys__n29778, ys__n29780, ys__n29781, ys__n29783, ys__n29784, ys__n29786,
    ys__n29787, ys__n29789, ys__n29790, ys__n29792, ys__n29793, ys__n29795,
    ys__n29796, ys__n29798, ys__n29799, ys__n29801, ys__n29802, ys__n29806,
    ys__n29808, ys__n29812, ys__n29846, ys__n29880, ys__n29881, ys__n29883,
    ys__n29884, ys__n29885, ys__n29886, ys__n29887, ys__n29888, ys__n29889,
    ys__n29890, ys__n29891, ys__n29892, ys__n29893, ys__n29894, ys__n29895,
    ys__n29896, ys__n29897, ys__n29898, ys__n29899, ys__n29900, ys__n29901,
    ys__n29902, ys__n29903, ys__n29904, ys__n29905, ys__n29906, ys__n29907,
    ys__n29908, ys__n29909, ys__n29910, ys__n29911, ys__n29912, ys__n29913,
    ys__n30011, ys__n30014, ys__n30016, ys__n30018, ys__n30020, ys__n30022,
    ys__n30024, ys__n30026, ys__n30028, ys__n30030, ys__n30032, ys__n30034,
    ys__n30036, ys__n30038, ys__n30040, ys__n30042, ys__n30044, ys__n30046,
    ys__n30048, ys__n30050, ys__n30052, ys__n30054, ys__n30056, ys__n30058,
    ys__n30060, ys__n30062, ys__n30064, ys__n30066, ys__n30068, ys__n30070,
    ys__n30072, ys__n30074, ys__n30214, ys__n30216, ys__n30217, ys__n30219,
    ys__n30220, ys__n30225, ys__n30230, ys__n30232, ys__n30333, ys__n30334,
    ys__n30553, ys__n30815, ys__n30816, ys__n30818, ys__n30819, ys__n30820,
    ys__n30837, ys__n30861, ys__n30862, ys__n30863, ys__n30865, ys__n30867,
    ys__n30869, ys__n30871, ys__n30877, ys__n30879, ys__n30881, ys__n30883,
    ys__n30885, ys__n30887, ys__n30889, ys__n30891, ys__n30893, ys__n30895,
    ys__n30897, ys__n30899, ys__n30901, ys__n30903, ys__n30905, ys__n30907,
    ys__n30909, ys__n30911, ys__n30913, ys__n30915, ys__n30917, ys__n30919,
    ys__n30921, ys__n30923, ys__n30925, ys__n30927, ys__n30929, ys__n30931,
    ys__n30933, ys__n30935, ys__n30937, ys__n30939, ys__n30941, ys__n30957,
    ys__n30960, ys__n30961, ys__n30962, ys__n30974, ys__n31031, ys__n33212,
    ys__n33214, ys__n33216, ys__n33218, ys__n33220, ys__n33222, ys__n33259,
    ys__n33261, ys__n33263, ys__n33265, ys__n33267, ys__n33269, ys__n33272,
    ys__n33274, ys__n33276, ys__n33278, ys__n33300, ys__n33309, ys__n33311,
    ys__n33313, ys__n33318, ys__n33320, ys__n33328, ys__n33330, ys__n33332,
    ys__n33334, ys__n33336, ys__n33338, ys__n33340, ys__n33342, ys__n33350,
    ys__n33352, ys__n33359, ys__n33364, ys__n33370, ys__n33375, ys__n33380,
    ys__n33384, ys__n33386, ys__n33389, ys__n33394, ys__n33396, ys__n33398,
    ys__n33403, ys__n33407, ys__n33409, ys__n33411, ys__n33423, ys__n33431,
    ys__n33442, ys__n33451, ys__n33464, ys__n33469, ys__n33471, ys__n33473,
    ys__n33475, ys__n33479, ys__n33481, ys__n33488, ys__n33491, ys__n33493,
    ys__n33495, ys__n33497, ys__n33499, ys__n33509, ys__n33511, ys__n33522,
    ys__n33532, ys__n33541, ys__n33545, ys__n33548, ys__n33552, ys__n33558,
    ys__n33563, ys__n33564, ys__n33566, ys__n33568, ys__n33570, ys__n33572,
    ys__n33574, ys__n33576, ys__n33579, ys__n33581, ys__n33614, ys__n33632,
    ys__n33634, ys__n33636, ys__n33638, ys__n33640, ys__n33642, ys__n33644,
    ys__n33646, ys__n33648, ys__n33650, ys__n33652, ys__n33654, ys__n33656,
    ys__n33658, ys__n33660, ys__n33662, ys__n33664, ys__n33666, ys__n33668,
    ys__n33670, ys__n33672, ys__n33674, ys__n33676, ys__n33678, ys__n33681,
    ys__n33683, ys__n33685, ys__n33687, ys__n33689, ys__n33691, ys__n33693,
    ys__n33695, ys__n33697, ys__n33699, ys__n33701, ys__n33703, ys__n33705,
    ys__n33707, ys__n33709, ys__n33711, ys__n33713, ys__n33715, ys__n33717,
    ys__n33719, ys__n33721, ys__n33723, ys__n33725, ys__n33727, ys__n33729,
    ys__n33731, ys__n33733, ys__n33735, ys__n33737, ys__n33739, ys__n33741,
    ys__n33743, ys__n33745, ys__n33747, ys__n33749, ys__n34666, ys__n34668,
    ys__n34670, ys__n34672, ys__n34674, ys__n34676, ys__n34678, ys__n34680,
    ys__n34682, ys__n34684, ys__n34686, ys__n34688, ys__n34690, ys__n34692,
    ys__n34694, ys__n34696, ys__n34698, ys__n34700, ys__n34702, ys__n34704,
    ys__n34706, ys__n34708, ys__n34710, ys__n34712, ys__n34714, ys__n34716,
    ys__n34718, ys__n34720, ys__n34722, ys__n34724, ys__n34726, ys__n34728,
    ys__n34730, ys__n34732, ys__n34734, ys__n34736, ys__n34738, ys__n34740,
    ys__n34742, ys__n34744, ys__n34746, ys__n34748, ys__n34750, ys__n34752,
    ys__n34754, ys__n34756, ys__n34758, ys__n34760, ys__n34762, ys__n34764,
    ys__n34766, ys__n34768, ys__n34770, ys__n34772, ys__n34774, ys__n34776,
    ys__n34778, ys__n34780, ys__n34782, ys__n34784, ys__n34786, ys__n34788,
    ys__n34790, ys__n34792, ys__n34794, ys__n34796, ys__n34798, ys__n34800,
    ys__n34802, ys__n34804, ys__n34806, ys__n34808, ys__n34810, ys__n34812,
    ys__n34814, ys__n34816, ys__n34818, ys__n34820, ys__n34822, ys__n34824,
    ys__n34826, ys__n34828, ys__n34830, ys__n34832, ys__n34834, ys__n34836,
    ys__n34838, ys__n34840, ys__n34842, ys__n34844, ys__n34846, ys__n34848,
    ys__n34850, ys__n34852, ys__n34854, ys__n34856, ys__n34858, ys__n34860,
    ys__n34862, ys__n34864, ys__n34866, ys__n34868, ys__n34870, ys__n34872,
    ys__n34874, ys__n34876, ys__n34878, ys__n34880, ys__n34882, ys__n34884,
    ys__n34886, ys__n34888, ys__n34890, ys__n34892, ys__n34894, ys__n34896,
    ys__n34898, ys__n34900, ys__n34902, ys__n34904, ys__n34906, ys__n34908,
    ys__n34910, ys__n34912, ys__n34914, ys__n34916, ys__n34918, ys__n34920,
    ys__n34922, ys__n34924, ys__n34926, ys__n34928, ys__n34930, ys__n34932,
    ys__n34934, ys__n34936, ys__n34938, ys__n34940, ys__n34942, ys__n34944,
    ys__n34946, ys__n34948, ys__n34950, ys__n34959, ys__n34966, ys__n34972,
    ys__n34976, ys__n34978, ys__n34984, ys__n34988, ys__n34990, ys__n34996,
    ys__n35000, ys__n35002, ys__n35008, ys__n35012, ys__n35014, ys__n35020,
    ys__n35024, ys__n35026, ys__n35028, ys__n35031, ys__n35033, ys__n35035,
    ys__n35037, ys__n35039, ys__n35041, ys__n35047, ys__n35049, ys__n35057,
    ys__n35059, ys__n35065, ys__n35076, ys__n35078, ys__n35080, ys__n35082,
    ys__n35084, ys__n35086, ys__n35088, ys__n35090, ys__n35092, ys__n35094,
    ys__n35096, ys__n35098, ys__n35102, ys__n35104, ys__n35106, ys__n35108,
    ys__n35110, ys__n35112, ys__n35114, ys__n35116, ys__n35118, ys__n35120,
    ys__n35122, ys__n35124, ys__n35413, ys__n35415, ys__n35417, ys__n35419,
    ys__n35421, ys__n35423, ys__n35426, ys__n35704, ys__n35717, ys__n35719,
    ys__n35721, ys__n35723, ys__n35725, ys__n35727, ys__n37668, ys__n37669,
    ys__n37670, ys__n37671, ys__n37672, ys__n37673, ys__n37674, ys__n37675,
    ys__n37678, ys__n37679, ys__n37682, ys__n37692, ys__n37694, ys__n37696,
    ys__n37710, ys__n37712, ys__n37713, ys__n37743, ys__n37744, ys__n37745,
    ys__n37746, ys__n37747, ys__n37748, ys__n37749, ys__n37750, ys__n37751,
    ys__n37752, ys__n37753, ys__n37754, ys__n37755, ys__n37756, ys__n37757,
    ys__n37758, ys__n37759, ys__n37760, ys__n37761, ys__n37762, ys__n37763,
    ys__n37764, ys__n37765, ys__n37766, ys__n37767, ys__n37768, ys__n37769,
    ys__n37770, ys__n37771, ys__n37772, ys__n37773, ys__n37774, ys__n37775,
    ys__n37776, ys__n37777, ys__n37778, ys__n37779, ys__n37780, ys__n37781,
    ys__n37782, ys__n37783, ys__n37784, ys__n37785, ys__n37786, ys__n37787,
    ys__n37788, ys__n37789, ys__n37790, ys__n37791, ys__n37792, ys__n37793,
    ys__n37794, ys__n37795, ys__n37796, ys__n37797, ys__n37798, ys__n37799,
    ys__n37800, ys__n37801, ys__n37802, ys__n37803, ys__n37804, ys__n37805,
    ys__n37806, ys__n37807, ys__n37808, ys__n37809, ys__n37810, ys__n37811,
    ys__n37812, ys__n37813, ys__n37814, ys__n37815, ys__n37816, ys__n37817,
    ys__n37818, ys__n37819, ys__n37820, ys__n37821, ys__n37822, ys__n37823,
    ys__n37824, ys__n37825, ys__n37826, ys__n37827, ys__n37828, ys__n37829,
    ys__n37830, ys__n37831, ys__n37832, ys__n37833, ys__n37834, ys__n37835,
    ys__n37836, ys__n37837, ys__n37838, ys__n37839, ys__n37840, ys__n37841,
    ys__n37842, ys__n37843, ys__n37844, ys__n37845, ys__n37846, ys__n37847,
    ys__n37848, ys__n37849, ys__n37850, ys__n37851, ys__n37852, ys__n37853,
    ys__n37854, ys__n37855, ys__n37856, ys__n37857, ys__n37858, ys__n37859,
    ys__n37860, ys__n37861, ys__n37862, ys__n37863, ys__n37864, ys__n37865,
    ys__n37866, ys__n37867, ys__n37868, ys__n37869, ys__n37870, ys__n37871,
    ys__n37872, ys__n37873, ys__n37874, ys__n37875, ys__n37876, ys__n37877,
    ys__n37878, ys__n37879, ys__n37880, ys__n37881, ys__n37882, ys__n37883,
    ys__n37884, ys__n37885, ys__n37886, ys__n37887, ys__n37888, ys__n37889,
    ys__n37890, ys__n37891, ys__n37892, ys__n37893, ys__n37894, ys__n37895,
    ys__n37896, ys__n37897, ys__n37898, ys__n37899, ys__n37900, ys__n37901,
    ys__n37902, ys__n37903, ys__n37904, ys__n37905, ys__n37906, ys__n37907,
    ys__n37908, ys__n37909, ys__n37910, ys__n37911, ys__n37912, ys__n37913,
    ys__n37914, ys__n37915, ys__n37916, ys__n37917, ys__n37918, ys__n37919,
    ys__n37920, ys__n37921, ys__n37922, ys__n37923, ys__n37924, ys__n37925,
    ys__n37926, ys__n37927, ys__n37928, ys__n37929, ys__n37930, ys__n37931,
    ys__n37932, ys__n37933, ys__n37934, ys__n37935, ys__n37936, ys__n37937,
    ys__n37938, ys__n37939, ys__n37940, ys__n37941, ys__n37942, ys__n37943,
    ys__n37944, ys__n37945, ys__n37946, ys__n37947, ys__n37948, ys__n37949,
    ys__n37950, ys__n37951, ys__n37952, ys__n37953, ys__n37954, ys__n37955,
    ys__n37956, ys__n37957, ys__n37958, ys__n37959, ys__n37960, ys__n37961,
    ys__n37962, ys__n37963, ys__n37964, ys__n37965, ys__n37966, ys__n37967,
    ys__n37968, ys__n37969, ys__n37970, ys__n37971, ys__n37972, ys__n37973,
    ys__n37974, ys__n37975, ys__n37976, ys__n37977, ys__n37978, ys__n37979,
    ys__n37980, ys__n37981, ys__n37982, ys__n37983, ys__n37984, ys__n37985,
    ys__n37986, ys__n37987, ys__n37988, ys__n37989, ys__n37990, ys__n37991,
    ys__n37992, ys__n37993, ys__n37994, ys__n37995, ys__n37996, ys__n37997,
    ys__n37998, ys__n37999, ys__n38000, ys__n38001, ys__n38002, ys__n38003,
    ys__n38004, ys__n38005, ys__n38006, ys__n38007, ys__n38008, ys__n38009,
    ys__n38010, ys__n38011, ys__n38012, ys__n38013, ys__n38014, ys__n38015,
    ys__n38016, ys__n38017, ys__n38018, ys__n38019, ys__n38020, ys__n38021,
    ys__n38022, ys__n38023, ys__n38024, ys__n38025, ys__n38026, ys__n38027,
    ys__n38028, ys__n38029, ys__n38030, ys__n38031, ys__n38032, ys__n38033,
    ys__n38034, ys__n38035, ys__n38036, ys__n38037, ys__n38038, ys__n38039,
    ys__n38040, ys__n38041, ys__n38042, ys__n38043, ys__n38044, ys__n38045,
    ys__n38046, ys__n38047, ys__n38048, ys__n38049, ys__n38050, ys__n38051,
    ys__n38052, ys__n38053, ys__n38054, ys__n38055, ys__n38056, ys__n38057,
    ys__n38058, ys__n38059, ys__n38060, ys__n38061, ys__n38062, ys__n38063,
    ys__n38064, ys__n38065, ys__n38066, ys__n38067, ys__n38068, ys__n38069,
    ys__n38070, ys__n38071, ys__n38072, ys__n38073, ys__n38074, ys__n38075,
    ys__n38076, ys__n38077, ys__n38078, ys__n38079, ys__n38080, ys__n38081,
    ys__n38082, ys__n38083, ys__n38084, ys__n38085, ys__n38086, ys__n38087,
    ys__n38088, ys__n38089, ys__n38090, ys__n38091, ys__n38092, ys__n38093,
    ys__n38094, ys__n38095, ys__n38096, ys__n38097, ys__n38098, ys__n38099,
    ys__n38100, ys__n38101, ys__n38102, ys__n38103, ys__n38104, ys__n38105,
    ys__n38106, ys__n38107, ys__n38108, ys__n38109, ys__n38110, ys__n38111,
    ys__n38112, ys__n38113, ys__n38114, ys__n38115, ys__n38116, ys__n38117,
    ys__n38118, ys__n38119, ys__n38120, ys__n38121, ys__n38122, ys__n38123,
    ys__n38124, ys__n38125, ys__n38126, ys__n38127, ys__n38128, ys__n38129,
    ys__n38130, ys__n38131, ys__n38132, ys__n38133, ys__n38134, ys__n38135,
    ys__n38136, ys__n38137, ys__n38138, ys__n38139, ys__n38140, ys__n38141,
    ys__n38142, ys__n38143, ys__n38144, ys__n38145, ys__n38146, ys__n38147,
    ys__n38148, ys__n38149, ys__n38150, ys__n38151, ys__n38152, ys__n38153,
    ys__n38154, ys__n38155, ys__n38156, ys__n38157, ys__n38158, ys__n38159,
    ys__n38160, ys__n38161, ys__n38162, ys__n38163, ys__n38164, ys__n38165,
    ys__n38166, ys__n38167, ys__n38168, ys__n38169, ys__n38170, ys__n38171,
    ys__n38172, ys__n38173, ys__n38174, ys__n38175, ys__n38176, ys__n38177,
    ys__n38178, ys__n38179, ys__n38183, ys__n38192, ys__n38193, ys__n38194,
    ys__n38195, ys__n38196, ys__n38197, ys__n38198, ys__n38199, ys__n38200,
    ys__n38201, ys__n38202, ys__n38203, ys__n38212, ys__n38215, ys__n38217,
    ys__n38219, ys__n38220, ys__n38221, ys__n38236, ys__n38237, ys__n38257,
    ys__n38259, ys__n38272, ys__n38277, ys__n38278, ys__n38279, ys__n38282,
    ys__n38283, ys__n38286, ys__n38288, ys__n38290, ys__n38291, ys__n38300,
    ys__n38304, ys__n38305, ys__n38307, ys__n38311, ys__n38315, ys__n38320,
    ys__n38323, ys__n38346, ys__n38361, ys__n38376, ys__n38378, ys__n38380,
    ys__n38382, ys__n38384, ys__n38386, ys__n38398, ys__n38407, ys__n38408,
    ys__n38413, ys__n38418, ys__n38420, ys__n38424, ys__n38427, ys__n38437,
    ys__n38438, ys__n38441, ys__n38443, ys__n38448, ys__n38449, ys__n38451,
    ys__n38473, ys__n38486, ys__n38487, ys__n38488, ys__n38489, ys__n38490,
    ys__n38491, ys__n38494, ys__n38495, ys__n38496, ys__n38497, ys__n38498,
    ys__n38499, ys__n38502, ys__n38503, ys__n38504, ys__n38505, ys__n38506,
    ys__n38507, ys__n38513, ys__n38522, ys__n38524, ys__n38526, ys__n38527,
    ys__n38528, ys__n38529, ys__n38553, ys__n38557, ys__n38561, ys__n38564,
    ys__n38565, ys__n38567, ys__n38568, ys__n38569, ys__n38585, ys__n38586,
    ys__n38587, ys__n38588, ys__n38589, ys__n38590, ys__n38591, ys__n38592,
    ys__n38593, ys__n38594, ys__n38595, ys__n38596, ys__n38597, ys__n38598,
    ys__n38599, ys__n38600, ys__n38601, ys__n38602, ys__n38603, ys__n38604,
    ys__n38605, ys__n38606, ys__n38607, ys__n38608, ys__n38609, ys__n38610,
    ys__n38611, ys__n38620, ys__n38624, ys__n38631, ys__n38649, ys__n38654,
    ys__n38670, ys__n38680, ys__n38693, ys__n38694, ys__n38695, ys__n38724,
    ys__n38776, ys__n38777, ys__n38805, ys__n38827, ys__n38828, ys__n38829,
    ys__n38830, ys__n38831, ys__n38832, ys__n38833, ys__n38834, ys__n38835,
    ys__n38836, ys__n38837, ys__n38838, ys__n38839, ys__n38840, ys__n38841,
    ys__n38842, ys__n38843, ys__n38844, ys__n38845, ys__n38846, ys__n38847,
    ys__n38848, ys__n38849, ys__n38850, ys__n38851, ys__n38852, ys__n38853,
    ys__n38854, ys__n38855, ys__n38856, ys__n38857, ys__n38858, ys__n38859,
    ys__n38861, ys__n38862, ys__n38863, ys__n38864, ys__n38865, ys__n38883,
    ys__n38885, ys__n38893, ys__n38894, ys__n38896, ys__n38897, ys__n38898,
    ys__n38902, ys__n38904, ys__n38906, ys__n38908, ys__n38910, ys__n38919,
    ys__n38922, ys__n38927, ys__n38928, ys__n38929, ys__n39167, ys__n39518,
    ys__n39520, ys__n39718, ys__n39720, ys__n39722, ys__n39724, ys__n39726,
    ys__n39728, ys__n39730, ys__n39732, ys__n39734, ys__n39736, ys__n39738,
    ys__n39740, ys__n39742, ys__n39744, ys__n39746, ys__n39748, ys__n39750,
    ys__n39752, ys__n39754, ys__n39756, ys__n39758, ys__n39760, ys__n39762,
    ys__n39764, ys__n39766, ys__n39768, ys__n39770, ys__n39772, ys__n39774,
    ys__n39776, ys__n39778, ys__n44833, ys__n44840, ys__n44842, ys__n44847,
    ys__n44849, ys__n44892, ys__n44906, ys__n44907, ys__n44908, ys__n44988,
    ys__n44989, ys__n44990, ys__n44991, ys__n44992, ys__n44993, ys__n44995,
    ys__n44996, ys__n44998, ys__n44999, ys__n45001, ys__n45002, ys__n45004,
    ys__n45005, ys__n45007, ys__n45008, ys__n45010, ys__n45011, ys__n45013,
    ys__n45014, ys__n45016, ys__n45017, ys__n45019, ys__n45020, ys__n45022,
    ys__n45023, ys__n45025, ys__n45026, ys__n45028, ys__n45029, ys__n45031,
    ys__n45032, ys__n45034, ys__n45035, ys__n45037, ys__n45038, ys__n45040,
    ys__n45041, ys__n45043, ys__n45044, ys__n45046, ys__n45047, ys__n45049,
    ys__n45050, ys__n45052, ys__n45053, ys__n45055, ys__n45056, ys__n45058,
    ys__n45059, ys__n45061, ys__n45062, ys__n45064, ys__n45065, ys__n45067,
    ys__n45068, ys__n45070, ys__n45071, ys__n45073, ys__n45074, ys__n45076,
    ys__n45077, ys__n45079, ys__n45080, ys__n45082, ys__n45083, ys__n45084,
    ys__n45085, ys__n45086, ys__n45087, ys__n45088, ys__n45089, ys__n45090,
    ys__n45091, ys__n45092, ys__n45093, ys__n45094, ys__n45095, ys__n45096,
    ys__n45097, ys__n45098, ys__n45099, ys__n45100, ys__n45101, ys__n45102,
    ys__n45103, ys__n45104, ys__n45105, ys__n45106, ys__n45107, ys__n45108,
    ys__n45109, ys__n45110, ys__n45111, ys__n45112, ys__n45113, ys__n45115,
    ys__n45116, ys__n45118, ys__n45119, ys__n45121, ys__n45122, ys__n45124,
    ys__n45125, ys__n45127, ys__n45128, ys__n45130, ys__n45131, ys__n45133,
    ys__n45134, ys__n45136, ys__n45137, ys__n45139, ys__n45140, ys__n45142,
    ys__n45143, ys__n45145, ys__n45146, ys__n45148, ys__n45149, ys__n45151,
    ys__n45152, ys__n45154, ys__n45155, ys__n45157, ys__n45158, ys__n45160,
    ys__n45161, ys__n45163, ys__n45164, ys__n45166, ys__n45167, ys__n45169,
    ys__n45170, ys__n45172, ys__n45173, ys__n45175, ys__n45176, ys__n45178,
    ys__n45179, ys__n45181, ys__n45182, ys__n45184, ys__n45185, ys__n45187,
    ys__n45188, ys__n45190, ys__n45191, ys__n45193, ys__n45194, ys__n45196,
    ys__n45197, ys__n45199, ys__n45200, ys__n45202, ys__n45203, ys__n45205,
    ys__n45206, ys__n45208, ys__n45209, ys__n45210, ys__n45211, ys__n45212,
    ys__n45214, ys__n45216, ys__n45218, ys__n45220, ys__n45222, ys__n45224,
    ys__n45226, ys__n45228, ys__n45230, ys__n45232, ys__n45234, ys__n45236,
    ys__n45238, ys__n45240, ys__n45242, ys__n45244, ys__n45246, ys__n45248,
    ys__n45250, ys__n45252, ys__n45254, ys__n45256, ys__n45258, ys__n45260,
    ys__n45262, ys__n45264, ys__n45266, ys__n45268, ys__n45270, ys__n45272,
    ys__n45274, ys__n45276, ys__n45277, ys__n45278, ys__n45279, ys__n45280,
    ys__n45281, ys__n45282, ys__n45283, ys__n45284, ys__n45285, ys__n45286,
    ys__n45287, ys__n45288, ys__n45289, ys__n45290, ys__n45291, ys__n45292,
    ys__n45293, ys__n45294, ys__n45295, ys__n45296, ys__n45297, ys__n45298,
    ys__n45299, ys__n45300, ys__n45301, ys__n45302, ys__n45303, ys__n45304,
    ys__n45305, ys__n45306, ys__n45308, ys__n45310, ys__n45312, ys__n45314,
    ys__n45316, ys__n45318, ys__n45320, ys__n45322, ys__n45324, ys__n45326,
    ys__n45328, ys__n45330, ys__n45332, ys__n45334, ys__n45336, ys__n45338,
    ys__n45340, ys__n45342, ys__n45344, ys__n45346, ys__n45348, ys__n45350,
    ys__n45352, ys__n45354, ys__n45356, ys__n45358, ys__n45360, ys__n45362,
    ys__n45364, ys__n45366, ys__n45368, ys__n45370, ys__n45371, ys__n45372,
    ys__n45373, ys__n45374, ys__n45377, ys__n45380, ys__n45382, ys__n45384,
    ys__n45386, ys__n45388, ys__n45390, ys__n45392, ys__n45394, ys__n45396,
    ys__n45398, ys__n45400, ys__n45402, ys__n45404, ys__n45406, ys__n45408,
    ys__n45410, ys__n45412, ys__n45414, ys__n45416, ys__n45418, ys__n45420,
    ys__n45422, ys__n45424, ys__n45426, ys__n45428, ys__n45430, ys__n45432,
    ys__n45434, ys__n45436, ys__n45438, ys__n45440, ys__n45441, ys__n45442,
    ys__n45443, ys__n45444, ys__n45445, ys__n45446, ys__n45447, ys__n45448,
    ys__n45449, ys__n45450, ys__n45451, ys__n45452, ys__n45453, ys__n45454,
    ys__n45455, ys__n45456, ys__n45457, ys__n45458, ys__n45459, ys__n45460,
    ys__n45461, ys__n45462, ys__n45463, ys__n45464, ys__n45465, ys__n45466,
    ys__n45467, ys__n45468, ys__n45469, ys__n45470, ys__n45472, ys__n45474,
    ys__n45476, ys__n45478, ys__n45480, ys__n45482, ys__n45484, ys__n45486,
    ys__n45488, ys__n45490, ys__n45492, ys__n45494, ys__n45496, ys__n45498,
    ys__n45500, ys__n45502, ys__n45504, ys__n45506, ys__n45508, ys__n45510,
    ys__n45512, ys__n45514, ys__n45516, ys__n45518, ys__n45520, ys__n45522,
    ys__n45524, ys__n45526, ys__n45528, ys__n45530, ys__n45532, ys__n45534,
    ys__n45535, ys__n45536, ys__n45537, ys__n45538, ys__n45541, ys__n45544,
    ys__n45546, ys__n45548, ys__n45550, ys__n45552, ys__n45554, ys__n45556,
    ys__n45558, ys__n45560, ys__n45562, ys__n45564, ys__n45566, ys__n45568,
    ys__n45570, ys__n45572, ys__n45574, ys__n45576, ys__n45578, ys__n45580,
    ys__n45582, ys__n45584, ys__n45586, ys__n45588, ys__n45590, ys__n45592,
    ys__n45594, ys__n45596, ys__n45598, ys__n45600, ys__n45602, ys__n45604,
    ys__n45605, ys__n45606, ys__n45607, ys__n45608, ys__n45609, ys__n45610,
    ys__n45611, ys__n45612, ys__n45613, ys__n45614, ys__n45615, ys__n45616,
    ys__n45617, ys__n45618, ys__n45619, ys__n45620, ys__n45621, ys__n45622,
    ys__n45623, ys__n45624, ys__n45625, ys__n45626, ys__n45627, ys__n45628,
    ys__n45629, ys__n45630, ys__n45631, ys__n45632, ys__n45633, ys__n45634,
    ys__n45636, ys__n45638, ys__n45640, ys__n45642, ys__n45644, ys__n45646,
    ys__n45648, ys__n45650, ys__n45652, ys__n45654, ys__n45656, ys__n45658,
    ys__n45660, ys__n45662, ys__n45664, ys__n45666, ys__n45668, ys__n45670,
    ys__n45672, ys__n45674, ys__n45676, ys__n45678, ys__n45680, ys__n45682,
    ys__n45684, ys__n45686, ys__n45688, ys__n45690, ys__n45692, ys__n45694,
    ys__n45696, ys__n45698, ys__n45699, ys__n45700, ys__n45701, ys__n45702,
    ys__n45704, ys__n45707, ys__n45708, ys__n45709, ys__n45710, ys__n45711,
    ys__n45712, ys__n45714, ys__n45715, ys__n45717, ys__n45718, ys__n45720,
    ys__n45721, ys__n45723, ys__n45724, ys__n45726, ys__n45727, ys__n45729,
    ys__n45730, ys__n45732, ys__n45733, ys__n45735, ys__n45736, ys__n45738,
    ys__n45739, ys__n45741, ys__n45742, ys__n45744, ys__n45745, ys__n45747,
    ys__n45748, ys__n45750, ys__n45751, ys__n45753, ys__n45754, ys__n45756,
    ys__n45757, ys__n45759, ys__n45760, ys__n45762, ys__n45763, ys__n45765,
    ys__n45766, ys__n45768, ys__n45769, ys__n45771, ys__n45772, ys__n45774,
    ys__n45775, ys__n45777, ys__n45778, ys__n45780, ys__n45781, ys__n45783,
    ys__n45784, ys__n45786, ys__n45787, ys__n45789, ys__n45790, ys__n45792,
    ys__n45793, ys__n45795, ys__n45796, ys__n45798, ys__n45799, ys__n45801,
    ys__n45802, ys__n45804, ys__n45805, ys__n45806, ys__n45807, ys__n45808,
    ys__n45809, ys__n45810, ys__n45811, ys__n45812, ys__n45813, ys__n45814,
    ys__n45815, ys__n45816, ys__n45817, ys__n45818, ys__n45819, ys__n45820,
    ys__n45821, ys__n45822, ys__n45823, ys__n45824, ys__n45825, ys__n45826,
    ys__n45827, ys__n45828, ys__n45829, ys__n45830, ys__n45831, ys__n45832,
    ys__n45833, ys__n45834, ys__n45835, ys__n45836, ys__n45838, ys__n45840,
    ys__n45842, ys__n45844, ys__n45846, ys__n45848, ys__n45850, ys__n45852,
    ys__n45854, ys__n45856, ys__n45858, ys__n45860, ys__n45862, ys__n45864,
    ys__n45866, ys__n45868, ys__n45870, ys__n45872, ys__n45874, ys__n45876,
    ys__n45878, ys__n45880, ys__n45882, ys__n45884, ys__n45886, ys__n45888,
    ys__n45890, ys__n45892, ys__n45894, ys__n45896, ys__n45898, ys__n45900,
    ys__n45901, ys__n45902, ys__n45903, ys__n45904, ys__n45905, ys__n45906,
    ys__n45907, ys__n45908, ys__n45909, ys__n45910, ys__n45911, ys__n45912,
    ys__n45913, ys__n45914, ys__n45915, ys__n45916, ys__n45917, ys__n45918,
    ys__n45919, ys__n45920, ys__n45921, ys__n45922, ys__n45923, ys__n45924,
    ys__n45925, ys__n45926, ys__n45927, ys__n45928, ys__n45929, ys__n45930,
    ys__n45931, ys__n45933, ys__n45936, ys__n45938, ys__n45940, ys__n45942,
    ys__n45944, ys__n45946, ys__n45948, ys__n45950, ys__n45952, ys__n45954,
    ys__n45956, ys__n45958, ys__n45960, ys__n45962, ys__n45964, ys__n45966,
    ys__n45968, ys__n45970, ys__n45972, ys__n45974, ys__n45976, ys__n45978,
    ys__n45980, ys__n45982, ys__n45984, ys__n45986, ys__n45988, ys__n45990,
    ys__n45992, ys__n45994, ys__n45996, ys__n45998, ys__n45999, ys__n46000,
    ys__n46001, ys__n46002, ys__n46003, ys__n46004, ys__n46005, ys__n46006,
    ys__n46007, ys__n46008, ys__n46009, ys__n46010, ys__n46011, ys__n46012,
    ys__n46013, ys__n46014, ys__n46015, ys__n46016, ys__n46017, ys__n46018,
    ys__n46019, ys__n46020, ys__n46021, ys__n46022, ys__n46023, ys__n46024,
    ys__n46025, ys__n46026, ys__n46027, ys__n46028, ys__n46029, ys__n46031,
    ys__n46034, ys__n46036, ys__n46038, ys__n46040, ys__n46042, ys__n46044,
    ys__n46046, ys__n46048, ys__n46050, ys__n46052, ys__n46054, ys__n46056,
    ys__n46058, ys__n46060, ys__n46062, ys__n46064, ys__n46066, ys__n46068,
    ys__n46070, ys__n46072, ys__n46074, ys__n46076, ys__n46078, ys__n46080,
    ys__n46082, ys__n46084, ys__n46086, ys__n46088, ys__n46090, ys__n46092,
    ys__n46094, ys__n46096, ys__n46097, ys__n46098, ys__n46099, ys__n46100,
    ys__n46101, ys__n46102, ys__n46103, ys__n46104, ys__n46105, ys__n46106,
    ys__n46107, ys__n46108, ys__n46109, ys__n46110, ys__n46111, ys__n46112,
    ys__n46113, ys__n46114, ys__n46115, ys__n46116, ys__n46117, ys__n46118,
    ys__n46119, ys__n46120, ys__n46121, ys__n46122, ys__n46123, ys__n46124,
    ys__n46125, ys__n46126, ys__n46127, ys__n46128, ys__n46130, ys__n46132,
    ys__n46134, ys__n46136, ys__n46141, ys__n46142, ys__n46150, ys__n46151,
    ys__n46152, ys__n46153, ys__n46166, ys__n46168, ys__n46169, ys__n46170,
    ys__n46171, ys__n46180, ys__n46184, ys__n46185, ys__n46186, ys__n46187,
    ys__n46198, ys__n46200, ys__n46201, ys__n46202, ys__n46203, ys__n46214,
    ys__n46216, ys__n46217, ys__n46218, ys__n46219, ys__n46230, ys__n46231,
    ys__n46238, ys__n46239, ys__n46240, ys__n46242, ys__n46244, ys__n46245,
    ys__n46247, ys__n46248, ys__n46252, ys__n46254, ys__n46256, ys__n46258,
    ys__n46260, ys__n46262, ys__n46264, ys__n46266, ys__n46268, ys__n46270,
    ys__n46272, ys__n46274, ys__n46276, ys__n46278, ys__n46280, ys__n46282,
    ys__n46284, ys__n46286, ys__n46288, ys__n46290, ys__n46292, ys__n46294,
    ys__n46296, ys__n46298, ys__n46300, ys__n46302, ys__n46304, ys__n46306,
    ys__n46308, ys__n46310, ys__n46312, ys__n46314, ys__n46315, ys__n46316,
    ys__n46317, ys__n46318, ys__n46319, ys__n46320, ys__n46321, ys__n46322,
    ys__n46323, ys__n46324, ys__n46325, ys__n46326, ys__n46327, ys__n46328,
    ys__n46329, ys__n46330, ys__n46331, ys__n46332, ys__n46333, ys__n46334,
    ys__n46335, ys__n46336, ys__n46337, ys__n46338, ys__n46339, ys__n46340,
    ys__n46341, ys__n46342, ys__n46343, ys__n46344, ys__n46345, ys__n46346,
    ys__n46348, ys__n46350, ys__n46352, ys__n46354, ys__n46356, ys__n46358,
    ys__n46360, ys__n46362, ys__n46364, ys__n46366, ys__n46368, ys__n46370,
    ys__n46372, ys__n46374, ys__n46376, ys__n46378, ys__n46380, ys__n46382,
    ys__n46384, ys__n46386, ys__n46388, ys__n46390, ys__n46392, ys__n46393,
    ys__n46394, ys__n46395, ys__n46396, ys__n46397, ys__n46398, ys__n46399,
    ys__n46400, ys__n46401, ys__n46402, ys__n46403, ys__n46404, ys__n46405,
    ys__n46406, ys__n46407, ys__n46408, ys__n46409, ys__n46410, ys__n46411,
    ys__n46412, ys__n46413, ys__n46414, ys__n46415, ys__n46416, ys__n46417,
    ys__n46418, ys__n46419, ys__n46420, ys__n46421, ys__n46422, ys__n46423,
    ys__n46428, ys__n46430, ys__n46432, ys__n46434, ys__n46436, ys__n46438,
    ys__n46440, ys__n46442, ys__n46444, ys__n46446, ys__n46448, ys__n46450,
    ys__n46452, ys__n46454, ys__n46456, ys__n46458, ys__n46460, ys__n46462,
    ys__n46464, ys__n46466, ys__n46468, ys__n46470, ys__n46472, ys__n46474,
    ys__n46476, ys__n46478, ys__n46480, ys__n46482, ys__n46484, ys__n46486,
    ys__n46488, ys__n46490, ys__n46491, ys__n46492, ys__n46493, ys__n46494,
    ys__n46495, ys__n46496, ys__n46497, ys__n46498, ys__n46499, ys__n46500,
    ys__n46501, ys__n46502, ys__n46503, ys__n46504, ys__n46505, ys__n46506,
    ys__n46507, ys__n46508, ys__n46509, ys__n46510, ys__n46511, ys__n46512,
    ys__n46513, ys__n46514, ys__n46515, ys__n46516, ys__n46517, ys__n46518,
    ys__n46519, ys__n46520, ys__n46521, ys__n46522, ys__n46524, ys__n46526,
    ys__n46528, ys__n46530, ys__n46532, ys__n46534, ys__n46536, ys__n46538,
    ys__n46540, ys__n46542, ys__n46544, ys__n46546, ys__n46548, ys__n46550,
    ys__n46552, ys__n46554, ys__n46556, ys__n46558, ys__n46560, ys__n46562,
    ys__n46564, ys__n46566, ys__n46568, ys__n46569, ys__n46570, ys__n46571,
    ys__n46572, ys__n46573, ys__n46574, ys__n46575, ys__n46576, ys__n46577,
    ys__n46578, ys__n46579, ys__n46580, ys__n46581, ys__n46582, ys__n46583,
    ys__n46584, ys__n46585, ys__n46586, ys__n46587, ys__n46588, ys__n46589,
    ys__n46590, ys__n46591, ys__n46592, ys__n46593, ys__n46594, ys__n46595,
    ys__n46596, ys__n46597, ys__n46598, ys__n46599, ys__n46604, ys__n46606,
    ys__n46608, ys__n46610, ys__n46612, ys__n46614, ys__n46616, ys__n46618,
    ys__n46620, ys__n46622, ys__n46624, ys__n46626, ys__n46628, ys__n46630,
    ys__n46632, ys__n46634, ys__n46636, ys__n46638, ys__n46640, ys__n46642,
    ys__n46644, ys__n46646, ys__n46648, ys__n46650, ys__n46652, ys__n46654,
    ys__n46656, ys__n46658, ys__n46660, ys__n46662, ys__n46664, ys__n46666,
    ys__n46667, ys__n46668, ys__n46669, ys__n46670, ys__n46671, ys__n46672,
    ys__n46673, ys__n46674, ys__n46675, ys__n46676, ys__n46677, ys__n46678,
    ys__n46679, ys__n46680, ys__n46681, ys__n46682, ys__n46683, ys__n46684,
    ys__n46685, ys__n46686, ys__n46687, ys__n46688, ys__n46689, ys__n46690,
    ys__n46691, ys__n46692, ys__n46693, ys__n46694, ys__n46695, ys__n46696,
    ys__n46697, ys__n46698, ys__n46700, ys__n46702, ys__n46704, ys__n46706,
    ys__n46708, ys__n46710, ys__n46712, ys__n46714, ys__n46716, ys__n46718,
    ys__n46720, ys__n46722, ys__n46724, ys__n46726, ys__n46728, ys__n46730,
    ys__n46732, ys__n46734, ys__n46736, ys__n46738, ys__n46740, ys__n46742,
    ys__n46744, ys__n46745, ys__n46746, ys__n46747, ys__n46748, ys__n46749,
    ys__n46750, ys__n46751, ys__n46752, ys__n46753, ys__n46754, ys__n46755,
    ys__n46756, ys__n46757, ys__n46758, ys__n46759, ys__n46760, ys__n46761,
    ys__n46762, ys__n46763, ys__n46764, ys__n46765, ys__n46766, ys__n46767,
    ys__n46768, ys__n46769, ys__n46770, ys__n46771, ys__n46772, ys__n46773,
    ys__n46774, ys__n46775, ys__n46780, ys__n46782, ys__n46784, ys__n46786,
    ys__n46788, ys__n46790, ys__n46792, ys__n46794, ys__n46796, ys__n46798,
    ys__n46800, ys__n46802, ys__n46804, ys__n46806, ys__n46808, ys__n46810,
    ys__n46812, ys__n46814, ys__n46816, ys__n46818, ys__n46820, ys__n46822,
    ys__n46824, ys__n46826, ys__n46828, ys__n46830, ys__n46832, ys__n46834,
    ys__n46836, ys__n46838, ys__n46840, ys__n46842, ys__n46843, ys__n46844,
    ys__n46845, ys__n46846, ys__n46847, ys__n46848, ys__n46849, ys__n46850,
    ys__n46851, ys__n46852, ys__n46853, ys__n46854, ys__n46855, ys__n46856,
    ys__n46857, ys__n46858, ys__n46859, ys__n46860, ys__n46861, ys__n46862,
    ys__n46863, ys__n46864, ys__n46865, ys__n46866, ys__n46867, ys__n46868,
    ys__n46869, ys__n46870, ys__n46871, ys__n46872, ys__n46873, ys__n46874,
    ys__n46876, ys__n46878, ys__n46880, ys__n46882, ys__n46884, ys__n46886,
    ys__n46888, ys__n46890, ys__n46892, ys__n46894, ys__n46896, ys__n46898,
    ys__n46900, ys__n46902, ys__n46904, ys__n46906, ys__n46908, ys__n46910,
    ys__n46912, ys__n46914, ys__n46916, ys__n46918, ys__n46920, ys__n46921,
    ys__n46922, ys__n46923, ys__n46924, ys__n46925, ys__n46926, ys__n46927,
    ys__n46928, ys__n46929, ys__n46930, ys__n46931, ys__n46932, ys__n46933,
    ys__n46934, ys__n46935, ys__n46936, ys__n46937, ys__n46938, ys__n46939,
    ys__n46940, ys__n46941, ys__n46942, ys__n46943, ys__n46944, ys__n46945,
    ys__n46946, ys__n46947, ys__n46948, ys__n46949, ys__n46950, ys__n46951,
    ys__n46954, ys__n46955, ys__n46956, ys__n46957, ys__n46958, ys__n46959,
    ys__n46960, ys__n46961, ys__n46962, ys__n46963, ys__n46964, ys__n46965,
    ys__n46966, ys__n46967, ys__n46968, ys__n46969, ys__n46970, ys__n46971,
    ys__n46972, ys__n46973, ys__n46974, ys__n46975, ys__n46976, ys__n46977,
    ys__n46978, ys__n46979, ys__n46980, ys__n46981, ys__n46982, ys__n46983,
    ys__n46984, ys__n46985, ys__n46986, ys__n46987, ys__n46988, ys__n46989,
    ys__n46990, ys__n46991, ys__n46992, ys__n46993, ys__n46994, ys__n46995,
    ys__n46996, ys__n46997, ys__n46998, ys__n46999, ys__n47000, ys__n47001,
    ys__n47002, ys__n47003, ys__n47004, ys__n47005, ys__n47006, ys__n47007,
    ys__n47008, ys__n47009, ys__n47010, ys__n47011, ys__n47012, ys__n47013,
    ys__n47014, ys__n47015, ys__n47016, ys__n47017, ys__n47018, ys__n47019,
    ys__n47020, ys__n47021, ys__n47022, ys__n47023, ys__n47024, ys__n47025,
    ys__n47026, ys__n47027, ys__n47028, ys__n47029, ys__n47030, ys__n47031,
    ys__n47032, ys__n47033, ys__n47034, ys__n47035, ys__n47036, ys__n47037,
    ys__n47038, ys__n47039, ys__n47040, ys__n47041, ys__n47074, ys__n47075,
    ys__n47076, ys__n47077, ys__n47078, ys__n47079, ys__n47080, ys__n47081,
    ys__n47082, ys__n47083, ys__n47084, ys__n47085, ys__n47086, ys__n47087,
    ys__n47088, ys__n47089, ys__n47090, ys__n47091, ys__n47092, ys__n47093,
    ys__n47094, ys__n47095, ys__n47096, ys__n47097, ys__n47098, ys__n47099,
    ys__n47100, ys__n47101, ys__n47102, ys__n47103, ys__n47104, ys__n47105,
    ys__n47106, ys__n47107, ys__n47108, ys__n47109, ys__n47110, ys__n47111,
    ys__n47112, ys__n47113, ys__n47114, ys__n47115, ys__n47116, ys__n47117,
    ys__n47118, ys__n47119, ys__n47184, ys__n47185, ys__n47186, ys__n47187,
    ys__n47188, ys__n47189, ys__n47190, ys__n47191, ys__n47192, ys__n47193,
    ys__n47194, ys__n47195, ys__n47196, ys__n47197, ys__n47198, ys__n47199,
    ys__n47200, ys__n47201, ys__n47202, ys__n47203, ys__n47204, ys__n47205,
    ys__n47206, ys__n47207, ys__n47208, ys__n47209, ys__n47210, ys__n47211,
    ys__n47212, ys__n47213, ys__n47214, ys__n47215, ys__n47216, ys__n47217,
    ys__n47218, ys__n47219, ys__n47220, ys__n47221, ys__n47222, ys__n47223,
    ys__n47224, ys__n47225, ys__n47226, ys__n47227, ys__n47228, ys__n47229,
    ys__n47230, ys__n47231, ys__n47232, ys__n47233, ys__n47234, ys__n47235,
    ys__n47236, ys__n47237, ys__n47238, ys__n47239, ys__n47240, ys__n47241,
    ys__n47242, ys__n47243, ys__n47244, ys__n47245, ys__n47246, ys__n47247,
    ys__n47248, ys__n47249, ys__n47250, ys__n47251, ys__n47252, ys__n47253,
    ys__n47254, ys__n47255, ys__n47256, ys__n47257, ys__n47258, ys__n47259,
    ys__n47260, ys__n47261, ys__n47262, ys__n47263, ys__n47264, ys__n47265,
    ys__n47266, ys__n47267, ys__n47268, ys__n47269, ys__n47270, ys__n47271,
    ys__n47272, ys__n47273, ys__n47274, ys__n47275, ys__n47276, ys__n47277,
    ys__n47278, ys__n47279, ys__n47280, ys__n47281, ys__n47282, ys__n47283,
    ys__n47284, ys__n47285, ys__n47286, ys__n47287, ys__n47288, ys__n47289,
    ys__n47290, ys__n47291, ys__n47292, ys__n47293, ys__n47294, ys__n47295,
    ys__n47296, ys__n47297, ys__n47298, ys__n47299, ys__n47300, ys__n47301,
    ys__n47302, ys__n47303, ys__n47305, ys__n47306, ys__n47307, ys__n47308,
    ys__n47309, ys__n47310, ys__n47311, ys__n47312, ys__n47313, ys__n47314,
    ys__n47315, ys__n47316, ys__n47317, ys__n47318, ys__n47319, ys__n47320,
    ys__n47321, ys__n47322, ys__n47323, ys__n47324, ys__n47325, ys__n47326,
    ys__n47327, ys__n47328, ys__n47329, ys__n47330, ys__n47331, ys__n47332,
    ys__n47333, ys__n47334, ys__n47335, ys__n47336, ys__n47337, ys__n47338,
    ys__n47339, ys__n47340, ys__n47341, ys__n47342, ys__n47343, ys__n47344,
    ys__n47345, ys__n47346, ys__n47347, ys__n47348, ys__n47349, ys__n47350,
    ys__n47351, ys__n47352, ys__n47353, ys__n47354, ys__n47355, ys__n47356,
    ys__n47357, ys__n47358, ys__n47359, ys__n47360, ys__n47361, ys__n47362,
    ys__n47363, ys__n47364, ys__n47365, ys__n47366, ys__n47367, ys__n47368,
    ys__n47369, ys__n47370, ys__n47371, ys__n47372, ys__n47373, ys__n47374,
    ys__n47375, ys__n47376, ys__n47377, ys__n47378, ys__n47379, ys__n47380,
    ys__n47381, ys__n47382, ys__n47383, ys__n47384, ys__n47385, ys__n47386,
    ys__n47387, ys__n47388, ys__n47389, ys__n47390, ys__n47391, ys__n47392,
    ys__n47393, ys__n47394, ys__n47395, ys__n47396, ys__n47397, ys__n47398,
    ys__n47399, ys__n47400, ys__n47401, ys__n47402, ys__n47403, ys__n47404,
    ys__n47405, ys__n47406, ys__n47407, ys__n47408, ys__n47409, ys__n47410,
    ys__n47411, ys__n47412, ys__n47413, ys__n47414, ys__n47415, ys__n47416,
    ys__n47417, ys__n47418, ys__n47419, ys__n47420, ys__n47421, ys__n47422,
    ys__n47423, ys__n47424, ys__n47425, ys__n47426, ys__n47427, ys__n47428,
    ys__n47429, ys__n47430, ys__n47431, ys__n47432, ys__n47433, ys__n47434,
    ys__n47435, ys__n47436, ys__n47437, ys__n47438, ys__n47439, ys__n47440,
    ys__n47441, ys__n47442, ys__n47443, ys__n47444, ys__n47445, ys__n47446,
    ys__n47447, ys__n47448, ys__n47449, ys__n47450, ys__n47451, ys__n47452,
    ys__n47453, ys__n47454, ys__n47455, ys__n47456, ys__n47457, ys__n47458,
    ys__n47459, ys__n47460, ys__n47461, ys__n47462, ys__n47463, ys__n47464,
    ys__n47465, ys__n47466, ys__n47467, ys__n47468, ys__n47469, ys__n47470,
    ys__n47471, ys__n47472, ys__n47473, ys__n47474, ys__n47475, ys__n47476,
    ys__n47477, ys__n47478, ys__n47479, ys__n47480, ys__n47481, ys__n47482,
    ys__n47483, ys__n47484, ys__n47485, ys__n47486, ys__n47487, ys__n47488,
    ys__n47489, ys__n47490, ys__n47491, ys__n47492, ys__n47493, ys__n47494,
    ys__n47495, ys__n47496, ys__n47497, ys__n47498, ys__n47499, ys__n47500,
    ys__n47501, ys__n47502, ys__n47503, ys__n47504, ys__n47505, ys__n47506,
    ys__n47507, ys__n47508, ys__n47509, ys__n47510, ys__n47511, ys__n47512,
    ys__n47513, ys__n47514, ys__n47515, ys__n47516, ys__n47517, ys__n47518,
    ys__n47519, ys__n47520, ys__n47521, ys__n47522, ys__n47523, ys__n47524,
    ys__n47525, ys__n47526, ys__n47527, ys__n47528, ys__n47529, ys__n47530,
    ys__n47531, ys__n47532, ys__n47533, ys__n47534, ys__n47535, ys__n47536,
    ys__n47537, ys__n47538, ys__n47539, ys__n47540, ys__n47541, ys__n47542,
    ys__n47543, ys__n47544, ys__n47545, ys__n47546, ys__n47547, ys__n47548,
    ys__n47549, ys__n47550, ys__n47551, ys__n47552, ys__n47553, ys__n47554,
    ys__n47555, ys__n47556, ys__n47557, ys__n47558, ys__n47559, ys__n47560,
    ys__n47561, ys__n47562, ys__n47563, ys__n47564, ys__n47565, ys__n47566,
    ys__n47567, ys__n47568, ys__n47569, ys__n47570, ys__n47571, ys__n47572,
    ys__n47573, ys__n47574, ys__n47575, ys__n47576, ys__n47577, ys__n47578,
    ys__n47579, ys__n47580, ys__n47581, ys__n47582, ys__n47583, ys__n47584,
    ys__n47585, ys__n47586, ys__n47587, ys__n47588, ys__n47589, ys__n47590,
    ys__n47591, ys__n47592, ys__n47593, ys__n47594, ys__n47595, ys__n47596,
    ys__n47597, ys__n47598, ys__n47599, ys__n47600, ys__n47601, ys__n47602,
    ys__n47603, ys__n47604, ys__n47605, ys__n47606, ys__n47607, ys__n47608,
    ys__n47609, ys__n47610, ys__n47611, ys__n47612, ys__n47613, ys__n47614,
    ys__n47615, ys__n47616, ys__n47617, ys__n47618, ys__n47619, ys__n47620,
    ys__n47621, ys__n47622, ys__n47623, ys__n47624, ys__n47625, ys__n47626,
    ys__n47627, ys__n47628, ys__n47629, ys__n47630, ys__n47631, ys__n47632,
    ys__n47633, ys__n47634, ys__n47635, ys__n47636, ys__n47637, ys__n47638,
    ys__n47639, ys__n47640, ys__n47641, ys__n47642, ys__n47643, ys__n47644,
    ys__n47645, ys__n47646, ys__n47647, ys__n47648, ys__n47649, ys__n47650,
    ys__n47651, ys__n47652, ys__n47653, ys__n47654, ys__n47655, ys__n47656,
    ys__n47657, ys__n47658, ys__n47659, ys__n47660, ys__n47661, ys__n47662,
    ys__n47663, ys__n47664, ys__n47665, ys__n47666, ys__n47667, ys__n47668,
    ys__n47669, ys__n47670, ys__n47671, ys__n47672, ys__n47673, ys__n47674,
    ys__n47675, ys__n47676, ys__n47677, ys__n47678, ys__n47679, ys__n47680,
    ys__n47681, ys__n47682, ys__n47683, ys__n47684, ys__n47685, ys__n47686,
    ys__n47687, ys__n47688, ys__n47689, ys__n47690, ys__n47691, ys__n47692,
    ys__n47693, ys__n47694, ys__n47695, ys__n47696, ys__n47697, ys__n47698,
    ys__n47699, ys__n47700, ys__n47701, ys__n47702, ys__n47703, ys__n47704,
    ys__n47705, ys__n47706, ys__n47707, ys__n47708, ys__n47709, ys__n47710,
    ys__n47711, ys__n47712, ys__n47713, ys__n47714, ys__n47715, ys__n47716,
    ys__n47717, ys__n47718, ys__n47719, ys__n47720, ys__n47721, ys__n47722,
    ys__n47723, ys__n47724, ys__n47725, ys__n47726, ys__n47727, ys__n47728,
    ys__n47729, ys__n47730, ys__n47731, ys__n47732, ys__n47733, ys__n47734,
    ys__n47735, ys__n47736, ys__n47737, ys__n47738, ys__n47739, ys__n47740,
    ys__n47741, ys__n47742, ys__n47743, ys__n47744, ys__n47745, ys__n47746,
    ys__n47747, ys__n47748, ys__n47749, ys__n47750, ys__n47751, ys__n47752,
    ys__n47753, ys__n47754, ys__n47755, ys__n47756, ys__n47757, ys__n47758,
    ys__n47759, ys__n47760, ys__n47761, ys__n47762, ys__n47763, ys__n47764,
    ys__n47765, ys__n47766, ys__n47767, ys__n47768, ys__n47769, ys__n47770,
    ys__n47771, ys__n47772, ys__n47773, ys__n47774, ys__n47775, ys__n47776,
    ys__n47777, ys__n47778, ys__n47779, ys__n47780, ys__n47781, ys__n47782,
    ys__n47783, ys__n47784, ys__n47785, ys__n47786, ys__n47787, ys__n47788,
    ys__n47789, ys__n47790, ys__n47791, ys__n47792, ys__n47793, ys__n47794,
    ys__n47795, ys__n47796, ys__n47797, ys__n47798, ys__n47799, ys__n47800,
    ys__n47801, ys__n47802, ys__n47803, ys__n47804, ys__n47805, ys__n47806,
    ys__n47807, ys__n47808, ys__n47809, ys__n47810, ys__n47811, ys__n47812,
    ys__n47813, ys__n47814, ys__n47815, ys__n47816, ys__n47817, ys__n47818,
    ys__n47819, ys__n47820, ys__n47821, ys__n47822, ys__n47823, ys__n47824,
    ys__n47825, ys__n47826, ys__n47827, ys__n47828, ys__n47829, ys__n47830,
    ys__n47831, ys__n47832, ys__n47833, ys__n47834, ys__n47835, ys__n47836,
    ys__n47837, ys__n47838, ys__n47839, ys__n47840, ys__n47841, ys__n47842,
    ys__n47843, ys__n47844, ys__n47845, ys__n47846, ys__n47847, ys__n47848,
    ys__n47849, ys__n47850, ys__n47851, ys__n47852, ys__n47853, ys__n47854,
    ys__n47855, ys__n47856, ys__n47857, ys__n47858, ys__n47859, ys__n47860,
    ys__n47861, ys__n47862, ys__n47863, ys__n47864, ys__n47865, ys__n47866,
    ys__n47867, ys__n47868, ys__n47869, ys__n47870, ys__n47871, ys__n47872,
    ys__n47873, ys__n47874, ys__n47875, ys__n47876, ys__n47877, ys__n47878,
    ys__n47879, ys__n47880, ys__n47881, ys__n47882, ys__n47883, ys__n47884,
    ys__n47885, ys__n47886, ys__n47887, ys__n47888, ys__n47889, ys__n47890,
    ys__n47891, ys__n47892, ys__n47893, ys__n47894, ys__n47895, ys__n47896,
    ys__n47897, ys__n47898, ys__n47899, ys__n47900, ys__n47901, ys__n47902,
    ys__n47903, ys__n47904, ys__n47905, ys__n47906, ys__n47907, ys__n47908,
    ys__n47909, ys__n47910, ys__n47911, ys__n47912, ys__n47913, ys__n47914,
    ys__n47915, ys__n47916, ys__n47917, ys__n47918, ys__n47919, ys__n47920,
    ys__n47921, ys__n47922, ys__n47923, ys__n47924, ys__n47925, ys__n47926,
    ys__n47927, ys__n47928, ys__n47929, ys__n47930, ys__n47931, ys__n47932,
    ys__n47933, ys__n47934, ys__n47935, ys__n47936, ys__n47937, ys__n47938,
    ys__n47939, ys__n47940, ys__n47941, ys__n47942, ys__n47943, ys__n47944,
    ys__n47945, ys__n47946, ys__n47947, ys__n47948, ys__n47949, ys__n47950,
    ys__n47951, ys__n47952, ys__n47953, ys__n47954, ys__n47955, ys__n47956,
    ys__n47957, ys__n47958, ys__n47959, ys__n47960, ys__n47961, ys__n47962,
    ys__n47963, ys__n47964, ys__n47965, ys__n47966, ys__n47967, ys__n47968,
    ys__n47969, ys__n47970, ys__n47971, ys__n47972, ys__n47973, ys__n47974,
    ys__n47975, ys__n47976, ys__n47977, ys__n47978, ys__n47979, ys__n47980,
    ys__n47981, ys__n47982, ys__n47983, ys__n47984, ys__n47985, ys__n47986,
    ys__n47987, ys__n47988, ys__n47989, ys__n47990, ys__n47991, ys__n47992,
    ys__n47993, ys__n47994, ys__n47995, ys__n47996, ys__n47997, ys__n47998,
    ys__n47999, ys__n48000, ys__n48001, ys__n48002, ys__n48003, ys__n48004,
    ys__n48005, ys__n48006, ys__n48007, ys__n48008, ys__n48009, ys__n48010,
    ys__n48011, ys__n48012, ys__n48013, ys__n48014, ys__n48015, ys__n48016,
    ys__n48017, ys__n48018, ys__n48019, ys__n48020, ys__n48021, ys__n48022,
    ys__n48023, ys__n48024, ys__n48025, ys__n48026, ys__n48027, ys__n48028,
    ys__n48029, ys__n48030, ys__n48031, ys__n48032, ys__n48033, ys__n48034,
    ys__n48035, ys__n48036, ys__n48037, ys__n48038, ys__n48039, ys__n48040,
    ys__n48041, ys__n48042, ys__n48043, ys__n48044, ys__n48045, ys__n48046,
    ys__n48047, ys__n48048, ys__n48049, ys__n48050, ys__n48051, ys__n48052,
    ys__n48053, ys__n48054, ys__n48055, ys__n48056, ys__n48057, ys__n48058,
    ys__n48059, ys__n48060, ys__n48061, ys__n48062, ys__n48063, ys__n48064,
    ys__n48065, ys__n48066, ys__n48067, ys__n48068, ys__n48069, ys__n48070,
    ys__n48071, ys__n48072, ys__n48073, ys__n48074, ys__n48075, ys__n48076,
    ys__n48077, ys__n48078, ys__n48079, ys__n48080, ys__n48081, ys__n48082,
    ys__n48083, ys__n48084, ys__n48085, ys__n48086, ys__n48087, ys__n48088,
    ys__n48089, ys__n48090, ys__n48091, ys__n48092, ys__n48093, ys__n48094,
    ys__n48095, ys__n48096, ys__n48097, ys__n48098, ys__n48099, ys__n48100,
    ys__n48101, ys__n48102, ys__n48103, ys__n48104, ys__n48105, ys__n48106,
    ys__n48107, ys__n48108, ys__n48109, ys__n48110, ys__n48111, ys__n48112,
    ys__n48113, ys__n48114, ys__n48115, ys__n48116, ys__n48117, ys__n48118,
    ys__n48119, ys__n48120, ys__n48121, ys__n48122, ys__n48123, ys__n48124,
    ys__n48125, ys__n48126, ys__n48127, ys__n48128, ys__n48129, ys__n48130,
    ys__n48131, ys__n48132, ys__n48133, ys__n48134, ys__n48135, ys__n48136,
    ys__n48137, ys__n48138, ys__n48139, ys__n48140, ys__n48141, ys__n48142,
    ys__n48143, ys__n48144, ys__n48145, ys__n48146, ys__n48147, ys__n48148,
    ys__n48149, ys__n48150, ys__n48151, ys__n48152, ys__n48153, ys__n48154,
    ys__n48155, ys__n48156, ys__n48157, ys__n48158, ys__n48159, ys__n48160,
    ys__n48161, ys__n48162, ys__n48163, ys__n48164, ys__n48165, ys__n48166,
    ys__n48167, ys__n48168, ys__n48169, ys__n48170, ys__n48171, ys__n48172,
    ys__n48173, ys__n48174, ys__n48175, ys__n48176, ys__n48177, ys__n48178,
    ys__n48179, ys__n48180, ys__n48181, ys__n48182, ys__n48183, ys__n48184,
    ys__n48185, ys__n48186, ys__n48187, ys__n48188, ys__n48189, ys__n48190,
    ys__n48191, ys__n48192, ys__n48193, ys__n48194, ys__n48195, ys__n48196,
    ys__n48197, ys__n48198, ys__n48199, ys__n48200, ys__n48201, ys__n48202,
    ys__n48203, ys__n48204, ys__n48205, ys__n48206, ys__n48207, ys__n48208,
    ys__n48209, ys__n48210, ys__n48211, ys__n48212, ys__n48213, ys__n48214,
    ys__n48215, ys__n48216, ys__n48217, ys__n48218, ys__n48219, ys__n48220,
    ys__n48221, ys__n48222, ys__n48223, ys__n48224, ys__n48225, ys__n48226,
    ys__n48227, ys__n48228, ys__n48229, ys__n48230, ys__n48231, ys__n48232,
    ys__n48233, ys__n48234, ys__n48235, ys__n48236, ys__n48237, ys__n48238,
    ys__n48239, ys__n48240, ys__n48241, ys__n48242, ys__n48243, ys__n48244,
    ys__n48245, ys__n48246, ys__n48247, ys__n48248, ys__n48249, ys__n48250,
    ys__n48251, ys__n48252, ys__n48253, ys__n48254, ys__n48255, ys__n48256,
    ys__n48257, ys__n48258, ys__n48259, ys__n48260, ys__n48261, ys__n48262,
    ys__n48263, ys__n48264, ys__n48265, ys__n48266, ys__n48267, ys__n48268,
    ys__n48269, ys__n48270, ys__n48271, ys__n48272, ys__n48273, ys__n48274,
    ys__n48275, ys__n48324, ys__n48325, ys__n48327, ys__n48330, ys__n48331,
    ys__n48332, ys__n48333, ys__n48334, ys__n48335,
    ys__n2, ys__n246, ys__n250, ys__n252, ys__n254, ys__n264, ys__n270,
    ys__n278, ys__n280, ys__n313, ys__n319, ys__n404, ys__n415, ys__n417,
    ys__n455, ys__n457, ys__n478, ys__n480, ys__n482, ys__n502, ys__n565,
    ys__n574, ys__n576, ys__n628, ys__n630, ys__n714, ys__n716, ys__n730,
    ys__n732, ys__n738, ys__n740, ys__n754, ys__n756, ys__n786, ys__n788,
    ys__n790, ys__n792, ys__n794, ys__n796, ys__n798, ys__n800, ys__n802,
    ys__n804, ys__n806, ys__n808, ys__n810, ys__n812, ys__n814, ys__n862,
    ys__n863, ys__n865, ys__n866, ys__n868, ys__n870, ys__n871, ys__n872,
    ys__n873, ys__n876, ys__n878, ys__n879, ys__n881, ys__n888, ys__n890,
    ys__n900, ys__n902, ys__n904, ys__n911, ys__n920, ys__n923, ys__n927,
    ys__n929, ys__n930, ys__n932, ys__n934, ys__n936, ys__n942, ys__n944,
    ys__n948, ys__n949, ys__n970, ys__n972, ys__n974, ys__n976, ys__n978,
    ys__n980, ys__n982, ys__n989, ys__n991, ys__n993, ys__n995, ys__n999,
    ys__n1001, ys__n1004, ys__n1007, ys__n1009, ys__n1013, ys__n1020,
    ys__n1028, ys__n1030, ys__n1031, ys__n1032, ys__n1037, ys__n1040,
    ys__n1043, ys__n1046, ys__n1047, ys__n1049, ys__n1060, ys__n1071,
    ys__n1073, ys__n1074, ys__n1075, ys__n1077, ys__n1079, ys__n1080,
    ys__n1083, ys__n1085, ys__n1087, ys__n1088, ys__n1089, ys__n1090,
    ys__n1091, ys__n1095, ys__n1103, ys__n1115, ys__n1125, ys__n1128,
    ys__n1135, ys__n1138, ys__n1141, ys__n1142, ys__n1143, ys__n1146,
    ys__n1148, ys__n1161, ys__n1163, ys__n1164, ys__n1165, ys__n1167,
    ys__n1170, ys__n1171, ys__n1183, ys__n1189, ys__n1195, ys__n1201,
    ys__n1207, ys__n1213, ys__n1219, ys__n1222, ys__n1228, ys__n1234,
    ys__n1240, ys__n1246, ys__n1252, ys__n1258, ys__n1261, ys__n1266,
    ys__n1272, ys__n1278, ys__n1284, ys__n1290, ys__n1296, ys__n1303,
    ys__n1377, ys__n1386, ys__n1445, ys__n1448, ys__n1470, ys__n1591,
    ys__n1598, ys__n1601, ys__n1616, ys__n1790, ys__n1802, ys__n1817,
    ys__n1835, ys__n1837, ys__n2152, ys__n2365, ys__n2400, ys__n2423,
    ys__n2491, ys__n2535, ys__n2536, ys__n2582, ys__n2635, ys__n2651,
    ys__n2653, ys__n2655, ys__n2674, ys__n2684, ys__n2733, ys__n2776,
    ys__n2778, ys__n2780, ys__n2782, ys__n2804, ys__n2806, ys__n2845,
    ys__n2855, ys__n3021, ys__n3024, ys__n3035, ys__n3039, ys__n3040,
    ys__n3051, ys__n3061, ys__n3068, ys__n3083, ys__n3085, ys__n3097,
    ys__n3106, ys__n3114, ys__n3115, ys__n3118, ys__n3121, ys__n3195,
    ys__n3249, ys__n3250, ys__n3252, ys__n4175, ys__n4189, ys__n4192,
    ys__n4320, ys__n4414, ys__n4521, ys__n4566, ys__n4588, ys__n4603,
    ys__n4615, ys__n4696, ys__n4764, ys__n4791, ys__n4793, ys__n4798,
    ys__n4817, ys__n4818, ys__n4820, ys__n4821, ys__n4824, ys__n4825,
    ys__n4839, ys__n4840, ys__n12455, ys__n12458, ys__n12461, ys__n12464,
    ys__n12467, ys__n12470, ys__n12473, ys__n12476, ys__n12479, ys__n12482,
    ys__n12485, ys__n12488, ys__n12491, ys__n12494, ys__n12497, ys__n12500,
    ys__n12503, ys__n12506, ys__n12509, ys__n12512, ys__n12515, ys__n12518,
    ys__n12521, ys__n12524, ys__n12527, ys__n12530, ys__n12533, ys__n12536,
    ys__n12539, ys__n12542, ys__n12545, ys__n12548, ys__n16188, ys__n16191,
    ys__n16412, ys__n16415, ys__n16424, ys__n16427, ys__n16706, ys__n16709,
    ys__n16718, ys__n16721, ys__n17692, ys__n17697, ys__n17780, ys__n18007,
    ys__n18009, ys__n18015, ys__n18019, ys__n18028, ys__n18078, ys__n18080,
    ys__n18082, ys__n18087, ys__n18088, ys__n18089, ys__n18120, ys__n18125,
    ys__n18128, ys__n18131, ys__n18133, ys__n18134, ys__n18136, ys__n18137,
    ys__n18154, ys__n18165, ys__n18166, ys__n18169, ys__n18170, ys__n18174,
    ys__n18176, ys__n18178, ys__n18210, ys__n18214, ys__n18216, ys__n18217,
    ys__n18218, ys__n18223, ys__n18227, ys__n18236, ys__n18238, ys__n18239,
    ys__n18241, ys__n18251, ys__n18268, ys__n18272, ys__n18273, ys__n18278,
    ys__n18281, ys__n18284, ys__n18287, ys__n18303, ys__n18321, ys__n18329,
    ys__n18331, ys__n18333, ys__n18335, ys__n18337, ys__n18339, ys__n18341,
    ys__n18343, ys__n18345, ys__n18347, ys__n18349, ys__n18351, ys__n18353,
    ys__n18355, ys__n18357, ys__n18360, ys__n18380, ys__n18383, ys__n18386,
    ys__n18391, ys__n18392, ys__n18394, ys__n18395, ys__n18396, ys__n18397,
    ys__n18398, ys__n18399, ys__n18400, ys__n18401, ys__n18402, ys__n18403,
    ys__n18404, ys__n18405, ys__n18406, ys__n18407, ys__n18408, ys__n18409,
    ys__n18410, ys__n18411, ys__n18412, ys__n18413, ys__n18414, ys__n18415,
    ys__n18416, ys__n18417, ys__n18418, ys__n18419, ys__n18420, ys__n18421,
    ys__n18422, ys__n18423, ys__n18424, ys__n18425, ys__n18426, ys__n18427,
    ys__n18428, ys__n18429, ys__n18430, ys__n18431, ys__n18432, ys__n18433,
    ys__n18434, ys__n18435, ys__n18436, ys__n18437, ys__n18438, ys__n18439,
    ys__n18440, ys__n18441, ys__n18442, ys__n18443, ys__n18444, ys__n18445,
    ys__n18449, ys__n18450, ys__n18452, ys__n18453, ys__n18455, ys__n18456,
    ys__n18458, ys__n18459, ys__n18461, ys__n18462, ys__n18464, ys__n18465,
    ys__n18467, ys__n18468, ys__n18470, ys__n18471, ys__n18473, ys__n18474,
    ys__n18476, ys__n18477, ys__n18479, ys__n18480, ys__n18482, ys__n18483,
    ys__n18485, ys__n18486, ys__n18488, ys__n18489, ys__n18491, ys__n18492,
    ys__n18494, ys__n18495, ys__n18497, ys__n18498, ys__n18500, ys__n18501,
    ys__n18503, ys__n18504, ys__n18506, ys__n18507, ys__n18509, ys__n18510,
    ys__n18512, ys__n18513, ys__n18515, ys__n18516, ys__n18518, ys__n18519,
    ys__n18521, ys__n18522, ys__n18524, ys__n18525, ys__n18527, ys__n18528,
    ys__n18530, ys__n18531, ys__n18533, ys__n18534, ys__n18536, ys__n18537,
    ys__n18539, ys__n18540, ys__n18542, ys__n18543, ys__n18545, ys__n18547,
    ys__n18548, ys__n18549, ys__n18550, ys__n18551, ys__n18553, ys__n18554,
    ys__n18555, ys__n18557, ys__n18559, ys__n18561, ys__n18564, ys__n18567,
    ys__n18570, ys__n18573, ys__n18576, ys__n18579, ys__n18582, ys__n18585,
    ys__n18588, ys__n18591, ys__n18594, ys__n18597, ys__n18600, ys__n18603,
    ys__n18606, ys__n18609, ys__n18612, ys__n18615, ys__n18618, ys__n18621,
    ys__n18624, ys__n18627, ys__n18629, ys__n18631, ys__n18633, ys__n18635,
    ys__n18637, ys__n18640, ys__n18643, ys__n18646, ys__n18649, ys__n18652,
    ys__n18654, ys__n18655, ys__n18657, ys__n18658, ys__n18660, ys__n18661,
    ys__n18663, ys__n18664, ys__n18666, ys__n18667, ys__n18669, ys__n18670,
    ys__n18672, ys__n18673, ys__n18675, ys__n18676, ys__n18678, ys__n18679,
    ys__n18681, ys__n18682, ys__n18684, ys__n18685, ys__n18687, ys__n18688,
    ys__n18690, ys__n18691, ys__n18693, ys__n18694, ys__n18696, ys__n18697,
    ys__n18699, ys__n18700, ys__n18702, ys__n18703, ys__n18705, ys__n18706,
    ys__n18708, ys__n18709, ys__n18711, ys__n18712, ys__n18714, ys__n18715,
    ys__n18717, ys__n18718, ys__n18720, ys__n18721, ys__n18723, ys__n18724,
    ys__n18726, ys__n18727, ys__n18729, ys__n18730, ys__n18732, ys__n18733,
    ys__n18735, ys__n18736, ys__n18738, ys__n18739, ys__n18741, ys__n18742,
    ys__n18744, ys__n18745, ys__n18747, ys__n18748, ys__n18750, ys__n18751,
    ys__n18753, ys__n18754, ys__n18757, ys__n18759, ys__n18760, ys__n18763,
    ys__n18764, ys__n18766, ys__n18768, ys__n18770, ys__n18772, ys__n18774,
    ys__n18776, ys__n18778, ys__n18780, ys__n18782, ys__n18784, ys__n18786,
    ys__n18788, ys__n18790, ys__n18792, ys__n18794, ys__n18796, ys__n18798,
    ys__n18800, ys__n18802, ys__n18804, ys__n18806, ys__n18808, ys__n18810,
    ys__n18812, ys__n18814, ys__n18816, ys__n18818, ys__n18820, ys__n18822,
    ys__n18824, ys__n18826, ys__n19149, ys__n19151, ys__n19159, ys__n19173,
    ys__n19177, ys__n19178, ys__n19183, ys__n19227, ys__n19229, ys__n19231,
    ys__n19233, ys__n19235, ys__n19239, ys__n19254, ys__n19256, ys__n19257,
    ys__n19264, ys__n19266, ys__n19878, ys__n19881, ys__n19884, ys__n19887,
    ys__n19890, ys__n19893, ys__n19896, ys__n19899, ys__n19902, ys__n19905,
    ys__n19908, ys__n19911, ys__n19914, ys__n19917, ys__n19920, ys__n19923,
    ys__n19926, ys__n19929, ys__n19932, ys__n19935, ys__n19938, ys__n19941,
    ys__n19944, ys__n19947, ys__n19950, ys__n19953, ys__n19956, ys__n19959,
    ys__n19962, ys__n19965, ys__n19968, ys__n19971, ys__n20006, ys__n20007,
    ys__n20008, ys__n20009, ys__n20010, ys__n20011, ys__n20012, ys__n20013,
    ys__n20014, ys__n20015, ys__n20016, ys__n20017, ys__n20018, ys__n20019,
    ys__n20020, ys__n20021, ys__n20022, ys__n20023, ys__n20024, ys__n20025,
    ys__n20026, ys__n20027, ys__n20028, ys__n20029, ys__n20030, ys__n20031,
    ys__n20032, ys__n20033, ys__n20034, ys__n20038, ys__n20040, ys__n20043,
    ys__n20045, ys__n20053, ys__n20059, ys__n20062, ys__n20065, ys__n20068,
    ys__n20071, ys__n20074, ys__n20077, ys__n20080, ys__n20082, ys__n20084,
    ys__n20086, ys__n20088, ys__n20090, ys__n20092, ys__n20094, ys__n20096,
    ys__n20098, ys__n20100, ys__n20102, ys__n20104, ys__n20106, ys__n20108,
    ys__n20110, ys__n20112, ys__n20114, ys__n20116, ys__n20118, ys__n20120,
    ys__n20122, ys__n20124, ys__n20126, ys__n20128, ys__n22466, ys__n22919,
    ys__n22922, ys__n22925, ys__n22928, ys__n22931, ys__n22934, ys__n22937,
    ys__n22940, ys__n22943, ys__n22946, ys__n22949, ys__n22952, ys__n22955,
    ys__n22958, ys__n22961, ys__n22964, ys__n22967, ys__n22970, ys__n22973,
    ys__n22976, ys__n22979, ys__n22982, ys__n22985, ys__n22988, ys__n22991,
    ys__n22994, ys__n22997, ys__n23000, ys__n23003, ys__n23006, ys__n23009,
    ys__n23012, ys__n23263, ys__n23264, ys__n23340, ys__n23483, ys__n23485,
    ys__n23487, ys__n23489, ys__n23491, ys__n23493, ys__n23495, ys__n23497,
    ys__n23499, ys__n23501, ys__n23503, ys__n23505, ys__n23507, ys__n23509,
    ys__n23511, ys__n23513, ys__n23515, ys__n23517, ys__n23519, ys__n23521,
    ys__n23523, ys__n23525, ys__n23527, ys__n23529, ys__n23531, ys__n23533,
    ys__n23535, ys__n23537, ys__n23539, ys__n23541, ys__n23543, ys__n23635,
    ys__n23636, ys__n23764, ys__n23795, ys__n23798, ys__n23801, ys__n23804,
    ys__n23807, ys__n23853, ys__n23865, ys__n23868, ys__n23871, ys__n23874,
    ys__n23877, ys__n23921, ys__n23933, ys__n23936, ys__n23939, ys__n23942,
    ys__n23945, ys__n24099, ys__n24101, ys__n24102, ys__n24104, ys__n24105,
    ys__n24116, ys__n24118, ys__n24120, ys__n24126, ys__n24130, ys__n24134,
    ys__n24140, ys__n24145, ys__n24149, ys__n24154, ys__n24160, ys__n24162,
    ys__n24163, ys__n24165, ys__n24166, ys__n24176, ys__n24179, ys__n24180,
    ys__n24182, ys__n24183, ys__n24185, ys__n24186, ys__n24188, ys__n24189,
    ys__n24191, ys__n24192, ys__n24194, ys__n24195, ys__n24222, ys__n24227,
    ys__n24231, ys__n24236, ys__n24240, ys__n24245, ys__n24250, ys__n24255,
    ys__n24256, ys__n24258, ys__n24259, ys__n24260, ys__n24262, ys__n24265,
    ys__n24268, ys__n24271, ys__n24272, ys__n24274, ys__n24275, ys__n24277,
    ys__n24278, ys__n24286, ys__n24289, ys__n24291, ys__n24293, ys__n24295,
    ys__n24297, ys__n24299, ys__n24301, ys__n24305, ys__n24307, ys__n24309,
    ys__n24311, ys__n24313, ys__n24315, ys__n24317, ys__n24319, ys__n24320,
    ys__n24323, ys__n24325, ys__n24327, ys__n24329, ys__n24331, ys__n24333,
    ys__n24335, ys__n24339, ys__n24341, ys__n24343, ys__n24345, ys__n24347,
    ys__n24349, ys__n24351, ys__n24353, ys__n24354, ys__n24357, ys__n24359,
    ys__n24361, ys__n24363, ys__n24365, ys__n24367, ys__n24369, ys__n24373,
    ys__n24375, ys__n24377, ys__n24379, ys__n24381, ys__n24383, ys__n24385,
    ys__n24387, ys__n24388, ys__n24392, ys__n24394, ys__n24396, ys__n24398,
    ys__n24400, ys__n24402, ys__n24404, ys__n24408, ys__n24410, ys__n24412,
    ys__n24414, ys__n24416, ys__n24418, ys__n24420, ys__n24422, ys__n24425,
    ys__n24430, ys__n24436, ys__n24440, ys__n24445, ys__n24447, ys__n24466,
    ys__n24470, ys__n24488, ys__n24499, ys__n24502, ys__n24522, ys__n24532,
    ys__n24541, ys__n24552, ys__n24570, ys__n24573, ys__n24577, ys__n24579,
    ys__n24581, ys__n24585, ys__n24604, ys__n24713, ys__n24714, ys__n24742,
    ys__n24745, ys__n24748, ys__n24751, ys__n24754, ys__n24757, ys__n24760,
    ys__n24763, ys__n24766, ys__n24769, ys__n24772, ys__n24775, ys__n24778,
    ys__n24781, ys__n24784, ys__n24787, ys__n24790, ys__n24793, ys__n24796,
    ys__n24799, ys__n24802, ys__n24805, ys__n24808, ys__n24811, ys__n24814,
    ys__n24817, ys__n24820, ys__n24823, ys__n24826, ys__n24829, ys__n24832,
    ys__n24835, ys__n24837, ys__n24839, ys__n24907, ys__n24910, ys__n24913,
    ys__n24916, ys__n24919, ys__n24922, ys__n24925, ys__n24928, ys__n24931,
    ys__n24934, ys__n24937, ys__n24940, ys__n24943, ys__n24946, ys__n24949,
    ys__n24952, ys__n24955, ys__n25294, ys__n25302, ys__n25304, ys__n25306,
    ys__n25308, ys__n25310, ys__n25385, ys__n25386, ys__n25387, ys__n25388,
    ys__n25390, ys__n25406, ys__n25421, ys__n25430, ys__n25431, ys__n25432,
    ys__n25433, ys__n25434, ys__n25435, ys__n25436, ys__n25438, ys__n25441,
    ys__n25449, ys__n25456, ys__n25461, ys__n25463, ys__n25465, ys__n25467,
    ys__n25469, ys__n25472, ys__n25486, ys__n25496, ys__n25504, ys__n25519,
    ys__n25522, ys__n25534, ys__n25550, ys__n25661, ys__n25663, ys__n25665,
    ys__n25667, ys__n25669, ys__n25671, ys__n25673, ys__n25675, ys__n25677,
    ys__n25679, ys__n25681, ys__n25683, ys__n25685, ys__n25687, ys__n25689,
    ys__n25691, ys__n25693, ys__n25695, ys__n25697, ys__n25699, ys__n25701,
    ys__n25703, ys__n25705, ys__n25707, ys__n25709, ys__n25711, ys__n25713,
    ys__n25715, ys__n25717, ys__n25719, ys__n25721, ys__n25723, ys__n25725,
    ys__n25830, ys__n25833, ys__n25836, ys__n25839, ys__n25842, ys__n25844,
    ys__n25846, ys__n25852, ys__n25957, ys__n25960, ys__n25963, ys__n25966,
    ys__n26118, ys__n26119, ys__n26120, ys__n26121, ys__n26122, ys__n26123,
    ys__n26124, ys__n26125, ys__n26126, ys__n26127, ys__n26128, ys__n26129,
    ys__n26130, ys__n26131, ys__n26132, ys__n26133, ys__n26134, ys__n26135,
    ys__n26136, ys__n26137, ys__n26138, ys__n26139, ys__n26141, ys__n26144,
    ys__n26146, ys__n26148, ys__n26150, ys__n26152, ys__n26154, ys__n26156,
    ys__n26158, ys__n26160, ys__n26220, ys__n26222, ys__n26224, ys__n26226,
    ys__n26228, ys__n26230, ys__n26232, ys__n26234, ys__n26236, ys__n26238,
    ys__n26240, ys__n26242, ys__n26244, ys__n26246, ys__n26248, ys__n26250,
    ys__n26252, ys__n26254, ys__n26256, ys__n26258, ys__n26260, ys__n26262,
    ys__n26264, ys__n26266, ys__n26268, ys__n26270, ys__n26272, ys__n26274,
    ys__n26276, ys__n26278, ys__n26282, ys__n26284, ys__n26286, ys__n26288,
    ys__n26291, ys__n26293, ys__n26294, ys__n26555, ys__n26566, ys__n26573,
    ys__n26607, ys__n26609, ys__n26611, ys__n26613, ys__n26615, ys__n26617,
    ys__n26619, ys__n26621, ys__n26623, ys__n26625, ys__n26627, ys__n26629,
    ys__n26631, ys__n26633, ys__n26635, ys__n26637, ys__n26639, ys__n26641,
    ys__n26643, ys__n26645, ys__n26647, ys__n26649, ys__n26651, ys__n26653,
    ys__n26655, ys__n26657, ys__n26659, ys__n26661, ys__n26663, ys__n26665,
    ys__n26667, ys__n26669, ys__n26671, ys__n26673, ys__n26675, ys__n26677,
    ys__n26679, ys__n26681, ys__n26683, ys__n26685, ys__n26687, ys__n26689,
    ys__n26691, ys__n26693, ys__n26695, ys__n26697, ys__n26699, ys__n26701,
    ys__n26703, ys__n26705, ys__n26707, ys__n26709, ys__n26711, ys__n26713,
    ys__n26715, ys__n26717, ys__n26719, ys__n26721, ys__n26723, ys__n26725,
    ys__n26727, ys__n26729, ys__n26731, ys__n26733, ys__n26734, ys__n26735,
    ys__n26736, ys__n26737, ys__n26738, ys__n26739, ys__n26740, ys__n26741,
    ys__n26742, ys__n26743, ys__n26744, ys__n26745, ys__n26746, ys__n26747,
    ys__n26748, ys__n26749, ys__n26750, ys__n26751, ys__n26752, ys__n26753,
    ys__n26754, ys__n26755, ys__n26756, ys__n26757, ys__n26758, ys__n26759,
    ys__n26760, ys__n26761, ys__n26762, ys__n26763, ys__n26764, ys__n26765,
    ys__n26802, ys__n26803, ys__n26804, ys__n26805, ys__n26806, ys__n26807,
    ys__n26808, ys__n26809, ys__n26810, ys__n26811, ys__n26812, ys__n26813,
    ys__n26814, ys__n26815, ys__n26816, ys__n26817, ys__n26818, ys__n26819,
    ys__n26820, ys__n26821, ys__n26822, ys__n26823, ys__n26824, ys__n26825,
    ys__n26826, ys__n26827, ys__n26828, ys__n26829, ys__n26830, ys__n26831,
    ys__n26832, ys__n26833, ys__n26834, ys__n26835, ys__n26836, ys__n26837,
    ys__n26838, ys__n26839, ys__n26840, ys__n26841, ys__n26842, ys__n26843,
    ys__n26844, ys__n26845, ys__n26846, ys__n26847, ys__n26848, ys__n26849,
    ys__n26850, ys__n26851, ys__n26852, ys__n26853, ys__n26854, ys__n26855,
    ys__n26856, ys__n26857, ys__n26858, ys__n26859, ys__n26860, ys__n26861,
    ys__n26862, ys__n26863, ys__n26864, ys__n26865, ys__n26866, ys__n26867,
    ys__n26868, ys__n26869, ys__n26870, ys__n26871, ys__n26872, ys__n26873,
    ys__n26874, ys__n26875, ys__n26876, ys__n26877, ys__n26878, ys__n26879,
    ys__n26880, ys__n26881, ys__n26882, ys__n26883, ys__n26884, ys__n26885,
    ys__n26886, ys__n26887, ys__n26888, ys__n26889, ys__n26890, ys__n26891,
    ys__n26892, ys__n26893, ys__n26894, ys__n26895, ys__n26896, ys__n26897,
    ys__n26898, ys__n26899, ys__n26900, ys__n26901, ys__n26902, ys__n26903,
    ys__n26904, ys__n26905, ys__n26906, ys__n26907, ys__n26908, ys__n26909,
    ys__n26910, ys__n26911, ys__n26912, ys__n26913, ys__n26914, ys__n26915,
    ys__n26916, ys__n26917, ys__n26918, ys__n26919, ys__n26920, ys__n26921,
    ys__n26922, ys__n26923, ys__n26924, ys__n26925, ys__n26926, ys__n26927,
    ys__n26928, ys__n26929, ys__n26930, ys__n26931, ys__n26932, ys__n26933,
    ys__n26934, ys__n26935, ys__n26936, ys__n26937, ys__n26938, ys__n26939,
    ys__n26940, ys__n26941, ys__n26942, ys__n26943, ys__n26944, ys__n26945,
    ys__n26946, ys__n26947, ys__n26948, ys__n26949, ys__n26950, ys__n26951,
    ys__n26952, ys__n26953, ys__n26954, ys__n26955, ys__n26956, ys__n26957,
    ys__n26958, ys__n26959, ys__n26960, ys__n26961, ys__n26962, ys__n26963,
    ys__n26964, ys__n26965, ys__n26966, ys__n26967, ys__n26968, ys__n26969,
    ys__n26970, ys__n26971, ys__n26972, ys__n26973, ys__n26974, ys__n26975,
    ys__n26976, ys__n26977, ys__n26978, ys__n26979, ys__n26980, ys__n26981,
    ys__n26982, ys__n26983, ys__n26984, ys__n26985, ys__n26986, ys__n26987,
    ys__n26988, ys__n26989, ys__n26990, ys__n26991, ys__n26992, ys__n26993,
    ys__n26994, ys__n26995, ys__n26996, ys__n26997, ys__n26998, ys__n26999,
    ys__n27000, ys__n27001, ys__n27002, ys__n27003, ys__n27004, ys__n27005,
    ys__n27006, ys__n27007, ys__n27008, ys__n27009, ys__n27010, ys__n27011,
    ys__n27012, ys__n27013, ys__n27014, ys__n27015, ys__n27016, ys__n27017,
    ys__n27018, ys__n27019, ys__n27020, ys__n27021, ys__n27022, ys__n27023,
    ys__n27024, ys__n27025, ys__n27026, ys__n27027, ys__n27028, ys__n27029,
    ys__n27030, ys__n27031, ys__n27032, ys__n27033, ys__n27034, ys__n27035,
    ys__n27036, ys__n27037, ys__n27038, ys__n27039, ys__n27040, ys__n27041,
    ys__n27042, ys__n27043, ys__n27044, ys__n27045, ys__n27046, ys__n27047,
    ys__n27048, ys__n27049, ys__n27050, ys__n27051, ys__n27052, ys__n27053,
    ys__n27054, ys__n27055, ys__n27056, ys__n27057, ys__n27058, ys__n27059,
    ys__n27060, ys__n27061, ys__n27062, ys__n27063, ys__n27064, ys__n27065,
    ys__n27066, ys__n27067, ys__n27068, ys__n27069, ys__n27070, ys__n27071,
    ys__n27072, ys__n27073, ys__n27074, ys__n27075, ys__n27076, ys__n27077,
    ys__n27078, ys__n27079, ys__n27080, ys__n27081, ys__n27082, ys__n27083,
    ys__n27084, ys__n27085, ys__n27086, ys__n27087, ys__n27088, ys__n27089,
    ys__n27090, ys__n27091, ys__n27092, ys__n27093, ys__n27094, ys__n27095,
    ys__n27096, ys__n27097, ys__n27098, ys__n27099, ys__n27100, ys__n27101,
    ys__n27102, ys__n27103, ys__n27104, ys__n27105, ys__n27106, ys__n27107,
    ys__n27108, ys__n27109, ys__n27110, ys__n27111, ys__n27112, ys__n27113,
    ys__n27114, ys__n27115, ys__n27116, ys__n27117, ys__n27118, ys__n27119,
    ys__n27120, ys__n27121, ys__n27122, ys__n27123, ys__n27124, ys__n27125,
    ys__n27126, ys__n27127, ys__n27128, ys__n27129, ys__n27130, ys__n27131,
    ys__n27132, ys__n27133, ys__n27134, ys__n27135, ys__n27136, ys__n27137,
    ys__n27138, ys__n27139, ys__n27140, ys__n27141, ys__n27142, ys__n27143,
    ys__n27144, ys__n27145, ys__n27146, ys__n27147, ys__n27148, ys__n27149,
    ys__n27150, ys__n27151, ys__n27152, ys__n27153, ys__n27154, ys__n27155,
    ys__n27156, ys__n27157, ys__n27158, ys__n27159, ys__n27160, ys__n27161,
    ys__n27162, ys__n27163, ys__n27164, ys__n27165, ys__n27166, ys__n27167,
    ys__n27168, ys__n27169, ys__n27170, ys__n27171, ys__n27172, ys__n27173,
    ys__n27174, ys__n27175, ys__n27176, ys__n27177, ys__n27178, ys__n27179,
    ys__n27180, ys__n27181, ys__n27182, ys__n27183, ys__n27184, ys__n27185,
    ys__n27186, ys__n27187, ys__n27188, ys__n27189, ys__n27190, ys__n27191,
    ys__n27192, ys__n27193, ys__n27194, ys__n27195, ys__n27196, ys__n27197,
    ys__n27198, ys__n27199, ys__n27200, ys__n27201, ys__n27202, ys__n27203,
    ys__n27204, ys__n27205, ys__n27206, ys__n27207, ys__n27208, ys__n27209,
    ys__n27210, ys__n27211, ys__n27212, ys__n27213, ys__n27214, ys__n27215,
    ys__n27216, ys__n27217, ys__n27218, ys__n27219, ys__n27220, ys__n27221,
    ys__n27222, ys__n27223, ys__n27224, ys__n27225, ys__n27226, ys__n27227,
    ys__n27228, ys__n27229, ys__n27230, ys__n27231, ys__n27232, ys__n27233,
    ys__n27234, ys__n27235, ys__n27236, ys__n27237, ys__n27238, ys__n27239,
    ys__n27240, ys__n27241, ys__n27242, ys__n27243, ys__n27244, ys__n27245,
    ys__n27246, ys__n27247, ys__n27248, ys__n27249, ys__n27250, ys__n27251,
    ys__n27252, ys__n27253, ys__n27254, ys__n27255, ys__n27256, ys__n27257,
    ys__n27258, ys__n27259, ys__n27260, ys__n27261, ys__n27262, ys__n27263,
    ys__n27264, ys__n27265, ys__n27266, ys__n27267, ys__n27268, ys__n27269,
    ys__n27270, ys__n27271, ys__n27272, ys__n27273, ys__n27274, ys__n27275,
    ys__n27276, ys__n27277, ys__n27278, ys__n27279, ys__n27280, ys__n27281,
    ys__n27282, ys__n27283, ys__n27284, ys__n27285, ys__n27286, ys__n27287,
    ys__n27288, ys__n27289, ys__n27290, ys__n27291, ys__n27292, ys__n27293,
    ys__n27294, ys__n27295, ys__n27296, ys__n27297, ys__n27298, ys__n27299,
    ys__n27300, ys__n27301, ys__n27302, ys__n27303, ys__n27304, ys__n27305,
    ys__n27306, ys__n27307, ys__n27308, ys__n27309, ys__n27310, ys__n27311,
    ys__n27312, ys__n27313, ys__n27314, ys__n27315, ys__n27316, ys__n27317,
    ys__n27318, ys__n27319, ys__n27320, ys__n27321, ys__n27322, ys__n27323,
    ys__n27324, ys__n27325, ys__n27326, ys__n27327, ys__n27328, ys__n27329,
    ys__n27330, ys__n27331, ys__n27332, ys__n27333, ys__n27334, ys__n27335,
    ys__n27336, ys__n27337, ys__n27338, ys__n27339, ys__n27340, ys__n27341,
    ys__n27342, ys__n27343, ys__n27344, ys__n27345, ys__n27346, ys__n27347,
    ys__n27348, ys__n27349, ys__n27350, ys__n27351, ys__n27352, ys__n27353,
    ys__n27354, ys__n27355, ys__n27356, ys__n27357, ys__n27358, ys__n27359,
    ys__n27360, ys__n27361, ys__n27362, ys__n27363, ys__n27364, ys__n27365,
    ys__n27366, ys__n27367, ys__n27368, ys__n27369, ys__n27370, ys__n27371,
    ys__n27372, ys__n27373, ys__n27374, ys__n27375, ys__n27376, ys__n27377,
    ys__n27378, ys__n27379, ys__n27380, ys__n27381, ys__n27382, ys__n27383,
    ys__n27384, ys__n27385, ys__n27386, ys__n27387, ys__n27388, ys__n27389,
    ys__n27390, ys__n27391, ys__n27392, ys__n27393, ys__n27394, ys__n27395,
    ys__n27396, ys__n27397, ys__n27398, ys__n27399, ys__n27400, ys__n27401,
    ys__n27402, ys__n27403, ys__n27404, ys__n27405, ys__n27406, ys__n27407,
    ys__n27408, ys__n27409, ys__n27410, ys__n27411, ys__n27412, ys__n27413,
    ys__n27414, ys__n27415, ys__n27416, ys__n27417, ys__n27418, ys__n27419,
    ys__n27420, ys__n27421, ys__n27422, ys__n27423, ys__n27424, ys__n27425,
    ys__n27426, ys__n27427, ys__n27428, ys__n27429, ys__n27430, ys__n27431,
    ys__n27432, ys__n27433, ys__n27434, ys__n27435, ys__n27436, ys__n27437,
    ys__n27484, ys__n27493, ys__n27504, ys__n27513, ys__n27515, ys__n27517,
    ys__n27550, ys__n27551, ys__n27598, ys__n27603, ys__n27605, ys__n27610,
    ys__n27613, ys__n27616, ys__n27619, ys__n27622, ys__n27625, ys__n27628,
    ys__n27631, ys__n27634, ys__n27637, ys__n27640, ys__n27643, ys__n27646,
    ys__n27649, ys__n27652, ys__n27655, ys__n27658, ys__n27661, ys__n27664,
    ys__n27667, ys__n27670, ys__n27673, ys__n27676, ys__n27679, ys__n27682,
    ys__n27685, ys__n27688, ys__n27691, ys__n27694, ys__n27697, ys__n27700,
    ys__n27703, ys__n27705, ys__n27706, ys__n27707, ys__n27708, ys__n27709,
    ys__n27710, ys__n27711, ys__n27712, ys__n27713, ys__n27714, ys__n27715,
    ys__n27716, ys__n27717, ys__n27718, ys__n27719, ys__n27720, ys__n27721,
    ys__n27722, ys__n27723, ys__n27724, ys__n27725, ys__n27726, ys__n27727,
    ys__n27728, ys__n27729, ys__n27730, ys__n27731, ys__n27732, ys__n27733,
    ys__n27734, ys__n27735, ys__n27736, ys__n27739, ys__n27741, ys__n28247,
    ys__n28249, ys__n28250, ys__n28251, ys__n28252, ys__n28254, ys__n28256,
    ys__n28258, ys__n28259, ys__n28261, ys__n28263, ys__n28265, ys__n28266,
    ys__n28268, ys__n28269, ys__n28270, ys__n28271, ys__n28272, ys__n28274,
    ys__n28276, ys__n28328, ys__n28330, ys__n28332, ys__n28334, ys__n28336,
    ys__n28343, ys__n28345, ys__n28347, ys__n28349, ys__n28351, ys__n28353,
    ys__n28355, ys__n28357, ys__n28359, ys__n28361, ys__n28363, ys__n28365,
    ys__n28367, ys__n28369, ys__n28371, ys__n28373, ys__n28375, ys__n28377,
    ys__n28379, ys__n28381, ys__n28383, ys__n28385, ys__n28387, ys__n28389,
    ys__n28391, ys__n28393, ys__n28395, ys__n28397, ys__n28399, ys__n28401,
    ys__n28403, ys__n28406, ys__n28409, ys__n28410, ys__n28411, ys__n28412,
    ys__n28413, ys__n28414, ys__n28415, ys__n28416, ys__n28417, ys__n28418,
    ys__n28419, ys__n28420, ys__n28421, ys__n28422, ys__n28423, ys__n28425,
    ys__n28427, ys__n28429, ys__n28431, ys__n28433, ys__n28435, ys__n28437,
    ys__n28439, ys__n28440, ys__n28441, ys__n28442, ys__n28443, ys__n28444,
    ys__n28445, ys__n28447, ys__n28448, ys__n28449, ys__n28450, ys__n28451,
    ys__n28452, ys__n28454, ys__n28456, ys__n28458, ys__n28460, ys__n28475,
    ys__n28476, ys__n28477, ys__n28478, ys__n28479, ys__n28480, ys__n28481,
    ys__n28482, ys__n28483, ys__n28484, ys__n28485, ys__n28486, ys__n28487,
    ys__n28488, ys__n28489, ys__n28490, ys__n28491, ys__n28492, ys__n28493,
    ys__n28494, ys__n28495, ys__n28496, ys__n28497, ys__n28498, ys__n28499,
    ys__n28500, ys__n28501, ys__n28502, ys__n28503, ys__n28504, ys__n28505,
    ys__n28506, ys__n28510, ys__n28513, ys__n28518, ys__n28533, ys__n28536,
    ys__n28539, ys__n28542, ys__n28545, ys__n28548, ys__n28551, ys__n28554,
    ys__n28557, ys__n28560, ys__n28563, ys__n28566, ys__n28569, ys__n28572,
    ys__n28575, ys__n28578, ys__n28581, ys__n28584, ys__n28587, ys__n28661,
    ys__n28662, ys__n28781, ys__n28782, ys__n28783, ys__n28784, ys__n28785,
    ys__n28786, ys__n28787, ys__n28788, ys__n28789, ys__n28790, ys__n28791,
    ys__n28792, ys__n28793, ys__n28794, ys__n28796, ys__n28798, ys__n28800,
    ys__n28802, ys__n28804, ys__n28806, ys__n28808, ys__n28810, ys__n28812,
    ys__n28814, ys__n28816, ys__n28818, ys__n28820, ys__n28822, ys__n28824,
    ys__n28826, ys__n28828, ys__n28830, ys__n28832, ys__n28834, ys__n28836,
    ys__n28838, ys__n28840, ys__n28842, ys__n28844, ys__n28846, ys__n28848,
    ys__n28850, ys__n28852, ys__n28854, ys__n28856, ys__n28858, ys__n29022,
    ys__n29025, ys__n29028, ys__n29031, ys__n29034, ys__n29037, ys__n29040,
    ys__n29043, ys__n29046, ys__n29049, ys__n29052, ys__n29055, ys__n29058,
    ys__n29061, ys__n29064, ys__n29067, ys__n29070, ys__n29073, ys__n29076,
    ys__n29079, ys__n29082, ys__n29085, ys__n29088, ys__n29091, ys__n29094,
    ys__n29097, ys__n29100, ys__n29103, ys__n29106, ys__n29109, ys__n29112,
    ys__n29115, ys__n29118, ys__n29122, ys__n29125, ys__n29128, ys__n29131,
    ys__n29134, ys__n29137, ys__n29140, ys__n29143, ys__n29146, ys__n29149,
    ys__n29152, ys__n29155, ys__n29158, ys__n29161, ys__n29164, ys__n29167,
    ys__n29170, ys__n29173, ys__n29176, ys__n29179, ys__n29182, ys__n29185,
    ys__n29188, ys__n29191, ys__n29194, ys__n29197, ys__n29200, ys__n29203,
    ys__n29206, ys__n29209, ys__n29212, ys__n29215, ys__n29217, ys__n29219,
    ys__n29221, ys__n29223, ys__n29225, ys__n29226, ys__n29227, ys__n29228,
    ys__n29229, ys__n29230, ys__n29231, ys__n29232, ys__n29233, ys__n29234,
    ys__n29235, ys__n29336, ys__n29339, ys__n29342, ys__n29345, ys__n29348,
    ys__n29351, ys__n29354, ys__n29357, ys__n29360, ys__n29363, ys__n29366,
    ys__n29369, ys__n29372, ys__n29375, ys__n29378, ys__n29381, ys__n29384,
    ys__n29387, ys__n29390, ys__n29393, ys__n29396, ys__n29399, ys__n29402,
    ys__n29405, ys__n29408, ys__n29411, ys__n29414, ys__n29417, ys__n29420,
    ys__n29423, ys__n29426, ys__n29429, ys__n29431, ys__n29435, ys__n29438,
    ys__n29441, ys__n29444, ys__n29447, ys__n29450, ys__n29453, ys__n29456,
    ys__n29459, ys__n29462, ys__n29465, ys__n29468, ys__n29471, ys__n29474,
    ys__n29477, ys__n29480, ys__n29483, ys__n29486, ys__n29489, ys__n29492,
    ys__n29495, ys__n29498, ys__n29501, ys__n29504, ys__n29507, ys__n29510,
    ys__n29513, ys__n29516, ys__n29519, ys__n29522, ys__n29525, ys__n29528,
    ys__n29530, ys__n29532, ys__n29534, ys__n29536, ys__n29538, ys__n29539,
    ys__n29540, ys__n29541, ys__n29542, ys__n29543, ys__n29544, ys__n29545,
    ys__n29546, ys__n29547, ys__n29548, ys__n29611, ys__n29614, ys__n29617,
    ys__n29620, ys__n29623, ys__n29626, ys__n29629, ys__n29632, ys__n29635,
    ys__n29638, ys__n29641, ys__n29644, ys__n29647, ys__n29650, ys__n29653,
    ys__n29656, ys__n29659, ys__n29662, ys__n29665, ys__n29668, ys__n29671,
    ys__n29674, ys__n29677, ys__n29680, ys__n29683, ys__n29686, ys__n29689,
    ys__n29692, ys__n29695, ys__n29698, ys__n29701, ys__n29704, ys__n29706,
    ys__n29710, ys__n29713, ys__n29716, ys__n29719, ys__n29722, ys__n29725,
    ys__n29728, ys__n29731, ys__n29734, ys__n29737, ys__n29740, ys__n29743,
    ys__n29746, ys__n29749, ys__n29752, ys__n29755, ys__n29758, ys__n29761,
    ys__n29764, ys__n29767, ys__n29770, ys__n29773, ys__n29776, ys__n29779,
    ys__n29782, ys__n29785, ys__n29788, ys__n29791, ys__n29794, ys__n29797,
    ys__n29800, ys__n29803, ys__n29805, ys__n29807, ys__n29809, ys__n29811,
    ys__n29813, ys__n29814, ys__n29815, ys__n29816, ys__n29817, ys__n29818,
    ys__n29819, ys__n29820, ys__n29821, ys__n29822, ys__n29823, ys__n29847,
    ys__n30010, ys__n30080, ys__n30081, ys__n30082, ys__n30083, ys__n30084,
    ys__n30085, ys__n30086, ys__n30087, ys__n30089, ys__n30090, ys__n30091,
    ys__n30092, ys__n30093, ys__n30094, ys__n30095, ys__n30096, ys__n30098,
    ys__n30099, ys__n30100, ys__n30101, ys__n30102, ys__n30103, ys__n30104,
    ys__n30105, ys__n30106, ys__n30107, ys__n30108, ys__n30109, ys__n30110,
    ys__n30111, ys__n30112, ys__n30113, ys__n30119, ys__n30122, ys__n30125,
    ys__n30128, ys__n30131, ys__n30134, ys__n30137, ys__n30140, ys__n30143,
    ys__n30146, ys__n30149, ys__n30152, ys__n30155, ys__n30158, ys__n30161,
    ys__n30164, ys__n30167, ys__n30170, ys__n30173, ys__n30176, ys__n30179,
    ys__n30182, ys__n30185, ys__n30188, ys__n30191, ys__n30194, ys__n30197,
    ys__n30200, ys__n30203, ys__n30206, ys__n30209, ys__n30212, ys__n30215,
    ys__n30223, ys__n30226, ys__n30235, ys__n30238, ys__n30241, ys__n30244,
    ys__n30247, ys__n30250, ys__n30253, ys__n30256, ys__n30259, ys__n30262,
    ys__n30265, ys__n30268, ys__n30271, ys__n30274, ys__n30277, ys__n30280,
    ys__n30283, ys__n30286, ys__n30289, ys__n30292, ys__n30295, ys__n30298,
    ys__n30301, ys__n30304, ys__n30307, ys__n30310, ys__n30313, ys__n30316,
    ys__n30319, ys__n30322, ys__n30325, ys__n30328, ys__n30330, ys__n30331,
    ys__n30616, ys__n30619, ys__n30622, ys__n30625, ys__n30628, ys__n30631,
    ys__n30634, ys__n30637, ys__n30640, ys__n30643, ys__n30646, ys__n30649,
    ys__n30652, ys__n30655, ys__n30658, ys__n30661, ys__n30664, ys__n30667,
    ys__n30668, ys__n30670, ys__n30797, ys__n30798, ys__n30799, ys__n30800,
    ys__n30801, ys__n30802, ys__n30803, ys__n30804, ys__n30805, ys__n30806,
    ys__n30807, ys__n30808, ys__n30809, ys__n30810, ys__n30811, ys__n30812,
    ys__n30813, ys__n30832, ys__n30833, ys__n30835, ys__n30836, ys__n30856,
    ys__n30858, ys__n30860, ys__n30864, ys__n30873, ys__n30874, ys__n30875,
    ys__n30876, ys__n30942, ys__n30943, ys__n30944, ys__n30945, ys__n30946,
    ys__n30947, ys__n30948, ys__n30949, ys__n30950, ys__n30951, ys__n30952,
    ys__n30953, ys__n30954, ys__n30955, ys__n30956, ys__n31202, ys__n31203,
    ys__n31207, ys__n31208, ys__n31209, ys__n31210, ys__n31211, ys__n31212,
    ys__n31213, ys__n31214, ys__n31215, ys__n31216, ys__n31217, ys__n31218,
    ys__n31219, ys__n31220, ys__n31221, ys__n31222, ys__n31223, ys__n31224,
    ys__n31225, ys__n31226, ys__n31227, ys__n31228, ys__n31229, ys__n31230,
    ys__n31231, ys__n31232, ys__n31233, ys__n31234, ys__n31235, ys__n31236,
    ys__n31237, ys__n31238, ys__n31326, ys__n31327, ys__n31328, ys__n31329,
    ys__n31330, ys__n31331, ys__n31332, ys__n31333, ys__n31334, ys__n31335,
    ys__n31336, ys__n31337, ys__n31338, ys__n31339, ys__n31340, ys__n31341,
    ys__n31342, ys__n31343, ys__n31344, ys__n31345, ys__n31346, ys__n31347,
    ys__n31348, ys__n31349, ys__n31350, ys__n31351, ys__n31352, ys__n31353,
    ys__n31354, ys__n31355, ys__n31356, ys__n31357, ys__n31358, ys__n31359,
    ys__n31360, ys__n31361, ys__n31362, ys__n31363, ys__n31364, ys__n31365,
    ys__n31366, ys__n31367, ys__n31368, ys__n31369, ys__n31370, ys__n31371,
    ys__n31372, ys__n31373, ys__n31374, ys__n31375, ys__n31376, ys__n31377,
    ys__n31378, ys__n31379, ys__n31380, ys__n31381, ys__n31382, ys__n31383,
    ys__n31384, ys__n31385, ys__n31386, ys__n31387, ys__n31388, ys__n31389,
    ys__n31390, ys__n31391, ys__n31392, ys__n31393, ys__n31394, ys__n31395,
    ys__n31397, ys__n31398, ys__n31399, ys__n31400, ys__n31401, ys__n31402,
    ys__n31403, ys__n31404, ys__n31405, ys__n31406, ys__n31407, ys__n31408,
    ys__n31409, ys__n31410, ys__n31411, ys__n31412, ys__n31413, ys__n31414,
    ys__n31415, ys__n31416, ys__n31417, ys__n31418, ys__n31419, ys__n31420,
    ys__n31421, ys__n31422, ys__n31423, ys__n31424, ys__n31425, ys__n31426,
    ys__n31427, ys__n31428, ys__n31429, ys__n31430, ys__n31431, ys__n31432,
    ys__n31433, ys__n31434, ys__n31435, ys__n31436, ys__n31437, ys__n31438,
    ys__n31439, ys__n31440, ys__n31441, ys__n31442, ys__n31443, ys__n31444,
    ys__n31445, ys__n31446, ys__n31447, ys__n31448, ys__n31449, ys__n31450,
    ys__n31451, ys__n31452, ys__n31453, ys__n31454, ys__n31455, ys__n31456,
    ys__n31457, ys__n31458, ys__n31459, ys__n31460, ys__n31461, ys__n31462,
    ys__n31463, ys__n31464, ys__n31465, ys__n31466, ys__n31467, ys__n31468,
    ys__n31469, ys__n31470, ys__n31471, ys__n31472, ys__n31473, ys__n31474,
    ys__n31475, ys__n31476, ys__n31477, ys__n31478, ys__n31479, ys__n31480,
    ys__n31481, ys__n31482, ys__n31483, ys__n31484, ys__n31485, ys__n31486,
    ys__n31487, ys__n31488, ys__n31489, ys__n31490, ys__n31491, ys__n31492,
    ys__n31493, ys__n31494, ys__n31495, ys__n31496, ys__n31497, ys__n31498,
    ys__n31499, ys__n31500, ys__n31501, ys__n31502, ys__n31503, ys__n31504,
    ys__n31505, ys__n31506, ys__n31507, ys__n31508, ys__n31509, ys__n31510,
    ys__n31511, ys__n31512, ys__n31513, ys__n31514, ys__n31515, ys__n31516,
    ys__n31517, ys__n31518, ys__n31519, ys__n31520, ys__n31521, ys__n31522,
    ys__n31523, ys__n31524, ys__n31525, ys__n31526, ys__n31527, ys__n31528,
    ys__n31529, ys__n31530, ys__n31531, ys__n31532, ys__n31533, ys__n31534,
    ys__n31535, ys__n31536, ys__n31537, ys__n31538, ys__n31539, ys__n31540,
    ys__n31541, ys__n31542, ys__n31543, ys__n31544, ys__n31559, ys__n31560,
    ys__n31562, ys__n31564, ys__n31567, ys__n31571, ys__n31740, ys__n31741,
    ys__n31742, ys__n31743, ys__n31744, ys__n31745, ys__n31746, ys__n31747,
    ys__n31748, ys__n31749, ys__n31750, ys__n31751, ys__n31752, ys__n31753,
    ys__n31754, ys__n31755, ys__n31756, ys__n31757, ys__n31758, ys__n31759,
    ys__n31760, ys__n31761, ys__n31762, ys__n31763, ys__n31764, ys__n31765,
    ys__n31766, ys__n31767, ys__n31768, ys__n31769, ys__n31770, ys__n31771,
    ys__n31772, ys__n31773, ys__n31774, ys__n31775, ys__n31776, ys__n31777,
    ys__n31778, ys__n31779, ys__n31780, ys__n31781, ys__n31782, ys__n31783,
    ys__n31784, ys__n31785, ys__n31786, ys__n31787, ys__n31788, ys__n31789,
    ys__n31790, ys__n31791, ys__n31792, ys__n31793, ys__n31794, ys__n31795,
    ys__n31796, ys__n31797, ys__n31798, ys__n31799, ys__n31800, ys__n31801,
    ys__n31802, ys__n31803, ys__n31804, ys__n31805, ys__n31806, ys__n31807,
    ys__n31808, ys__n31809, ys__n31810, ys__n31811, ys__n31812, ys__n31813,
    ys__n31814, ys__n31815, ys__n31816, ys__n31817, ys__n31818, ys__n31819,
    ys__n31820, ys__n31821, ys__n31822, ys__n31823, ys__n31824, ys__n31825,
    ys__n31826, ys__n31827, ys__n31828, ys__n31829, ys__n31830, ys__n31831,
    ys__n31832, ys__n31833, ys__n31834, ys__n31835, ys__n31836, ys__n31837,
    ys__n31838, ys__n31839, ys__n31840, ys__n31841, ys__n31842, ys__n31843,
    ys__n31844, ys__n31845, ys__n31846, ys__n31847, ys__n31848, ys__n31849,
    ys__n31850, ys__n31851, ys__n31852, ys__n31853, ys__n31854, ys__n31855,
    ys__n31856, ys__n31857, ys__n31858, ys__n31859, ys__n31860, ys__n31861,
    ys__n31862, ys__n31863, ys__n31864, ys__n31865, ys__n31866, ys__n31867,
    ys__n31868, ys__n31869, ys__n31870, ys__n31871, ys__n31872, ys__n31873,
    ys__n31874, ys__n31875, ys__n31876, ys__n31877, ys__n31878, ys__n31879,
    ys__n31880, ys__n31881, ys__n31882, ys__n31883, ys__n31884, ys__n31885,
    ys__n31886, ys__n31887, ys__n31888, ys__n31889, ys__n31890, ys__n31891,
    ys__n31892, ys__n31893, ys__n31894, ys__n31895, ys__n31896, ys__n31897,
    ys__n31898, ys__n31899, ys__n31900, ys__n31901, ys__n31902, ys__n31903,
    ys__n31904, ys__n31905, ys__n31906, ys__n31907, ys__n31908, ys__n31909,
    ys__n31910, ys__n31911, ys__n31912, ys__n31913, ys__n31914, ys__n31915,
    ys__n31916, ys__n31917, ys__n31918, ys__n31919, ys__n31920, ys__n31921,
    ys__n31922, ys__n31923, ys__n31924, ys__n31925, ys__n31926, ys__n31927,
    ys__n31928, ys__n31929, ys__n31930, ys__n31931, ys__n31932, ys__n31933,
    ys__n31934, ys__n31935, ys__n31936, ys__n31937, ys__n31938, ys__n31939,
    ys__n31940, ys__n31941, ys__n31942, ys__n31943, ys__n31944, ys__n31945,
    ys__n31946, ys__n31947, ys__n31948, ys__n31949, ys__n31950, ys__n31953,
    ys__n31954, ys__n31955, ys__n31965, ys__n31971, ys__n31973, ys__n31975,
    ys__n31976, ys__n31978, ys__n31979, ys__n31984, ys__n31986, ys__n31988,
    ys__n31990, ys__n31992, ys__n31994, ys__n31996, ys__n31998, ys__n32000,
    ys__n32002, ys__n32004, ys__n32006, ys__n32007, ys__n32008, ys__n32010,
    ys__n32012, ys__n32014, ys__n32016, ys__n32018, ys__n32022, ys__n32023,
    ys__n32024, ys__n32025, ys__n32026, ys__n32027, ys__n32028, ys__n32029,
    ys__n32030, ys__n32031, ys__n32032, ys__n32033, ys__n32034, ys__n32035,
    ys__n32036, ys__n32037, ys__n32038, ys__n32039, ys__n32040, ys__n32041,
    ys__n32042, ys__n32043, ys__n32044, ys__n32045, ys__n32046, ys__n32047,
    ys__n32048, ys__n32049, ys__n32050, ys__n32051, ys__n32052, ys__n32053,
    ys__n32054, ys__n32055, ys__n32056, ys__n32057, ys__n32058, ys__n32059,
    ys__n32060, ys__n32061, ys__n32062, ys__n32063, ys__n32064, ys__n32065,
    ys__n32066, ys__n32067, ys__n32068, ys__n32069, ys__n32070, ys__n32071,
    ys__n32072, ys__n32073, ys__n32074, ys__n32075, ys__n32076, ys__n32077,
    ys__n32078, ys__n32079, ys__n32080, ys__n32081, ys__n32082, ys__n32083,
    ys__n32084, ys__n32085, ys__n32086, ys__n32087, ys__n32088, ys__n32124,
    ys__n32125, ys__n32126, ys__n32127, ys__n32128, ys__n32129, ys__n32130,
    ys__n32131, ys__n32132, ys__n32133, ys__n32134, ys__n32135, ys__n32136,
    ys__n32137, ys__n32138, ys__n32139, ys__n32140, ys__n32141, ys__n32142,
    ys__n32143, ys__n32144, ys__n32145, ys__n32146, ys__n32147, ys__n32148,
    ys__n32149, ys__n32150, ys__n32151, ys__n32152, ys__n32153, ys__n32154,
    ys__n32155, ys__n32158, ys__n32159, ys__n32160, ys__n32161, ys__n32162,
    ys__n32163, ys__n32164, ys__n32165, ys__n32166, ys__n32167, ys__n32168,
    ys__n32169, ys__n32170, ys__n32171, ys__n32172, ys__n32173, ys__n32174,
    ys__n32175, ys__n32176, ys__n32177, ys__n32178, ys__n32179, ys__n32180,
    ys__n32181, ys__n32182, ys__n32183, ys__n32184, ys__n32185, ys__n32186,
    ys__n32187, ys__n32188, ys__n32189, ys__n32190, ys__n32191, ys__n32192,
    ys__n32193, ys__n32194, ys__n32195, ys__n32196, ys__n32197, ys__n32198,
    ys__n32199, ys__n32200, ys__n32201, ys__n32202, ys__n32203, ys__n32204,
    ys__n32205, ys__n32206, ys__n32207, ys__n32208, ys__n32209, ys__n32210,
    ys__n32211, ys__n32212, ys__n32213, ys__n32214, ys__n32215, ys__n32216,
    ys__n32217, ys__n32218, ys__n32219, ys__n32220, ys__n32221, ys__n32222,
    ys__n32223, ys__n32224, ys__n32225, ys__n32226, ys__n32227, ys__n32228,
    ys__n32229, ys__n32230, ys__n32231, ys__n32232, ys__n32233, ys__n32234,
    ys__n32235, ys__n32236, ys__n32237, ys__n32238, ys__n32239, ys__n32240,
    ys__n32241, ys__n32242, ys__n32243, ys__n32244, ys__n32245, ys__n32246,
    ys__n32247, ys__n32248, ys__n32249, ys__n32250, ys__n32251, ys__n32252,
    ys__n32253, ys__n32254, ys__n32255, ys__n32256, ys__n32257, ys__n32258,
    ys__n32259, ys__n32260, ys__n32261, ys__n32262, ys__n32263, ys__n32264,
    ys__n32265, ys__n32266, ys__n32267, ys__n32268, ys__n32269, ys__n32270,
    ys__n32271, ys__n32272, ys__n32273, ys__n32274, ys__n32275, ys__n32276,
    ys__n32277, ys__n32278, ys__n32279, ys__n32280, ys__n32281, ys__n32282,
    ys__n32283, ys__n32284, ys__n32285, ys__n32286, ys__n32287, ys__n32288,
    ys__n32289, ys__n32290, ys__n32291, ys__n32292, ys__n32293, ys__n32294,
    ys__n32295, ys__n32296, ys__n32297, ys__n32298, ys__n32299, ys__n32300,
    ys__n32301, ys__n32302, ys__n32303, ys__n32304, ys__n32305, ys__n32306,
    ys__n32307, ys__n32308, ys__n32309, ys__n32310, ys__n32311, ys__n32312,
    ys__n32313, ys__n32314, ys__n32315, ys__n32316, ys__n32317, ys__n32318,
    ys__n32319, ys__n32320, ys__n32321, ys__n32322, ys__n32323, ys__n32324,
    ys__n32325, ys__n32326, ys__n32327, ys__n32328, ys__n32329, ys__n32330,
    ys__n32331, ys__n32332, ys__n32333, ys__n32334, ys__n32335, ys__n32336,
    ys__n32337, ys__n32338, ys__n32339, ys__n32340, ys__n32341, ys__n32342,
    ys__n32343, ys__n32344, ys__n32345, ys__n32346, ys__n32347, ys__n32348,
    ys__n32349, ys__n32350, ys__n32351, ys__n32352, ys__n32353, ys__n32354,
    ys__n32355, ys__n32356, ys__n32357, ys__n32358, ys__n32359, ys__n32360,
    ys__n32361, ys__n32362, ys__n32363, ys__n32364, ys__n32365, ys__n32366,
    ys__n32367, ys__n32368, ys__n32369, ys__n32370, ys__n32371, ys__n32372,
    ys__n32373, ys__n32374, ys__n32375, ys__n32376, ys__n32377, ys__n32378,
    ys__n32379, ys__n32380, ys__n32381, ys__n32382, ys__n32383, ys__n32384,
    ys__n32385, ys__n32386, ys__n32387, ys__n32388, ys__n32389, ys__n32390,
    ys__n32391, ys__n32392, ys__n32393, ys__n32394, ys__n32395, ys__n32396,
    ys__n32397, ys__n32398, ys__n32399, ys__n32400, ys__n32401, ys__n32402,
    ys__n32403, ys__n32404, ys__n32405, ys__n32406, ys__n32407, ys__n32408,
    ys__n32409, ys__n32410, ys__n32411, ys__n32412, ys__n32413, ys__n32414,
    ys__n32415, ys__n32416, ys__n32417, ys__n32418, ys__n32419, ys__n32420,
    ys__n32421, ys__n32422, ys__n32423, ys__n32424, ys__n32425, ys__n32426,
    ys__n32427, ys__n32428, ys__n32429, ys__n32430, ys__n32431, ys__n32432,
    ys__n32433, ys__n32434, ys__n32435, ys__n32436, ys__n32437, ys__n32438,
    ys__n32439, ys__n32440, ys__n32441, ys__n32442, ys__n32443, ys__n32444,
    ys__n32445, ys__n32446, ys__n32447, ys__n32448, ys__n32449, ys__n32450,
    ys__n32451, ys__n32452, ys__n32453, ys__n32454, ys__n32455, ys__n32456,
    ys__n32457, ys__n32458, ys__n32459, ys__n32460, ys__n32461, ys__n32462,
    ys__n32463, ys__n32464, ys__n32465, ys__n32466, ys__n32467, ys__n32468,
    ys__n32469, ys__n32470, ys__n32471, ys__n32472, ys__n32473, ys__n32474,
    ys__n32475, ys__n32476, ys__n32477, ys__n32478, ys__n32479, ys__n32480,
    ys__n32481, ys__n32482, ys__n32483, ys__n32484, ys__n32485, ys__n32486,
    ys__n32487, ys__n32488, ys__n32489, ys__n32490, ys__n32491, ys__n32492,
    ys__n32493, ys__n32494, ys__n32495, ys__n32496, ys__n32497, ys__n32498,
    ys__n32499, ys__n32500, ys__n32501, ys__n32502, ys__n32503, ys__n32504,
    ys__n32505, ys__n32506, ys__n32507, ys__n32508, ys__n32509, ys__n32510,
    ys__n32511, ys__n32512, ys__n32513, ys__n32514, ys__n32515, ys__n32516,
    ys__n32517, ys__n32518, ys__n32519, ys__n32520, ys__n32521, ys__n32522,
    ys__n32523, ys__n32524, ys__n32525, ys__n32526, ys__n32527, ys__n32528,
    ys__n32529, ys__n32530, ys__n32531, ys__n32532, ys__n32533, ys__n32534,
    ys__n32535, ys__n32536, ys__n32537, ys__n32538, ys__n32539, ys__n32540,
    ys__n32541, ys__n32542, ys__n32543, ys__n32544, ys__n32545, ys__n32546,
    ys__n32547, ys__n32548, ys__n32549, ys__n32550, ys__n32551, ys__n32552,
    ys__n32553, ys__n32554, ys__n32555, ys__n32556, ys__n32557, ys__n32558,
    ys__n32559, ys__n32560, ys__n32561, ys__n32562, ys__n32563, ys__n32564,
    ys__n32565, ys__n32566, ys__n32567, ys__n32568, ys__n32569, ys__n32570,
    ys__n32571, ys__n32572, ys__n32573, ys__n32574, ys__n32575, ys__n32576,
    ys__n32577, ys__n32578, ys__n32579, ys__n32580, ys__n32581, ys__n32582,
    ys__n32583, ys__n32584, ys__n32585, ys__n32586, ys__n32587, ys__n32588,
    ys__n32589, ys__n32590, ys__n32591, ys__n32592, ys__n32593, ys__n32594,
    ys__n32595, ys__n32596, ys__n32597, ys__n32598, ys__n32599, ys__n32600,
    ys__n32601, ys__n32602, ys__n32603, ys__n32604, ys__n32605, ys__n32606,
    ys__n32607, ys__n32608, ys__n32609, ys__n32610, ys__n32611, ys__n32612,
    ys__n32613, ys__n32614, ys__n32615, ys__n32616, ys__n32617, ys__n32618,
    ys__n32619, ys__n32620, ys__n32621, ys__n32622, ys__n32623, ys__n32624,
    ys__n32625, ys__n32626, ys__n32627, ys__n32628, ys__n32629, ys__n32630,
    ys__n32631, ys__n32632, ys__n32633, ys__n32634, ys__n32635, ys__n32636,
    ys__n32637, ys__n32638, ys__n32639, ys__n32640, ys__n32641, ys__n32642,
    ys__n32643, ys__n32644, ys__n32645, ys__n32646, ys__n32647, ys__n32648,
    ys__n32649, ys__n32650, ys__n32651, ys__n32652, ys__n32653, ys__n32654,
    ys__n32655, ys__n32656, ys__n32657, ys__n32658, ys__n32659, ys__n32660,
    ys__n32661, ys__n32662, ys__n32663, ys__n32664, ys__n32665, ys__n32666,
    ys__n32667, ys__n32668, ys__n32669, ys__n32670, ys__n32671, ys__n32672,
    ys__n32673, ys__n32674, ys__n32675, ys__n32676, ys__n32677, ys__n32678,
    ys__n32679, ys__n32680, ys__n32681, ys__n32682, ys__n32683, ys__n32684,
    ys__n32685, ys__n32686, ys__n32687, ys__n32688, ys__n32689, ys__n32690,
    ys__n32691, ys__n32692, ys__n32693, ys__n32694, ys__n32695, ys__n32696,
    ys__n32697, ys__n32698, ys__n32699, ys__n32700, ys__n32701, ys__n32702,
    ys__n32703, ys__n32704, ys__n32705, ys__n32706, ys__n32707, ys__n32708,
    ys__n32709, ys__n32710, ys__n32711, ys__n32712, ys__n32713, ys__n32714,
    ys__n32715, ys__n32716, ys__n32717, ys__n32718, ys__n32719, ys__n32720,
    ys__n32721, ys__n32722, ys__n32723, ys__n32724, ys__n32725, ys__n32726,
    ys__n32727, ys__n32728, ys__n32729, ys__n32730, ys__n32731, ys__n32732,
    ys__n32733, ys__n32734, ys__n32735, ys__n32736, ys__n32737, ys__n32738,
    ys__n32739, ys__n32740, ys__n32741, ys__n32742, ys__n32743, ys__n32744,
    ys__n32745, ys__n32746, ys__n32747, ys__n32748, ys__n32749, ys__n32750,
    ys__n32751, ys__n32752, ys__n32753, ys__n32754, ys__n32755, ys__n32756,
    ys__n32757, ys__n32758, ys__n32759, ys__n32760, ys__n32761, ys__n32762,
    ys__n32763, ys__n32764, ys__n32765, ys__n32766, ys__n32767, ys__n32768,
    ys__n32769, ys__n32770, ys__n32771, ys__n32772, ys__n32773, ys__n32774,
    ys__n32775, ys__n32776, ys__n32777, ys__n32778, ys__n32779, ys__n32780,
    ys__n32781, ys__n32782, ys__n32783, ys__n32784, ys__n32785, ys__n32786,
    ys__n32787, ys__n32788, ys__n32789, ys__n32790, ys__n32791, ys__n32792,
    ys__n32793, ys__n32794, ys__n32795, ys__n32796, ys__n32797, ys__n32798,
    ys__n32799, ys__n32800, ys__n32801, ys__n32802, ys__n32803, ys__n32804,
    ys__n32805, ys__n32806, ys__n32807, ys__n32808, ys__n32809, ys__n32810,
    ys__n32811, ys__n32812, ys__n32813, ys__n32814, ys__n32815, ys__n32816,
    ys__n32817, ys__n32818, ys__n32819, ys__n32820, ys__n32821, ys__n32822,
    ys__n32823, ys__n32824, ys__n32825, ys__n32826, ys__n32827, ys__n32828,
    ys__n32829, ys__n32830, ys__n32831, ys__n32832, ys__n32833, ys__n32834,
    ys__n32835, ys__n32836, ys__n32837, ys__n32838, ys__n32839, ys__n32840,
    ys__n32841, ys__n32842, ys__n32843, ys__n32844, ys__n32845, ys__n32846,
    ys__n32847, ys__n32848, ys__n32849, ys__n32850, ys__n32851, ys__n32852,
    ys__n32853, ys__n32854, ys__n32855, ys__n32856, ys__n32857, ys__n32858,
    ys__n32859, ys__n32860, ys__n32861, ys__n32862, ys__n32863, ys__n32864,
    ys__n32865, ys__n32866, ys__n32867, ys__n32868, ys__n32869, ys__n32870,
    ys__n32871, ys__n32872, ys__n32873, ys__n32874, ys__n32875, ys__n32876,
    ys__n32877, ys__n32878, ys__n32879, ys__n32880, ys__n32881, ys__n32882,
    ys__n32883, ys__n32884, ys__n32885, ys__n32886, ys__n32887, ys__n32888,
    ys__n32889, ys__n32890, ys__n32891, ys__n32892, ys__n32893, ys__n32894,
    ys__n32895, ys__n32896, ys__n32897, ys__n32898, ys__n32899, ys__n32900,
    ys__n32901, ys__n32902, ys__n32903, ys__n32904, ys__n32905, ys__n32906,
    ys__n32907, ys__n32908, ys__n32909, ys__n32910, ys__n32911, ys__n32912,
    ys__n32913, ys__n32914, ys__n32915, ys__n32916, ys__n32917, ys__n32918,
    ys__n32919, ys__n32920, ys__n32921, ys__n32922, ys__n32923, ys__n32924,
    ys__n32925, ys__n32926, ys__n32927, ys__n32928, ys__n32929, ys__n32930,
    ys__n32931, ys__n32932, ys__n32933, ys__n32934, ys__n32935, ys__n32936,
    ys__n32937, ys__n32938, ys__n32939, ys__n32940, ys__n32941, ys__n32942,
    ys__n32943, ys__n32944, ys__n32945, ys__n32946, ys__n32947, ys__n32948,
    ys__n32949, ys__n32950, ys__n32951, ys__n32952, ys__n32953, ys__n32954,
    ys__n32955, ys__n32956, ys__n32957, ys__n32958, ys__n32959, ys__n32960,
    ys__n32961, ys__n32962, ys__n32963, ys__n32964, ys__n32965, ys__n32966,
    ys__n32967, ys__n32968, ys__n32969, ys__n32970, ys__n32971, ys__n32972,
    ys__n32973, ys__n32974, ys__n32975, ys__n32976, ys__n32977, ys__n32978,
    ys__n32979, ys__n32980, ys__n32981, ys__n32982, ys__n32983, ys__n32984,
    ys__n32985, ys__n32986, ys__n32987, ys__n32988, ys__n32989, ys__n32990,
    ys__n32991, ys__n32992, ys__n32993, ys__n32994, ys__n32995, ys__n32996,
    ys__n32997, ys__n32998, ys__n33007, ys__n33008, ys__n33009, ys__n33014,
    ys__n33015, ys__n33016, ys__n33017, ys__n33018, ys__n33019, ys__n33020,
    ys__n33021, ys__n33022, ys__n33023, ys__n33024, ys__n33025, ys__n33026,
    ys__n33027, ys__n33028, ys__n33029, ys__n33030, ys__n33031, ys__n33032,
    ys__n33033, ys__n33034, ys__n33035, ys__n33036, ys__n33037, ys__n33038,
    ys__n33039, ys__n33040, ys__n33041, ys__n33042, ys__n33043, ys__n33044,
    ys__n33045, ys__n33046, ys__n33047, ys__n33048, ys__n33049, ys__n33050,
    ys__n33051, ys__n33052, ys__n33053, ys__n33054, ys__n33055, ys__n33056,
    ys__n33058, ys__n33059, ys__n33060, ys__n33061, ys__n33062, ys__n33063,
    ys__n33064, ys__n33065, ys__n33066, ys__n33067, ys__n33068, ys__n33069,
    ys__n33070, ys__n33071, ys__n33072, ys__n33073, ys__n33074, ys__n33075,
    ys__n33076, ys__n33077, ys__n33078, ys__n33079, ys__n33080, ys__n33081,
    ys__n33082, ys__n33083, ys__n33084, ys__n33085, ys__n33086, ys__n33087,
    ys__n33088, ys__n33089, ys__n33090, ys__n33091, ys__n33092, ys__n33093,
    ys__n33094, ys__n33095, ys__n33096, ys__n33097, ys__n33098, ys__n33099,
    ys__n33100, ys__n33101, ys__n33102, ys__n33103, ys__n33104, ys__n33105,
    ys__n33106, ys__n33107, ys__n33108, ys__n33109, ys__n33110, ys__n33111,
    ys__n33178, ys__n33179, ys__n33180, ys__n33181, ys__n33182, ys__n33183,
    ys__n33184, ys__n33185, ys__n33186, ys__n33187, ys__n33188, ys__n33189,
    ys__n33190, ys__n33191, ys__n33192, ys__n33193, ys__n33194, ys__n33195,
    ys__n33196, ys__n33197, ys__n33198, ys__n33199, ys__n33200, ys__n33201,
    ys__n33202, ys__n33203, ys__n33204, ys__n33205, ys__n33206, ys__n33207,
    ys__n33208, ys__n33209, ys__n33211, ys__n33317, ys__n33324, ys__n33329,
    ys__n33331, ys__n33333, ys__n33335, ys__n33337, ys__n33339, ys__n33357,
    ys__n33366, ys__n33414, ys__n33420, ys__n33437, ys__n33438, ys__n33439,
    ys__n33453, ys__n33454, ys__n33455, ys__n33456, ys__n33457, ys__n33513,
    ys__n33514, ys__n33515, ys__n33521, ys__n33535, ys__n34952, ys__n34953,
    ys__n34962, ys__n35052, ys__n35144, ys__n35146, ys__n35148, ys__n35150,
    ys__n35152, ys__n35154, ys__n35156, ys__n35158, ys__n35160, ys__n35162,
    ys__n35164, ys__n35166, ys__n35168, ys__n35170, ys__n35172, ys__n35174,
    ys__n35176, ys__n35178, ys__n35180, ys__n35182, ys__n35184, ys__n35186,
    ys__n35188, ys__n35190, ys__n35192, ys__n35194, ys__n35196, ys__n35198,
    ys__n35200, ys__n35202, ys__n35204, ys__n35206, ys__n35402, ys__n35404,
    ys__n35406, ys__n35408, ys__n35410, ys__n35412, ys__n35425, ys__n35705,
    ys__n35706, ys__n35708, ys__n35710, ys__n35712, ys__n35714, ys__n35716,
    ys__n37676, ys__n37687, ys__n37695, ys__n37697, ys__n37699, ys__n37702,
    ys__n37703, ys__n37707, ys__n37714, ys__n37731, ys__n37732, ys__n37733,
    ys__n37738, ys__n37739, ys__n37741, ys__n37742, ys__n38180, ys__n38182,
    ys__n38184, ys__n38185, ys__n38186, ys__n38188, ys__n38191, ys__n38205,
    ys__n38207, ys__n38209, ys__n38211, ys__n38213, ys__n38214, ys__n38216,
    ys__n38218, ys__n38222, ys__n38224, ys__n38246, ys__n38247, ys__n38248,
    ys__n38250, ys__n38252, ys__n38263, ys__n38266, ys__n38281, ys__n38285,
    ys__n38287, ys__n38289, ys__n38292, ys__n38294, ys__n38296, ys__n38303,
    ys__n38325, ys__n38326, ys__n38327, ys__n38328, ys__n38330, ys__n38331,
    ys__n38332, ys__n38334, ys__n38336, ys__n38337, ys__n38338, ys__n38339,
    ys__n38340, ys__n38341, ys__n38342, ys__n38343, ys__n38344, ys__n38345,
    ys__n38347, ys__n38349, ys__n38351, ys__n38352, ys__n38353, ys__n38354,
    ys__n38355, ys__n38356, ys__n38357, ys__n38359, ys__n38360, ys__n38362,
    ys__n38364, ys__n38365, ys__n38366, ys__n38367, ys__n38368, ys__n38369,
    ys__n38370, ys__n38371, ys__n38372, ys__n38373, ys__n38374, ys__n38375,
    ys__n38377, ys__n38379, ys__n38381, ys__n38383, ys__n38385, ys__n38387,
    ys__n38388, ys__n38389, ys__n38390, ys__n38391, ys__n38392, ys__n38393,
    ys__n38394, ys__n38396, ys__n38397, ys__n38417, ys__n38453, ys__n38456,
    ys__n38508, ys__n38509, ys__n38510, ys__n38515, ys__n38518, ys__n38520,
    ys__n38521, ys__n38523, ys__n38525, ys__n38552, ys__n38555, ys__n38556,
    ys__n38563, ys__n38566, ys__n38615, ys__n38623, ys__n38628, ys__n38633,
    ys__n38650, ys__n38662, ys__n38668, ys__n38669, ys__n38672, ys__n38674,
    ys__n38677, ys__n38689, ys__n38742, ys__n38768, ys__n38795, ys__n38799,
    ys__n38801, ys__n38884, ys__n38886, ys__n38887, ys__n38900, ys__n38912,
    ys__n38913, ys__n38914, ys__n38915, ys__n38917, ys__n38923, ys__n38925,
    ys__n38930, ys__n39392, ys__n39393, ys__n39395, ys__n39396, ys__n39397,
    ys__n39398, ys__n39399, ys__n39400, ys__n39401, ys__n39402, ys__n39403,
    ys__n39404, ys__n39405, ys__n39406, ys__n39407, ys__n39408, ys__n39409,
    ys__n39410, ys__n39411, ys__n39412, ys__n39413, ys__n39414, ys__n39415,
    ys__n39416, ys__n39417, ys__n39418, ys__n40052, ys__n42129, ys__n42153,
    ys__n42189, ys__n42194, ys__n42229, ys__n42234, ys__n42270, ys__n42275,
    ys__n42311, ys__n42316, ys__n42352, ys__n42357, ys__n42393, ys__n42398,
    ys__n42434, ys__n42439, ys__n42488, ys__n42493, ys__n42541, ys__n42546,
    ys__n42594, ys__n42599, ys__n42647, ys__n42652, ys__n42701, ys__n42706,
    ys__n42755, ys__n42760, ys__n42809, ys__n42814, ys__n42863, ys__n42868,
    ys__n42917, ys__n42922, ys__n42971, ys__n42976, ys__n43025, ys__n43030,
    ys__n43079, ys__n43084, ys__n43133, ys__n43138, ys__n43187, ys__n43192,
    ys__n43241, ys__n43246, ys__n43295, ys__n43300, ys__n43349, ys__n43354,
    ys__n43403, ys__n43408, ys__n43457, ys__n43462, ys__n43511, ys__n43516,
    ys__n43565, ys__n43570, ys__n43619, ys__n43624, ys__n43673, ys__n43678,
    ys__n43727, ys__n43732, ys__n43781, ys__n43786, ys__n43835, ys__n43840,
    ys__n43889, ys__n43894, ys__n43932, ys__n43937, ys__n43975, ys__n43980,
    ys__n44018, ys__n44023, ys__n44048, ys__n44053, ys__n44089, ys__n44094,
    ys__n44119, ys__n44122, ys__n44136, ys__n44139, ys__n44155, ys__n44160,
    ys__n44183, ys__n44186, ys__n44189, ys__n44192, ys__n44195, ys__n44198,
    ys__n44205, ys__n44213, ys__n44216, ys__n44219, ys__n44836, ys__n44838,
    ys__n44841, ys__n44843, ys__n44844, ys__n44845, ys__n44846, ys__n44848,
    ys__n44850, ys__n44851, ys__n44852, ys__n44853, ys__n44854, ys__n44855,
    ys__n44858, ys__n44948, ys__n44949, ys__n44950, ys__n44952, ys__n44953,
    ys__n44954, ys__n44955, ys__n44956, ys__n44957, ys__n44958, ys__n44959,
    ys__n44960, ys__n44961, ys__n44962, ys__n44963, ys__n44964, ys__n44965,
    ys__n44966, ys__n44967, ys__n44968, ys__n44969, ys__n44970, ys__n44971,
    ys__n44972, ys__n44973, ys__n44974, ys__n44975, ys__n44976, ys__n44977,
    ys__n44978, ys__n44979, ys__n44980, ys__n44981, ys__n44982, ys__n44983,
    ys__n44985, ys__n44987, ys__n46131, ys__n46133, ys__n46135, ys__n46137,
    ys__n46143, ys__n46146, ys__n46154, ys__n46155, ys__n46158, ys__n46159,
    ys__n46162, ys__n46163, ys__n46172, ys__n46173, ys__n46176, ys__n46179,
    ys__n46188, ys__n46189, ys__n46192, ys__n46195, ys__n46204, ys__n46205,
    ys__n46208, ys__n46211, ys__n46220, ys__n46221, ys__n46224, ys__n46227,
    ys__n46233, ys__n46234, ys__n48339, ys__n48340, ys__n48341, ys__n48342,
    ys__n48343, ys__n48344, ys__n48348, ys__n48349, ys__n48350, ys__n48351,
    ys__n48352, ys__n48353, ys__n48354, ys__n48355, ys__n48356, ys__n48357,
    ys__n48358, ys__n48359, ys__n48360, ys__n48361, ys__n48362  );
  input  ys__n14, ys__n16, ys__n22, ys__n24, ys__n26, ys__n28, ys__n30,
    ys__n32, ys__n34, ys__n36, ys__n38, ys__n40, ys__n42, ys__n44, ys__n46,
    ys__n48, ys__n50, ys__n52, ys__n54, ys__n56, ys__n58, ys__n60, ys__n62,
    ys__n66, ys__n70, ys__n72, ys__n74, ys__n76, ys__n78, ys__n80, ys__n82,
    ys__n84, ys__n86, ys__n88, ys__n90, ys__n96, ys__n98, ys__n100,
    ys__n108, ys__n110, ys__n112, ys__n114, ys__n116, ys__n118, ys__n120,
    ys__n122, ys__n124, ys__n126, ys__n128, ys__n130, ys__n132, ys__n134,
    ys__n136, ys__n138, ys__n140, ys__n142, ys__n148, ys__n150, ys__n152,
    ys__n156, ys__n158, ys__n160, ys__n162, ys__n164, ys__n166, ys__n168,
    ys__n170, ys__n172, ys__n174, ys__n176, ys__n178, ys__n182, ys__n184,
    ys__n186, ys__n190, ys__n192, ys__n194, ys__n196, ys__n198, ys__n202,
    ys__n204, ys__n206, ys__n208, ys__n210, ys__n212, ys__n214, ys__n216,
    ys__n218, ys__n220, ys__n222, ys__n226, ys__n232, ys__n238, ys__n240,
    ys__n242, ys__n244, ys__n248, ys__n256, ys__n258, ys__n262, ys__n290,
    ys__n294, ys__n296, ys__n298, ys__n300, ys__n302, ys__n304, ys__n306,
    ys__n308, ys__n310, ys__n312, ys__n314, ys__n316, ys__n318, ys__n326,
    ys__n328, ys__n330, ys__n332, ys__n336, ys__n338, ys__n340, ys__n342,
    ys__n344, ys__n346, ys__n348, ys__n350, ys__n352, ys__n354, ys__n356,
    ys__n358, ys__n360, ys__n362, ys__n364, ys__n366, ys__n368, ys__n370,
    ys__n372, ys__n374, ys__n376, ys__n378, ys__n380, ys__n382, ys__n384,
    ys__n386, ys__n392, ys__n394, ys__n396, ys__n398, ys__n402, ys__n408,
    ys__n414, ys__n416, ys__n418, ys__n420, ys__n422, ys__n424, ys__n426,
    ys__n428, ys__n430, ys__n432, ys__n434, ys__n436, ys__n438, ys__n440,
    ys__n442, ys__n444, ys__n446, ys__n448, ys__n450, ys__n452, ys__n454,
    ys__n456, ys__n464, ys__n488, ys__n490, ys__n500, ys__n504, ys__n512,
    ys__n514, ys__n516, ys__n518, ys__n520, ys__n522, ys__n524, ys__n526,
    ys__n528, ys__n530, ys__n532, ys__n536, ys__n538, ys__n544, ys__n546,
    ys__n548, ys__n550, ys__n556, ys__n558, ys__n562, ys__n564, ys__n566,
    ys__n568, ys__n570, ys__n572, ys__n580, ys__n582, ys__n584, ys__n586,
    ys__n588, ys__n598, ys__n600, ys__n602, ys__n604, ys__n606, ys__n608,
    ys__n610, ys__n612, ys__n614, ys__n616, ys__n618, ys__n620, ys__n622,
    ys__n624, ys__n626, ys__n632, ys__n634, ys__n636, ys__n638, ys__n640,
    ys__n642, ys__n644, ys__n646, ys__n648, ys__n650, ys__n652, ys__n654,
    ys__n656, ys__n658, ys__n660, ys__n662, ys__n664, ys__n666, ys__n668,
    ys__n670, ys__n672, ys__n674, ys__n676, ys__n678, ys__n680, ys__n682,
    ys__n684, ys__n686, ys__n688, ys__n690, ys__n692, ys__n694, ys__n696,
    ys__n698, ys__n700, ys__n702, ys__n704, ys__n706, ys__n708, ys__n710,
    ys__n712, ys__n718, ys__n720, ys__n722, ys__n724, ys__n726, ys__n728,
    ys__n736, ys__n742, ys__n744, ys__n746, ys__n748, ys__n750, ys__n752,
    ys__n758, ys__n760, ys__n762, ys__n764, ys__n766, ys__n768, ys__n770,
    ys__n772, ys__n774, ys__n776, ys__n778, ys__n780, ys__n782, ys__n784,
    ys__n816, ys__n818, ys__n820, ys__n822, ys__n824, ys__n826, ys__n828,
    ys__n830, ys__n832, ys__n834, ys__n836, ys__n838, ys__n840, ys__n842,
    ys__n844, ys__n846, ys__n848, ys__n850, ys__n852, ys__n854, ys__n856,
    ys__n858, ys__n860, ys__n874, ys__n889, ys__n935, ys__n1029, ys__n1036,
    ys__n1038, ys__n1048, ys__n1072, ys__n1076, ys__n1078, ys__n1084,
    ys__n1094, ys__n1098, ys__n1099, ys__n1106, ys__n1107, ys__n1109,
    ys__n1110, ys__n1116, ys__n1117, ys__n1119, ys__n1120, ys__n1129,
    ys__n1147, ys__n1151, ys__n1153, ys__n1154, ys__n1156, ys__n1157,
    ys__n1301, ys__n1309, ys__n1489, ys__n1490, ys__n1492, ys__n1493,
    ys__n1495, ys__n1496, ys__n1498, ys__n1499, ys__n1502, ys__n1503,
    ys__n1505, ys__n1506, ys__n1508, ys__n1509, ys__n1511, ys__n1535,
    ys__n2024, ys__n2233, ys__n2239, ys__n2245, ys__n2247, ys__n2251,
    ys__n2276, ys__n2282, ys__n2306, ys__n2308, ys__n2312, ys__n2427,
    ys__n2429, ys__n2433, ys__n2644, ys__n2652, ys__n2693, ys__n2716,
    ys__n2779, ys__n2830, ys__n2924, ys__n3214, ys__n4168, ys__n4176,
    ys__n4177, ys__n4184, ys__n4185, ys__n4190, ys__n4291, ys__n4292,
    ys__n4294, ys__n4296, ys__n4297, ys__n4299, ys__n4300, ys__n4305,
    ys__n4340, ys__n4448, ys__n4449, ys__n4451, ys__n4452, ys__n4454,
    ys__n4455, ys__n4457, ys__n4458, ys__n4460, ys__n4461, ys__n4465,
    ys__n4478, ys__n4480, ys__n4488, ys__n4494, ys__n4496, ys__n4613,
    ys__n4625, ys__n4627, ys__n4688, ys__n4698, ys__n4736, ys__n4744,
    ys__n4746, ys__n4750, ys__n4751, ys__n4753, ys__n4754, ys__n4756,
    ys__n4757, ys__n4759, ys__n4761, ys__n4783, ys__n4784, ys__n4810,
    ys__n4826, ys__n4832, ys__n4833, ys__n4836, ys__n4837, ys__n6112,
    ys__n6113, ys__n6115, ys__n6118, ys__n6119, ys__n6120, ys__n6121,
    ys__n6123, ys__n6124, ys__n6126, ys__n6127, ys__n6129, ys__n6130,
    ys__n6133, ys__n6134, ys__n17803, ys__n17804, ys__n17806, ys__n17807,
    ys__n17809, ys__n17810, ys__n17812, ys__n17813, ys__n17815, ys__n17816,
    ys__n17818, ys__n17819, ys__n17821, ys__n17822, ys__n17824, ys__n17825,
    ys__n17827, ys__n17828, ys__n17830, ys__n17831, ys__n17833, ys__n17834,
    ys__n17836, ys__n17837, ys__n17839, ys__n17840, ys__n17842, ys__n17843,
    ys__n17845, ys__n17846, ys__n17848, ys__n17849, ys__n17866, ys__n17867,
    ys__n17869, ys__n17870, ys__n17872, ys__n17873, ys__n17875, ys__n17876,
    ys__n17878, ys__n17879, ys__n17881, ys__n17882, ys__n17884, ys__n17885,
    ys__n17887, ys__n17888, ys__n17890, ys__n17891, ys__n17893, ys__n17894,
    ys__n17896, ys__n17897, ys__n17899, ys__n17900, ys__n17902, ys__n17903,
    ys__n17905, ys__n17906, ys__n17908, ys__n17909, ys__n17911, ys__n17912,
    ys__n17941, ys__n17943, ys__n18041, ys__n18043, ys__n18045, ys__n18047,
    ys__n18049, ys__n18051, ys__n18053, ys__n18055, ys__n18057, ys__n18059,
    ys__n18061, ys__n18063, ys__n18065, ys__n18067, ys__n18070, ys__n18071,
    ys__n18090, ys__n18101, ys__n18105, ys__n18106, ys__n18109, ys__n18111,
    ys__n18112, ys__n18114, ys__n18116, ys__n18118, ys__n18121, ys__n18122,
    ys__n18124, ys__n18143, ys__n18149, ys__n18150, ys__n18156, ys__n18173,
    ys__n18208, ys__n18226, ys__n18229, ys__n18231, ys__n18240, ys__n18242,
    ys__n18243, ys__n18270, ys__n18271, ys__n18277, ys__n18280, ys__n18283,
    ys__n18286, ys__n18317, ys__n18378, ys__n18381, ys__n18384, ys__n18389,
    ys__n18393, ys__n18448, ys__n18451, ys__n18454, ys__n18457, ys__n18460,
    ys__n18463, ys__n18466, ys__n18469, ys__n18472, ys__n18475, ys__n18478,
    ys__n18481, ys__n18484, ys__n18487, ys__n18490, ys__n18493, ys__n18496,
    ys__n18499, ys__n18502, ys__n18505, ys__n18508, ys__n18511, ys__n18514,
    ys__n18517, ys__n18520, ys__n18523, ys__n18526, ys__n18529, ys__n18532,
    ys__n18535, ys__n18538, ys__n18541, ys__n18544, ys__n18546, ys__n18556,
    ys__n18558, ys__n18560, ys__n18562, ys__n18565, ys__n18568, ys__n18569,
    ys__n18571, ys__n18572, ys__n18574, ys__n18575, ys__n18577, ys__n18578,
    ys__n18580, ys__n18581, ys__n18583, ys__n18584, ys__n18586, ys__n18587,
    ys__n18589, ys__n18590, ys__n18592, ys__n18593, ys__n18595, ys__n18596,
    ys__n18598, ys__n18599, ys__n18601, ys__n18602, ys__n18604, ys__n18605,
    ys__n18607, ys__n18608, ys__n18610, ys__n18611, ys__n18613, ys__n18614,
    ys__n18616, ys__n18617, ys__n18619, ys__n18620, ys__n18622, ys__n18623,
    ys__n18625, ys__n18626, ys__n18628, ys__n18630, ys__n18632, ys__n18634,
    ys__n18636, ys__n18638, ys__n18639, ys__n18641, ys__n18642, ys__n18644,
    ys__n18645, ys__n18647, ys__n18650, ys__n18651, ys__n18749, ys__n18752,
    ys__n18755, ys__n18758, ys__n18761, ys__n18762, ys__n18765, ys__n18767,
    ys__n18769, ys__n18771, ys__n18773, ys__n18775, ys__n18777, ys__n18779,
    ys__n18781, ys__n18783, ys__n18785, ys__n18787, ys__n18789, ys__n18791,
    ys__n18793, ys__n18795, ys__n18797, ys__n18799, ys__n18801, ys__n18803,
    ys__n18805, ys__n18807, ys__n18809, ys__n18811, ys__n18813, ys__n18815,
    ys__n18817, ys__n18819, ys__n18821, ys__n18823, ys__n18825, ys__n18827,
    ys__n18829, ys__n18831, ys__n18833, ys__n18835, ys__n18837, ys__n18839,
    ys__n18841, ys__n18843, ys__n18845, ys__n18847, ys__n18849, ys__n18851,
    ys__n18853, ys__n18855, ys__n18857, ys__n18859, ys__n18861, ys__n18863,
    ys__n18865, ys__n18867, ys__n18869, ys__n18871, ys__n18873, ys__n18875,
    ys__n18877, ys__n18879, ys__n18881, ys__n18883, ys__n18885, ys__n18887,
    ys__n18889, ys__n18891, ys__n18956, ys__n18957, ys__n18958, ys__n18959,
    ys__n18960, ys__n18961, ys__n18962, ys__n18963, ys__n18964, ys__n18965,
    ys__n18966, ys__n18967, ys__n18968, ys__n18969, ys__n18970, ys__n18971,
    ys__n18972, ys__n18973, ys__n18974, ys__n18975, ys__n18976, ys__n18977,
    ys__n18978, ys__n18979, ys__n18980, ys__n18981, ys__n18982, ys__n18983,
    ys__n18984, ys__n18985, ys__n18986, ys__n18987, ys__n18989, ys__n18991,
    ys__n18993, ys__n18995, ys__n18997, ys__n18999, ys__n19001, ys__n19003,
    ys__n19005, ys__n19007, ys__n19009, ys__n19011, ys__n19013, ys__n19015,
    ys__n19017, ys__n19019, ys__n19021, ys__n19023, ys__n19025, ys__n19027,
    ys__n19029, ys__n19031, ys__n19033, ys__n19035, ys__n19037, ys__n19039,
    ys__n19041, ys__n19043, ys__n19045, ys__n19047, ys__n19049, ys__n19051,
    ys__n19116, ys__n19117, ys__n19118, ys__n19119, ys__n19120, ys__n19121,
    ys__n19122, ys__n19123, ys__n19124, ys__n19125, ys__n19126, ys__n19127,
    ys__n19128, ys__n19129, ys__n19130, ys__n19131, ys__n19132, ys__n19133,
    ys__n19134, ys__n19135, ys__n19136, ys__n19137, ys__n19138, ys__n19139,
    ys__n19140, ys__n19141, ys__n19142, ys__n19143, ys__n19144, ys__n19145,
    ys__n19146, ys__n19147, ys__n19156, ys__n19157, ys__n19166, ys__n19171,
    ys__n19203, ys__n19215, ys__n19245, ys__n19251, ys__n19253, ys__n19259,
    ys__n19261, ys__n19263, ys__n19843, ys__n19844, ys__n19845, ys__n19846,
    ys__n19847, ys__n19848, ys__n19849, ys__n19850, ys__n19851, ys__n19852,
    ys__n19853, ys__n19854, ys__n19855, ys__n19856, ys__n19857, ys__n19858,
    ys__n19859, ys__n19860, ys__n19861, ys__n19862, ys__n19863, ys__n19864,
    ys__n19865, ys__n19866, ys__n19867, ys__n19868, ys__n19869, ys__n19870,
    ys__n19871, ys__n19872, ys__n19873, ys__n19874, ys__n19875, ys__n19972,
    ys__n19973, ys__n19974, ys__n19975, ys__n19976, ys__n19977, ys__n19978,
    ys__n19979, ys__n19980, ys__n19981, ys__n19982, ys__n19983, ys__n19984,
    ys__n19985, ys__n19986, ys__n19987, ys__n19988, ys__n19989, ys__n19990,
    ys__n19991, ys__n19992, ys__n19993, ys__n19994, ys__n19995, ys__n19996,
    ys__n19997, ys__n19998, ys__n19999, ys__n20000, ys__n20001, ys__n20002,
    ys__n20003, ys__n20004, ys__n20035, ys__n20058, ys__n20061, ys__n20064,
    ys__n20067, ys__n20070, ys__n20073, ys__n20076, ys__n20079, ys__n20138,
    ys__n20140, ys__n20142, ys__n20144, ys__n20146, ys__n20148, ys__n20150,
    ys__n20152, ys__n20186, ys__n20188, ys__n20190, ys__n20192, ys__n20194,
    ys__n20196, ys__n20198, ys__n20200, ys__n20202, ys__n20204, ys__n20206,
    ys__n20208, ys__n20210, ys__n20212, ys__n20214, ys__n20216, ys__n20273,
    ys__n20279, ys__n20280, ys__n20540, ys__n20542, ys__n20544, ys__n20546,
    ys__n20548, ys__n20550, ys__n20552, ys__n20554, ys__n20556, ys__n20558,
    ys__n20560, ys__n20562, ys__n20564, ys__n20566, ys__n20568, ys__n20570,
    ys__n20572, ys__n20574, ys__n20576, ys__n20578, ys__n20580, ys__n20582,
    ys__n20584, ys__n20586, ys__n20588, ys__n20590, ys__n20592, ys__n20594,
    ys__n20596, ys__n20598, ys__n20600, ys__n20602, ys__n20604, ys__n20606,
    ys__n20608, ys__n20610, ys__n20612, ys__n20614, ys__n20616, ys__n20618,
    ys__n20620, ys__n20622, ys__n20624, ys__n20626, ys__n20628, ys__n20630,
    ys__n20632, ys__n20634, ys__n20636, ys__n20638, ys__n20640, ys__n20642,
    ys__n20644, ys__n20646, ys__n20648, ys__n20650, ys__n20652, ys__n20654,
    ys__n20656, ys__n20658, ys__n20660, ys__n20662, ys__n20664, ys__n20666,
    ys__n20668, ys__n20670, ys__n20672, ys__n20674, ys__n20676, ys__n20678,
    ys__n20680, ys__n20682, ys__n20684, ys__n20686, ys__n20688, ys__n20690,
    ys__n20692, ys__n20694, ys__n20696, ys__n20698, ys__n20700, ys__n20702,
    ys__n20704, ys__n20706, ys__n20708, ys__n20710, ys__n20712, ys__n20714,
    ys__n20716, ys__n20718, ys__n20720, ys__n20722, ys__n20724, ys__n20726,
    ys__n20728, ys__n20730, ys__n20732, ys__n20734, ys__n20736, ys__n20738,
    ys__n20740, ys__n20742, ys__n20744, ys__n20746, ys__n20748, ys__n20750,
    ys__n20752, ys__n20754, ys__n20756, ys__n20758, ys__n20760, ys__n20762,
    ys__n20764, ys__n20766, ys__n20768, ys__n20770, ys__n20772, ys__n20774,
    ys__n20776, ys__n20778, ys__n20780, ys__n20782, ys__n20784, ys__n20786,
    ys__n20788, ys__n20790, ys__n20792, ys__n20794, ys__n20796, ys__n20798,
    ys__n20800, ys__n20802, ys__n20804, ys__n20806, ys__n20808, ys__n20810,
    ys__n20812, ys__n20814, ys__n20816, ys__n20818, ys__n20820, ys__n20822,
    ys__n20824, ys__n20826, ys__n20828, ys__n20830, ys__n20832, ys__n20834,
    ys__n20836, ys__n20838, ys__n20840, ys__n20842, ys__n20844, ys__n20846,
    ys__n20848, ys__n20850, ys__n20852, ys__n20854, ys__n20856, ys__n20858,
    ys__n20860, ys__n20862, ys__n20864, ys__n20866, ys__n20868, ys__n20870,
    ys__n20872, ys__n20874, ys__n20876, ys__n20878, ys__n20880, ys__n20882,
    ys__n20884, ys__n20886, ys__n20888, ys__n20890, ys__n20892, ys__n20894,
    ys__n20896, ys__n20898, ys__n20900, ys__n20902, ys__n20904, ys__n20906,
    ys__n20908, ys__n20910, ys__n20912, ys__n20914, ys__n20916, ys__n20918,
    ys__n20920, ys__n20922, ys__n20924, ys__n20925, ys__n20926, ys__n20927,
    ys__n20928, ys__n20929, ys__n20930, ys__n20931, ys__n20932, ys__n20933,
    ys__n20934, ys__n20935, ys__n20936, ys__n20937, ys__n20938, ys__n20939,
    ys__n20940, ys__n20941, ys__n20942, ys__n20943, ys__n20944, ys__n20945,
    ys__n20946, ys__n20947, ys__n20948, ys__n20949, ys__n20950, ys__n20951,
    ys__n20952, ys__n20953, ys__n20954, ys__n20955, ys__n20956, ys__n20958,
    ys__n20960, ys__n20962, ys__n20964, ys__n20966, ys__n20968, ys__n20970,
    ys__n20972, ys__n20974, ys__n20976, ys__n20978, ys__n20980, ys__n20982,
    ys__n20984, ys__n20986, ys__n20988, ys__n20990, ys__n20992, ys__n20994,
    ys__n20996, ys__n20998, ys__n21000, ys__n21002, ys__n21004, ys__n21006,
    ys__n21008, ys__n21010, ys__n21012, ys__n21014, ys__n21016, ys__n21018,
    ys__n21020, ys__n21022, ys__n21024, ys__n21026, ys__n21028, ys__n21030,
    ys__n21032, ys__n21034, ys__n21036, ys__n21038, ys__n21040, ys__n21042,
    ys__n21044, ys__n21046, ys__n21048, ys__n21050, ys__n21052, ys__n21054,
    ys__n21056, ys__n21058, ys__n21060, ys__n21062, ys__n21064, ys__n21066,
    ys__n21068, ys__n21070, ys__n21072, ys__n21074, ys__n21076, ys__n21078,
    ys__n21080, ys__n21082, ys__n21084, ys__n21086, ys__n21088, ys__n21090,
    ys__n21092, ys__n21094, ys__n21096, ys__n21098, ys__n21100, ys__n21102,
    ys__n21104, ys__n21106, ys__n21108, ys__n21110, ys__n21112, ys__n21114,
    ys__n21116, ys__n21118, ys__n21120, ys__n21122, ys__n21124, ys__n21126,
    ys__n21128, ys__n21130, ys__n21132, ys__n21134, ys__n21136, ys__n21138,
    ys__n21140, ys__n21142, ys__n21144, ys__n21146, ys__n21148, ys__n21150,
    ys__n21152, ys__n21154, ys__n21156, ys__n21158, ys__n21160, ys__n21162,
    ys__n21164, ys__n21166, ys__n21168, ys__n21170, ys__n21172, ys__n21174,
    ys__n21176, ys__n21178, ys__n21180, ys__n21182, ys__n21184, ys__n21186,
    ys__n21188, ys__n21190, ys__n21192, ys__n21194, ys__n21196, ys__n21198,
    ys__n21200, ys__n21202, ys__n21204, ys__n21206, ys__n21208, ys__n21210,
    ys__n21212, ys__n21214, ys__n21216, ys__n21218, ys__n21220, ys__n21222,
    ys__n21224, ys__n21226, ys__n21228, ys__n21230, ys__n21232, ys__n21234,
    ys__n21236, ys__n21238, ys__n21240, ys__n21242, ys__n21244, ys__n21246,
    ys__n21248, ys__n21250, ys__n21252, ys__n21254, ys__n21256, ys__n21258,
    ys__n21260, ys__n21262, ys__n21264, ys__n21266, ys__n21268, ys__n21270,
    ys__n21272, ys__n21274, ys__n21276, ys__n21278, ys__n21280, ys__n21282,
    ys__n21284, ys__n21286, ys__n21288, ys__n21290, ys__n21292, ys__n21294,
    ys__n21296, ys__n21298, ys__n21300, ys__n21302, ys__n21304, ys__n21306,
    ys__n21308, ys__n21310, ys__n21312, ys__n21314, ys__n21316, ys__n21318,
    ys__n21320, ys__n21322, ys__n21324, ys__n21326, ys__n21328, ys__n21330,
    ys__n21332, ys__n21334, ys__n21336, ys__n21338, ys__n21340, ys__n21342,
    ys__n21344, ys__n21346, ys__n21348, ys__n21350, ys__n21352, ys__n21354,
    ys__n21356, ys__n21358, ys__n21360, ys__n21362, ys__n21364, ys__n21366,
    ys__n21368, ys__n21370, ys__n21372, ys__n21374, ys__n21376, ys__n21378,
    ys__n21380, ys__n21382, ys__n21384, ys__n21386, ys__n21388, ys__n21390,
    ys__n21392, ys__n21394, ys__n21396, ys__n21398, ys__n21400, ys__n21402,
    ys__n21404, ys__n21405, ys__n21406, ys__n21407, ys__n21408, ys__n21409,
    ys__n21410, ys__n21411, ys__n21412, ys__n21413, ys__n21414, ys__n21415,
    ys__n21416, ys__n21417, ys__n21418, ys__n21419, ys__n21420, ys__n21421,
    ys__n21422, ys__n21423, ys__n21424, ys__n21425, ys__n21426, ys__n21427,
    ys__n21428, ys__n21429, ys__n21430, ys__n21431, ys__n21432, ys__n21433,
    ys__n21434, ys__n21435, ys__n21500, ys__n21502, ys__n21504, ys__n21506,
    ys__n21508, ys__n21510, ys__n21512, ys__n21514, ys__n21516, ys__n21518,
    ys__n21520, ys__n21522, ys__n21524, ys__n21526, ys__n21528, ys__n21530,
    ys__n21532, ys__n21534, ys__n21536, ys__n21538, ys__n21540, ys__n21542,
    ys__n21544, ys__n21546, ys__n21548, ys__n21550, ys__n21552, ys__n21554,
    ys__n21556, ys__n21558, ys__n21560, ys__n21562, ys__n21564, ys__n21566,
    ys__n21568, ys__n21570, ys__n21572, ys__n21574, ys__n21576, ys__n21578,
    ys__n21580, ys__n21582, ys__n21584, ys__n21586, ys__n21588, ys__n21590,
    ys__n21592, ys__n21594, ys__n21596, ys__n21598, ys__n21600, ys__n21602,
    ys__n21604, ys__n21606, ys__n21608, ys__n21610, ys__n21612, ys__n21614,
    ys__n21616, ys__n21618, ys__n21620, ys__n21622, ys__n21624, ys__n21626,
    ys__n21628, ys__n21630, ys__n21632, ys__n21634, ys__n21636, ys__n21638,
    ys__n21640, ys__n21642, ys__n21644, ys__n21646, ys__n21648, ys__n21650,
    ys__n21652, ys__n21654, ys__n21656, ys__n21658, ys__n21660, ys__n21662,
    ys__n21664, ys__n21666, ys__n21668, ys__n21670, ys__n21672, ys__n21674,
    ys__n21676, ys__n21678, ys__n21680, ys__n21682, ys__n21684, ys__n21686,
    ys__n21688, ys__n21690, ys__n21692, ys__n21694, ys__n21696, ys__n21698,
    ys__n21700, ys__n21702, ys__n21704, ys__n21706, ys__n21708, ys__n21710,
    ys__n21712, ys__n21714, ys__n21716, ys__n21718, ys__n21720, ys__n21722,
    ys__n21724, ys__n21726, ys__n21728, ys__n21730, ys__n21732, ys__n21734,
    ys__n21736, ys__n21738, ys__n21740, ys__n21742, ys__n21744, ys__n21746,
    ys__n21748, ys__n21750, ys__n21752, ys__n21754, ys__n21756, ys__n21758,
    ys__n21760, ys__n21762, ys__n21764, ys__n21766, ys__n21768, ys__n21770,
    ys__n21772, ys__n21774, ys__n21776, ys__n21778, ys__n21780, ys__n21782,
    ys__n21784, ys__n21786, ys__n21788, ys__n21790, ys__n21792, ys__n21794,
    ys__n21796, ys__n21798, ys__n21800, ys__n21802, ys__n21804, ys__n21806,
    ys__n21808, ys__n21810, ys__n21812, ys__n21814, ys__n21816, ys__n21818,
    ys__n21820, ys__n21822, ys__n21824, ys__n21826, ys__n21828, ys__n21830,
    ys__n21832, ys__n21834, ys__n21836, ys__n21838, ys__n21840, ys__n21842,
    ys__n21844, ys__n21846, ys__n21848, ys__n21850, ys__n21852, ys__n21854,
    ys__n21856, ys__n21858, ys__n21860, ys__n21862, ys__n21864, ys__n21866,
    ys__n21868, ys__n21870, ys__n21872, ys__n21874, ys__n21876, ys__n21878,
    ys__n21880, ys__n21882, ys__n21884, ys__n21886, ys__n21888, ys__n21890,
    ys__n21892, ys__n21894, ys__n21896, ys__n21898, ys__n21900, ys__n21902,
    ys__n21904, ys__n21906, ys__n21908, ys__n21910, ys__n21912, ys__n21914,
    ys__n21916, ys__n21918, ys__n21920, ys__n21922, ys__n21924, ys__n21926,
    ys__n21928, ys__n21930, ys__n21932, ys__n21934, ys__n21936, ys__n21938,
    ys__n21940, ys__n21942, ys__n21944, ys__n21946, ys__n21948, ys__n21949,
    ys__n21950, ys__n21951, ys__n21952, ys__n21953, ys__n21954, ys__n21955,
    ys__n21956, ys__n21957, ys__n21958, ys__n21959, ys__n21960, ys__n21961,
    ys__n21962, ys__n21963, ys__n21964, ys__n21965, ys__n21966, ys__n21967,
    ys__n21968, ys__n21969, ys__n21970, ys__n21971, ys__n21972, ys__n21973,
    ys__n21974, ys__n21975, ys__n21976, ys__n21977, ys__n21978, ys__n21979,
    ys__n21980, ys__n21982, ys__n21984, ys__n21986, ys__n21988, ys__n21990,
    ys__n21992, ys__n21994, ys__n21996, ys__n21998, ys__n22000, ys__n22002,
    ys__n22004, ys__n22006, ys__n22008, ys__n22010, ys__n22012, ys__n22014,
    ys__n22016, ys__n22018, ys__n22020, ys__n22022, ys__n22024, ys__n22026,
    ys__n22028, ys__n22030, ys__n22032, ys__n22034, ys__n22036, ys__n22038,
    ys__n22040, ys__n22042, ys__n22044, ys__n22046, ys__n22048, ys__n22050,
    ys__n22052, ys__n22054, ys__n22056, ys__n22058, ys__n22060, ys__n22062,
    ys__n22064, ys__n22066, ys__n22068, ys__n22070, ys__n22072, ys__n22074,
    ys__n22076, ys__n22078, ys__n22080, ys__n22082, ys__n22084, ys__n22086,
    ys__n22088, ys__n22090, ys__n22092, ys__n22094, ys__n22096, ys__n22098,
    ys__n22100, ys__n22102, ys__n22104, ys__n22106, ys__n22108, ys__n22110,
    ys__n22112, ys__n22114, ys__n22116, ys__n22118, ys__n22120, ys__n22122,
    ys__n22124, ys__n22126, ys__n22128, ys__n22130, ys__n22132, ys__n22134,
    ys__n22136, ys__n22138, ys__n22140, ys__n22142, ys__n22144, ys__n22146,
    ys__n22148, ys__n22150, ys__n22152, ys__n22154, ys__n22156, ys__n22158,
    ys__n22160, ys__n22162, ys__n22164, ys__n22166, ys__n22168, ys__n22170,
    ys__n22172, ys__n22174, ys__n22176, ys__n22178, ys__n22180, ys__n22182,
    ys__n22184, ys__n22186, ys__n22188, ys__n22190, ys__n22192, ys__n22194,
    ys__n22196, ys__n22198, ys__n22200, ys__n22202, ys__n22204, ys__n22206,
    ys__n22208, ys__n22210, ys__n22212, ys__n22214, ys__n22216, ys__n22218,
    ys__n22220, ys__n22222, ys__n22224, ys__n22226, ys__n22228, ys__n22230,
    ys__n22232, ys__n22234, ys__n22236, ys__n22238, ys__n22240, ys__n22242,
    ys__n22244, ys__n22246, ys__n22248, ys__n22250, ys__n22252, ys__n22254,
    ys__n22256, ys__n22258, ys__n22260, ys__n22262, ys__n22264, ys__n22266,
    ys__n22268, ys__n22270, ys__n22272, ys__n22274, ys__n22276, ys__n22278,
    ys__n22280, ys__n22282, ys__n22284, ys__n22286, ys__n22288, ys__n22290,
    ys__n22292, ys__n22294, ys__n22296, ys__n22298, ys__n22300, ys__n22302,
    ys__n22304, ys__n22306, ys__n22308, ys__n22310, ys__n22312, ys__n22314,
    ys__n22316, ys__n22318, ys__n22320, ys__n22322, ys__n22324, ys__n22326,
    ys__n22328, ys__n22330, ys__n22332, ys__n22334, ys__n22336, ys__n22338,
    ys__n22340, ys__n22342, ys__n22344, ys__n22346, ys__n22348, ys__n22350,
    ys__n22352, ys__n22354, ys__n22356, ys__n22358, ys__n22360, ys__n22362,
    ys__n22364, ys__n22366, ys__n22368, ys__n22370, ys__n22372, ys__n22374,
    ys__n22376, ys__n22378, ys__n22380, ys__n22382, ys__n22384, ys__n22386,
    ys__n22388, ys__n22390, ys__n22392, ys__n22394, ys__n22396, ys__n22398,
    ys__n22400, ys__n22402, ys__n22404, ys__n22406, ys__n22408, ys__n22410,
    ys__n22412, ys__n22414, ys__n22416, ys__n22418, ys__n22420, ys__n22422,
    ys__n22424, ys__n22426, ys__n22428, ys__n22429, ys__n22430, ys__n22431,
    ys__n22432, ys__n22433, ys__n22434, ys__n22435, ys__n22436, ys__n22437,
    ys__n22438, ys__n22439, ys__n22440, ys__n22441, ys__n22442, ys__n22443,
    ys__n22444, ys__n22445, ys__n22446, ys__n22447, ys__n22448, ys__n22449,
    ys__n22450, ys__n22451, ys__n22452, ys__n22453, ys__n22454, ys__n22455,
    ys__n22456, ys__n22457, ys__n22458, ys__n22459, ys__n22464, ys__n22465,
    ys__n22564, ys__n22566, ys__n22568, ys__n22570, ys__n22572, ys__n22574,
    ys__n22576, ys__n22578, ys__n22580, ys__n22582, ys__n22584, ys__n22586,
    ys__n22588, ys__n22590, ys__n22592, ys__n22594, ys__n22596, ys__n22598,
    ys__n22600, ys__n22602, ys__n22604, ys__n22606, ys__n22608, ys__n22610,
    ys__n22612, ys__n22614, ys__n22616, ys__n22618, ys__n22620, ys__n22622,
    ys__n22624, ys__n22626, ys__n22630, ys__n22632, ys__n22634, ys__n22636,
    ys__n22640, ys__n22642, ys__n22644, ys__n22646, ys__n22648, ys__n22650,
    ys__n22652, ys__n22654, ys__n22668, ys__n22670, ys__n22673, ys__n22675,
    ys__n22677, ys__n22679, ys__n22681, ys__n22683, ys__n22685, ys__n22687,
    ys__n22689, ys__n22715, ys__n22717, ys__n22719, ys__n22721, ys__n22723,
    ys__n22725, ys__n22727, ys__n22729, ys__n22731, ys__n22733, ys__n22735,
    ys__n22737, ys__n22739, ys__n22741, ys__n22743, ys__n22745, ys__n22747,
    ys__n22749, ys__n22751, ys__n22753, ys__n22755, ys__n22757, ys__n22759,
    ys__n22761, ys__n22763, ys__n22765, ys__n22767, ys__n22769, ys__n22771,
    ys__n22773, ys__n22775, ys__n22777, ys__n22779, ys__n22781, ys__n22783,
    ys__n22785, ys__n22787, ys__n22789, ys__n22792, ys__n22794, ys__n22799,
    ys__n22818, ys__n22820, ys__n22822, ys__n22824, ys__n22826, ys__n22828,
    ys__n22830, ys__n22832, ys__n22834, ys__n22836, ys__n22838, ys__n22840,
    ys__n22842, ys__n22844, ys__n22846, ys__n22848, ys__n22850, ys__n22852,
    ys__n22854, ys__n22856, ys__n22858, ys__n22860, ys__n22862, ys__n22864,
    ys__n22866, ys__n22868, ys__n22870, ys__n22872, ys__n22874, ys__n22876,
    ys__n22878, ys__n22880, ys__n22882, ys__n22884, ys__n22885, ys__n22886,
    ys__n22887, ys__n22888, ys__n22889, ys__n22890, ys__n22891, ys__n22892,
    ys__n22893, ys__n22894, ys__n22895, ys__n22896, ys__n22897, ys__n22898,
    ys__n22899, ys__n22900, ys__n22901, ys__n22902, ys__n22903, ys__n22904,
    ys__n22905, ys__n22906, ys__n22907, ys__n22908, ys__n22909, ys__n22910,
    ys__n22911, ys__n22912, ys__n22913, ys__n22914, ys__n22915, ys__n22916,
    ys__n22918, ys__n22921, ys__n22924, ys__n22927, ys__n22930, ys__n22933,
    ys__n22936, ys__n22939, ys__n22942, ys__n22945, ys__n22948, ys__n22951,
    ys__n22954, ys__n22957, ys__n22960, ys__n22963, ys__n22966, ys__n22969,
    ys__n22972, ys__n22975, ys__n22978, ys__n22981, ys__n22984, ys__n22987,
    ys__n22990, ys__n22993, ys__n22996, ys__n22999, ys__n23002, ys__n23005,
    ys__n23008, ys__n23011, ys__n23014, ys__n23016, ys__n23018, ys__n23020,
    ys__n23022, ys__n23024, ys__n23026, ys__n23028, ys__n23030, ys__n23032,
    ys__n23034, ys__n23036, ys__n23038, ys__n23040, ys__n23042, ys__n23044,
    ys__n23046, ys__n23048, ys__n23050, ys__n23052, ys__n23054, ys__n23056,
    ys__n23058, ys__n23060, ys__n23062, ys__n23064, ys__n23066, ys__n23068,
    ys__n23070, ys__n23072, ys__n23074, ys__n23076, ys__n23077, ys__n23078,
    ys__n23079, ys__n23080, ys__n23081, ys__n23082, ys__n23083, ys__n23084,
    ys__n23085, ys__n23086, ys__n23087, ys__n23088, ys__n23089, ys__n23090,
    ys__n23091, ys__n23092, ys__n23093, ys__n23094, ys__n23095, ys__n23096,
    ys__n23097, ys__n23098, ys__n23099, ys__n23100, ys__n23101, ys__n23102,
    ys__n23103, ys__n23104, ys__n23105, ys__n23106, ys__n23107, ys__n23108,
    ys__n23111, ys__n23114, ys__n23117, ys__n23120, ys__n23123, ys__n23126,
    ys__n23129, ys__n23132, ys__n23135, ys__n23138, ys__n23141, ys__n23144,
    ys__n23147, ys__n23150, ys__n23153, ys__n23156, ys__n23159, ys__n23162,
    ys__n23165, ys__n23168, ys__n23171, ys__n23174, ys__n23177, ys__n23180,
    ys__n23183, ys__n23186, ys__n23189, ys__n23192, ys__n23195, ys__n23198,
    ys__n23203, ys__n23205, ys__n23207, ys__n23209, ys__n23211, ys__n23213,
    ys__n23215, ys__n23217, ys__n23219, ys__n23221, ys__n23223, ys__n23225,
    ys__n23227, ys__n23229, ys__n23231, ys__n23233, ys__n23235, ys__n23237,
    ys__n23239, ys__n23241, ys__n23243, ys__n23245, ys__n23247, ys__n23249,
    ys__n23251, ys__n23253, ys__n23255, ys__n23257, ys__n23259, ys__n23261,
    ys__n23269, ys__n23271, ys__n23272, ys__n23274, ys__n23276, ys__n23278,
    ys__n23280, ys__n23282, ys__n23284, ys__n23286, ys__n23288, ys__n23290,
    ys__n23292, ys__n23294, ys__n23296, ys__n23298, ys__n23300, ys__n23302,
    ys__n23304, ys__n23306, ys__n23308, ys__n23310, ys__n23312, ys__n23314,
    ys__n23316, ys__n23318, ys__n23320, ys__n23322, ys__n23324, ys__n23326,
    ys__n23328, ys__n23330, ys__n23332, ys__n23335, ys__n23339, ys__n23480,
    ys__n23548, ys__n23550, ys__n23552, ys__n23554, ys__n23556, ys__n23558,
    ys__n23560, ys__n23562, ys__n23564, ys__n23566, ys__n23568, ys__n23570,
    ys__n23572, ys__n23574, ys__n23627, ys__n23629, ys__n23641, ys__n23644,
    ys__n23645, ys__n23647, ys__n23650, ys__n23652, ys__n23655, ys__n23658,
    ys__n23661, ys__n23663, ys__n23705, ys__n23706, ys__n23707, ys__n23708,
    ys__n23709, ys__n23710, ys__n23711, ys__n23712, ys__n23713, ys__n23714,
    ys__n23715, ys__n23717, ys__n23729, ys__n23730, ys__n23763, ys__n23818,
    ys__n23819, ys__n23820, ys__n23821, ys__n23822, ys__n23834, ys__n23836,
    ys__n23838, ys__n23840, ys__n23842, ys__n23850, ys__n23888, ys__n23889,
    ys__n23890, ys__n23891, ys__n23892, ys__n23904, ys__n23906, ys__n23908,
    ys__n23910, ys__n23912, ys__n23956, ys__n23957, ys__n23958, ys__n23959,
    ys__n23960, ys__n23977, ys__n23979, ys__n23981, ys__n23983, ys__n23985,
    ys__n24106, ys__n24107, ys__n24108, ys__n24112, ys__n24123, ys__n24124,
    ys__n24131, ys__n24143, ys__n24158, ys__n24167, ys__n24168, ys__n24177,
    ys__n24197, ys__n24199, ys__n24201, ys__n24203, ys__n24205, ys__n24207,
    ys__n24209, ys__n24211, ys__n24213, ys__n24215, ys__n24217, ys__n24219,
    ys__n24228, ys__n24233, ys__n24235, ys__n24243, ys__n24248, ys__n24279,
    ys__n24280, ys__n24303, ys__n24306, ys__n24308, ys__n24310, ys__n24312,
    ys__n24314, ys__n24316, ys__n24318, ys__n24337, ys__n24340, ys__n24342,
    ys__n24344, ys__n24346, ys__n24348, ys__n24350, ys__n24352, ys__n24371,
    ys__n24374, ys__n24376, ys__n24378, ys__n24380, ys__n24382, ys__n24384,
    ys__n24386, ys__n24389, ys__n24406, ys__n24409, ys__n24411, ys__n24413,
    ys__n24415, ys__n24417, ys__n24419, ys__n24421, ys__n24427, ys__n24433,
    ys__n24434, ys__n24461, ys__n24463, ys__n24464, ys__n24483, ys__n24485,
    ys__n24506, ys__n24519, ys__n24567, ys__n24575, ys__n24578, ys__n24590,
    ys__n24591, ys__n24615, ys__n24616, ys__n24617, ys__n24618, ys__n24619,
    ys__n24620, ys__n24621, ys__n24622, ys__n24623, ys__n24624, ys__n24625,
    ys__n24626, ys__n24627, ys__n24628, ys__n24629, ys__n24630, ys__n24631,
    ys__n24632, ys__n24633, ys__n24634, ys__n24635, ys__n24636, ys__n24637,
    ys__n24638, ys__n24639, ys__n24640, ys__n24641, ys__n24642, ys__n24643,
    ys__n24644, ys__n24645, ys__n24646, ys__n24647, ys__n24648, ys__n24649,
    ys__n24650, ys__n24651, ys__n24652, ys__n24653, ys__n24654, ys__n24655,
    ys__n24656, ys__n24657, ys__n24658, ys__n24659, ys__n24660, ys__n24661,
    ys__n24662, ys__n24663, ys__n24664, ys__n24665, ys__n24666, ys__n24667,
    ys__n24668, ys__n24669, ys__n24670, ys__n24671, ys__n24672, ys__n24673,
    ys__n24674, ys__n24675, ys__n24677, ys__n24679, ys__n24681, ys__n24683,
    ys__n24684, ys__n24685, ys__n24686, ys__n24687, ys__n24688, ys__n24689,
    ys__n24690, ys__n24691, ys__n24692, ys__n24693, ys__n24694, ys__n24695,
    ys__n24696, ys__n24697, ys__n24698, ys__n24699, ys__n24700, ys__n24701,
    ys__n24702, ys__n24703, ys__n24704, ys__n24705, ys__n24706, ys__n24707,
    ys__n24708, ys__n24709, ys__n24710, ys__n24711, ys__n24712, ys__n24741,
    ys__n24744, ys__n24747, ys__n24750, ys__n24753, ys__n24756, ys__n24759,
    ys__n24762, ys__n24765, ys__n24768, ys__n24771, ys__n24774, ys__n24777,
    ys__n24780, ys__n24783, ys__n24786, ys__n24789, ys__n24792, ys__n24795,
    ys__n24798, ys__n24801, ys__n24804, ys__n24807, ys__n24810, ys__n24813,
    ys__n24816, ys__n24819, ys__n24822, ys__n24825, ys__n24828, ys__n24831,
    ys__n24834, ys__n25292, ys__n25300, ys__n25381, ys__n25382, ys__n25383,
    ys__n25384, ys__n25470, ys__n25564, ys__n25567, ys__n25570, ys__n25573,
    ys__n25576, ys__n25579, ys__n25582, ys__n25585, ys__n25588, ys__n25591,
    ys__n25594, ys__n25597, ys__n25600, ys__n25603, ys__n25606, ys__n25609,
    ys__n25612, ys__n25615, ys__n25618, ys__n25621, ys__n25624, ys__n25627,
    ys__n25630, ys__n25633, ys__n25636, ys__n25639, ys__n25642, ys__n25645,
    ys__n25648, ys__n25651, ys__n25654, ys__n25657, ys__n25727, ys__n25730,
    ys__n25733, ys__n25736, ys__n25853, ys__n25856, ys__n25859, ys__n25862,
    ys__n25980, ys__n25984, ys__n25987, ys__n25990, ys__n25993, ys__n25996,
    ys__n25999, ys__n26002, ys__n26005, ys__n26008, ys__n26011, ys__n26014,
    ys__n26017, ys__n26020, ys__n26023, ys__n26026, ys__n26029, ys__n26032,
    ys__n26035, ys__n26038, ys__n26041, ys__n26044, ys__n26047, ys__n26050,
    ys__n26053, ys__n26056, ys__n26059, ys__n26062, ys__n26065, ys__n26068,
    ys__n26071, ys__n26074, ys__n26143, ys__n26145, ys__n26147, ys__n26149,
    ys__n26151, ys__n26153, ys__n26155, ys__n26157, ys__n26159, ys__n26161,
    ys__n26162, ys__n26164, ys__n26166, ys__n26168, ys__n26170, ys__n26172,
    ys__n26174, ys__n26176, ys__n26178, ys__n26180, ys__n26182, ys__n26184,
    ys__n26186, ys__n26188, ys__n26190, ys__n26192, ys__n26194, ys__n26196,
    ys__n26198, ys__n26200, ys__n26202, ys__n26204, ys__n26206, ys__n26208,
    ys__n26210, ys__n26212, ys__n26214, ys__n26216, ys__n26218, ys__n26279,
    ys__n26285, ys__n26359, ys__n26362, ys__n26425, ys__n26428, ys__n26431,
    ys__n26434, ys__n26437, ys__n26440, ys__n26443, ys__n26446, ys__n26449,
    ys__n26452, ys__n26455, ys__n26460, ys__n26463, ys__n26466, ys__n26469,
    ys__n26472, ys__n26475, ys__n26478, ys__n26481, ys__n26484, ys__n26487,
    ys__n26490, ys__n26493, ys__n26496, ys__n26499, ys__n26502, ys__n26505,
    ys__n26508, ys__n26511, ys__n26514, ys__n26517, ys__n26552, ys__n26553,
    ys__n26554, ys__n26556, ys__n26557, ys__n26558, ys__n26559, ys__n26560,
    ys__n26561, ys__n26562, ys__n26563, ys__n26564, ys__n26565, ys__n26567,
    ys__n26568, ys__n26569, ys__n26570, ys__n26571, ys__n26572, ys__n26766,
    ys__n26768, ys__n26770, ys__n26772, ys__n27479, ys__n27481, ys__n27485,
    ys__n27488, ys__n27496, ys__n27498, ys__n27499, ys__n27507, ys__n27509,
    ys__n27510, ys__n27518, ys__n27520, ys__n27607, ys__n27608, ys__n27611,
    ys__n27612, ys__n27614, ys__n27615, ys__n27617, ys__n27618, ys__n27620,
    ys__n27621, ys__n27623, ys__n27624, ys__n27626, ys__n27627, ys__n27629,
    ys__n27630, ys__n27632, ys__n27633, ys__n27635, ys__n27636, ys__n27638,
    ys__n27639, ys__n27641, ys__n27642, ys__n27644, ys__n27645, ys__n27647,
    ys__n27648, ys__n27650, ys__n27651, ys__n27653, ys__n27654, ys__n27656,
    ys__n27657, ys__n27659, ys__n27660, ys__n27662, ys__n27663, ys__n27665,
    ys__n27666, ys__n27668, ys__n27669, ys__n27671, ys__n27672, ys__n27674,
    ys__n27675, ys__n27677, ys__n27678, ys__n27680, ys__n27681, ys__n27683,
    ys__n27684, ys__n27686, ys__n27687, ys__n27689, ys__n27690, ys__n27692,
    ys__n27693, ys__n27695, ys__n27696, ys__n27698, ys__n27699, ys__n27701,
    ys__n27702, ys__n27737, ys__n27738, ys__n27740, ys__n27743, ys__n27747,
    ys__n27750, ys__n27753, ys__n27756, ys__n27759, ys__n27762, ys__n27765,
    ys__n27768, ys__n27771, ys__n27774, ys__n27777, ys__n27780, ys__n27783,
    ys__n27786, ys__n27789, ys__n27792, ys__n27795, ys__n27798, ys__n27801,
    ys__n27804, ys__n27807, ys__n27810, ys__n27813, ys__n27816, ys__n27819,
    ys__n27822, ys__n27825, ys__n27828, ys__n27831, ys__n27834, ys__n27837,
    ys__n27855, ys__n27857, ys__n27859, ys__n27861, ys__n27863, ys__n27865,
    ys__n27867, ys__n27869, ys__n27871, ys__n27873, ys__n27875, ys__n27877,
    ys__n27879, ys__n27881, ys__n27883, ys__n27885, ys__n28015, ys__n28016,
    ys__n28017, ys__n28018, ys__n28019, ys__n28020, ys__n28021, ys__n28022,
    ys__n28023, ys__n28024, ys__n28025, ys__n28026, ys__n28027, ys__n28028,
    ys__n28029, ys__n28030, ys__n28243, ys__n28287, ys__n28288, ys__n28290,
    ys__n28292, ys__n28294, ys__n28296, ys__n28424, ys__n28426, ys__n28428,
    ys__n28430, ys__n28432, ys__n28434, ys__n28436, ys__n28438, ys__n28446,
    ys__n28453, ys__n28455, ys__n28457, ys__n28459, ys__n28462, ys__n28464,
    ys__n28466, ys__n28468, ys__n28470, ys__n28472, ys__n28632, ys__n28633,
    ys__n28634, ys__n28635, ys__n28636, ys__n28637, ys__n28638, ys__n28639,
    ys__n28640, ys__n28641, ys__n28718, ys__n28719, ys__n28720, ys__n28859,
    ys__n28863, ys__n28866, ys__n28869, ys__n28872, ys__n28875, ys__n28878,
    ys__n28881, ys__n28884, ys__n28887, ys__n28890, ys__n28893, ys__n28896,
    ys__n28899, ys__n28902, ys__n28905, ys__n28908, ys__n28911, ys__n28914,
    ys__n28917, ys__n28920, ys__n28923, ys__n28926, ys__n28929, ys__n28932,
    ys__n28935, ys__n28938, ys__n28941, ys__n28944, ys__n28947, ys__n28950,
    ys__n28953, ys__n29117, ys__n29119, ys__n29120, ys__n29121, ys__n29123,
    ys__n29124, ys__n29126, ys__n29127, ys__n29129, ys__n29130, ys__n29132,
    ys__n29133, ys__n29135, ys__n29136, ys__n29138, ys__n29139, ys__n29141,
    ys__n29142, ys__n29144, ys__n29145, ys__n29147, ys__n29148, ys__n29150,
    ys__n29151, ys__n29153, ys__n29154, ys__n29156, ys__n29157, ys__n29159,
    ys__n29160, ys__n29162, ys__n29163, ys__n29165, ys__n29166, ys__n29168,
    ys__n29169, ys__n29171, ys__n29172, ys__n29174, ys__n29175, ys__n29177,
    ys__n29178, ys__n29180, ys__n29181, ys__n29183, ys__n29184, ys__n29186,
    ys__n29187, ys__n29189, ys__n29190, ys__n29192, ys__n29193, ys__n29195,
    ys__n29196, ys__n29198, ys__n29199, ys__n29201, ys__n29202, ys__n29204,
    ys__n29205, ys__n29207, ys__n29208, ys__n29210, ys__n29211, ys__n29213,
    ys__n29214, ys__n29218, ys__n29220, ys__n29224, ys__n29237, ys__n29240,
    ys__n29242, ys__n29244, ys__n29246, ys__n29248, ys__n29250, ys__n29252,
    ys__n29254, ys__n29256, ys__n29258, ys__n29260, ys__n29262, ys__n29264,
    ys__n29266, ys__n29268, ys__n29270, ys__n29272, ys__n29274, ys__n29276,
    ys__n29278, ys__n29280, ys__n29282, ys__n29284, ys__n29286, ys__n29288,
    ys__n29290, ys__n29292, ys__n29294, ys__n29296, ys__n29298, ys__n29300,
    ys__n29432, ys__n29433, ys__n29434, ys__n29436, ys__n29437, ys__n29439,
    ys__n29440, ys__n29442, ys__n29443, ys__n29445, ys__n29446, ys__n29448,
    ys__n29449, ys__n29451, ys__n29452, ys__n29454, ys__n29455, ys__n29457,
    ys__n29458, ys__n29460, ys__n29461, ys__n29463, ys__n29464, ys__n29466,
    ys__n29467, ys__n29469, ys__n29470, ys__n29472, ys__n29473, ys__n29475,
    ys__n29476, ys__n29478, ys__n29479, ys__n29481, ys__n29482, ys__n29484,
    ys__n29485, ys__n29487, ys__n29488, ys__n29490, ys__n29491, ys__n29493,
    ys__n29494, ys__n29496, ys__n29497, ys__n29499, ys__n29500, ys__n29502,
    ys__n29503, ys__n29505, ys__n29506, ys__n29508, ys__n29509, ys__n29511,
    ys__n29512, ys__n29514, ys__n29515, ys__n29517, ys__n29518, ys__n29520,
    ys__n29521, ys__n29523, ys__n29524, ys__n29526, ys__n29527, ys__n29531,
    ys__n29533, ys__n29537, ys__n29550, ys__n29552, ys__n29553, ys__n29554,
    ys__n29555, ys__n29556, ys__n29557, ys__n29558, ys__n29559, ys__n29560,
    ys__n29561, ys__n29562, ys__n29563, ys__n29564, ys__n29565, ys__n29566,
    ys__n29567, ys__n29568, ys__n29569, ys__n29570, ys__n29571, ys__n29572,
    ys__n29573, ys__n29574, ys__n29575, ys__n29576, ys__n29577, ys__n29578,
    ys__n29579, ys__n29580, ys__n29581, ys__n29582, ys__n29583, ys__n29584,
    ys__n29585, ys__n29586, ys__n29587, ys__n29588, ys__n29589, ys__n29590,
    ys__n29591, ys__n29592, ys__n29593, ys__n29594, ys__n29595, ys__n29596,
    ys__n29597, ys__n29598, ys__n29599, ys__n29600, ys__n29601, ys__n29602,
    ys__n29603, ys__n29604, ys__n29605, ys__n29606, ys__n29607, ys__n29608,
    ys__n29707, ys__n29708, ys__n29709, ys__n29711, ys__n29712, ys__n29714,
    ys__n29715, ys__n29717, ys__n29718, ys__n29720, ys__n29721, ys__n29723,
    ys__n29724, ys__n29726, ys__n29727, ys__n29729, ys__n29730, ys__n29732,
    ys__n29733, ys__n29735, ys__n29736, ys__n29738, ys__n29739, ys__n29741,
    ys__n29742, ys__n29744, ys__n29745, ys__n29747, ys__n29748, ys__n29750,
    ys__n29751, ys__n29753, ys__n29754, ys__n29756, ys__n29757, ys__n29759,
    ys__n29760, ys__n29762, ys__n29763, ys__n29765, ys__n29766, ys__n29768,
    ys__n29769, ys__n29771, ys__n29772, ys__n29774, ys__n29775, ys__n29777,
    ys__n29778, ys__n29780, ys__n29781, ys__n29783, ys__n29784, ys__n29786,
    ys__n29787, ys__n29789, ys__n29790, ys__n29792, ys__n29793, ys__n29795,
    ys__n29796, ys__n29798, ys__n29799, ys__n29801, ys__n29802, ys__n29806,
    ys__n29808, ys__n29812, ys__n29846, ys__n29880, ys__n29881, ys__n29883,
    ys__n29884, ys__n29885, ys__n29886, ys__n29887, ys__n29888, ys__n29889,
    ys__n29890, ys__n29891, ys__n29892, ys__n29893, ys__n29894, ys__n29895,
    ys__n29896, ys__n29897, ys__n29898, ys__n29899, ys__n29900, ys__n29901,
    ys__n29902, ys__n29903, ys__n29904, ys__n29905, ys__n29906, ys__n29907,
    ys__n29908, ys__n29909, ys__n29910, ys__n29911, ys__n29912, ys__n29913,
    ys__n30011, ys__n30014, ys__n30016, ys__n30018, ys__n30020, ys__n30022,
    ys__n30024, ys__n30026, ys__n30028, ys__n30030, ys__n30032, ys__n30034,
    ys__n30036, ys__n30038, ys__n30040, ys__n30042, ys__n30044, ys__n30046,
    ys__n30048, ys__n30050, ys__n30052, ys__n30054, ys__n30056, ys__n30058,
    ys__n30060, ys__n30062, ys__n30064, ys__n30066, ys__n30068, ys__n30070,
    ys__n30072, ys__n30074, ys__n30214, ys__n30216, ys__n30217, ys__n30219,
    ys__n30220, ys__n30225, ys__n30230, ys__n30232, ys__n30333, ys__n30334,
    ys__n30553, ys__n30815, ys__n30816, ys__n30818, ys__n30819, ys__n30820,
    ys__n30837, ys__n30861, ys__n30862, ys__n30863, ys__n30865, ys__n30867,
    ys__n30869, ys__n30871, ys__n30877, ys__n30879, ys__n30881, ys__n30883,
    ys__n30885, ys__n30887, ys__n30889, ys__n30891, ys__n30893, ys__n30895,
    ys__n30897, ys__n30899, ys__n30901, ys__n30903, ys__n30905, ys__n30907,
    ys__n30909, ys__n30911, ys__n30913, ys__n30915, ys__n30917, ys__n30919,
    ys__n30921, ys__n30923, ys__n30925, ys__n30927, ys__n30929, ys__n30931,
    ys__n30933, ys__n30935, ys__n30937, ys__n30939, ys__n30941, ys__n30957,
    ys__n30960, ys__n30961, ys__n30962, ys__n30974, ys__n31031, ys__n33212,
    ys__n33214, ys__n33216, ys__n33218, ys__n33220, ys__n33222, ys__n33259,
    ys__n33261, ys__n33263, ys__n33265, ys__n33267, ys__n33269, ys__n33272,
    ys__n33274, ys__n33276, ys__n33278, ys__n33300, ys__n33309, ys__n33311,
    ys__n33313, ys__n33318, ys__n33320, ys__n33328, ys__n33330, ys__n33332,
    ys__n33334, ys__n33336, ys__n33338, ys__n33340, ys__n33342, ys__n33350,
    ys__n33352, ys__n33359, ys__n33364, ys__n33370, ys__n33375, ys__n33380,
    ys__n33384, ys__n33386, ys__n33389, ys__n33394, ys__n33396, ys__n33398,
    ys__n33403, ys__n33407, ys__n33409, ys__n33411, ys__n33423, ys__n33431,
    ys__n33442, ys__n33451, ys__n33464, ys__n33469, ys__n33471, ys__n33473,
    ys__n33475, ys__n33479, ys__n33481, ys__n33488, ys__n33491, ys__n33493,
    ys__n33495, ys__n33497, ys__n33499, ys__n33509, ys__n33511, ys__n33522,
    ys__n33532, ys__n33541, ys__n33545, ys__n33548, ys__n33552, ys__n33558,
    ys__n33563, ys__n33564, ys__n33566, ys__n33568, ys__n33570, ys__n33572,
    ys__n33574, ys__n33576, ys__n33579, ys__n33581, ys__n33614, ys__n33632,
    ys__n33634, ys__n33636, ys__n33638, ys__n33640, ys__n33642, ys__n33644,
    ys__n33646, ys__n33648, ys__n33650, ys__n33652, ys__n33654, ys__n33656,
    ys__n33658, ys__n33660, ys__n33662, ys__n33664, ys__n33666, ys__n33668,
    ys__n33670, ys__n33672, ys__n33674, ys__n33676, ys__n33678, ys__n33681,
    ys__n33683, ys__n33685, ys__n33687, ys__n33689, ys__n33691, ys__n33693,
    ys__n33695, ys__n33697, ys__n33699, ys__n33701, ys__n33703, ys__n33705,
    ys__n33707, ys__n33709, ys__n33711, ys__n33713, ys__n33715, ys__n33717,
    ys__n33719, ys__n33721, ys__n33723, ys__n33725, ys__n33727, ys__n33729,
    ys__n33731, ys__n33733, ys__n33735, ys__n33737, ys__n33739, ys__n33741,
    ys__n33743, ys__n33745, ys__n33747, ys__n33749, ys__n34666, ys__n34668,
    ys__n34670, ys__n34672, ys__n34674, ys__n34676, ys__n34678, ys__n34680,
    ys__n34682, ys__n34684, ys__n34686, ys__n34688, ys__n34690, ys__n34692,
    ys__n34694, ys__n34696, ys__n34698, ys__n34700, ys__n34702, ys__n34704,
    ys__n34706, ys__n34708, ys__n34710, ys__n34712, ys__n34714, ys__n34716,
    ys__n34718, ys__n34720, ys__n34722, ys__n34724, ys__n34726, ys__n34728,
    ys__n34730, ys__n34732, ys__n34734, ys__n34736, ys__n34738, ys__n34740,
    ys__n34742, ys__n34744, ys__n34746, ys__n34748, ys__n34750, ys__n34752,
    ys__n34754, ys__n34756, ys__n34758, ys__n34760, ys__n34762, ys__n34764,
    ys__n34766, ys__n34768, ys__n34770, ys__n34772, ys__n34774, ys__n34776,
    ys__n34778, ys__n34780, ys__n34782, ys__n34784, ys__n34786, ys__n34788,
    ys__n34790, ys__n34792, ys__n34794, ys__n34796, ys__n34798, ys__n34800,
    ys__n34802, ys__n34804, ys__n34806, ys__n34808, ys__n34810, ys__n34812,
    ys__n34814, ys__n34816, ys__n34818, ys__n34820, ys__n34822, ys__n34824,
    ys__n34826, ys__n34828, ys__n34830, ys__n34832, ys__n34834, ys__n34836,
    ys__n34838, ys__n34840, ys__n34842, ys__n34844, ys__n34846, ys__n34848,
    ys__n34850, ys__n34852, ys__n34854, ys__n34856, ys__n34858, ys__n34860,
    ys__n34862, ys__n34864, ys__n34866, ys__n34868, ys__n34870, ys__n34872,
    ys__n34874, ys__n34876, ys__n34878, ys__n34880, ys__n34882, ys__n34884,
    ys__n34886, ys__n34888, ys__n34890, ys__n34892, ys__n34894, ys__n34896,
    ys__n34898, ys__n34900, ys__n34902, ys__n34904, ys__n34906, ys__n34908,
    ys__n34910, ys__n34912, ys__n34914, ys__n34916, ys__n34918, ys__n34920,
    ys__n34922, ys__n34924, ys__n34926, ys__n34928, ys__n34930, ys__n34932,
    ys__n34934, ys__n34936, ys__n34938, ys__n34940, ys__n34942, ys__n34944,
    ys__n34946, ys__n34948, ys__n34950, ys__n34959, ys__n34966, ys__n34972,
    ys__n34976, ys__n34978, ys__n34984, ys__n34988, ys__n34990, ys__n34996,
    ys__n35000, ys__n35002, ys__n35008, ys__n35012, ys__n35014, ys__n35020,
    ys__n35024, ys__n35026, ys__n35028, ys__n35031, ys__n35033, ys__n35035,
    ys__n35037, ys__n35039, ys__n35041, ys__n35047, ys__n35049, ys__n35057,
    ys__n35059, ys__n35065, ys__n35076, ys__n35078, ys__n35080, ys__n35082,
    ys__n35084, ys__n35086, ys__n35088, ys__n35090, ys__n35092, ys__n35094,
    ys__n35096, ys__n35098, ys__n35102, ys__n35104, ys__n35106, ys__n35108,
    ys__n35110, ys__n35112, ys__n35114, ys__n35116, ys__n35118, ys__n35120,
    ys__n35122, ys__n35124, ys__n35413, ys__n35415, ys__n35417, ys__n35419,
    ys__n35421, ys__n35423, ys__n35426, ys__n35704, ys__n35717, ys__n35719,
    ys__n35721, ys__n35723, ys__n35725, ys__n35727, ys__n37668, ys__n37669,
    ys__n37670, ys__n37671, ys__n37672, ys__n37673, ys__n37674, ys__n37675,
    ys__n37678, ys__n37679, ys__n37682, ys__n37692, ys__n37694, ys__n37696,
    ys__n37710, ys__n37712, ys__n37713, ys__n37743, ys__n37744, ys__n37745,
    ys__n37746, ys__n37747, ys__n37748, ys__n37749, ys__n37750, ys__n37751,
    ys__n37752, ys__n37753, ys__n37754, ys__n37755, ys__n37756, ys__n37757,
    ys__n37758, ys__n37759, ys__n37760, ys__n37761, ys__n37762, ys__n37763,
    ys__n37764, ys__n37765, ys__n37766, ys__n37767, ys__n37768, ys__n37769,
    ys__n37770, ys__n37771, ys__n37772, ys__n37773, ys__n37774, ys__n37775,
    ys__n37776, ys__n37777, ys__n37778, ys__n37779, ys__n37780, ys__n37781,
    ys__n37782, ys__n37783, ys__n37784, ys__n37785, ys__n37786, ys__n37787,
    ys__n37788, ys__n37789, ys__n37790, ys__n37791, ys__n37792, ys__n37793,
    ys__n37794, ys__n37795, ys__n37796, ys__n37797, ys__n37798, ys__n37799,
    ys__n37800, ys__n37801, ys__n37802, ys__n37803, ys__n37804, ys__n37805,
    ys__n37806, ys__n37807, ys__n37808, ys__n37809, ys__n37810, ys__n37811,
    ys__n37812, ys__n37813, ys__n37814, ys__n37815, ys__n37816, ys__n37817,
    ys__n37818, ys__n37819, ys__n37820, ys__n37821, ys__n37822, ys__n37823,
    ys__n37824, ys__n37825, ys__n37826, ys__n37827, ys__n37828, ys__n37829,
    ys__n37830, ys__n37831, ys__n37832, ys__n37833, ys__n37834, ys__n37835,
    ys__n37836, ys__n37837, ys__n37838, ys__n37839, ys__n37840, ys__n37841,
    ys__n37842, ys__n37843, ys__n37844, ys__n37845, ys__n37846, ys__n37847,
    ys__n37848, ys__n37849, ys__n37850, ys__n37851, ys__n37852, ys__n37853,
    ys__n37854, ys__n37855, ys__n37856, ys__n37857, ys__n37858, ys__n37859,
    ys__n37860, ys__n37861, ys__n37862, ys__n37863, ys__n37864, ys__n37865,
    ys__n37866, ys__n37867, ys__n37868, ys__n37869, ys__n37870, ys__n37871,
    ys__n37872, ys__n37873, ys__n37874, ys__n37875, ys__n37876, ys__n37877,
    ys__n37878, ys__n37879, ys__n37880, ys__n37881, ys__n37882, ys__n37883,
    ys__n37884, ys__n37885, ys__n37886, ys__n37887, ys__n37888, ys__n37889,
    ys__n37890, ys__n37891, ys__n37892, ys__n37893, ys__n37894, ys__n37895,
    ys__n37896, ys__n37897, ys__n37898, ys__n37899, ys__n37900, ys__n37901,
    ys__n37902, ys__n37903, ys__n37904, ys__n37905, ys__n37906, ys__n37907,
    ys__n37908, ys__n37909, ys__n37910, ys__n37911, ys__n37912, ys__n37913,
    ys__n37914, ys__n37915, ys__n37916, ys__n37917, ys__n37918, ys__n37919,
    ys__n37920, ys__n37921, ys__n37922, ys__n37923, ys__n37924, ys__n37925,
    ys__n37926, ys__n37927, ys__n37928, ys__n37929, ys__n37930, ys__n37931,
    ys__n37932, ys__n37933, ys__n37934, ys__n37935, ys__n37936, ys__n37937,
    ys__n37938, ys__n37939, ys__n37940, ys__n37941, ys__n37942, ys__n37943,
    ys__n37944, ys__n37945, ys__n37946, ys__n37947, ys__n37948, ys__n37949,
    ys__n37950, ys__n37951, ys__n37952, ys__n37953, ys__n37954, ys__n37955,
    ys__n37956, ys__n37957, ys__n37958, ys__n37959, ys__n37960, ys__n37961,
    ys__n37962, ys__n37963, ys__n37964, ys__n37965, ys__n37966, ys__n37967,
    ys__n37968, ys__n37969, ys__n37970, ys__n37971, ys__n37972, ys__n37973,
    ys__n37974, ys__n37975, ys__n37976, ys__n37977, ys__n37978, ys__n37979,
    ys__n37980, ys__n37981, ys__n37982, ys__n37983, ys__n37984, ys__n37985,
    ys__n37986, ys__n37987, ys__n37988, ys__n37989, ys__n37990, ys__n37991,
    ys__n37992, ys__n37993, ys__n37994, ys__n37995, ys__n37996, ys__n37997,
    ys__n37998, ys__n37999, ys__n38000, ys__n38001, ys__n38002, ys__n38003,
    ys__n38004, ys__n38005, ys__n38006, ys__n38007, ys__n38008, ys__n38009,
    ys__n38010, ys__n38011, ys__n38012, ys__n38013, ys__n38014, ys__n38015,
    ys__n38016, ys__n38017, ys__n38018, ys__n38019, ys__n38020, ys__n38021,
    ys__n38022, ys__n38023, ys__n38024, ys__n38025, ys__n38026, ys__n38027,
    ys__n38028, ys__n38029, ys__n38030, ys__n38031, ys__n38032, ys__n38033,
    ys__n38034, ys__n38035, ys__n38036, ys__n38037, ys__n38038, ys__n38039,
    ys__n38040, ys__n38041, ys__n38042, ys__n38043, ys__n38044, ys__n38045,
    ys__n38046, ys__n38047, ys__n38048, ys__n38049, ys__n38050, ys__n38051,
    ys__n38052, ys__n38053, ys__n38054, ys__n38055, ys__n38056, ys__n38057,
    ys__n38058, ys__n38059, ys__n38060, ys__n38061, ys__n38062, ys__n38063,
    ys__n38064, ys__n38065, ys__n38066, ys__n38067, ys__n38068, ys__n38069,
    ys__n38070, ys__n38071, ys__n38072, ys__n38073, ys__n38074, ys__n38075,
    ys__n38076, ys__n38077, ys__n38078, ys__n38079, ys__n38080, ys__n38081,
    ys__n38082, ys__n38083, ys__n38084, ys__n38085, ys__n38086, ys__n38087,
    ys__n38088, ys__n38089, ys__n38090, ys__n38091, ys__n38092, ys__n38093,
    ys__n38094, ys__n38095, ys__n38096, ys__n38097, ys__n38098, ys__n38099,
    ys__n38100, ys__n38101, ys__n38102, ys__n38103, ys__n38104, ys__n38105,
    ys__n38106, ys__n38107, ys__n38108, ys__n38109, ys__n38110, ys__n38111,
    ys__n38112, ys__n38113, ys__n38114, ys__n38115, ys__n38116, ys__n38117,
    ys__n38118, ys__n38119, ys__n38120, ys__n38121, ys__n38122, ys__n38123,
    ys__n38124, ys__n38125, ys__n38126, ys__n38127, ys__n38128, ys__n38129,
    ys__n38130, ys__n38131, ys__n38132, ys__n38133, ys__n38134, ys__n38135,
    ys__n38136, ys__n38137, ys__n38138, ys__n38139, ys__n38140, ys__n38141,
    ys__n38142, ys__n38143, ys__n38144, ys__n38145, ys__n38146, ys__n38147,
    ys__n38148, ys__n38149, ys__n38150, ys__n38151, ys__n38152, ys__n38153,
    ys__n38154, ys__n38155, ys__n38156, ys__n38157, ys__n38158, ys__n38159,
    ys__n38160, ys__n38161, ys__n38162, ys__n38163, ys__n38164, ys__n38165,
    ys__n38166, ys__n38167, ys__n38168, ys__n38169, ys__n38170, ys__n38171,
    ys__n38172, ys__n38173, ys__n38174, ys__n38175, ys__n38176, ys__n38177,
    ys__n38178, ys__n38179, ys__n38183, ys__n38192, ys__n38193, ys__n38194,
    ys__n38195, ys__n38196, ys__n38197, ys__n38198, ys__n38199, ys__n38200,
    ys__n38201, ys__n38202, ys__n38203, ys__n38212, ys__n38215, ys__n38217,
    ys__n38219, ys__n38220, ys__n38221, ys__n38236, ys__n38237, ys__n38257,
    ys__n38259, ys__n38272, ys__n38277, ys__n38278, ys__n38279, ys__n38282,
    ys__n38283, ys__n38286, ys__n38288, ys__n38290, ys__n38291, ys__n38300,
    ys__n38304, ys__n38305, ys__n38307, ys__n38311, ys__n38315, ys__n38320,
    ys__n38323, ys__n38346, ys__n38361, ys__n38376, ys__n38378, ys__n38380,
    ys__n38382, ys__n38384, ys__n38386, ys__n38398, ys__n38407, ys__n38408,
    ys__n38413, ys__n38418, ys__n38420, ys__n38424, ys__n38427, ys__n38437,
    ys__n38438, ys__n38441, ys__n38443, ys__n38448, ys__n38449, ys__n38451,
    ys__n38473, ys__n38486, ys__n38487, ys__n38488, ys__n38489, ys__n38490,
    ys__n38491, ys__n38494, ys__n38495, ys__n38496, ys__n38497, ys__n38498,
    ys__n38499, ys__n38502, ys__n38503, ys__n38504, ys__n38505, ys__n38506,
    ys__n38507, ys__n38513, ys__n38522, ys__n38524, ys__n38526, ys__n38527,
    ys__n38528, ys__n38529, ys__n38553, ys__n38557, ys__n38561, ys__n38564,
    ys__n38565, ys__n38567, ys__n38568, ys__n38569, ys__n38585, ys__n38586,
    ys__n38587, ys__n38588, ys__n38589, ys__n38590, ys__n38591, ys__n38592,
    ys__n38593, ys__n38594, ys__n38595, ys__n38596, ys__n38597, ys__n38598,
    ys__n38599, ys__n38600, ys__n38601, ys__n38602, ys__n38603, ys__n38604,
    ys__n38605, ys__n38606, ys__n38607, ys__n38608, ys__n38609, ys__n38610,
    ys__n38611, ys__n38620, ys__n38624, ys__n38631, ys__n38649, ys__n38654,
    ys__n38670, ys__n38680, ys__n38693, ys__n38694, ys__n38695, ys__n38724,
    ys__n38776, ys__n38777, ys__n38805, ys__n38827, ys__n38828, ys__n38829,
    ys__n38830, ys__n38831, ys__n38832, ys__n38833, ys__n38834, ys__n38835,
    ys__n38836, ys__n38837, ys__n38838, ys__n38839, ys__n38840, ys__n38841,
    ys__n38842, ys__n38843, ys__n38844, ys__n38845, ys__n38846, ys__n38847,
    ys__n38848, ys__n38849, ys__n38850, ys__n38851, ys__n38852, ys__n38853,
    ys__n38854, ys__n38855, ys__n38856, ys__n38857, ys__n38858, ys__n38859,
    ys__n38861, ys__n38862, ys__n38863, ys__n38864, ys__n38865, ys__n38883,
    ys__n38885, ys__n38893, ys__n38894, ys__n38896, ys__n38897, ys__n38898,
    ys__n38902, ys__n38904, ys__n38906, ys__n38908, ys__n38910, ys__n38919,
    ys__n38922, ys__n38927, ys__n38928, ys__n38929, ys__n39167, ys__n39518,
    ys__n39520, ys__n39718, ys__n39720, ys__n39722, ys__n39724, ys__n39726,
    ys__n39728, ys__n39730, ys__n39732, ys__n39734, ys__n39736, ys__n39738,
    ys__n39740, ys__n39742, ys__n39744, ys__n39746, ys__n39748, ys__n39750,
    ys__n39752, ys__n39754, ys__n39756, ys__n39758, ys__n39760, ys__n39762,
    ys__n39764, ys__n39766, ys__n39768, ys__n39770, ys__n39772, ys__n39774,
    ys__n39776, ys__n39778, ys__n44833, ys__n44840, ys__n44842, ys__n44847,
    ys__n44849, ys__n44892, ys__n44906, ys__n44907, ys__n44908, ys__n44988,
    ys__n44989, ys__n44990, ys__n44991, ys__n44992, ys__n44993, ys__n44995,
    ys__n44996, ys__n44998, ys__n44999, ys__n45001, ys__n45002, ys__n45004,
    ys__n45005, ys__n45007, ys__n45008, ys__n45010, ys__n45011, ys__n45013,
    ys__n45014, ys__n45016, ys__n45017, ys__n45019, ys__n45020, ys__n45022,
    ys__n45023, ys__n45025, ys__n45026, ys__n45028, ys__n45029, ys__n45031,
    ys__n45032, ys__n45034, ys__n45035, ys__n45037, ys__n45038, ys__n45040,
    ys__n45041, ys__n45043, ys__n45044, ys__n45046, ys__n45047, ys__n45049,
    ys__n45050, ys__n45052, ys__n45053, ys__n45055, ys__n45056, ys__n45058,
    ys__n45059, ys__n45061, ys__n45062, ys__n45064, ys__n45065, ys__n45067,
    ys__n45068, ys__n45070, ys__n45071, ys__n45073, ys__n45074, ys__n45076,
    ys__n45077, ys__n45079, ys__n45080, ys__n45082, ys__n45083, ys__n45084,
    ys__n45085, ys__n45086, ys__n45087, ys__n45088, ys__n45089, ys__n45090,
    ys__n45091, ys__n45092, ys__n45093, ys__n45094, ys__n45095, ys__n45096,
    ys__n45097, ys__n45098, ys__n45099, ys__n45100, ys__n45101, ys__n45102,
    ys__n45103, ys__n45104, ys__n45105, ys__n45106, ys__n45107, ys__n45108,
    ys__n45109, ys__n45110, ys__n45111, ys__n45112, ys__n45113, ys__n45115,
    ys__n45116, ys__n45118, ys__n45119, ys__n45121, ys__n45122, ys__n45124,
    ys__n45125, ys__n45127, ys__n45128, ys__n45130, ys__n45131, ys__n45133,
    ys__n45134, ys__n45136, ys__n45137, ys__n45139, ys__n45140, ys__n45142,
    ys__n45143, ys__n45145, ys__n45146, ys__n45148, ys__n45149, ys__n45151,
    ys__n45152, ys__n45154, ys__n45155, ys__n45157, ys__n45158, ys__n45160,
    ys__n45161, ys__n45163, ys__n45164, ys__n45166, ys__n45167, ys__n45169,
    ys__n45170, ys__n45172, ys__n45173, ys__n45175, ys__n45176, ys__n45178,
    ys__n45179, ys__n45181, ys__n45182, ys__n45184, ys__n45185, ys__n45187,
    ys__n45188, ys__n45190, ys__n45191, ys__n45193, ys__n45194, ys__n45196,
    ys__n45197, ys__n45199, ys__n45200, ys__n45202, ys__n45203, ys__n45205,
    ys__n45206, ys__n45208, ys__n45209, ys__n45210, ys__n45211, ys__n45212,
    ys__n45214, ys__n45216, ys__n45218, ys__n45220, ys__n45222, ys__n45224,
    ys__n45226, ys__n45228, ys__n45230, ys__n45232, ys__n45234, ys__n45236,
    ys__n45238, ys__n45240, ys__n45242, ys__n45244, ys__n45246, ys__n45248,
    ys__n45250, ys__n45252, ys__n45254, ys__n45256, ys__n45258, ys__n45260,
    ys__n45262, ys__n45264, ys__n45266, ys__n45268, ys__n45270, ys__n45272,
    ys__n45274, ys__n45276, ys__n45277, ys__n45278, ys__n45279, ys__n45280,
    ys__n45281, ys__n45282, ys__n45283, ys__n45284, ys__n45285, ys__n45286,
    ys__n45287, ys__n45288, ys__n45289, ys__n45290, ys__n45291, ys__n45292,
    ys__n45293, ys__n45294, ys__n45295, ys__n45296, ys__n45297, ys__n45298,
    ys__n45299, ys__n45300, ys__n45301, ys__n45302, ys__n45303, ys__n45304,
    ys__n45305, ys__n45306, ys__n45308, ys__n45310, ys__n45312, ys__n45314,
    ys__n45316, ys__n45318, ys__n45320, ys__n45322, ys__n45324, ys__n45326,
    ys__n45328, ys__n45330, ys__n45332, ys__n45334, ys__n45336, ys__n45338,
    ys__n45340, ys__n45342, ys__n45344, ys__n45346, ys__n45348, ys__n45350,
    ys__n45352, ys__n45354, ys__n45356, ys__n45358, ys__n45360, ys__n45362,
    ys__n45364, ys__n45366, ys__n45368, ys__n45370, ys__n45371, ys__n45372,
    ys__n45373, ys__n45374, ys__n45377, ys__n45380, ys__n45382, ys__n45384,
    ys__n45386, ys__n45388, ys__n45390, ys__n45392, ys__n45394, ys__n45396,
    ys__n45398, ys__n45400, ys__n45402, ys__n45404, ys__n45406, ys__n45408,
    ys__n45410, ys__n45412, ys__n45414, ys__n45416, ys__n45418, ys__n45420,
    ys__n45422, ys__n45424, ys__n45426, ys__n45428, ys__n45430, ys__n45432,
    ys__n45434, ys__n45436, ys__n45438, ys__n45440, ys__n45441, ys__n45442,
    ys__n45443, ys__n45444, ys__n45445, ys__n45446, ys__n45447, ys__n45448,
    ys__n45449, ys__n45450, ys__n45451, ys__n45452, ys__n45453, ys__n45454,
    ys__n45455, ys__n45456, ys__n45457, ys__n45458, ys__n45459, ys__n45460,
    ys__n45461, ys__n45462, ys__n45463, ys__n45464, ys__n45465, ys__n45466,
    ys__n45467, ys__n45468, ys__n45469, ys__n45470, ys__n45472, ys__n45474,
    ys__n45476, ys__n45478, ys__n45480, ys__n45482, ys__n45484, ys__n45486,
    ys__n45488, ys__n45490, ys__n45492, ys__n45494, ys__n45496, ys__n45498,
    ys__n45500, ys__n45502, ys__n45504, ys__n45506, ys__n45508, ys__n45510,
    ys__n45512, ys__n45514, ys__n45516, ys__n45518, ys__n45520, ys__n45522,
    ys__n45524, ys__n45526, ys__n45528, ys__n45530, ys__n45532, ys__n45534,
    ys__n45535, ys__n45536, ys__n45537, ys__n45538, ys__n45541, ys__n45544,
    ys__n45546, ys__n45548, ys__n45550, ys__n45552, ys__n45554, ys__n45556,
    ys__n45558, ys__n45560, ys__n45562, ys__n45564, ys__n45566, ys__n45568,
    ys__n45570, ys__n45572, ys__n45574, ys__n45576, ys__n45578, ys__n45580,
    ys__n45582, ys__n45584, ys__n45586, ys__n45588, ys__n45590, ys__n45592,
    ys__n45594, ys__n45596, ys__n45598, ys__n45600, ys__n45602, ys__n45604,
    ys__n45605, ys__n45606, ys__n45607, ys__n45608, ys__n45609, ys__n45610,
    ys__n45611, ys__n45612, ys__n45613, ys__n45614, ys__n45615, ys__n45616,
    ys__n45617, ys__n45618, ys__n45619, ys__n45620, ys__n45621, ys__n45622,
    ys__n45623, ys__n45624, ys__n45625, ys__n45626, ys__n45627, ys__n45628,
    ys__n45629, ys__n45630, ys__n45631, ys__n45632, ys__n45633, ys__n45634,
    ys__n45636, ys__n45638, ys__n45640, ys__n45642, ys__n45644, ys__n45646,
    ys__n45648, ys__n45650, ys__n45652, ys__n45654, ys__n45656, ys__n45658,
    ys__n45660, ys__n45662, ys__n45664, ys__n45666, ys__n45668, ys__n45670,
    ys__n45672, ys__n45674, ys__n45676, ys__n45678, ys__n45680, ys__n45682,
    ys__n45684, ys__n45686, ys__n45688, ys__n45690, ys__n45692, ys__n45694,
    ys__n45696, ys__n45698, ys__n45699, ys__n45700, ys__n45701, ys__n45702,
    ys__n45704, ys__n45707, ys__n45708, ys__n45709, ys__n45710, ys__n45711,
    ys__n45712, ys__n45714, ys__n45715, ys__n45717, ys__n45718, ys__n45720,
    ys__n45721, ys__n45723, ys__n45724, ys__n45726, ys__n45727, ys__n45729,
    ys__n45730, ys__n45732, ys__n45733, ys__n45735, ys__n45736, ys__n45738,
    ys__n45739, ys__n45741, ys__n45742, ys__n45744, ys__n45745, ys__n45747,
    ys__n45748, ys__n45750, ys__n45751, ys__n45753, ys__n45754, ys__n45756,
    ys__n45757, ys__n45759, ys__n45760, ys__n45762, ys__n45763, ys__n45765,
    ys__n45766, ys__n45768, ys__n45769, ys__n45771, ys__n45772, ys__n45774,
    ys__n45775, ys__n45777, ys__n45778, ys__n45780, ys__n45781, ys__n45783,
    ys__n45784, ys__n45786, ys__n45787, ys__n45789, ys__n45790, ys__n45792,
    ys__n45793, ys__n45795, ys__n45796, ys__n45798, ys__n45799, ys__n45801,
    ys__n45802, ys__n45804, ys__n45805, ys__n45806, ys__n45807, ys__n45808,
    ys__n45809, ys__n45810, ys__n45811, ys__n45812, ys__n45813, ys__n45814,
    ys__n45815, ys__n45816, ys__n45817, ys__n45818, ys__n45819, ys__n45820,
    ys__n45821, ys__n45822, ys__n45823, ys__n45824, ys__n45825, ys__n45826,
    ys__n45827, ys__n45828, ys__n45829, ys__n45830, ys__n45831, ys__n45832,
    ys__n45833, ys__n45834, ys__n45835, ys__n45836, ys__n45838, ys__n45840,
    ys__n45842, ys__n45844, ys__n45846, ys__n45848, ys__n45850, ys__n45852,
    ys__n45854, ys__n45856, ys__n45858, ys__n45860, ys__n45862, ys__n45864,
    ys__n45866, ys__n45868, ys__n45870, ys__n45872, ys__n45874, ys__n45876,
    ys__n45878, ys__n45880, ys__n45882, ys__n45884, ys__n45886, ys__n45888,
    ys__n45890, ys__n45892, ys__n45894, ys__n45896, ys__n45898, ys__n45900,
    ys__n45901, ys__n45902, ys__n45903, ys__n45904, ys__n45905, ys__n45906,
    ys__n45907, ys__n45908, ys__n45909, ys__n45910, ys__n45911, ys__n45912,
    ys__n45913, ys__n45914, ys__n45915, ys__n45916, ys__n45917, ys__n45918,
    ys__n45919, ys__n45920, ys__n45921, ys__n45922, ys__n45923, ys__n45924,
    ys__n45925, ys__n45926, ys__n45927, ys__n45928, ys__n45929, ys__n45930,
    ys__n45931, ys__n45933, ys__n45936, ys__n45938, ys__n45940, ys__n45942,
    ys__n45944, ys__n45946, ys__n45948, ys__n45950, ys__n45952, ys__n45954,
    ys__n45956, ys__n45958, ys__n45960, ys__n45962, ys__n45964, ys__n45966,
    ys__n45968, ys__n45970, ys__n45972, ys__n45974, ys__n45976, ys__n45978,
    ys__n45980, ys__n45982, ys__n45984, ys__n45986, ys__n45988, ys__n45990,
    ys__n45992, ys__n45994, ys__n45996, ys__n45998, ys__n45999, ys__n46000,
    ys__n46001, ys__n46002, ys__n46003, ys__n46004, ys__n46005, ys__n46006,
    ys__n46007, ys__n46008, ys__n46009, ys__n46010, ys__n46011, ys__n46012,
    ys__n46013, ys__n46014, ys__n46015, ys__n46016, ys__n46017, ys__n46018,
    ys__n46019, ys__n46020, ys__n46021, ys__n46022, ys__n46023, ys__n46024,
    ys__n46025, ys__n46026, ys__n46027, ys__n46028, ys__n46029, ys__n46031,
    ys__n46034, ys__n46036, ys__n46038, ys__n46040, ys__n46042, ys__n46044,
    ys__n46046, ys__n46048, ys__n46050, ys__n46052, ys__n46054, ys__n46056,
    ys__n46058, ys__n46060, ys__n46062, ys__n46064, ys__n46066, ys__n46068,
    ys__n46070, ys__n46072, ys__n46074, ys__n46076, ys__n46078, ys__n46080,
    ys__n46082, ys__n46084, ys__n46086, ys__n46088, ys__n46090, ys__n46092,
    ys__n46094, ys__n46096, ys__n46097, ys__n46098, ys__n46099, ys__n46100,
    ys__n46101, ys__n46102, ys__n46103, ys__n46104, ys__n46105, ys__n46106,
    ys__n46107, ys__n46108, ys__n46109, ys__n46110, ys__n46111, ys__n46112,
    ys__n46113, ys__n46114, ys__n46115, ys__n46116, ys__n46117, ys__n46118,
    ys__n46119, ys__n46120, ys__n46121, ys__n46122, ys__n46123, ys__n46124,
    ys__n46125, ys__n46126, ys__n46127, ys__n46128, ys__n46130, ys__n46132,
    ys__n46134, ys__n46136, ys__n46141, ys__n46142, ys__n46150, ys__n46151,
    ys__n46152, ys__n46153, ys__n46166, ys__n46168, ys__n46169, ys__n46170,
    ys__n46171, ys__n46180, ys__n46184, ys__n46185, ys__n46186, ys__n46187,
    ys__n46198, ys__n46200, ys__n46201, ys__n46202, ys__n46203, ys__n46214,
    ys__n46216, ys__n46217, ys__n46218, ys__n46219, ys__n46230, ys__n46231,
    ys__n46238, ys__n46239, ys__n46240, ys__n46242, ys__n46244, ys__n46245,
    ys__n46247, ys__n46248, ys__n46252, ys__n46254, ys__n46256, ys__n46258,
    ys__n46260, ys__n46262, ys__n46264, ys__n46266, ys__n46268, ys__n46270,
    ys__n46272, ys__n46274, ys__n46276, ys__n46278, ys__n46280, ys__n46282,
    ys__n46284, ys__n46286, ys__n46288, ys__n46290, ys__n46292, ys__n46294,
    ys__n46296, ys__n46298, ys__n46300, ys__n46302, ys__n46304, ys__n46306,
    ys__n46308, ys__n46310, ys__n46312, ys__n46314, ys__n46315, ys__n46316,
    ys__n46317, ys__n46318, ys__n46319, ys__n46320, ys__n46321, ys__n46322,
    ys__n46323, ys__n46324, ys__n46325, ys__n46326, ys__n46327, ys__n46328,
    ys__n46329, ys__n46330, ys__n46331, ys__n46332, ys__n46333, ys__n46334,
    ys__n46335, ys__n46336, ys__n46337, ys__n46338, ys__n46339, ys__n46340,
    ys__n46341, ys__n46342, ys__n46343, ys__n46344, ys__n46345, ys__n46346,
    ys__n46348, ys__n46350, ys__n46352, ys__n46354, ys__n46356, ys__n46358,
    ys__n46360, ys__n46362, ys__n46364, ys__n46366, ys__n46368, ys__n46370,
    ys__n46372, ys__n46374, ys__n46376, ys__n46378, ys__n46380, ys__n46382,
    ys__n46384, ys__n46386, ys__n46388, ys__n46390, ys__n46392, ys__n46393,
    ys__n46394, ys__n46395, ys__n46396, ys__n46397, ys__n46398, ys__n46399,
    ys__n46400, ys__n46401, ys__n46402, ys__n46403, ys__n46404, ys__n46405,
    ys__n46406, ys__n46407, ys__n46408, ys__n46409, ys__n46410, ys__n46411,
    ys__n46412, ys__n46413, ys__n46414, ys__n46415, ys__n46416, ys__n46417,
    ys__n46418, ys__n46419, ys__n46420, ys__n46421, ys__n46422, ys__n46423,
    ys__n46428, ys__n46430, ys__n46432, ys__n46434, ys__n46436, ys__n46438,
    ys__n46440, ys__n46442, ys__n46444, ys__n46446, ys__n46448, ys__n46450,
    ys__n46452, ys__n46454, ys__n46456, ys__n46458, ys__n46460, ys__n46462,
    ys__n46464, ys__n46466, ys__n46468, ys__n46470, ys__n46472, ys__n46474,
    ys__n46476, ys__n46478, ys__n46480, ys__n46482, ys__n46484, ys__n46486,
    ys__n46488, ys__n46490, ys__n46491, ys__n46492, ys__n46493, ys__n46494,
    ys__n46495, ys__n46496, ys__n46497, ys__n46498, ys__n46499, ys__n46500,
    ys__n46501, ys__n46502, ys__n46503, ys__n46504, ys__n46505, ys__n46506,
    ys__n46507, ys__n46508, ys__n46509, ys__n46510, ys__n46511, ys__n46512,
    ys__n46513, ys__n46514, ys__n46515, ys__n46516, ys__n46517, ys__n46518,
    ys__n46519, ys__n46520, ys__n46521, ys__n46522, ys__n46524, ys__n46526,
    ys__n46528, ys__n46530, ys__n46532, ys__n46534, ys__n46536, ys__n46538,
    ys__n46540, ys__n46542, ys__n46544, ys__n46546, ys__n46548, ys__n46550,
    ys__n46552, ys__n46554, ys__n46556, ys__n46558, ys__n46560, ys__n46562,
    ys__n46564, ys__n46566, ys__n46568, ys__n46569, ys__n46570, ys__n46571,
    ys__n46572, ys__n46573, ys__n46574, ys__n46575, ys__n46576, ys__n46577,
    ys__n46578, ys__n46579, ys__n46580, ys__n46581, ys__n46582, ys__n46583,
    ys__n46584, ys__n46585, ys__n46586, ys__n46587, ys__n46588, ys__n46589,
    ys__n46590, ys__n46591, ys__n46592, ys__n46593, ys__n46594, ys__n46595,
    ys__n46596, ys__n46597, ys__n46598, ys__n46599, ys__n46604, ys__n46606,
    ys__n46608, ys__n46610, ys__n46612, ys__n46614, ys__n46616, ys__n46618,
    ys__n46620, ys__n46622, ys__n46624, ys__n46626, ys__n46628, ys__n46630,
    ys__n46632, ys__n46634, ys__n46636, ys__n46638, ys__n46640, ys__n46642,
    ys__n46644, ys__n46646, ys__n46648, ys__n46650, ys__n46652, ys__n46654,
    ys__n46656, ys__n46658, ys__n46660, ys__n46662, ys__n46664, ys__n46666,
    ys__n46667, ys__n46668, ys__n46669, ys__n46670, ys__n46671, ys__n46672,
    ys__n46673, ys__n46674, ys__n46675, ys__n46676, ys__n46677, ys__n46678,
    ys__n46679, ys__n46680, ys__n46681, ys__n46682, ys__n46683, ys__n46684,
    ys__n46685, ys__n46686, ys__n46687, ys__n46688, ys__n46689, ys__n46690,
    ys__n46691, ys__n46692, ys__n46693, ys__n46694, ys__n46695, ys__n46696,
    ys__n46697, ys__n46698, ys__n46700, ys__n46702, ys__n46704, ys__n46706,
    ys__n46708, ys__n46710, ys__n46712, ys__n46714, ys__n46716, ys__n46718,
    ys__n46720, ys__n46722, ys__n46724, ys__n46726, ys__n46728, ys__n46730,
    ys__n46732, ys__n46734, ys__n46736, ys__n46738, ys__n46740, ys__n46742,
    ys__n46744, ys__n46745, ys__n46746, ys__n46747, ys__n46748, ys__n46749,
    ys__n46750, ys__n46751, ys__n46752, ys__n46753, ys__n46754, ys__n46755,
    ys__n46756, ys__n46757, ys__n46758, ys__n46759, ys__n46760, ys__n46761,
    ys__n46762, ys__n46763, ys__n46764, ys__n46765, ys__n46766, ys__n46767,
    ys__n46768, ys__n46769, ys__n46770, ys__n46771, ys__n46772, ys__n46773,
    ys__n46774, ys__n46775, ys__n46780, ys__n46782, ys__n46784, ys__n46786,
    ys__n46788, ys__n46790, ys__n46792, ys__n46794, ys__n46796, ys__n46798,
    ys__n46800, ys__n46802, ys__n46804, ys__n46806, ys__n46808, ys__n46810,
    ys__n46812, ys__n46814, ys__n46816, ys__n46818, ys__n46820, ys__n46822,
    ys__n46824, ys__n46826, ys__n46828, ys__n46830, ys__n46832, ys__n46834,
    ys__n46836, ys__n46838, ys__n46840, ys__n46842, ys__n46843, ys__n46844,
    ys__n46845, ys__n46846, ys__n46847, ys__n46848, ys__n46849, ys__n46850,
    ys__n46851, ys__n46852, ys__n46853, ys__n46854, ys__n46855, ys__n46856,
    ys__n46857, ys__n46858, ys__n46859, ys__n46860, ys__n46861, ys__n46862,
    ys__n46863, ys__n46864, ys__n46865, ys__n46866, ys__n46867, ys__n46868,
    ys__n46869, ys__n46870, ys__n46871, ys__n46872, ys__n46873, ys__n46874,
    ys__n46876, ys__n46878, ys__n46880, ys__n46882, ys__n46884, ys__n46886,
    ys__n46888, ys__n46890, ys__n46892, ys__n46894, ys__n46896, ys__n46898,
    ys__n46900, ys__n46902, ys__n46904, ys__n46906, ys__n46908, ys__n46910,
    ys__n46912, ys__n46914, ys__n46916, ys__n46918, ys__n46920, ys__n46921,
    ys__n46922, ys__n46923, ys__n46924, ys__n46925, ys__n46926, ys__n46927,
    ys__n46928, ys__n46929, ys__n46930, ys__n46931, ys__n46932, ys__n46933,
    ys__n46934, ys__n46935, ys__n46936, ys__n46937, ys__n46938, ys__n46939,
    ys__n46940, ys__n46941, ys__n46942, ys__n46943, ys__n46944, ys__n46945,
    ys__n46946, ys__n46947, ys__n46948, ys__n46949, ys__n46950, ys__n46951,
    ys__n46954, ys__n46955, ys__n46956, ys__n46957, ys__n46958, ys__n46959,
    ys__n46960, ys__n46961, ys__n46962, ys__n46963, ys__n46964, ys__n46965,
    ys__n46966, ys__n46967, ys__n46968, ys__n46969, ys__n46970, ys__n46971,
    ys__n46972, ys__n46973, ys__n46974, ys__n46975, ys__n46976, ys__n46977,
    ys__n46978, ys__n46979, ys__n46980, ys__n46981, ys__n46982, ys__n46983,
    ys__n46984, ys__n46985, ys__n46986, ys__n46987, ys__n46988, ys__n46989,
    ys__n46990, ys__n46991, ys__n46992, ys__n46993, ys__n46994, ys__n46995,
    ys__n46996, ys__n46997, ys__n46998, ys__n46999, ys__n47000, ys__n47001,
    ys__n47002, ys__n47003, ys__n47004, ys__n47005, ys__n47006, ys__n47007,
    ys__n47008, ys__n47009, ys__n47010, ys__n47011, ys__n47012, ys__n47013,
    ys__n47014, ys__n47015, ys__n47016, ys__n47017, ys__n47018, ys__n47019,
    ys__n47020, ys__n47021, ys__n47022, ys__n47023, ys__n47024, ys__n47025,
    ys__n47026, ys__n47027, ys__n47028, ys__n47029, ys__n47030, ys__n47031,
    ys__n47032, ys__n47033, ys__n47034, ys__n47035, ys__n47036, ys__n47037,
    ys__n47038, ys__n47039, ys__n47040, ys__n47041, ys__n47074, ys__n47075,
    ys__n47076, ys__n47077, ys__n47078, ys__n47079, ys__n47080, ys__n47081,
    ys__n47082, ys__n47083, ys__n47084, ys__n47085, ys__n47086, ys__n47087,
    ys__n47088, ys__n47089, ys__n47090, ys__n47091, ys__n47092, ys__n47093,
    ys__n47094, ys__n47095, ys__n47096, ys__n47097, ys__n47098, ys__n47099,
    ys__n47100, ys__n47101, ys__n47102, ys__n47103, ys__n47104, ys__n47105,
    ys__n47106, ys__n47107, ys__n47108, ys__n47109, ys__n47110, ys__n47111,
    ys__n47112, ys__n47113, ys__n47114, ys__n47115, ys__n47116, ys__n47117,
    ys__n47118, ys__n47119, ys__n47184, ys__n47185, ys__n47186, ys__n47187,
    ys__n47188, ys__n47189, ys__n47190, ys__n47191, ys__n47192, ys__n47193,
    ys__n47194, ys__n47195, ys__n47196, ys__n47197, ys__n47198, ys__n47199,
    ys__n47200, ys__n47201, ys__n47202, ys__n47203, ys__n47204, ys__n47205,
    ys__n47206, ys__n47207, ys__n47208, ys__n47209, ys__n47210, ys__n47211,
    ys__n47212, ys__n47213, ys__n47214, ys__n47215, ys__n47216, ys__n47217,
    ys__n47218, ys__n47219, ys__n47220, ys__n47221, ys__n47222, ys__n47223,
    ys__n47224, ys__n47225, ys__n47226, ys__n47227, ys__n47228, ys__n47229,
    ys__n47230, ys__n47231, ys__n47232, ys__n47233, ys__n47234, ys__n47235,
    ys__n47236, ys__n47237, ys__n47238, ys__n47239, ys__n47240, ys__n47241,
    ys__n47242, ys__n47243, ys__n47244, ys__n47245, ys__n47246, ys__n47247,
    ys__n47248, ys__n47249, ys__n47250, ys__n47251, ys__n47252, ys__n47253,
    ys__n47254, ys__n47255, ys__n47256, ys__n47257, ys__n47258, ys__n47259,
    ys__n47260, ys__n47261, ys__n47262, ys__n47263, ys__n47264, ys__n47265,
    ys__n47266, ys__n47267, ys__n47268, ys__n47269, ys__n47270, ys__n47271,
    ys__n47272, ys__n47273, ys__n47274, ys__n47275, ys__n47276, ys__n47277,
    ys__n47278, ys__n47279, ys__n47280, ys__n47281, ys__n47282, ys__n47283,
    ys__n47284, ys__n47285, ys__n47286, ys__n47287, ys__n47288, ys__n47289,
    ys__n47290, ys__n47291, ys__n47292, ys__n47293, ys__n47294, ys__n47295,
    ys__n47296, ys__n47297, ys__n47298, ys__n47299, ys__n47300, ys__n47301,
    ys__n47302, ys__n47303, ys__n47305, ys__n47306, ys__n47307, ys__n47308,
    ys__n47309, ys__n47310, ys__n47311, ys__n47312, ys__n47313, ys__n47314,
    ys__n47315, ys__n47316, ys__n47317, ys__n47318, ys__n47319, ys__n47320,
    ys__n47321, ys__n47322, ys__n47323, ys__n47324, ys__n47325, ys__n47326,
    ys__n47327, ys__n47328, ys__n47329, ys__n47330, ys__n47331, ys__n47332,
    ys__n47333, ys__n47334, ys__n47335, ys__n47336, ys__n47337, ys__n47338,
    ys__n47339, ys__n47340, ys__n47341, ys__n47342, ys__n47343, ys__n47344,
    ys__n47345, ys__n47346, ys__n47347, ys__n47348, ys__n47349, ys__n47350,
    ys__n47351, ys__n47352, ys__n47353, ys__n47354, ys__n47355, ys__n47356,
    ys__n47357, ys__n47358, ys__n47359, ys__n47360, ys__n47361, ys__n47362,
    ys__n47363, ys__n47364, ys__n47365, ys__n47366, ys__n47367, ys__n47368,
    ys__n47369, ys__n47370, ys__n47371, ys__n47372, ys__n47373, ys__n47374,
    ys__n47375, ys__n47376, ys__n47377, ys__n47378, ys__n47379, ys__n47380,
    ys__n47381, ys__n47382, ys__n47383, ys__n47384, ys__n47385, ys__n47386,
    ys__n47387, ys__n47388, ys__n47389, ys__n47390, ys__n47391, ys__n47392,
    ys__n47393, ys__n47394, ys__n47395, ys__n47396, ys__n47397, ys__n47398,
    ys__n47399, ys__n47400, ys__n47401, ys__n47402, ys__n47403, ys__n47404,
    ys__n47405, ys__n47406, ys__n47407, ys__n47408, ys__n47409, ys__n47410,
    ys__n47411, ys__n47412, ys__n47413, ys__n47414, ys__n47415, ys__n47416,
    ys__n47417, ys__n47418, ys__n47419, ys__n47420, ys__n47421, ys__n47422,
    ys__n47423, ys__n47424, ys__n47425, ys__n47426, ys__n47427, ys__n47428,
    ys__n47429, ys__n47430, ys__n47431, ys__n47432, ys__n47433, ys__n47434,
    ys__n47435, ys__n47436, ys__n47437, ys__n47438, ys__n47439, ys__n47440,
    ys__n47441, ys__n47442, ys__n47443, ys__n47444, ys__n47445, ys__n47446,
    ys__n47447, ys__n47448, ys__n47449, ys__n47450, ys__n47451, ys__n47452,
    ys__n47453, ys__n47454, ys__n47455, ys__n47456, ys__n47457, ys__n47458,
    ys__n47459, ys__n47460, ys__n47461, ys__n47462, ys__n47463, ys__n47464,
    ys__n47465, ys__n47466, ys__n47467, ys__n47468, ys__n47469, ys__n47470,
    ys__n47471, ys__n47472, ys__n47473, ys__n47474, ys__n47475, ys__n47476,
    ys__n47477, ys__n47478, ys__n47479, ys__n47480, ys__n47481, ys__n47482,
    ys__n47483, ys__n47484, ys__n47485, ys__n47486, ys__n47487, ys__n47488,
    ys__n47489, ys__n47490, ys__n47491, ys__n47492, ys__n47493, ys__n47494,
    ys__n47495, ys__n47496, ys__n47497, ys__n47498, ys__n47499, ys__n47500,
    ys__n47501, ys__n47502, ys__n47503, ys__n47504, ys__n47505, ys__n47506,
    ys__n47507, ys__n47508, ys__n47509, ys__n47510, ys__n47511, ys__n47512,
    ys__n47513, ys__n47514, ys__n47515, ys__n47516, ys__n47517, ys__n47518,
    ys__n47519, ys__n47520, ys__n47521, ys__n47522, ys__n47523, ys__n47524,
    ys__n47525, ys__n47526, ys__n47527, ys__n47528, ys__n47529, ys__n47530,
    ys__n47531, ys__n47532, ys__n47533, ys__n47534, ys__n47535, ys__n47536,
    ys__n47537, ys__n47538, ys__n47539, ys__n47540, ys__n47541, ys__n47542,
    ys__n47543, ys__n47544, ys__n47545, ys__n47546, ys__n47547, ys__n47548,
    ys__n47549, ys__n47550, ys__n47551, ys__n47552, ys__n47553, ys__n47554,
    ys__n47555, ys__n47556, ys__n47557, ys__n47558, ys__n47559, ys__n47560,
    ys__n47561, ys__n47562, ys__n47563, ys__n47564, ys__n47565, ys__n47566,
    ys__n47567, ys__n47568, ys__n47569, ys__n47570, ys__n47571, ys__n47572,
    ys__n47573, ys__n47574, ys__n47575, ys__n47576, ys__n47577, ys__n47578,
    ys__n47579, ys__n47580, ys__n47581, ys__n47582, ys__n47583, ys__n47584,
    ys__n47585, ys__n47586, ys__n47587, ys__n47588, ys__n47589, ys__n47590,
    ys__n47591, ys__n47592, ys__n47593, ys__n47594, ys__n47595, ys__n47596,
    ys__n47597, ys__n47598, ys__n47599, ys__n47600, ys__n47601, ys__n47602,
    ys__n47603, ys__n47604, ys__n47605, ys__n47606, ys__n47607, ys__n47608,
    ys__n47609, ys__n47610, ys__n47611, ys__n47612, ys__n47613, ys__n47614,
    ys__n47615, ys__n47616, ys__n47617, ys__n47618, ys__n47619, ys__n47620,
    ys__n47621, ys__n47622, ys__n47623, ys__n47624, ys__n47625, ys__n47626,
    ys__n47627, ys__n47628, ys__n47629, ys__n47630, ys__n47631, ys__n47632,
    ys__n47633, ys__n47634, ys__n47635, ys__n47636, ys__n47637, ys__n47638,
    ys__n47639, ys__n47640, ys__n47641, ys__n47642, ys__n47643, ys__n47644,
    ys__n47645, ys__n47646, ys__n47647, ys__n47648, ys__n47649, ys__n47650,
    ys__n47651, ys__n47652, ys__n47653, ys__n47654, ys__n47655, ys__n47656,
    ys__n47657, ys__n47658, ys__n47659, ys__n47660, ys__n47661, ys__n47662,
    ys__n47663, ys__n47664, ys__n47665, ys__n47666, ys__n47667, ys__n47668,
    ys__n47669, ys__n47670, ys__n47671, ys__n47672, ys__n47673, ys__n47674,
    ys__n47675, ys__n47676, ys__n47677, ys__n47678, ys__n47679, ys__n47680,
    ys__n47681, ys__n47682, ys__n47683, ys__n47684, ys__n47685, ys__n47686,
    ys__n47687, ys__n47688, ys__n47689, ys__n47690, ys__n47691, ys__n47692,
    ys__n47693, ys__n47694, ys__n47695, ys__n47696, ys__n47697, ys__n47698,
    ys__n47699, ys__n47700, ys__n47701, ys__n47702, ys__n47703, ys__n47704,
    ys__n47705, ys__n47706, ys__n47707, ys__n47708, ys__n47709, ys__n47710,
    ys__n47711, ys__n47712, ys__n47713, ys__n47714, ys__n47715, ys__n47716,
    ys__n47717, ys__n47718, ys__n47719, ys__n47720, ys__n47721, ys__n47722,
    ys__n47723, ys__n47724, ys__n47725, ys__n47726, ys__n47727, ys__n47728,
    ys__n47729, ys__n47730, ys__n47731, ys__n47732, ys__n47733, ys__n47734,
    ys__n47735, ys__n47736, ys__n47737, ys__n47738, ys__n47739, ys__n47740,
    ys__n47741, ys__n47742, ys__n47743, ys__n47744, ys__n47745, ys__n47746,
    ys__n47747, ys__n47748, ys__n47749, ys__n47750, ys__n47751, ys__n47752,
    ys__n47753, ys__n47754, ys__n47755, ys__n47756, ys__n47757, ys__n47758,
    ys__n47759, ys__n47760, ys__n47761, ys__n47762, ys__n47763, ys__n47764,
    ys__n47765, ys__n47766, ys__n47767, ys__n47768, ys__n47769, ys__n47770,
    ys__n47771, ys__n47772, ys__n47773, ys__n47774, ys__n47775, ys__n47776,
    ys__n47777, ys__n47778, ys__n47779, ys__n47780, ys__n47781, ys__n47782,
    ys__n47783, ys__n47784, ys__n47785, ys__n47786, ys__n47787, ys__n47788,
    ys__n47789, ys__n47790, ys__n47791, ys__n47792, ys__n47793, ys__n47794,
    ys__n47795, ys__n47796, ys__n47797, ys__n47798, ys__n47799, ys__n47800,
    ys__n47801, ys__n47802, ys__n47803, ys__n47804, ys__n47805, ys__n47806,
    ys__n47807, ys__n47808, ys__n47809, ys__n47810, ys__n47811, ys__n47812,
    ys__n47813, ys__n47814, ys__n47815, ys__n47816, ys__n47817, ys__n47818,
    ys__n47819, ys__n47820, ys__n47821, ys__n47822, ys__n47823, ys__n47824,
    ys__n47825, ys__n47826, ys__n47827, ys__n47828, ys__n47829, ys__n47830,
    ys__n47831, ys__n47832, ys__n47833, ys__n47834, ys__n47835, ys__n47836,
    ys__n47837, ys__n47838, ys__n47839, ys__n47840, ys__n47841, ys__n47842,
    ys__n47843, ys__n47844, ys__n47845, ys__n47846, ys__n47847, ys__n47848,
    ys__n47849, ys__n47850, ys__n47851, ys__n47852, ys__n47853, ys__n47854,
    ys__n47855, ys__n47856, ys__n47857, ys__n47858, ys__n47859, ys__n47860,
    ys__n47861, ys__n47862, ys__n47863, ys__n47864, ys__n47865, ys__n47866,
    ys__n47867, ys__n47868, ys__n47869, ys__n47870, ys__n47871, ys__n47872,
    ys__n47873, ys__n47874, ys__n47875, ys__n47876, ys__n47877, ys__n47878,
    ys__n47879, ys__n47880, ys__n47881, ys__n47882, ys__n47883, ys__n47884,
    ys__n47885, ys__n47886, ys__n47887, ys__n47888, ys__n47889, ys__n47890,
    ys__n47891, ys__n47892, ys__n47893, ys__n47894, ys__n47895, ys__n47896,
    ys__n47897, ys__n47898, ys__n47899, ys__n47900, ys__n47901, ys__n47902,
    ys__n47903, ys__n47904, ys__n47905, ys__n47906, ys__n47907, ys__n47908,
    ys__n47909, ys__n47910, ys__n47911, ys__n47912, ys__n47913, ys__n47914,
    ys__n47915, ys__n47916, ys__n47917, ys__n47918, ys__n47919, ys__n47920,
    ys__n47921, ys__n47922, ys__n47923, ys__n47924, ys__n47925, ys__n47926,
    ys__n47927, ys__n47928, ys__n47929, ys__n47930, ys__n47931, ys__n47932,
    ys__n47933, ys__n47934, ys__n47935, ys__n47936, ys__n47937, ys__n47938,
    ys__n47939, ys__n47940, ys__n47941, ys__n47942, ys__n47943, ys__n47944,
    ys__n47945, ys__n47946, ys__n47947, ys__n47948, ys__n47949, ys__n47950,
    ys__n47951, ys__n47952, ys__n47953, ys__n47954, ys__n47955, ys__n47956,
    ys__n47957, ys__n47958, ys__n47959, ys__n47960, ys__n47961, ys__n47962,
    ys__n47963, ys__n47964, ys__n47965, ys__n47966, ys__n47967, ys__n47968,
    ys__n47969, ys__n47970, ys__n47971, ys__n47972, ys__n47973, ys__n47974,
    ys__n47975, ys__n47976, ys__n47977, ys__n47978, ys__n47979, ys__n47980,
    ys__n47981, ys__n47982, ys__n47983, ys__n47984, ys__n47985, ys__n47986,
    ys__n47987, ys__n47988, ys__n47989, ys__n47990, ys__n47991, ys__n47992,
    ys__n47993, ys__n47994, ys__n47995, ys__n47996, ys__n47997, ys__n47998,
    ys__n47999, ys__n48000, ys__n48001, ys__n48002, ys__n48003, ys__n48004,
    ys__n48005, ys__n48006, ys__n48007, ys__n48008, ys__n48009, ys__n48010,
    ys__n48011, ys__n48012, ys__n48013, ys__n48014, ys__n48015, ys__n48016,
    ys__n48017, ys__n48018, ys__n48019, ys__n48020, ys__n48021, ys__n48022,
    ys__n48023, ys__n48024, ys__n48025, ys__n48026, ys__n48027, ys__n48028,
    ys__n48029, ys__n48030, ys__n48031, ys__n48032, ys__n48033, ys__n48034,
    ys__n48035, ys__n48036, ys__n48037, ys__n48038, ys__n48039, ys__n48040,
    ys__n48041, ys__n48042, ys__n48043, ys__n48044, ys__n48045, ys__n48046,
    ys__n48047, ys__n48048, ys__n48049, ys__n48050, ys__n48051, ys__n48052,
    ys__n48053, ys__n48054, ys__n48055, ys__n48056, ys__n48057, ys__n48058,
    ys__n48059, ys__n48060, ys__n48061, ys__n48062, ys__n48063, ys__n48064,
    ys__n48065, ys__n48066, ys__n48067, ys__n48068, ys__n48069, ys__n48070,
    ys__n48071, ys__n48072, ys__n48073, ys__n48074, ys__n48075, ys__n48076,
    ys__n48077, ys__n48078, ys__n48079, ys__n48080, ys__n48081, ys__n48082,
    ys__n48083, ys__n48084, ys__n48085, ys__n48086, ys__n48087, ys__n48088,
    ys__n48089, ys__n48090, ys__n48091, ys__n48092, ys__n48093, ys__n48094,
    ys__n48095, ys__n48096, ys__n48097, ys__n48098, ys__n48099, ys__n48100,
    ys__n48101, ys__n48102, ys__n48103, ys__n48104, ys__n48105, ys__n48106,
    ys__n48107, ys__n48108, ys__n48109, ys__n48110, ys__n48111, ys__n48112,
    ys__n48113, ys__n48114, ys__n48115, ys__n48116, ys__n48117, ys__n48118,
    ys__n48119, ys__n48120, ys__n48121, ys__n48122, ys__n48123, ys__n48124,
    ys__n48125, ys__n48126, ys__n48127, ys__n48128, ys__n48129, ys__n48130,
    ys__n48131, ys__n48132, ys__n48133, ys__n48134, ys__n48135, ys__n48136,
    ys__n48137, ys__n48138, ys__n48139, ys__n48140, ys__n48141, ys__n48142,
    ys__n48143, ys__n48144, ys__n48145, ys__n48146, ys__n48147, ys__n48148,
    ys__n48149, ys__n48150, ys__n48151, ys__n48152, ys__n48153, ys__n48154,
    ys__n48155, ys__n48156, ys__n48157, ys__n48158, ys__n48159, ys__n48160,
    ys__n48161, ys__n48162, ys__n48163, ys__n48164, ys__n48165, ys__n48166,
    ys__n48167, ys__n48168, ys__n48169, ys__n48170, ys__n48171, ys__n48172,
    ys__n48173, ys__n48174, ys__n48175, ys__n48176, ys__n48177, ys__n48178,
    ys__n48179, ys__n48180, ys__n48181, ys__n48182, ys__n48183, ys__n48184,
    ys__n48185, ys__n48186, ys__n48187, ys__n48188, ys__n48189, ys__n48190,
    ys__n48191, ys__n48192, ys__n48193, ys__n48194, ys__n48195, ys__n48196,
    ys__n48197, ys__n48198, ys__n48199, ys__n48200, ys__n48201, ys__n48202,
    ys__n48203, ys__n48204, ys__n48205, ys__n48206, ys__n48207, ys__n48208,
    ys__n48209, ys__n48210, ys__n48211, ys__n48212, ys__n48213, ys__n48214,
    ys__n48215, ys__n48216, ys__n48217, ys__n48218, ys__n48219, ys__n48220,
    ys__n48221, ys__n48222, ys__n48223, ys__n48224, ys__n48225, ys__n48226,
    ys__n48227, ys__n48228, ys__n48229, ys__n48230, ys__n48231, ys__n48232,
    ys__n48233, ys__n48234, ys__n48235, ys__n48236, ys__n48237, ys__n48238,
    ys__n48239, ys__n48240, ys__n48241, ys__n48242, ys__n48243, ys__n48244,
    ys__n48245, ys__n48246, ys__n48247, ys__n48248, ys__n48249, ys__n48250,
    ys__n48251, ys__n48252, ys__n48253, ys__n48254, ys__n48255, ys__n48256,
    ys__n48257, ys__n48258, ys__n48259, ys__n48260, ys__n48261, ys__n48262,
    ys__n48263, ys__n48264, ys__n48265, ys__n48266, ys__n48267, ys__n48268,
    ys__n48269, ys__n48270, ys__n48271, ys__n48272, ys__n48273, ys__n48274,
    ys__n48275, ys__n48324, ys__n48325, ys__n48327, ys__n48330, ys__n48331,
    ys__n48332, ys__n48333, ys__n48334, ys__n48335;
  output ys__n2, ys__n246, ys__n250, ys__n252, ys__n254, ys__n264, ys__n270,
    ys__n278, ys__n280, ys__n313, ys__n319, ys__n404, ys__n415, ys__n417,
    ys__n455, ys__n457, ys__n478, ys__n480, ys__n482, ys__n502, ys__n565,
    ys__n574, ys__n576, ys__n628, ys__n630, ys__n714, ys__n716, ys__n730,
    ys__n732, ys__n738, ys__n740, ys__n754, ys__n756, ys__n786, ys__n788,
    ys__n790, ys__n792, ys__n794, ys__n796, ys__n798, ys__n800, ys__n802,
    ys__n804, ys__n806, ys__n808, ys__n810, ys__n812, ys__n814, ys__n862,
    ys__n863, ys__n865, ys__n866, ys__n868, ys__n870, ys__n871, ys__n872,
    ys__n873, ys__n876, ys__n878, ys__n879, ys__n881, ys__n888, ys__n890,
    ys__n900, ys__n902, ys__n904, ys__n911, ys__n920, ys__n923, ys__n927,
    ys__n929, ys__n930, ys__n932, ys__n934, ys__n936, ys__n942, ys__n944,
    ys__n948, ys__n949, ys__n970, ys__n972, ys__n974, ys__n976, ys__n978,
    ys__n980, ys__n982, ys__n989, ys__n991, ys__n993, ys__n995, ys__n999,
    ys__n1001, ys__n1004, ys__n1007, ys__n1009, ys__n1013, ys__n1020,
    ys__n1028, ys__n1030, ys__n1031, ys__n1032, ys__n1037, ys__n1040,
    ys__n1043, ys__n1046, ys__n1047, ys__n1049, ys__n1060, ys__n1071,
    ys__n1073, ys__n1074, ys__n1075, ys__n1077, ys__n1079, ys__n1080,
    ys__n1083, ys__n1085, ys__n1087, ys__n1088, ys__n1089, ys__n1090,
    ys__n1091, ys__n1095, ys__n1103, ys__n1115, ys__n1125, ys__n1128,
    ys__n1135, ys__n1138, ys__n1141, ys__n1142, ys__n1143, ys__n1146,
    ys__n1148, ys__n1161, ys__n1163, ys__n1164, ys__n1165, ys__n1167,
    ys__n1170, ys__n1171, ys__n1183, ys__n1189, ys__n1195, ys__n1201,
    ys__n1207, ys__n1213, ys__n1219, ys__n1222, ys__n1228, ys__n1234,
    ys__n1240, ys__n1246, ys__n1252, ys__n1258, ys__n1261, ys__n1266,
    ys__n1272, ys__n1278, ys__n1284, ys__n1290, ys__n1296, ys__n1303,
    ys__n1377, ys__n1386, ys__n1445, ys__n1448, ys__n1470, ys__n1591,
    ys__n1598, ys__n1601, ys__n1616, ys__n1790, ys__n1802, ys__n1817,
    ys__n1835, ys__n1837, ys__n2152, ys__n2365, ys__n2400, ys__n2423,
    ys__n2491, ys__n2535, ys__n2536, ys__n2582, ys__n2635, ys__n2651,
    ys__n2653, ys__n2655, ys__n2674, ys__n2684, ys__n2733, ys__n2776,
    ys__n2778, ys__n2780, ys__n2782, ys__n2804, ys__n2806, ys__n2845,
    ys__n2855, ys__n3021, ys__n3024, ys__n3035, ys__n3039, ys__n3040,
    ys__n3051, ys__n3061, ys__n3068, ys__n3083, ys__n3085, ys__n3097,
    ys__n3106, ys__n3114, ys__n3115, ys__n3118, ys__n3121, ys__n3195,
    ys__n3249, ys__n3250, ys__n3252, ys__n4175, ys__n4189, ys__n4192,
    ys__n4320, ys__n4414, ys__n4521, ys__n4566, ys__n4588, ys__n4603,
    ys__n4615, ys__n4696, ys__n4764, ys__n4791, ys__n4793, ys__n4798,
    ys__n4817, ys__n4818, ys__n4820, ys__n4821, ys__n4824, ys__n4825,
    ys__n4839, ys__n4840, ys__n12455, ys__n12458, ys__n12461, ys__n12464,
    ys__n12467, ys__n12470, ys__n12473, ys__n12476, ys__n12479, ys__n12482,
    ys__n12485, ys__n12488, ys__n12491, ys__n12494, ys__n12497, ys__n12500,
    ys__n12503, ys__n12506, ys__n12509, ys__n12512, ys__n12515, ys__n12518,
    ys__n12521, ys__n12524, ys__n12527, ys__n12530, ys__n12533, ys__n12536,
    ys__n12539, ys__n12542, ys__n12545, ys__n12548, ys__n16188, ys__n16191,
    ys__n16412, ys__n16415, ys__n16424, ys__n16427, ys__n16706, ys__n16709,
    ys__n16718, ys__n16721, ys__n17692, ys__n17697, ys__n17780, ys__n18007,
    ys__n18009, ys__n18015, ys__n18019, ys__n18028, ys__n18078, ys__n18080,
    ys__n18082, ys__n18087, ys__n18088, ys__n18089, ys__n18120, ys__n18125,
    ys__n18128, ys__n18131, ys__n18133, ys__n18134, ys__n18136, ys__n18137,
    ys__n18154, ys__n18165, ys__n18166, ys__n18169, ys__n18170, ys__n18174,
    ys__n18176, ys__n18178, ys__n18210, ys__n18214, ys__n18216, ys__n18217,
    ys__n18218, ys__n18223, ys__n18227, ys__n18236, ys__n18238, ys__n18239,
    ys__n18241, ys__n18251, ys__n18268, ys__n18272, ys__n18273, ys__n18278,
    ys__n18281, ys__n18284, ys__n18287, ys__n18303, ys__n18321, ys__n18329,
    ys__n18331, ys__n18333, ys__n18335, ys__n18337, ys__n18339, ys__n18341,
    ys__n18343, ys__n18345, ys__n18347, ys__n18349, ys__n18351, ys__n18353,
    ys__n18355, ys__n18357, ys__n18360, ys__n18380, ys__n18383, ys__n18386,
    ys__n18391, ys__n18392, ys__n18394, ys__n18395, ys__n18396, ys__n18397,
    ys__n18398, ys__n18399, ys__n18400, ys__n18401, ys__n18402, ys__n18403,
    ys__n18404, ys__n18405, ys__n18406, ys__n18407, ys__n18408, ys__n18409,
    ys__n18410, ys__n18411, ys__n18412, ys__n18413, ys__n18414, ys__n18415,
    ys__n18416, ys__n18417, ys__n18418, ys__n18419, ys__n18420, ys__n18421,
    ys__n18422, ys__n18423, ys__n18424, ys__n18425, ys__n18426, ys__n18427,
    ys__n18428, ys__n18429, ys__n18430, ys__n18431, ys__n18432, ys__n18433,
    ys__n18434, ys__n18435, ys__n18436, ys__n18437, ys__n18438, ys__n18439,
    ys__n18440, ys__n18441, ys__n18442, ys__n18443, ys__n18444, ys__n18445,
    ys__n18449, ys__n18450, ys__n18452, ys__n18453, ys__n18455, ys__n18456,
    ys__n18458, ys__n18459, ys__n18461, ys__n18462, ys__n18464, ys__n18465,
    ys__n18467, ys__n18468, ys__n18470, ys__n18471, ys__n18473, ys__n18474,
    ys__n18476, ys__n18477, ys__n18479, ys__n18480, ys__n18482, ys__n18483,
    ys__n18485, ys__n18486, ys__n18488, ys__n18489, ys__n18491, ys__n18492,
    ys__n18494, ys__n18495, ys__n18497, ys__n18498, ys__n18500, ys__n18501,
    ys__n18503, ys__n18504, ys__n18506, ys__n18507, ys__n18509, ys__n18510,
    ys__n18512, ys__n18513, ys__n18515, ys__n18516, ys__n18518, ys__n18519,
    ys__n18521, ys__n18522, ys__n18524, ys__n18525, ys__n18527, ys__n18528,
    ys__n18530, ys__n18531, ys__n18533, ys__n18534, ys__n18536, ys__n18537,
    ys__n18539, ys__n18540, ys__n18542, ys__n18543, ys__n18545, ys__n18547,
    ys__n18548, ys__n18549, ys__n18550, ys__n18551, ys__n18553, ys__n18554,
    ys__n18555, ys__n18557, ys__n18559, ys__n18561, ys__n18564, ys__n18567,
    ys__n18570, ys__n18573, ys__n18576, ys__n18579, ys__n18582, ys__n18585,
    ys__n18588, ys__n18591, ys__n18594, ys__n18597, ys__n18600, ys__n18603,
    ys__n18606, ys__n18609, ys__n18612, ys__n18615, ys__n18618, ys__n18621,
    ys__n18624, ys__n18627, ys__n18629, ys__n18631, ys__n18633, ys__n18635,
    ys__n18637, ys__n18640, ys__n18643, ys__n18646, ys__n18649, ys__n18652,
    ys__n18654, ys__n18655, ys__n18657, ys__n18658, ys__n18660, ys__n18661,
    ys__n18663, ys__n18664, ys__n18666, ys__n18667, ys__n18669, ys__n18670,
    ys__n18672, ys__n18673, ys__n18675, ys__n18676, ys__n18678, ys__n18679,
    ys__n18681, ys__n18682, ys__n18684, ys__n18685, ys__n18687, ys__n18688,
    ys__n18690, ys__n18691, ys__n18693, ys__n18694, ys__n18696, ys__n18697,
    ys__n18699, ys__n18700, ys__n18702, ys__n18703, ys__n18705, ys__n18706,
    ys__n18708, ys__n18709, ys__n18711, ys__n18712, ys__n18714, ys__n18715,
    ys__n18717, ys__n18718, ys__n18720, ys__n18721, ys__n18723, ys__n18724,
    ys__n18726, ys__n18727, ys__n18729, ys__n18730, ys__n18732, ys__n18733,
    ys__n18735, ys__n18736, ys__n18738, ys__n18739, ys__n18741, ys__n18742,
    ys__n18744, ys__n18745, ys__n18747, ys__n18748, ys__n18750, ys__n18751,
    ys__n18753, ys__n18754, ys__n18757, ys__n18759, ys__n18760, ys__n18763,
    ys__n18764, ys__n18766, ys__n18768, ys__n18770, ys__n18772, ys__n18774,
    ys__n18776, ys__n18778, ys__n18780, ys__n18782, ys__n18784, ys__n18786,
    ys__n18788, ys__n18790, ys__n18792, ys__n18794, ys__n18796, ys__n18798,
    ys__n18800, ys__n18802, ys__n18804, ys__n18806, ys__n18808, ys__n18810,
    ys__n18812, ys__n18814, ys__n18816, ys__n18818, ys__n18820, ys__n18822,
    ys__n18824, ys__n18826, ys__n19149, ys__n19151, ys__n19159, ys__n19173,
    ys__n19177, ys__n19178, ys__n19183, ys__n19227, ys__n19229, ys__n19231,
    ys__n19233, ys__n19235, ys__n19239, ys__n19254, ys__n19256, ys__n19257,
    ys__n19264, ys__n19266, ys__n19878, ys__n19881, ys__n19884, ys__n19887,
    ys__n19890, ys__n19893, ys__n19896, ys__n19899, ys__n19902, ys__n19905,
    ys__n19908, ys__n19911, ys__n19914, ys__n19917, ys__n19920, ys__n19923,
    ys__n19926, ys__n19929, ys__n19932, ys__n19935, ys__n19938, ys__n19941,
    ys__n19944, ys__n19947, ys__n19950, ys__n19953, ys__n19956, ys__n19959,
    ys__n19962, ys__n19965, ys__n19968, ys__n19971, ys__n20006, ys__n20007,
    ys__n20008, ys__n20009, ys__n20010, ys__n20011, ys__n20012, ys__n20013,
    ys__n20014, ys__n20015, ys__n20016, ys__n20017, ys__n20018, ys__n20019,
    ys__n20020, ys__n20021, ys__n20022, ys__n20023, ys__n20024, ys__n20025,
    ys__n20026, ys__n20027, ys__n20028, ys__n20029, ys__n20030, ys__n20031,
    ys__n20032, ys__n20033, ys__n20034, ys__n20038, ys__n20040, ys__n20043,
    ys__n20045, ys__n20053, ys__n20059, ys__n20062, ys__n20065, ys__n20068,
    ys__n20071, ys__n20074, ys__n20077, ys__n20080, ys__n20082, ys__n20084,
    ys__n20086, ys__n20088, ys__n20090, ys__n20092, ys__n20094, ys__n20096,
    ys__n20098, ys__n20100, ys__n20102, ys__n20104, ys__n20106, ys__n20108,
    ys__n20110, ys__n20112, ys__n20114, ys__n20116, ys__n20118, ys__n20120,
    ys__n20122, ys__n20124, ys__n20126, ys__n20128, ys__n22466, ys__n22919,
    ys__n22922, ys__n22925, ys__n22928, ys__n22931, ys__n22934, ys__n22937,
    ys__n22940, ys__n22943, ys__n22946, ys__n22949, ys__n22952, ys__n22955,
    ys__n22958, ys__n22961, ys__n22964, ys__n22967, ys__n22970, ys__n22973,
    ys__n22976, ys__n22979, ys__n22982, ys__n22985, ys__n22988, ys__n22991,
    ys__n22994, ys__n22997, ys__n23000, ys__n23003, ys__n23006, ys__n23009,
    ys__n23012, ys__n23263, ys__n23264, ys__n23340, ys__n23483, ys__n23485,
    ys__n23487, ys__n23489, ys__n23491, ys__n23493, ys__n23495, ys__n23497,
    ys__n23499, ys__n23501, ys__n23503, ys__n23505, ys__n23507, ys__n23509,
    ys__n23511, ys__n23513, ys__n23515, ys__n23517, ys__n23519, ys__n23521,
    ys__n23523, ys__n23525, ys__n23527, ys__n23529, ys__n23531, ys__n23533,
    ys__n23535, ys__n23537, ys__n23539, ys__n23541, ys__n23543, ys__n23635,
    ys__n23636, ys__n23764, ys__n23795, ys__n23798, ys__n23801, ys__n23804,
    ys__n23807, ys__n23853, ys__n23865, ys__n23868, ys__n23871, ys__n23874,
    ys__n23877, ys__n23921, ys__n23933, ys__n23936, ys__n23939, ys__n23942,
    ys__n23945, ys__n24099, ys__n24101, ys__n24102, ys__n24104, ys__n24105,
    ys__n24116, ys__n24118, ys__n24120, ys__n24126, ys__n24130, ys__n24134,
    ys__n24140, ys__n24145, ys__n24149, ys__n24154, ys__n24160, ys__n24162,
    ys__n24163, ys__n24165, ys__n24166, ys__n24176, ys__n24179, ys__n24180,
    ys__n24182, ys__n24183, ys__n24185, ys__n24186, ys__n24188, ys__n24189,
    ys__n24191, ys__n24192, ys__n24194, ys__n24195, ys__n24222, ys__n24227,
    ys__n24231, ys__n24236, ys__n24240, ys__n24245, ys__n24250, ys__n24255,
    ys__n24256, ys__n24258, ys__n24259, ys__n24260, ys__n24262, ys__n24265,
    ys__n24268, ys__n24271, ys__n24272, ys__n24274, ys__n24275, ys__n24277,
    ys__n24278, ys__n24286, ys__n24289, ys__n24291, ys__n24293, ys__n24295,
    ys__n24297, ys__n24299, ys__n24301, ys__n24305, ys__n24307, ys__n24309,
    ys__n24311, ys__n24313, ys__n24315, ys__n24317, ys__n24319, ys__n24320,
    ys__n24323, ys__n24325, ys__n24327, ys__n24329, ys__n24331, ys__n24333,
    ys__n24335, ys__n24339, ys__n24341, ys__n24343, ys__n24345, ys__n24347,
    ys__n24349, ys__n24351, ys__n24353, ys__n24354, ys__n24357, ys__n24359,
    ys__n24361, ys__n24363, ys__n24365, ys__n24367, ys__n24369, ys__n24373,
    ys__n24375, ys__n24377, ys__n24379, ys__n24381, ys__n24383, ys__n24385,
    ys__n24387, ys__n24388, ys__n24392, ys__n24394, ys__n24396, ys__n24398,
    ys__n24400, ys__n24402, ys__n24404, ys__n24408, ys__n24410, ys__n24412,
    ys__n24414, ys__n24416, ys__n24418, ys__n24420, ys__n24422, ys__n24425,
    ys__n24430, ys__n24436, ys__n24440, ys__n24445, ys__n24447, ys__n24466,
    ys__n24470, ys__n24488, ys__n24499, ys__n24502, ys__n24522, ys__n24532,
    ys__n24541, ys__n24552, ys__n24570, ys__n24573, ys__n24577, ys__n24579,
    ys__n24581, ys__n24585, ys__n24604, ys__n24713, ys__n24714, ys__n24742,
    ys__n24745, ys__n24748, ys__n24751, ys__n24754, ys__n24757, ys__n24760,
    ys__n24763, ys__n24766, ys__n24769, ys__n24772, ys__n24775, ys__n24778,
    ys__n24781, ys__n24784, ys__n24787, ys__n24790, ys__n24793, ys__n24796,
    ys__n24799, ys__n24802, ys__n24805, ys__n24808, ys__n24811, ys__n24814,
    ys__n24817, ys__n24820, ys__n24823, ys__n24826, ys__n24829, ys__n24832,
    ys__n24835, ys__n24837, ys__n24839, ys__n24907, ys__n24910, ys__n24913,
    ys__n24916, ys__n24919, ys__n24922, ys__n24925, ys__n24928, ys__n24931,
    ys__n24934, ys__n24937, ys__n24940, ys__n24943, ys__n24946, ys__n24949,
    ys__n24952, ys__n24955, ys__n25294, ys__n25302, ys__n25304, ys__n25306,
    ys__n25308, ys__n25310, ys__n25385, ys__n25386, ys__n25387, ys__n25388,
    ys__n25390, ys__n25406, ys__n25421, ys__n25430, ys__n25431, ys__n25432,
    ys__n25433, ys__n25434, ys__n25435, ys__n25436, ys__n25438, ys__n25441,
    ys__n25449, ys__n25456, ys__n25461, ys__n25463, ys__n25465, ys__n25467,
    ys__n25469, ys__n25472, ys__n25486, ys__n25496, ys__n25504, ys__n25519,
    ys__n25522, ys__n25534, ys__n25550, ys__n25661, ys__n25663, ys__n25665,
    ys__n25667, ys__n25669, ys__n25671, ys__n25673, ys__n25675, ys__n25677,
    ys__n25679, ys__n25681, ys__n25683, ys__n25685, ys__n25687, ys__n25689,
    ys__n25691, ys__n25693, ys__n25695, ys__n25697, ys__n25699, ys__n25701,
    ys__n25703, ys__n25705, ys__n25707, ys__n25709, ys__n25711, ys__n25713,
    ys__n25715, ys__n25717, ys__n25719, ys__n25721, ys__n25723, ys__n25725,
    ys__n25830, ys__n25833, ys__n25836, ys__n25839, ys__n25842, ys__n25844,
    ys__n25846, ys__n25852, ys__n25957, ys__n25960, ys__n25963, ys__n25966,
    ys__n26118, ys__n26119, ys__n26120, ys__n26121, ys__n26122, ys__n26123,
    ys__n26124, ys__n26125, ys__n26126, ys__n26127, ys__n26128, ys__n26129,
    ys__n26130, ys__n26131, ys__n26132, ys__n26133, ys__n26134, ys__n26135,
    ys__n26136, ys__n26137, ys__n26138, ys__n26139, ys__n26141, ys__n26144,
    ys__n26146, ys__n26148, ys__n26150, ys__n26152, ys__n26154, ys__n26156,
    ys__n26158, ys__n26160, ys__n26220, ys__n26222, ys__n26224, ys__n26226,
    ys__n26228, ys__n26230, ys__n26232, ys__n26234, ys__n26236, ys__n26238,
    ys__n26240, ys__n26242, ys__n26244, ys__n26246, ys__n26248, ys__n26250,
    ys__n26252, ys__n26254, ys__n26256, ys__n26258, ys__n26260, ys__n26262,
    ys__n26264, ys__n26266, ys__n26268, ys__n26270, ys__n26272, ys__n26274,
    ys__n26276, ys__n26278, ys__n26282, ys__n26284, ys__n26286, ys__n26288,
    ys__n26291, ys__n26293, ys__n26294, ys__n26555, ys__n26566, ys__n26573,
    ys__n26607, ys__n26609, ys__n26611, ys__n26613, ys__n26615, ys__n26617,
    ys__n26619, ys__n26621, ys__n26623, ys__n26625, ys__n26627, ys__n26629,
    ys__n26631, ys__n26633, ys__n26635, ys__n26637, ys__n26639, ys__n26641,
    ys__n26643, ys__n26645, ys__n26647, ys__n26649, ys__n26651, ys__n26653,
    ys__n26655, ys__n26657, ys__n26659, ys__n26661, ys__n26663, ys__n26665,
    ys__n26667, ys__n26669, ys__n26671, ys__n26673, ys__n26675, ys__n26677,
    ys__n26679, ys__n26681, ys__n26683, ys__n26685, ys__n26687, ys__n26689,
    ys__n26691, ys__n26693, ys__n26695, ys__n26697, ys__n26699, ys__n26701,
    ys__n26703, ys__n26705, ys__n26707, ys__n26709, ys__n26711, ys__n26713,
    ys__n26715, ys__n26717, ys__n26719, ys__n26721, ys__n26723, ys__n26725,
    ys__n26727, ys__n26729, ys__n26731, ys__n26733, ys__n26734, ys__n26735,
    ys__n26736, ys__n26737, ys__n26738, ys__n26739, ys__n26740, ys__n26741,
    ys__n26742, ys__n26743, ys__n26744, ys__n26745, ys__n26746, ys__n26747,
    ys__n26748, ys__n26749, ys__n26750, ys__n26751, ys__n26752, ys__n26753,
    ys__n26754, ys__n26755, ys__n26756, ys__n26757, ys__n26758, ys__n26759,
    ys__n26760, ys__n26761, ys__n26762, ys__n26763, ys__n26764, ys__n26765,
    ys__n26802, ys__n26803, ys__n26804, ys__n26805, ys__n26806, ys__n26807,
    ys__n26808, ys__n26809, ys__n26810, ys__n26811, ys__n26812, ys__n26813,
    ys__n26814, ys__n26815, ys__n26816, ys__n26817, ys__n26818, ys__n26819,
    ys__n26820, ys__n26821, ys__n26822, ys__n26823, ys__n26824, ys__n26825,
    ys__n26826, ys__n26827, ys__n26828, ys__n26829, ys__n26830, ys__n26831,
    ys__n26832, ys__n26833, ys__n26834, ys__n26835, ys__n26836, ys__n26837,
    ys__n26838, ys__n26839, ys__n26840, ys__n26841, ys__n26842, ys__n26843,
    ys__n26844, ys__n26845, ys__n26846, ys__n26847, ys__n26848, ys__n26849,
    ys__n26850, ys__n26851, ys__n26852, ys__n26853, ys__n26854, ys__n26855,
    ys__n26856, ys__n26857, ys__n26858, ys__n26859, ys__n26860, ys__n26861,
    ys__n26862, ys__n26863, ys__n26864, ys__n26865, ys__n26866, ys__n26867,
    ys__n26868, ys__n26869, ys__n26870, ys__n26871, ys__n26872, ys__n26873,
    ys__n26874, ys__n26875, ys__n26876, ys__n26877, ys__n26878, ys__n26879,
    ys__n26880, ys__n26881, ys__n26882, ys__n26883, ys__n26884, ys__n26885,
    ys__n26886, ys__n26887, ys__n26888, ys__n26889, ys__n26890, ys__n26891,
    ys__n26892, ys__n26893, ys__n26894, ys__n26895, ys__n26896, ys__n26897,
    ys__n26898, ys__n26899, ys__n26900, ys__n26901, ys__n26902, ys__n26903,
    ys__n26904, ys__n26905, ys__n26906, ys__n26907, ys__n26908, ys__n26909,
    ys__n26910, ys__n26911, ys__n26912, ys__n26913, ys__n26914, ys__n26915,
    ys__n26916, ys__n26917, ys__n26918, ys__n26919, ys__n26920, ys__n26921,
    ys__n26922, ys__n26923, ys__n26924, ys__n26925, ys__n26926, ys__n26927,
    ys__n26928, ys__n26929, ys__n26930, ys__n26931, ys__n26932, ys__n26933,
    ys__n26934, ys__n26935, ys__n26936, ys__n26937, ys__n26938, ys__n26939,
    ys__n26940, ys__n26941, ys__n26942, ys__n26943, ys__n26944, ys__n26945,
    ys__n26946, ys__n26947, ys__n26948, ys__n26949, ys__n26950, ys__n26951,
    ys__n26952, ys__n26953, ys__n26954, ys__n26955, ys__n26956, ys__n26957,
    ys__n26958, ys__n26959, ys__n26960, ys__n26961, ys__n26962, ys__n26963,
    ys__n26964, ys__n26965, ys__n26966, ys__n26967, ys__n26968, ys__n26969,
    ys__n26970, ys__n26971, ys__n26972, ys__n26973, ys__n26974, ys__n26975,
    ys__n26976, ys__n26977, ys__n26978, ys__n26979, ys__n26980, ys__n26981,
    ys__n26982, ys__n26983, ys__n26984, ys__n26985, ys__n26986, ys__n26987,
    ys__n26988, ys__n26989, ys__n26990, ys__n26991, ys__n26992, ys__n26993,
    ys__n26994, ys__n26995, ys__n26996, ys__n26997, ys__n26998, ys__n26999,
    ys__n27000, ys__n27001, ys__n27002, ys__n27003, ys__n27004, ys__n27005,
    ys__n27006, ys__n27007, ys__n27008, ys__n27009, ys__n27010, ys__n27011,
    ys__n27012, ys__n27013, ys__n27014, ys__n27015, ys__n27016, ys__n27017,
    ys__n27018, ys__n27019, ys__n27020, ys__n27021, ys__n27022, ys__n27023,
    ys__n27024, ys__n27025, ys__n27026, ys__n27027, ys__n27028, ys__n27029,
    ys__n27030, ys__n27031, ys__n27032, ys__n27033, ys__n27034, ys__n27035,
    ys__n27036, ys__n27037, ys__n27038, ys__n27039, ys__n27040, ys__n27041,
    ys__n27042, ys__n27043, ys__n27044, ys__n27045, ys__n27046, ys__n27047,
    ys__n27048, ys__n27049, ys__n27050, ys__n27051, ys__n27052, ys__n27053,
    ys__n27054, ys__n27055, ys__n27056, ys__n27057, ys__n27058, ys__n27059,
    ys__n27060, ys__n27061, ys__n27062, ys__n27063, ys__n27064, ys__n27065,
    ys__n27066, ys__n27067, ys__n27068, ys__n27069, ys__n27070, ys__n27071,
    ys__n27072, ys__n27073, ys__n27074, ys__n27075, ys__n27076, ys__n27077,
    ys__n27078, ys__n27079, ys__n27080, ys__n27081, ys__n27082, ys__n27083,
    ys__n27084, ys__n27085, ys__n27086, ys__n27087, ys__n27088, ys__n27089,
    ys__n27090, ys__n27091, ys__n27092, ys__n27093, ys__n27094, ys__n27095,
    ys__n27096, ys__n27097, ys__n27098, ys__n27099, ys__n27100, ys__n27101,
    ys__n27102, ys__n27103, ys__n27104, ys__n27105, ys__n27106, ys__n27107,
    ys__n27108, ys__n27109, ys__n27110, ys__n27111, ys__n27112, ys__n27113,
    ys__n27114, ys__n27115, ys__n27116, ys__n27117, ys__n27118, ys__n27119,
    ys__n27120, ys__n27121, ys__n27122, ys__n27123, ys__n27124, ys__n27125,
    ys__n27126, ys__n27127, ys__n27128, ys__n27129, ys__n27130, ys__n27131,
    ys__n27132, ys__n27133, ys__n27134, ys__n27135, ys__n27136, ys__n27137,
    ys__n27138, ys__n27139, ys__n27140, ys__n27141, ys__n27142, ys__n27143,
    ys__n27144, ys__n27145, ys__n27146, ys__n27147, ys__n27148, ys__n27149,
    ys__n27150, ys__n27151, ys__n27152, ys__n27153, ys__n27154, ys__n27155,
    ys__n27156, ys__n27157, ys__n27158, ys__n27159, ys__n27160, ys__n27161,
    ys__n27162, ys__n27163, ys__n27164, ys__n27165, ys__n27166, ys__n27167,
    ys__n27168, ys__n27169, ys__n27170, ys__n27171, ys__n27172, ys__n27173,
    ys__n27174, ys__n27175, ys__n27176, ys__n27177, ys__n27178, ys__n27179,
    ys__n27180, ys__n27181, ys__n27182, ys__n27183, ys__n27184, ys__n27185,
    ys__n27186, ys__n27187, ys__n27188, ys__n27189, ys__n27190, ys__n27191,
    ys__n27192, ys__n27193, ys__n27194, ys__n27195, ys__n27196, ys__n27197,
    ys__n27198, ys__n27199, ys__n27200, ys__n27201, ys__n27202, ys__n27203,
    ys__n27204, ys__n27205, ys__n27206, ys__n27207, ys__n27208, ys__n27209,
    ys__n27210, ys__n27211, ys__n27212, ys__n27213, ys__n27214, ys__n27215,
    ys__n27216, ys__n27217, ys__n27218, ys__n27219, ys__n27220, ys__n27221,
    ys__n27222, ys__n27223, ys__n27224, ys__n27225, ys__n27226, ys__n27227,
    ys__n27228, ys__n27229, ys__n27230, ys__n27231, ys__n27232, ys__n27233,
    ys__n27234, ys__n27235, ys__n27236, ys__n27237, ys__n27238, ys__n27239,
    ys__n27240, ys__n27241, ys__n27242, ys__n27243, ys__n27244, ys__n27245,
    ys__n27246, ys__n27247, ys__n27248, ys__n27249, ys__n27250, ys__n27251,
    ys__n27252, ys__n27253, ys__n27254, ys__n27255, ys__n27256, ys__n27257,
    ys__n27258, ys__n27259, ys__n27260, ys__n27261, ys__n27262, ys__n27263,
    ys__n27264, ys__n27265, ys__n27266, ys__n27267, ys__n27268, ys__n27269,
    ys__n27270, ys__n27271, ys__n27272, ys__n27273, ys__n27274, ys__n27275,
    ys__n27276, ys__n27277, ys__n27278, ys__n27279, ys__n27280, ys__n27281,
    ys__n27282, ys__n27283, ys__n27284, ys__n27285, ys__n27286, ys__n27287,
    ys__n27288, ys__n27289, ys__n27290, ys__n27291, ys__n27292, ys__n27293,
    ys__n27294, ys__n27295, ys__n27296, ys__n27297, ys__n27298, ys__n27299,
    ys__n27300, ys__n27301, ys__n27302, ys__n27303, ys__n27304, ys__n27305,
    ys__n27306, ys__n27307, ys__n27308, ys__n27309, ys__n27310, ys__n27311,
    ys__n27312, ys__n27313, ys__n27314, ys__n27315, ys__n27316, ys__n27317,
    ys__n27318, ys__n27319, ys__n27320, ys__n27321, ys__n27322, ys__n27323,
    ys__n27324, ys__n27325, ys__n27326, ys__n27327, ys__n27328, ys__n27329,
    ys__n27330, ys__n27331, ys__n27332, ys__n27333, ys__n27334, ys__n27335,
    ys__n27336, ys__n27337, ys__n27338, ys__n27339, ys__n27340, ys__n27341,
    ys__n27342, ys__n27343, ys__n27344, ys__n27345, ys__n27346, ys__n27347,
    ys__n27348, ys__n27349, ys__n27350, ys__n27351, ys__n27352, ys__n27353,
    ys__n27354, ys__n27355, ys__n27356, ys__n27357, ys__n27358, ys__n27359,
    ys__n27360, ys__n27361, ys__n27362, ys__n27363, ys__n27364, ys__n27365,
    ys__n27366, ys__n27367, ys__n27368, ys__n27369, ys__n27370, ys__n27371,
    ys__n27372, ys__n27373, ys__n27374, ys__n27375, ys__n27376, ys__n27377,
    ys__n27378, ys__n27379, ys__n27380, ys__n27381, ys__n27382, ys__n27383,
    ys__n27384, ys__n27385, ys__n27386, ys__n27387, ys__n27388, ys__n27389,
    ys__n27390, ys__n27391, ys__n27392, ys__n27393, ys__n27394, ys__n27395,
    ys__n27396, ys__n27397, ys__n27398, ys__n27399, ys__n27400, ys__n27401,
    ys__n27402, ys__n27403, ys__n27404, ys__n27405, ys__n27406, ys__n27407,
    ys__n27408, ys__n27409, ys__n27410, ys__n27411, ys__n27412, ys__n27413,
    ys__n27414, ys__n27415, ys__n27416, ys__n27417, ys__n27418, ys__n27419,
    ys__n27420, ys__n27421, ys__n27422, ys__n27423, ys__n27424, ys__n27425,
    ys__n27426, ys__n27427, ys__n27428, ys__n27429, ys__n27430, ys__n27431,
    ys__n27432, ys__n27433, ys__n27434, ys__n27435, ys__n27436, ys__n27437,
    ys__n27484, ys__n27493, ys__n27504, ys__n27513, ys__n27515, ys__n27517,
    ys__n27550, ys__n27551, ys__n27598, ys__n27603, ys__n27605, ys__n27610,
    ys__n27613, ys__n27616, ys__n27619, ys__n27622, ys__n27625, ys__n27628,
    ys__n27631, ys__n27634, ys__n27637, ys__n27640, ys__n27643, ys__n27646,
    ys__n27649, ys__n27652, ys__n27655, ys__n27658, ys__n27661, ys__n27664,
    ys__n27667, ys__n27670, ys__n27673, ys__n27676, ys__n27679, ys__n27682,
    ys__n27685, ys__n27688, ys__n27691, ys__n27694, ys__n27697, ys__n27700,
    ys__n27703, ys__n27705, ys__n27706, ys__n27707, ys__n27708, ys__n27709,
    ys__n27710, ys__n27711, ys__n27712, ys__n27713, ys__n27714, ys__n27715,
    ys__n27716, ys__n27717, ys__n27718, ys__n27719, ys__n27720, ys__n27721,
    ys__n27722, ys__n27723, ys__n27724, ys__n27725, ys__n27726, ys__n27727,
    ys__n27728, ys__n27729, ys__n27730, ys__n27731, ys__n27732, ys__n27733,
    ys__n27734, ys__n27735, ys__n27736, ys__n27739, ys__n27741, ys__n28247,
    ys__n28249, ys__n28250, ys__n28251, ys__n28252, ys__n28254, ys__n28256,
    ys__n28258, ys__n28259, ys__n28261, ys__n28263, ys__n28265, ys__n28266,
    ys__n28268, ys__n28269, ys__n28270, ys__n28271, ys__n28272, ys__n28274,
    ys__n28276, ys__n28328, ys__n28330, ys__n28332, ys__n28334, ys__n28336,
    ys__n28343, ys__n28345, ys__n28347, ys__n28349, ys__n28351, ys__n28353,
    ys__n28355, ys__n28357, ys__n28359, ys__n28361, ys__n28363, ys__n28365,
    ys__n28367, ys__n28369, ys__n28371, ys__n28373, ys__n28375, ys__n28377,
    ys__n28379, ys__n28381, ys__n28383, ys__n28385, ys__n28387, ys__n28389,
    ys__n28391, ys__n28393, ys__n28395, ys__n28397, ys__n28399, ys__n28401,
    ys__n28403, ys__n28406, ys__n28409, ys__n28410, ys__n28411, ys__n28412,
    ys__n28413, ys__n28414, ys__n28415, ys__n28416, ys__n28417, ys__n28418,
    ys__n28419, ys__n28420, ys__n28421, ys__n28422, ys__n28423, ys__n28425,
    ys__n28427, ys__n28429, ys__n28431, ys__n28433, ys__n28435, ys__n28437,
    ys__n28439, ys__n28440, ys__n28441, ys__n28442, ys__n28443, ys__n28444,
    ys__n28445, ys__n28447, ys__n28448, ys__n28449, ys__n28450, ys__n28451,
    ys__n28452, ys__n28454, ys__n28456, ys__n28458, ys__n28460, ys__n28475,
    ys__n28476, ys__n28477, ys__n28478, ys__n28479, ys__n28480, ys__n28481,
    ys__n28482, ys__n28483, ys__n28484, ys__n28485, ys__n28486, ys__n28487,
    ys__n28488, ys__n28489, ys__n28490, ys__n28491, ys__n28492, ys__n28493,
    ys__n28494, ys__n28495, ys__n28496, ys__n28497, ys__n28498, ys__n28499,
    ys__n28500, ys__n28501, ys__n28502, ys__n28503, ys__n28504, ys__n28505,
    ys__n28506, ys__n28510, ys__n28513, ys__n28518, ys__n28533, ys__n28536,
    ys__n28539, ys__n28542, ys__n28545, ys__n28548, ys__n28551, ys__n28554,
    ys__n28557, ys__n28560, ys__n28563, ys__n28566, ys__n28569, ys__n28572,
    ys__n28575, ys__n28578, ys__n28581, ys__n28584, ys__n28587, ys__n28661,
    ys__n28662, ys__n28781, ys__n28782, ys__n28783, ys__n28784, ys__n28785,
    ys__n28786, ys__n28787, ys__n28788, ys__n28789, ys__n28790, ys__n28791,
    ys__n28792, ys__n28793, ys__n28794, ys__n28796, ys__n28798, ys__n28800,
    ys__n28802, ys__n28804, ys__n28806, ys__n28808, ys__n28810, ys__n28812,
    ys__n28814, ys__n28816, ys__n28818, ys__n28820, ys__n28822, ys__n28824,
    ys__n28826, ys__n28828, ys__n28830, ys__n28832, ys__n28834, ys__n28836,
    ys__n28838, ys__n28840, ys__n28842, ys__n28844, ys__n28846, ys__n28848,
    ys__n28850, ys__n28852, ys__n28854, ys__n28856, ys__n28858, ys__n29022,
    ys__n29025, ys__n29028, ys__n29031, ys__n29034, ys__n29037, ys__n29040,
    ys__n29043, ys__n29046, ys__n29049, ys__n29052, ys__n29055, ys__n29058,
    ys__n29061, ys__n29064, ys__n29067, ys__n29070, ys__n29073, ys__n29076,
    ys__n29079, ys__n29082, ys__n29085, ys__n29088, ys__n29091, ys__n29094,
    ys__n29097, ys__n29100, ys__n29103, ys__n29106, ys__n29109, ys__n29112,
    ys__n29115, ys__n29118, ys__n29122, ys__n29125, ys__n29128, ys__n29131,
    ys__n29134, ys__n29137, ys__n29140, ys__n29143, ys__n29146, ys__n29149,
    ys__n29152, ys__n29155, ys__n29158, ys__n29161, ys__n29164, ys__n29167,
    ys__n29170, ys__n29173, ys__n29176, ys__n29179, ys__n29182, ys__n29185,
    ys__n29188, ys__n29191, ys__n29194, ys__n29197, ys__n29200, ys__n29203,
    ys__n29206, ys__n29209, ys__n29212, ys__n29215, ys__n29217, ys__n29219,
    ys__n29221, ys__n29223, ys__n29225, ys__n29226, ys__n29227, ys__n29228,
    ys__n29229, ys__n29230, ys__n29231, ys__n29232, ys__n29233, ys__n29234,
    ys__n29235, ys__n29336, ys__n29339, ys__n29342, ys__n29345, ys__n29348,
    ys__n29351, ys__n29354, ys__n29357, ys__n29360, ys__n29363, ys__n29366,
    ys__n29369, ys__n29372, ys__n29375, ys__n29378, ys__n29381, ys__n29384,
    ys__n29387, ys__n29390, ys__n29393, ys__n29396, ys__n29399, ys__n29402,
    ys__n29405, ys__n29408, ys__n29411, ys__n29414, ys__n29417, ys__n29420,
    ys__n29423, ys__n29426, ys__n29429, ys__n29431, ys__n29435, ys__n29438,
    ys__n29441, ys__n29444, ys__n29447, ys__n29450, ys__n29453, ys__n29456,
    ys__n29459, ys__n29462, ys__n29465, ys__n29468, ys__n29471, ys__n29474,
    ys__n29477, ys__n29480, ys__n29483, ys__n29486, ys__n29489, ys__n29492,
    ys__n29495, ys__n29498, ys__n29501, ys__n29504, ys__n29507, ys__n29510,
    ys__n29513, ys__n29516, ys__n29519, ys__n29522, ys__n29525, ys__n29528,
    ys__n29530, ys__n29532, ys__n29534, ys__n29536, ys__n29538, ys__n29539,
    ys__n29540, ys__n29541, ys__n29542, ys__n29543, ys__n29544, ys__n29545,
    ys__n29546, ys__n29547, ys__n29548, ys__n29611, ys__n29614, ys__n29617,
    ys__n29620, ys__n29623, ys__n29626, ys__n29629, ys__n29632, ys__n29635,
    ys__n29638, ys__n29641, ys__n29644, ys__n29647, ys__n29650, ys__n29653,
    ys__n29656, ys__n29659, ys__n29662, ys__n29665, ys__n29668, ys__n29671,
    ys__n29674, ys__n29677, ys__n29680, ys__n29683, ys__n29686, ys__n29689,
    ys__n29692, ys__n29695, ys__n29698, ys__n29701, ys__n29704, ys__n29706,
    ys__n29710, ys__n29713, ys__n29716, ys__n29719, ys__n29722, ys__n29725,
    ys__n29728, ys__n29731, ys__n29734, ys__n29737, ys__n29740, ys__n29743,
    ys__n29746, ys__n29749, ys__n29752, ys__n29755, ys__n29758, ys__n29761,
    ys__n29764, ys__n29767, ys__n29770, ys__n29773, ys__n29776, ys__n29779,
    ys__n29782, ys__n29785, ys__n29788, ys__n29791, ys__n29794, ys__n29797,
    ys__n29800, ys__n29803, ys__n29805, ys__n29807, ys__n29809, ys__n29811,
    ys__n29813, ys__n29814, ys__n29815, ys__n29816, ys__n29817, ys__n29818,
    ys__n29819, ys__n29820, ys__n29821, ys__n29822, ys__n29823, ys__n29847,
    ys__n30010, ys__n30080, ys__n30081, ys__n30082, ys__n30083, ys__n30084,
    ys__n30085, ys__n30086, ys__n30087, ys__n30089, ys__n30090, ys__n30091,
    ys__n30092, ys__n30093, ys__n30094, ys__n30095, ys__n30096, ys__n30098,
    ys__n30099, ys__n30100, ys__n30101, ys__n30102, ys__n30103, ys__n30104,
    ys__n30105, ys__n30106, ys__n30107, ys__n30108, ys__n30109, ys__n30110,
    ys__n30111, ys__n30112, ys__n30113, ys__n30119, ys__n30122, ys__n30125,
    ys__n30128, ys__n30131, ys__n30134, ys__n30137, ys__n30140, ys__n30143,
    ys__n30146, ys__n30149, ys__n30152, ys__n30155, ys__n30158, ys__n30161,
    ys__n30164, ys__n30167, ys__n30170, ys__n30173, ys__n30176, ys__n30179,
    ys__n30182, ys__n30185, ys__n30188, ys__n30191, ys__n30194, ys__n30197,
    ys__n30200, ys__n30203, ys__n30206, ys__n30209, ys__n30212, ys__n30215,
    ys__n30223, ys__n30226, ys__n30235, ys__n30238, ys__n30241, ys__n30244,
    ys__n30247, ys__n30250, ys__n30253, ys__n30256, ys__n30259, ys__n30262,
    ys__n30265, ys__n30268, ys__n30271, ys__n30274, ys__n30277, ys__n30280,
    ys__n30283, ys__n30286, ys__n30289, ys__n30292, ys__n30295, ys__n30298,
    ys__n30301, ys__n30304, ys__n30307, ys__n30310, ys__n30313, ys__n30316,
    ys__n30319, ys__n30322, ys__n30325, ys__n30328, ys__n30330, ys__n30331,
    ys__n30616, ys__n30619, ys__n30622, ys__n30625, ys__n30628, ys__n30631,
    ys__n30634, ys__n30637, ys__n30640, ys__n30643, ys__n30646, ys__n30649,
    ys__n30652, ys__n30655, ys__n30658, ys__n30661, ys__n30664, ys__n30667,
    ys__n30668, ys__n30670, ys__n30797, ys__n30798, ys__n30799, ys__n30800,
    ys__n30801, ys__n30802, ys__n30803, ys__n30804, ys__n30805, ys__n30806,
    ys__n30807, ys__n30808, ys__n30809, ys__n30810, ys__n30811, ys__n30812,
    ys__n30813, ys__n30832, ys__n30833, ys__n30835, ys__n30836, ys__n30856,
    ys__n30858, ys__n30860, ys__n30864, ys__n30873, ys__n30874, ys__n30875,
    ys__n30876, ys__n30942, ys__n30943, ys__n30944, ys__n30945, ys__n30946,
    ys__n30947, ys__n30948, ys__n30949, ys__n30950, ys__n30951, ys__n30952,
    ys__n30953, ys__n30954, ys__n30955, ys__n30956, ys__n31202, ys__n31203,
    ys__n31207, ys__n31208, ys__n31209, ys__n31210, ys__n31211, ys__n31212,
    ys__n31213, ys__n31214, ys__n31215, ys__n31216, ys__n31217, ys__n31218,
    ys__n31219, ys__n31220, ys__n31221, ys__n31222, ys__n31223, ys__n31224,
    ys__n31225, ys__n31226, ys__n31227, ys__n31228, ys__n31229, ys__n31230,
    ys__n31231, ys__n31232, ys__n31233, ys__n31234, ys__n31235, ys__n31236,
    ys__n31237, ys__n31238, ys__n31326, ys__n31327, ys__n31328, ys__n31329,
    ys__n31330, ys__n31331, ys__n31332, ys__n31333, ys__n31334, ys__n31335,
    ys__n31336, ys__n31337, ys__n31338, ys__n31339, ys__n31340, ys__n31341,
    ys__n31342, ys__n31343, ys__n31344, ys__n31345, ys__n31346, ys__n31347,
    ys__n31348, ys__n31349, ys__n31350, ys__n31351, ys__n31352, ys__n31353,
    ys__n31354, ys__n31355, ys__n31356, ys__n31357, ys__n31358, ys__n31359,
    ys__n31360, ys__n31361, ys__n31362, ys__n31363, ys__n31364, ys__n31365,
    ys__n31366, ys__n31367, ys__n31368, ys__n31369, ys__n31370, ys__n31371,
    ys__n31372, ys__n31373, ys__n31374, ys__n31375, ys__n31376, ys__n31377,
    ys__n31378, ys__n31379, ys__n31380, ys__n31381, ys__n31382, ys__n31383,
    ys__n31384, ys__n31385, ys__n31386, ys__n31387, ys__n31388, ys__n31389,
    ys__n31390, ys__n31391, ys__n31392, ys__n31393, ys__n31394, ys__n31395,
    ys__n31397, ys__n31398, ys__n31399, ys__n31400, ys__n31401, ys__n31402,
    ys__n31403, ys__n31404, ys__n31405, ys__n31406, ys__n31407, ys__n31408,
    ys__n31409, ys__n31410, ys__n31411, ys__n31412, ys__n31413, ys__n31414,
    ys__n31415, ys__n31416, ys__n31417, ys__n31418, ys__n31419, ys__n31420,
    ys__n31421, ys__n31422, ys__n31423, ys__n31424, ys__n31425, ys__n31426,
    ys__n31427, ys__n31428, ys__n31429, ys__n31430, ys__n31431, ys__n31432,
    ys__n31433, ys__n31434, ys__n31435, ys__n31436, ys__n31437, ys__n31438,
    ys__n31439, ys__n31440, ys__n31441, ys__n31442, ys__n31443, ys__n31444,
    ys__n31445, ys__n31446, ys__n31447, ys__n31448, ys__n31449, ys__n31450,
    ys__n31451, ys__n31452, ys__n31453, ys__n31454, ys__n31455, ys__n31456,
    ys__n31457, ys__n31458, ys__n31459, ys__n31460, ys__n31461, ys__n31462,
    ys__n31463, ys__n31464, ys__n31465, ys__n31466, ys__n31467, ys__n31468,
    ys__n31469, ys__n31470, ys__n31471, ys__n31472, ys__n31473, ys__n31474,
    ys__n31475, ys__n31476, ys__n31477, ys__n31478, ys__n31479, ys__n31480,
    ys__n31481, ys__n31482, ys__n31483, ys__n31484, ys__n31485, ys__n31486,
    ys__n31487, ys__n31488, ys__n31489, ys__n31490, ys__n31491, ys__n31492,
    ys__n31493, ys__n31494, ys__n31495, ys__n31496, ys__n31497, ys__n31498,
    ys__n31499, ys__n31500, ys__n31501, ys__n31502, ys__n31503, ys__n31504,
    ys__n31505, ys__n31506, ys__n31507, ys__n31508, ys__n31509, ys__n31510,
    ys__n31511, ys__n31512, ys__n31513, ys__n31514, ys__n31515, ys__n31516,
    ys__n31517, ys__n31518, ys__n31519, ys__n31520, ys__n31521, ys__n31522,
    ys__n31523, ys__n31524, ys__n31525, ys__n31526, ys__n31527, ys__n31528,
    ys__n31529, ys__n31530, ys__n31531, ys__n31532, ys__n31533, ys__n31534,
    ys__n31535, ys__n31536, ys__n31537, ys__n31538, ys__n31539, ys__n31540,
    ys__n31541, ys__n31542, ys__n31543, ys__n31544, ys__n31559, ys__n31560,
    ys__n31562, ys__n31564, ys__n31567, ys__n31571, ys__n31740, ys__n31741,
    ys__n31742, ys__n31743, ys__n31744, ys__n31745, ys__n31746, ys__n31747,
    ys__n31748, ys__n31749, ys__n31750, ys__n31751, ys__n31752, ys__n31753,
    ys__n31754, ys__n31755, ys__n31756, ys__n31757, ys__n31758, ys__n31759,
    ys__n31760, ys__n31761, ys__n31762, ys__n31763, ys__n31764, ys__n31765,
    ys__n31766, ys__n31767, ys__n31768, ys__n31769, ys__n31770, ys__n31771,
    ys__n31772, ys__n31773, ys__n31774, ys__n31775, ys__n31776, ys__n31777,
    ys__n31778, ys__n31779, ys__n31780, ys__n31781, ys__n31782, ys__n31783,
    ys__n31784, ys__n31785, ys__n31786, ys__n31787, ys__n31788, ys__n31789,
    ys__n31790, ys__n31791, ys__n31792, ys__n31793, ys__n31794, ys__n31795,
    ys__n31796, ys__n31797, ys__n31798, ys__n31799, ys__n31800, ys__n31801,
    ys__n31802, ys__n31803, ys__n31804, ys__n31805, ys__n31806, ys__n31807,
    ys__n31808, ys__n31809, ys__n31810, ys__n31811, ys__n31812, ys__n31813,
    ys__n31814, ys__n31815, ys__n31816, ys__n31817, ys__n31818, ys__n31819,
    ys__n31820, ys__n31821, ys__n31822, ys__n31823, ys__n31824, ys__n31825,
    ys__n31826, ys__n31827, ys__n31828, ys__n31829, ys__n31830, ys__n31831,
    ys__n31832, ys__n31833, ys__n31834, ys__n31835, ys__n31836, ys__n31837,
    ys__n31838, ys__n31839, ys__n31840, ys__n31841, ys__n31842, ys__n31843,
    ys__n31844, ys__n31845, ys__n31846, ys__n31847, ys__n31848, ys__n31849,
    ys__n31850, ys__n31851, ys__n31852, ys__n31853, ys__n31854, ys__n31855,
    ys__n31856, ys__n31857, ys__n31858, ys__n31859, ys__n31860, ys__n31861,
    ys__n31862, ys__n31863, ys__n31864, ys__n31865, ys__n31866, ys__n31867,
    ys__n31868, ys__n31869, ys__n31870, ys__n31871, ys__n31872, ys__n31873,
    ys__n31874, ys__n31875, ys__n31876, ys__n31877, ys__n31878, ys__n31879,
    ys__n31880, ys__n31881, ys__n31882, ys__n31883, ys__n31884, ys__n31885,
    ys__n31886, ys__n31887, ys__n31888, ys__n31889, ys__n31890, ys__n31891,
    ys__n31892, ys__n31893, ys__n31894, ys__n31895, ys__n31896, ys__n31897,
    ys__n31898, ys__n31899, ys__n31900, ys__n31901, ys__n31902, ys__n31903,
    ys__n31904, ys__n31905, ys__n31906, ys__n31907, ys__n31908, ys__n31909,
    ys__n31910, ys__n31911, ys__n31912, ys__n31913, ys__n31914, ys__n31915,
    ys__n31916, ys__n31917, ys__n31918, ys__n31919, ys__n31920, ys__n31921,
    ys__n31922, ys__n31923, ys__n31924, ys__n31925, ys__n31926, ys__n31927,
    ys__n31928, ys__n31929, ys__n31930, ys__n31931, ys__n31932, ys__n31933,
    ys__n31934, ys__n31935, ys__n31936, ys__n31937, ys__n31938, ys__n31939,
    ys__n31940, ys__n31941, ys__n31942, ys__n31943, ys__n31944, ys__n31945,
    ys__n31946, ys__n31947, ys__n31948, ys__n31949, ys__n31950, ys__n31953,
    ys__n31954, ys__n31955, ys__n31965, ys__n31971, ys__n31973, ys__n31975,
    ys__n31976, ys__n31978, ys__n31979, ys__n31984, ys__n31986, ys__n31988,
    ys__n31990, ys__n31992, ys__n31994, ys__n31996, ys__n31998, ys__n32000,
    ys__n32002, ys__n32004, ys__n32006, ys__n32007, ys__n32008, ys__n32010,
    ys__n32012, ys__n32014, ys__n32016, ys__n32018, ys__n32022, ys__n32023,
    ys__n32024, ys__n32025, ys__n32026, ys__n32027, ys__n32028, ys__n32029,
    ys__n32030, ys__n32031, ys__n32032, ys__n32033, ys__n32034, ys__n32035,
    ys__n32036, ys__n32037, ys__n32038, ys__n32039, ys__n32040, ys__n32041,
    ys__n32042, ys__n32043, ys__n32044, ys__n32045, ys__n32046, ys__n32047,
    ys__n32048, ys__n32049, ys__n32050, ys__n32051, ys__n32052, ys__n32053,
    ys__n32054, ys__n32055, ys__n32056, ys__n32057, ys__n32058, ys__n32059,
    ys__n32060, ys__n32061, ys__n32062, ys__n32063, ys__n32064, ys__n32065,
    ys__n32066, ys__n32067, ys__n32068, ys__n32069, ys__n32070, ys__n32071,
    ys__n32072, ys__n32073, ys__n32074, ys__n32075, ys__n32076, ys__n32077,
    ys__n32078, ys__n32079, ys__n32080, ys__n32081, ys__n32082, ys__n32083,
    ys__n32084, ys__n32085, ys__n32086, ys__n32087, ys__n32088, ys__n32124,
    ys__n32125, ys__n32126, ys__n32127, ys__n32128, ys__n32129, ys__n32130,
    ys__n32131, ys__n32132, ys__n32133, ys__n32134, ys__n32135, ys__n32136,
    ys__n32137, ys__n32138, ys__n32139, ys__n32140, ys__n32141, ys__n32142,
    ys__n32143, ys__n32144, ys__n32145, ys__n32146, ys__n32147, ys__n32148,
    ys__n32149, ys__n32150, ys__n32151, ys__n32152, ys__n32153, ys__n32154,
    ys__n32155, ys__n32158, ys__n32159, ys__n32160, ys__n32161, ys__n32162,
    ys__n32163, ys__n32164, ys__n32165, ys__n32166, ys__n32167, ys__n32168,
    ys__n32169, ys__n32170, ys__n32171, ys__n32172, ys__n32173, ys__n32174,
    ys__n32175, ys__n32176, ys__n32177, ys__n32178, ys__n32179, ys__n32180,
    ys__n32181, ys__n32182, ys__n32183, ys__n32184, ys__n32185, ys__n32186,
    ys__n32187, ys__n32188, ys__n32189, ys__n32190, ys__n32191, ys__n32192,
    ys__n32193, ys__n32194, ys__n32195, ys__n32196, ys__n32197, ys__n32198,
    ys__n32199, ys__n32200, ys__n32201, ys__n32202, ys__n32203, ys__n32204,
    ys__n32205, ys__n32206, ys__n32207, ys__n32208, ys__n32209, ys__n32210,
    ys__n32211, ys__n32212, ys__n32213, ys__n32214, ys__n32215, ys__n32216,
    ys__n32217, ys__n32218, ys__n32219, ys__n32220, ys__n32221, ys__n32222,
    ys__n32223, ys__n32224, ys__n32225, ys__n32226, ys__n32227, ys__n32228,
    ys__n32229, ys__n32230, ys__n32231, ys__n32232, ys__n32233, ys__n32234,
    ys__n32235, ys__n32236, ys__n32237, ys__n32238, ys__n32239, ys__n32240,
    ys__n32241, ys__n32242, ys__n32243, ys__n32244, ys__n32245, ys__n32246,
    ys__n32247, ys__n32248, ys__n32249, ys__n32250, ys__n32251, ys__n32252,
    ys__n32253, ys__n32254, ys__n32255, ys__n32256, ys__n32257, ys__n32258,
    ys__n32259, ys__n32260, ys__n32261, ys__n32262, ys__n32263, ys__n32264,
    ys__n32265, ys__n32266, ys__n32267, ys__n32268, ys__n32269, ys__n32270,
    ys__n32271, ys__n32272, ys__n32273, ys__n32274, ys__n32275, ys__n32276,
    ys__n32277, ys__n32278, ys__n32279, ys__n32280, ys__n32281, ys__n32282,
    ys__n32283, ys__n32284, ys__n32285, ys__n32286, ys__n32287, ys__n32288,
    ys__n32289, ys__n32290, ys__n32291, ys__n32292, ys__n32293, ys__n32294,
    ys__n32295, ys__n32296, ys__n32297, ys__n32298, ys__n32299, ys__n32300,
    ys__n32301, ys__n32302, ys__n32303, ys__n32304, ys__n32305, ys__n32306,
    ys__n32307, ys__n32308, ys__n32309, ys__n32310, ys__n32311, ys__n32312,
    ys__n32313, ys__n32314, ys__n32315, ys__n32316, ys__n32317, ys__n32318,
    ys__n32319, ys__n32320, ys__n32321, ys__n32322, ys__n32323, ys__n32324,
    ys__n32325, ys__n32326, ys__n32327, ys__n32328, ys__n32329, ys__n32330,
    ys__n32331, ys__n32332, ys__n32333, ys__n32334, ys__n32335, ys__n32336,
    ys__n32337, ys__n32338, ys__n32339, ys__n32340, ys__n32341, ys__n32342,
    ys__n32343, ys__n32344, ys__n32345, ys__n32346, ys__n32347, ys__n32348,
    ys__n32349, ys__n32350, ys__n32351, ys__n32352, ys__n32353, ys__n32354,
    ys__n32355, ys__n32356, ys__n32357, ys__n32358, ys__n32359, ys__n32360,
    ys__n32361, ys__n32362, ys__n32363, ys__n32364, ys__n32365, ys__n32366,
    ys__n32367, ys__n32368, ys__n32369, ys__n32370, ys__n32371, ys__n32372,
    ys__n32373, ys__n32374, ys__n32375, ys__n32376, ys__n32377, ys__n32378,
    ys__n32379, ys__n32380, ys__n32381, ys__n32382, ys__n32383, ys__n32384,
    ys__n32385, ys__n32386, ys__n32387, ys__n32388, ys__n32389, ys__n32390,
    ys__n32391, ys__n32392, ys__n32393, ys__n32394, ys__n32395, ys__n32396,
    ys__n32397, ys__n32398, ys__n32399, ys__n32400, ys__n32401, ys__n32402,
    ys__n32403, ys__n32404, ys__n32405, ys__n32406, ys__n32407, ys__n32408,
    ys__n32409, ys__n32410, ys__n32411, ys__n32412, ys__n32413, ys__n32414,
    ys__n32415, ys__n32416, ys__n32417, ys__n32418, ys__n32419, ys__n32420,
    ys__n32421, ys__n32422, ys__n32423, ys__n32424, ys__n32425, ys__n32426,
    ys__n32427, ys__n32428, ys__n32429, ys__n32430, ys__n32431, ys__n32432,
    ys__n32433, ys__n32434, ys__n32435, ys__n32436, ys__n32437, ys__n32438,
    ys__n32439, ys__n32440, ys__n32441, ys__n32442, ys__n32443, ys__n32444,
    ys__n32445, ys__n32446, ys__n32447, ys__n32448, ys__n32449, ys__n32450,
    ys__n32451, ys__n32452, ys__n32453, ys__n32454, ys__n32455, ys__n32456,
    ys__n32457, ys__n32458, ys__n32459, ys__n32460, ys__n32461, ys__n32462,
    ys__n32463, ys__n32464, ys__n32465, ys__n32466, ys__n32467, ys__n32468,
    ys__n32469, ys__n32470, ys__n32471, ys__n32472, ys__n32473, ys__n32474,
    ys__n32475, ys__n32476, ys__n32477, ys__n32478, ys__n32479, ys__n32480,
    ys__n32481, ys__n32482, ys__n32483, ys__n32484, ys__n32485, ys__n32486,
    ys__n32487, ys__n32488, ys__n32489, ys__n32490, ys__n32491, ys__n32492,
    ys__n32493, ys__n32494, ys__n32495, ys__n32496, ys__n32497, ys__n32498,
    ys__n32499, ys__n32500, ys__n32501, ys__n32502, ys__n32503, ys__n32504,
    ys__n32505, ys__n32506, ys__n32507, ys__n32508, ys__n32509, ys__n32510,
    ys__n32511, ys__n32512, ys__n32513, ys__n32514, ys__n32515, ys__n32516,
    ys__n32517, ys__n32518, ys__n32519, ys__n32520, ys__n32521, ys__n32522,
    ys__n32523, ys__n32524, ys__n32525, ys__n32526, ys__n32527, ys__n32528,
    ys__n32529, ys__n32530, ys__n32531, ys__n32532, ys__n32533, ys__n32534,
    ys__n32535, ys__n32536, ys__n32537, ys__n32538, ys__n32539, ys__n32540,
    ys__n32541, ys__n32542, ys__n32543, ys__n32544, ys__n32545, ys__n32546,
    ys__n32547, ys__n32548, ys__n32549, ys__n32550, ys__n32551, ys__n32552,
    ys__n32553, ys__n32554, ys__n32555, ys__n32556, ys__n32557, ys__n32558,
    ys__n32559, ys__n32560, ys__n32561, ys__n32562, ys__n32563, ys__n32564,
    ys__n32565, ys__n32566, ys__n32567, ys__n32568, ys__n32569, ys__n32570,
    ys__n32571, ys__n32572, ys__n32573, ys__n32574, ys__n32575, ys__n32576,
    ys__n32577, ys__n32578, ys__n32579, ys__n32580, ys__n32581, ys__n32582,
    ys__n32583, ys__n32584, ys__n32585, ys__n32586, ys__n32587, ys__n32588,
    ys__n32589, ys__n32590, ys__n32591, ys__n32592, ys__n32593, ys__n32594,
    ys__n32595, ys__n32596, ys__n32597, ys__n32598, ys__n32599, ys__n32600,
    ys__n32601, ys__n32602, ys__n32603, ys__n32604, ys__n32605, ys__n32606,
    ys__n32607, ys__n32608, ys__n32609, ys__n32610, ys__n32611, ys__n32612,
    ys__n32613, ys__n32614, ys__n32615, ys__n32616, ys__n32617, ys__n32618,
    ys__n32619, ys__n32620, ys__n32621, ys__n32622, ys__n32623, ys__n32624,
    ys__n32625, ys__n32626, ys__n32627, ys__n32628, ys__n32629, ys__n32630,
    ys__n32631, ys__n32632, ys__n32633, ys__n32634, ys__n32635, ys__n32636,
    ys__n32637, ys__n32638, ys__n32639, ys__n32640, ys__n32641, ys__n32642,
    ys__n32643, ys__n32644, ys__n32645, ys__n32646, ys__n32647, ys__n32648,
    ys__n32649, ys__n32650, ys__n32651, ys__n32652, ys__n32653, ys__n32654,
    ys__n32655, ys__n32656, ys__n32657, ys__n32658, ys__n32659, ys__n32660,
    ys__n32661, ys__n32662, ys__n32663, ys__n32664, ys__n32665, ys__n32666,
    ys__n32667, ys__n32668, ys__n32669, ys__n32670, ys__n32671, ys__n32672,
    ys__n32673, ys__n32674, ys__n32675, ys__n32676, ys__n32677, ys__n32678,
    ys__n32679, ys__n32680, ys__n32681, ys__n32682, ys__n32683, ys__n32684,
    ys__n32685, ys__n32686, ys__n32687, ys__n32688, ys__n32689, ys__n32690,
    ys__n32691, ys__n32692, ys__n32693, ys__n32694, ys__n32695, ys__n32696,
    ys__n32697, ys__n32698, ys__n32699, ys__n32700, ys__n32701, ys__n32702,
    ys__n32703, ys__n32704, ys__n32705, ys__n32706, ys__n32707, ys__n32708,
    ys__n32709, ys__n32710, ys__n32711, ys__n32712, ys__n32713, ys__n32714,
    ys__n32715, ys__n32716, ys__n32717, ys__n32718, ys__n32719, ys__n32720,
    ys__n32721, ys__n32722, ys__n32723, ys__n32724, ys__n32725, ys__n32726,
    ys__n32727, ys__n32728, ys__n32729, ys__n32730, ys__n32731, ys__n32732,
    ys__n32733, ys__n32734, ys__n32735, ys__n32736, ys__n32737, ys__n32738,
    ys__n32739, ys__n32740, ys__n32741, ys__n32742, ys__n32743, ys__n32744,
    ys__n32745, ys__n32746, ys__n32747, ys__n32748, ys__n32749, ys__n32750,
    ys__n32751, ys__n32752, ys__n32753, ys__n32754, ys__n32755, ys__n32756,
    ys__n32757, ys__n32758, ys__n32759, ys__n32760, ys__n32761, ys__n32762,
    ys__n32763, ys__n32764, ys__n32765, ys__n32766, ys__n32767, ys__n32768,
    ys__n32769, ys__n32770, ys__n32771, ys__n32772, ys__n32773, ys__n32774,
    ys__n32775, ys__n32776, ys__n32777, ys__n32778, ys__n32779, ys__n32780,
    ys__n32781, ys__n32782, ys__n32783, ys__n32784, ys__n32785, ys__n32786,
    ys__n32787, ys__n32788, ys__n32789, ys__n32790, ys__n32791, ys__n32792,
    ys__n32793, ys__n32794, ys__n32795, ys__n32796, ys__n32797, ys__n32798,
    ys__n32799, ys__n32800, ys__n32801, ys__n32802, ys__n32803, ys__n32804,
    ys__n32805, ys__n32806, ys__n32807, ys__n32808, ys__n32809, ys__n32810,
    ys__n32811, ys__n32812, ys__n32813, ys__n32814, ys__n32815, ys__n32816,
    ys__n32817, ys__n32818, ys__n32819, ys__n32820, ys__n32821, ys__n32822,
    ys__n32823, ys__n32824, ys__n32825, ys__n32826, ys__n32827, ys__n32828,
    ys__n32829, ys__n32830, ys__n32831, ys__n32832, ys__n32833, ys__n32834,
    ys__n32835, ys__n32836, ys__n32837, ys__n32838, ys__n32839, ys__n32840,
    ys__n32841, ys__n32842, ys__n32843, ys__n32844, ys__n32845, ys__n32846,
    ys__n32847, ys__n32848, ys__n32849, ys__n32850, ys__n32851, ys__n32852,
    ys__n32853, ys__n32854, ys__n32855, ys__n32856, ys__n32857, ys__n32858,
    ys__n32859, ys__n32860, ys__n32861, ys__n32862, ys__n32863, ys__n32864,
    ys__n32865, ys__n32866, ys__n32867, ys__n32868, ys__n32869, ys__n32870,
    ys__n32871, ys__n32872, ys__n32873, ys__n32874, ys__n32875, ys__n32876,
    ys__n32877, ys__n32878, ys__n32879, ys__n32880, ys__n32881, ys__n32882,
    ys__n32883, ys__n32884, ys__n32885, ys__n32886, ys__n32887, ys__n32888,
    ys__n32889, ys__n32890, ys__n32891, ys__n32892, ys__n32893, ys__n32894,
    ys__n32895, ys__n32896, ys__n32897, ys__n32898, ys__n32899, ys__n32900,
    ys__n32901, ys__n32902, ys__n32903, ys__n32904, ys__n32905, ys__n32906,
    ys__n32907, ys__n32908, ys__n32909, ys__n32910, ys__n32911, ys__n32912,
    ys__n32913, ys__n32914, ys__n32915, ys__n32916, ys__n32917, ys__n32918,
    ys__n32919, ys__n32920, ys__n32921, ys__n32922, ys__n32923, ys__n32924,
    ys__n32925, ys__n32926, ys__n32927, ys__n32928, ys__n32929, ys__n32930,
    ys__n32931, ys__n32932, ys__n32933, ys__n32934, ys__n32935, ys__n32936,
    ys__n32937, ys__n32938, ys__n32939, ys__n32940, ys__n32941, ys__n32942,
    ys__n32943, ys__n32944, ys__n32945, ys__n32946, ys__n32947, ys__n32948,
    ys__n32949, ys__n32950, ys__n32951, ys__n32952, ys__n32953, ys__n32954,
    ys__n32955, ys__n32956, ys__n32957, ys__n32958, ys__n32959, ys__n32960,
    ys__n32961, ys__n32962, ys__n32963, ys__n32964, ys__n32965, ys__n32966,
    ys__n32967, ys__n32968, ys__n32969, ys__n32970, ys__n32971, ys__n32972,
    ys__n32973, ys__n32974, ys__n32975, ys__n32976, ys__n32977, ys__n32978,
    ys__n32979, ys__n32980, ys__n32981, ys__n32982, ys__n32983, ys__n32984,
    ys__n32985, ys__n32986, ys__n32987, ys__n32988, ys__n32989, ys__n32990,
    ys__n32991, ys__n32992, ys__n32993, ys__n32994, ys__n32995, ys__n32996,
    ys__n32997, ys__n32998, ys__n33007, ys__n33008, ys__n33009, ys__n33014,
    ys__n33015, ys__n33016, ys__n33017, ys__n33018, ys__n33019, ys__n33020,
    ys__n33021, ys__n33022, ys__n33023, ys__n33024, ys__n33025, ys__n33026,
    ys__n33027, ys__n33028, ys__n33029, ys__n33030, ys__n33031, ys__n33032,
    ys__n33033, ys__n33034, ys__n33035, ys__n33036, ys__n33037, ys__n33038,
    ys__n33039, ys__n33040, ys__n33041, ys__n33042, ys__n33043, ys__n33044,
    ys__n33045, ys__n33046, ys__n33047, ys__n33048, ys__n33049, ys__n33050,
    ys__n33051, ys__n33052, ys__n33053, ys__n33054, ys__n33055, ys__n33056,
    ys__n33058, ys__n33059, ys__n33060, ys__n33061, ys__n33062, ys__n33063,
    ys__n33064, ys__n33065, ys__n33066, ys__n33067, ys__n33068, ys__n33069,
    ys__n33070, ys__n33071, ys__n33072, ys__n33073, ys__n33074, ys__n33075,
    ys__n33076, ys__n33077, ys__n33078, ys__n33079, ys__n33080, ys__n33081,
    ys__n33082, ys__n33083, ys__n33084, ys__n33085, ys__n33086, ys__n33087,
    ys__n33088, ys__n33089, ys__n33090, ys__n33091, ys__n33092, ys__n33093,
    ys__n33094, ys__n33095, ys__n33096, ys__n33097, ys__n33098, ys__n33099,
    ys__n33100, ys__n33101, ys__n33102, ys__n33103, ys__n33104, ys__n33105,
    ys__n33106, ys__n33107, ys__n33108, ys__n33109, ys__n33110, ys__n33111,
    ys__n33178, ys__n33179, ys__n33180, ys__n33181, ys__n33182, ys__n33183,
    ys__n33184, ys__n33185, ys__n33186, ys__n33187, ys__n33188, ys__n33189,
    ys__n33190, ys__n33191, ys__n33192, ys__n33193, ys__n33194, ys__n33195,
    ys__n33196, ys__n33197, ys__n33198, ys__n33199, ys__n33200, ys__n33201,
    ys__n33202, ys__n33203, ys__n33204, ys__n33205, ys__n33206, ys__n33207,
    ys__n33208, ys__n33209, ys__n33211, ys__n33317, ys__n33324, ys__n33329,
    ys__n33331, ys__n33333, ys__n33335, ys__n33337, ys__n33339, ys__n33357,
    ys__n33366, ys__n33414, ys__n33420, ys__n33437, ys__n33438, ys__n33439,
    ys__n33453, ys__n33454, ys__n33455, ys__n33456, ys__n33457, ys__n33513,
    ys__n33514, ys__n33515, ys__n33521, ys__n33535, ys__n34952, ys__n34953,
    ys__n34962, ys__n35052, ys__n35144, ys__n35146, ys__n35148, ys__n35150,
    ys__n35152, ys__n35154, ys__n35156, ys__n35158, ys__n35160, ys__n35162,
    ys__n35164, ys__n35166, ys__n35168, ys__n35170, ys__n35172, ys__n35174,
    ys__n35176, ys__n35178, ys__n35180, ys__n35182, ys__n35184, ys__n35186,
    ys__n35188, ys__n35190, ys__n35192, ys__n35194, ys__n35196, ys__n35198,
    ys__n35200, ys__n35202, ys__n35204, ys__n35206, ys__n35402, ys__n35404,
    ys__n35406, ys__n35408, ys__n35410, ys__n35412, ys__n35425, ys__n35705,
    ys__n35706, ys__n35708, ys__n35710, ys__n35712, ys__n35714, ys__n35716,
    ys__n37676, ys__n37687, ys__n37695, ys__n37697, ys__n37699, ys__n37702,
    ys__n37703, ys__n37707, ys__n37714, ys__n37731, ys__n37732, ys__n37733,
    ys__n37738, ys__n37739, ys__n37741, ys__n37742, ys__n38180, ys__n38182,
    ys__n38184, ys__n38185, ys__n38186, ys__n38188, ys__n38191, ys__n38205,
    ys__n38207, ys__n38209, ys__n38211, ys__n38213, ys__n38214, ys__n38216,
    ys__n38218, ys__n38222, ys__n38224, ys__n38246, ys__n38247, ys__n38248,
    ys__n38250, ys__n38252, ys__n38263, ys__n38266, ys__n38281, ys__n38285,
    ys__n38287, ys__n38289, ys__n38292, ys__n38294, ys__n38296, ys__n38303,
    ys__n38325, ys__n38326, ys__n38327, ys__n38328, ys__n38330, ys__n38331,
    ys__n38332, ys__n38334, ys__n38336, ys__n38337, ys__n38338, ys__n38339,
    ys__n38340, ys__n38341, ys__n38342, ys__n38343, ys__n38344, ys__n38345,
    ys__n38347, ys__n38349, ys__n38351, ys__n38352, ys__n38353, ys__n38354,
    ys__n38355, ys__n38356, ys__n38357, ys__n38359, ys__n38360, ys__n38362,
    ys__n38364, ys__n38365, ys__n38366, ys__n38367, ys__n38368, ys__n38369,
    ys__n38370, ys__n38371, ys__n38372, ys__n38373, ys__n38374, ys__n38375,
    ys__n38377, ys__n38379, ys__n38381, ys__n38383, ys__n38385, ys__n38387,
    ys__n38388, ys__n38389, ys__n38390, ys__n38391, ys__n38392, ys__n38393,
    ys__n38394, ys__n38396, ys__n38397, ys__n38417, ys__n38453, ys__n38456,
    ys__n38508, ys__n38509, ys__n38510, ys__n38515, ys__n38518, ys__n38520,
    ys__n38521, ys__n38523, ys__n38525, ys__n38552, ys__n38555, ys__n38556,
    ys__n38563, ys__n38566, ys__n38615, ys__n38623, ys__n38628, ys__n38633,
    ys__n38650, ys__n38662, ys__n38668, ys__n38669, ys__n38672, ys__n38674,
    ys__n38677, ys__n38689, ys__n38742, ys__n38768, ys__n38795, ys__n38799,
    ys__n38801, ys__n38884, ys__n38886, ys__n38887, ys__n38900, ys__n38912,
    ys__n38913, ys__n38914, ys__n38915, ys__n38917, ys__n38923, ys__n38925,
    ys__n38930, ys__n39392, ys__n39393, ys__n39395, ys__n39396, ys__n39397,
    ys__n39398, ys__n39399, ys__n39400, ys__n39401, ys__n39402, ys__n39403,
    ys__n39404, ys__n39405, ys__n39406, ys__n39407, ys__n39408, ys__n39409,
    ys__n39410, ys__n39411, ys__n39412, ys__n39413, ys__n39414, ys__n39415,
    ys__n39416, ys__n39417, ys__n39418, ys__n40052, ys__n42129, ys__n42153,
    ys__n42189, ys__n42194, ys__n42229, ys__n42234, ys__n42270, ys__n42275,
    ys__n42311, ys__n42316, ys__n42352, ys__n42357, ys__n42393, ys__n42398,
    ys__n42434, ys__n42439, ys__n42488, ys__n42493, ys__n42541, ys__n42546,
    ys__n42594, ys__n42599, ys__n42647, ys__n42652, ys__n42701, ys__n42706,
    ys__n42755, ys__n42760, ys__n42809, ys__n42814, ys__n42863, ys__n42868,
    ys__n42917, ys__n42922, ys__n42971, ys__n42976, ys__n43025, ys__n43030,
    ys__n43079, ys__n43084, ys__n43133, ys__n43138, ys__n43187, ys__n43192,
    ys__n43241, ys__n43246, ys__n43295, ys__n43300, ys__n43349, ys__n43354,
    ys__n43403, ys__n43408, ys__n43457, ys__n43462, ys__n43511, ys__n43516,
    ys__n43565, ys__n43570, ys__n43619, ys__n43624, ys__n43673, ys__n43678,
    ys__n43727, ys__n43732, ys__n43781, ys__n43786, ys__n43835, ys__n43840,
    ys__n43889, ys__n43894, ys__n43932, ys__n43937, ys__n43975, ys__n43980,
    ys__n44018, ys__n44023, ys__n44048, ys__n44053, ys__n44089, ys__n44094,
    ys__n44119, ys__n44122, ys__n44136, ys__n44139, ys__n44155, ys__n44160,
    ys__n44183, ys__n44186, ys__n44189, ys__n44192, ys__n44195, ys__n44198,
    ys__n44205, ys__n44213, ys__n44216, ys__n44219, ys__n44836, ys__n44838,
    ys__n44841, ys__n44843, ys__n44844, ys__n44845, ys__n44846, ys__n44848,
    ys__n44850, ys__n44851, ys__n44852, ys__n44853, ys__n44854, ys__n44855,
    ys__n44858, ys__n44948, ys__n44949, ys__n44950, ys__n44952, ys__n44953,
    ys__n44954, ys__n44955, ys__n44956, ys__n44957, ys__n44958, ys__n44959,
    ys__n44960, ys__n44961, ys__n44962, ys__n44963, ys__n44964, ys__n44965,
    ys__n44966, ys__n44967, ys__n44968, ys__n44969, ys__n44970, ys__n44971,
    ys__n44972, ys__n44973, ys__n44974, ys__n44975, ys__n44976, ys__n44977,
    ys__n44978, ys__n44979, ys__n44980, ys__n44981, ys__n44982, ys__n44983,
    ys__n44985, ys__n44987, ys__n46131, ys__n46133, ys__n46135, ys__n46137,
    ys__n46143, ys__n46146, ys__n46154, ys__n46155, ys__n46158, ys__n46159,
    ys__n46162, ys__n46163, ys__n46172, ys__n46173, ys__n46176, ys__n46179,
    ys__n46188, ys__n46189, ys__n46192, ys__n46195, ys__n46204, ys__n46205,
    ys__n46208, ys__n46211, ys__n46220, ys__n46221, ys__n46224, ys__n46227,
    ys__n46233, ys__n46234, ys__n48339, ys__n48340, ys__n48341, ys__n48342,
    ys__n48343, ys__n48344, ys__n48348, ys__n48349, ys__n48350, ys__n48351,
    ys__n48352, ys__n48353, ys__n48354, ys__n48355, ys__n48356, ys__n48357,
    ys__n48358, ys__n48359, ys__n48360, ys__n48361, ys__n48362;
  wire new_n11532_, new_n11533_, new_n11534_, new_n11535_, new_n11536_,
    new_n11537_, new_n11538_, new_n11539_, new_n11540_, new_n11541_,
    new_n11542_, new_n11543_, new_n11544_, new_n11545_, new_n11546_,
    new_n11547_, new_n11548_, new_n11549_, new_n11550_, new_n11551_,
    new_n11552_, new_n11553_, new_n11554_, new_n11555_, new_n11556_,
    new_n11557_, new_n11558_, new_n11559_, new_n11560_, new_n11561_,
    new_n11562_, new_n11563_, new_n11564_, new_n11565_, new_n11566_,
    new_n11567_, new_n11568_, new_n11569_, new_n11570_, new_n11571_,
    new_n11572_, new_n11573_, new_n11574_, new_n11575_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11749_, new_n11750_, new_n11752_, new_n11753_, new_n11754_,
    new_n11755_, new_n11756_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11964_, new_n11965_, new_n11966_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11979_,
    new_n11980_, new_n11981_, new_n11982_, new_n11983_, new_n11984_,
    new_n11985_, new_n11986_, new_n11987_, new_n11988_, new_n11989_,
    new_n11990_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12008_, new_n12009_, new_n12010_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12024_,
    new_n12025_, new_n12026_, new_n12027_, new_n12028_, new_n12029_,
    new_n12030_, new_n12031_, new_n12032_, new_n12033_, new_n12034_,
    new_n12035_, new_n12036_, new_n12037_, new_n12038_, new_n12039_,
    new_n12040_, new_n12041_, new_n12042_, new_n12043_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12075_, new_n12076_,
    new_n12077_, new_n12078_, new_n12079_, new_n12081_, new_n12082_,
    new_n12083_, new_n12084_, new_n12085_, new_n12086_, new_n12087_,
    new_n12088_, new_n12089_, new_n12090_, new_n12091_, new_n12092_,
    new_n12093_, new_n12094_, new_n12095_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12101_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12116_,
    new_n12117_, new_n12118_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12142_, new_n12143_,
    new_n12144_, new_n12145_, new_n12146_, new_n12147_, new_n12148_,
    new_n12149_, new_n12150_, new_n12151_, new_n12152_, new_n12153_,
    new_n12154_, new_n12155_, new_n12156_, new_n12157_, new_n12158_,
    new_n12159_, new_n12160_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12197_, new_n12198_, new_n12199_, new_n12200_, new_n12201_,
    new_n12202_, new_n12203_, new_n12204_, new_n12205_, new_n12206_,
    new_n12207_, new_n12208_, new_n12209_, new_n12210_, new_n12211_,
    new_n12212_, new_n12213_, new_n12214_, new_n12215_, new_n12216_,
    new_n12217_, new_n12218_, new_n12219_, new_n12220_, new_n12221_,
    new_n12222_, new_n12223_, new_n12224_, new_n12225_, new_n12226_,
    new_n12227_, new_n12228_, new_n12229_, new_n12230_, new_n12231_,
    new_n12232_, new_n12233_, new_n12234_, new_n12235_, new_n12236_,
    new_n12237_, new_n12238_, new_n12239_, new_n12240_, new_n12241_,
    new_n12242_, new_n12243_, new_n12245_, new_n12246_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12253_, new_n12254_,
    new_n12255_, new_n12256_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12271_,
    new_n12272_, new_n12274_, new_n12275_, new_n12276_, new_n12277_,
    new_n12278_, new_n12279_, new_n12280_, new_n12281_, new_n12282_,
    new_n12283_, new_n12284_, new_n12285_, new_n12286_, new_n12287_,
    new_n12288_, new_n12289_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12297_, new_n12298_, new_n12299_,
    new_n12300_, new_n12301_, new_n12302_, new_n12303_, new_n12304_,
    new_n12305_, new_n12306_, new_n12307_, new_n12308_, new_n12309_,
    new_n12310_, new_n12311_, new_n12312_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12454_, new_n12455_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12787_, new_n12788_, new_n12789_, new_n12790_, new_n12791_,
    new_n12792_, new_n12793_, new_n12794_, new_n12795_, new_n12796_,
    new_n12797_, new_n12798_, new_n12799_, new_n12800_, new_n12801_,
    new_n12802_, new_n12803_, new_n12805_, new_n12806_, new_n12807_,
    new_n12808_, new_n12809_, new_n12810_, new_n12811_, new_n12812_,
    new_n12813_, new_n12814_, new_n12815_, new_n12816_, new_n12817_,
    new_n12818_, new_n12819_, new_n12820_, new_n12821_, new_n12822_,
    new_n12823_, new_n12824_, new_n12825_, new_n12826_, new_n12827_,
    new_n12828_, new_n12829_, new_n12830_, new_n12831_, new_n12832_,
    new_n12833_, new_n12834_, new_n12835_, new_n12836_, new_n12837_,
    new_n12838_, new_n12839_, new_n12840_, new_n12842_, new_n12843_,
    new_n12844_, new_n12845_, new_n12846_, new_n12847_, new_n12848_,
    new_n12849_, new_n12850_, new_n12851_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12869_, new_n12870_,
    new_n12871_, new_n12873_, new_n12874_, new_n12875_, new_n12877_,
    new_n12879_, new_n12880_, new_n12881_, new_n12882_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12905_, new_n12906_,
    new_n12907_, new_n12908_, new_n12909_, new_n12910_, new_n12911_,
    new_n12912_, new_n12913_, new_n12915_, new_n12916_, new_n12917_,
    new_n12918_, new_n12919_, new_n12920_, new_n12921_, new_n12923_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12948_, new_n12949_, new_n12950_, new_n12951_,
    new_n12953_, new_n12954_, new_n12955_, new_n12956_, new_n12957_,
    new_n12958_, new_n12960_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12970_,
    new_n12971_, new_n12972_, new_n12974_, new_n12975_, new_n12976_,
    new_n12977_, new_n12978_, new_n12979_, new_n12980_, new_n12982_,
    new_n12983_, new_n12985_, new_n12986_, new_n12987_, new_n12988_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12997_, new_n12999_, new_n13000_, new_n13001_,
    new_n13002_, new_n13003_, new_n13005_, new_n13006_, new_n13007_,
    new_n13008_, new_n13010_, new_n13011_, new_n13012_, new_n13013_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13022_, new_n13024_, new_n13025_, new_n13026_,
    new_n13027_, new_n13028_, new_n13030_, new_n13031_, new_n13032_,
    new_n13033_, new_n13035_, new_n13036_, new_n13037_, new_n13038_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13047_, new_n13049_, new_n13050_, new_n13051_,
    new_n13052_, new_n13053_, new_n13055_, new_n13056_, new_n13057_,
    new_n13058_, new_n13060_, new_n13061_, new_n13062_, new_n13063_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13072_, new_n13074_, new_n13075_, new_n13076_,
    new_n13077_, new_n13078_, new_n13080_, new_n13081_, new_n13082_,
    new_n13083_, new_n13085_, new_n13086_, new_n13087_, new_n13088_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13097_, new_n13099_, new_n13100_, new_n13101_,
    new_n13102_, new_n13103_, new_n13105_, new_n13106_, new_n13107_,
    new_n13108_, new_n13110_, new_n13111_, new_n13112_, new_n13113_,
    new_n13115_, new_n13116_, new_n13117_, new_n13118_, new_n13119_,
    new_n13120_, new_n13122_, new_n13124_, new_n13125_, new_n13126_,
    new_n13127_, new_n13128_, new_n13130_, new_n13131_, new_n13132_,
    new_n13133_, new_n13135_, new_n13136_, new_n13137_, new_n13138_,
    new_n13140_, new_n13141_, new_n13142_, new_n13143_, new_n13144_,
    new_n13145_, new_n13147_, new_n13149_, new_n13150_, new_n13151_,
    new_n13152_, new_n13153_, new_n13155_, new_n13156_, new_n13157_,
    new_n13158_, new_n13160_, new_n13161_, new_n13162_, new_n13163_,
    new_n13165_, new_n13166_, new_n13167_, new_n13168_, new_n13169_,
    new_n13170_, new_n13172_, new_n13174_, new_n13175_, new_n13176_,
    new_n13177_, new_n13178_, new_n13180_, new_n13181_, new_n13182_,
    new_n13183_, new_n13185_, new_n13187_, new_n13188_, new_n13189_,
    new_n13190_, new_n13191_, new_n13192_, new_n13193_, new_n13194_,
    new_n13195_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13206_,
    new_n13207_, new_n13208_, new_n13209_, new_n13210_, new_n13211_,
    new_n13212_, new_n13213_, new_n13214_, new_n13215_, new_n13216_,
    new_n13217_, new_n13218_, new_n13219_, new_n13220_, new_n13221_,
    new_n13222_, new_n13223_, new_n13224_, new_n13226_, new_n13227_,
    new_n13228_, new_n13229_, new_n13230_, new_n13231_, new_n13232_,
    new_n13233_, new_n13234_, new_n13235_, new_n13236_, new_n13237_,
    new_n13238_, new_n13239_, new_n13240_, new_n13242_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13258_, new_n13259_, new_n13260_, new_n13261_,
    new_n13263_, new_n13264_, new_n13265_, new_n13266_, new_n13267_,
    new_n13268_, new_n13269_, new_n13270_, new_n13271_, new_n13272_,
    new_n13274_, new_n13275_, new_n13276_, new_n13277_, new_n13278_,
    new_n13280_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13293_, new_n13294_, new_n13295_, new_n13296_,
    new_n13297_, new_n13298_, new_n13299_, new_n13300_, new_n13301_,
    new_n13302_, new_n13304_, new_n13305_, new_n13306_, new_n13307_,
    new_n13308_, new_n13309_, new_n13310_, new_n13311_, new_n13312_,
    new_n13313_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13326_, new_n13327_, new_n13328_, new_n13329_,
    new_n13330_, new_n13331_, new_n13332_, new_n13333_, new_n13334_,
    new_n13335_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13348_, new_n13349_, new_n13350_, new_n13351_,
    new_n13352_, new_n13353_, new_n13355_, new_n13356_, new_n13357_,
    new_n13358_, new_n13359_, new_n13360_, new_n13361_, new_n13362_,
    new_n13366_, new_n13368_, new_n13369_, new_n13370_, new_n13371_,
    new_n13372_, new_n13374_, new_n13375_, new_n13376_, new_n13377_,
    new_n13378_, new_n13379_, new_n13380_, new_n13381_, new_n13382_,
    new_n13383_, new_n13384_, new_n13385_, new_n13386_, new_n13387_,
    new_n13388_, new_n13389_, new_n13390_, new_n13391_, new_n13393_,
    new_n13394_, new_n13395_, new_n13396_, new_n13397_, new_n13398_,
    new_n13399_, new_n13400_, new_n13401_, new_n13402_, new_n13403_,
    new_n13404_, new_n13405_, new_n13406_, new_n13407_, new_n13408_,
    new_n13409_, new_n13410_, new_n13411_, new_n13412_, new_n13413_,
    new_n13414_, new_n13415_, new_n13416_, new_n13417_, new_n13418_,
    new_n13419_, new_n13420_, new_n13421_, new_n13423_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13431_, new_n13432_,
    new_n13434_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13451_,
    new_n13452_, new_n13453_, new_n13454_, new_n13455_, new_n13456_,
    new_n13457_, new_n13458_, new_n13459_, new_n13460_, new_n13461_,
    new_n13462_, new_n13463_, new_n13465_, new_n13466_, new_n13467_,
    new_n13470_, new_n13471_, new_n13472_, new_n13473_, new_n13474_,
    new_n13475_, new_n13476_, new_n13477_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13507_,
    new_n13508_, new_n13509_, new_n13511_, new_n13512_, new_n13513_,
    new_n13514_, new_n13516_, new_n13517_, new_n13519_, new_n13520_,
    new_n13522_, new_n13523_, new_n13525_, new_n13526_, new_n13527_,
    new_n13528_, new_n13529_, new_n13530_, new_n13531_, new_n13534_,
    new_n13535_, new_n13537_, new_n13538_, new_n13540_, new_n13541_,
    new_n13542_, new_n13544_, new_n13545_, new_n13547_, new_n13548_,
    new_n13550_, new_n13551_, new_n13553_, new_n13554_, new_n13556_,
    new_n13557_, new_n13559_, new_n13560_, new_n13562_, new_n13563_,
    new_n13564_, new_n13565_, new_n13566_, new_n13568_, new_n13573_,
    new_n13577_, new_n13581_, new_n13582_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13589_, new_n13590_, new_n13592_,
    new_n13593_, new_n13594_, new_n13595_, new_n13606_, new_n13607_,
    new_n13609_, new_n13610_, new_n13611_, new_n13617_, new_n13618_,
    new_n13619_, new_n13620_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13639_, new_n13641_, new_n13643_,
    new_n13644_, new_n13651_, new_n13652_, new_n13653_, new_n13655_,
    new_n13660_, new_n13662_, new_n13687_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13696_,
    new_n13698_, new_n13699_, new_n13700_, new_n13701_, new_n13702_,
    new_n13703_, new_n13707_, new_n13708_, new_n13709_, new_n13713_,
    new_n13714_, new_n13715_, new_n13716_, new_n13717_, new_n13718_,
    new_n13719_, new_n13720_, new_n13722_, new_n13723_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13744_, new_n13746_, new_n13747_, new_n13748_,
    new_n13749_, new_n13750_, new_n13751_, new_n13752_, new_n13753_,
    new_n13754_, new_n13755_, new_n13756_, new_n13757_, new_n13758_,
    new_n13759_, new_n13760_, new_n13761_, new_n13763_, new_n13765_,
    new_n13767_, new_n13769_, new_n13771_, new_n13772_, new_n13773_,
    new_n13774_, new_n13775_, new_n13776_, new_n13777_, new_n13778_,
    new_n13779_, new_n13780_, new_n13781_, new_n13782_, new_n13783_,
    new_n13784_, new_n13785_, new_n13786_, new_n13787_, new_n13788_,
    new_n13789_, new_n13790_, new_n13791_, new_n13792_, new_n13793_,
    new_n13794_, new_n13795_, new_n13796_, new_n13797_, new_n13798_,
    new_n13799_, new_n13800_, new_n13801_, new_n13802_, new_n13803_,
    new_n13804_, new_n13805_, new_n13806_, new_n13807_, new_n13808_,
    new_n13809_, new_n13810_, new_n13811_, new_n13812_, new_n13813_,
    new_n13814_, new_n13815_, new_n13816_, new_n13817_, new_n13818_,
    new_n13819_, new_n13820_, new_n13821_, new_n13822_, new_n13823_,
    new_n13824_, new_n13825_, new_n13826_, new_n13827_, new_n13828_,
    new_n13829_, new_n13830_, new_n13831_, new_n13832_, new_n13833_,
    new_n13834_, new_n13835_, new_n13836_, new_n13837_, new_n13838_,
    new_n13839_, new_n13840_, new_n13841_, new_n13842_, new_n13843_,
    new_n13844_, new_n13845_, new_n13846_, new_n13847_, new_n13848_,
    new_n13849_, new_n13850_, new_n13851_, new_n13852_, new_n13853_,
    new_n13854_, new_n13855_, new_n13856_, new_n13857_, new_n13858_,
    new_n13859_, new_n13860_, new_n13861_, new_n13862_, new_n13863_,
    new_n13864_, new_n13865_, new_n13866_, new_n13867_, new_n13868_,
    new_n13869_, new_n13870_, new_n13871_, new_n13872_, new_n13873_,
    new_n13874_, new_n13875_, new_n13876_, new_n13877_, new_n13878_,
    new_n13879_, new_n13880_, new_n13881_, new_n13882_, new_n13883_,
    new_n13884_, new_n13885_, new_n13886_, new_n13887_, new_n13888_,
    new_n13889_, new_n13890_, new_n13891_, new_n13892_, new_n13893_,
    new_n13894_, new_n13895_, new_n13896_, new_n13897_, new_n13898_,
    new_n13899_, new_n13900_, new_n13901_, new_n13902_, new_n13903_,
    new_n13904_, new_n13905_, new_n13906_, new_n13907_, new_n13908_,
    new_n13909_, new_n13910_, new_n13911_, new_n13912_, new_n13913_,
    new_n13914_, new_n13915_, new_n13916_, new_n13917_, new_n13918_,
    new_n13919_, new_n13920_, new_n13921_, new_n13922_, new_n13923_,
    new_n13924_, new_n13925_, new_n13926_, new_n13927_, new_n13928_,
    new_n13929_, new_n13930_, new_n13931_, new_n13932_, new_n13933_,
    new_n13934_, new_n13935_, new_n13936_, new_n13937_, new_n13938_,
    new_n13939_, new_n13940_, new_n13941_, new_n13942_, new_n13943_,
    new_n13944_, new_n13945_, new_n13946_, new_n13947_, new_n13948_,
    new_n13949_, new_n13950_, new_n13951_, new_n13952_, new_n13953_,
    new_n13954_, new_n13955_, new_n13956_, new_n13957_, new_n13958_,
    new_n13959_, new_n13960_, new_n13961_, new_n13962_, new_n13963_,
    new_n13964_, new_n13965_, new_n13966_, new_n13967_, new_n13968_,
    new_n13969_, new_n13970_, new_n13971_, new_n13972_, new_n13973_,
    new_n13974_, new_n13975_, new_n13976_, new_n13977_, new_n13978_,
    new_n13979_, new_n13980_, new_n13981_, new_n13982_, new_n13983_,
    new_n13984_, new_n13985_, new_n13986_, new_n13987_, new_n13988_,
    new_n13989_, new_n13990_, new_n13991_, new_n13992_, new_n13993_,
    new_n13994_, new_n13995_, new_n13996_, new_n13997_, new_n13998_,
    new_n13999_, new_n14000_, new_n14001_, new_n14002_, new_n14003_,
    new_n14004_, new_n14005_, new_n14006_, new_n14007_, new_n14008_,
    new_n14009_, new_n14010_, new_n14011_, new_n14012_, new_n14013_,
    new_n14014_, new_n14015_, new_n14016_, new_n14017_, new_n14018_,
    new_n14019_, new_n14020_, new_n14021_, new_n14022_, new_n14023_,
    new_n14024_, new_n14025_, new_n14026_, new_n14027_, new_n14028_,
    new_n14029_, new_n14030_, new_n14031_, new_n14032_, new_n14033_,
    new_n14034_, new_n14035_, new_n14036_, new_n14037_, new_n14038_,
    new_n14039_, new_n14040_, new_n14041_, new_n14042_, new_n14043_,
    new_n14044_, new_n14045_, new_n14046_, new_n14047_, new_n14048_,
    new_n14049_, new_n14050_, new_n14051_, new_n14052_, new_n14053_,
    new_n14054_, new_n14055_, new_n14056_, new_n14057_, new_n14058_,
    new_n14059_, new_n14060_, new_n14061_, new_n14062_, new_n14063_,
    new_n14064_, new_n14065_, new_n14066_, new_n14067_, new_n14068_,
    new_n14069_, new_n14070_, new_n14071_, new_n14072_, new_n14073_,
    new_n14074_, new_n14075_, new_n14076_, new_n14077_, new_n14078_,
    new_n14079_, new_n14080_, new_n14081_, new_n14082_, new_n14083_,
    new_n14084_, new_n14085_, new_n14086_, new_n14087_, new_n14088_,
    new_n14089_, new_n14090_, new_n14091_, new_n14092_, new_n14093_,
    new_n14094_, new_n14095_, new_n14096_, new_n14097_, new_n14098_,
    new_n14099_, new_n14100_, new_n14101_, new_n14102_, new_n14103_,
    new_n14104_, new_n14105_, new_n14106_, new_n14107_, new_n14108_,
    new_n14109_, new_n14110_, new_n14111_, new_n14112_, new_n14113_,
    new_n14114_, new_n14115_, new_n14116_, new_n14117_, new_n14118_,
    new_n14119_, new_n14120_, new_n14121_, new_n14122_, new_n14123_,
    new_n14124_, new_n14125_, new_n14126_, new_n14127_, new_n14128_,
    new_n14129_, new_n14130_, new_n14131_, new_n14132_, new_n14133_,
    new_n14134_, new_n14135_, new_n14136_, new_n14137_, new_n14138_,
    new_n14139_, new_n14140_, new_n14141_, new_n14142_, new_n14143_,
    new_n14144_, new_n14145_, new_n14146_, new_n14147_, new_n14148_,
    new_n14149_, new_n14150_, new_n14151_, new_n14152_, new_n14153_,
    new_n14154_, new_n14155_, new_n14156_, new_n14157_, new_n14158_,
    new_n14159_, new_n14160_, new_n14161_, new_n14162_, new_n14163_,
    new_n14164_, new_n14165_, new_n14166_, new_n14167_, new_n14168_,
    new_n14169_, new_n14170_, new_n14171_, new_n14172_, new_n14173_,
    new_n14174_, new_n14175_, new_n14176_, new_n14177_, new_n14178_,
    new_n14179_, new_n14180_, new_n14181_, new_n14182_, new_n14183_,
    new_n14184_, new_n14185_, new_n14186_, new_n14187_, new_n14188_,
    new_n14189_, new_n14190_, new_n14191_, new_n14192_, new_n14193_,
    new_n14194_, new_n14195_, new_n14196_, new_n14197_, new_n14198_,
    new_n14199_, new_n14200_, new_n14201_, new_n14202_, new_n14203_,
    new_n14204_, new_n14205_, new_n14206_, new_n14207_, new_n14208_,
    new_n14209_, new_n14210_, new_n14211_, new_n14212_, new_n14213_,
    new_n14214_, new_n14215_, new_n14216_, new_n14217_, new_n14218_,
    new_n14219_, new_n14220_, new_n14221_, new_n14222_, new_n14223_,
    new_n14224_, new_n14225_, new_n14226_, new_n14227_, new_n14228_,
    new_n14229_, new_n14230_, new_n14231_, new_n14232_, new_n14233_,
    new_n14234_, new_n14235_, new_n14236_, new_n14237_, new_n14238_,
    new_n14239_, new_n14240_, new_n14241_, new_n14242_, new_n14243_,
    new_n14244_, new_n14245_, new_n14246_, new_n14247_, new_n14248_,
    new_n14249_, new_n14250_, new_n14251_, new_n14252_, new_n14253_,
    new_n14254_, new_n14255_, new_n14256_, new_n14257_, new_n14258_,
    new_n14259_, new_n14260_, new_n14261_, new_n14262_, new_n14263_,
    new_n14264_, new_n14265_, new_n14266_, new_n14267_, new_n14268_,
    new_n14269_, new_n14270_, new_n14271_, new_n14272_, new_n14273_,
    new_n14274_, new_n14275_, new_n14276_, new_n14277_, new_n14278_,
    new_n14279_, new_n14280_, new_n14281_, new_n14282_, new_n14283_,
    new_n14284_, new_n14285_, new_n14286_, new_n14287_, new_n14288_,
    new_n14289_, new_n14290_, new_n14291_, new_n14292_, new_n14293_,
    new_n14294_, new_n14295_, new_n14296_, new_n14297_, new_n14298_,
    new_n14299_, new_n14300_, new_n14301_, new_n14302_, new_n14303_,
    new_n14304_, new_n14305_, new_n14306_, new_n14307_, new_n14308_,
    new_n14309_, new_n14310_, new_n14311_, new_n14312_, new_n14313_,
    new_n14314_, new_n14315_, new_n14316_, new_n14317_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14324_, new_n14325_, new_n14326_, new_n14327_, new_n14328_,
    new_n14329_, new_n14330_, new_n14331_, new_n14332_, new_n14333_,
    new_n14334_, new_n14335_, new_n14336_, new_n14337_, new_n14338_,
    new_n14339_, new_n14340_, new_n14341_, new_n14342_, new_n14343_,
    new_n14344_, new_n14345_, new_n14346_, new_n14347_, new_n14348_,
    new_n14349_, new_n14350_, new_n14351_, new_n14352_, new_n14353_,
    new_n14354_, new_n14355_, new_n14356_, new_n14357_, new_n14358_,
    new_n14359_, new_n14360_, new_n14361_, new_n14362_, new_n14363_,
    new_n14364_, new_n14365_, new_n14366_, new_n14367_, new_n14368_,
    new_n14369_, new_n14370_, new_n14371_, new_n14372_, new_n14373_,
    new_n14374_, new_n14375_, new_n14376_, new_n14377_, new_n14378_,
    new_n14379_, new_n14380_, new_n14381_, new_n14382_, new_n14383_,
    new_n14384_, new_n14385_, new_n14386_, new_n14387_, new_n14388_,
    new_n14389_, new_n14390_, new_n14391_, new_n14392_, new_n14393_,
    new_n14394_, new_n14395_, new_n14396_, new_n14397_, new_n14398_,
    new_n14399_, new_n14400_, new_n14401_, new_n14402_, new_n14403_,
    new_n14404_, new_n14405_, new_n14406_, new_n14407_, new_n14408_,
    new_n14409_, new_n14410_, new_n14411_, new_n14412_, new_n14413_,
    new_n14414_, new_n14415_, new_n14416_, new_n14417_, new_n14418_,
    new_n14419_, new_n14420_, new_n14421_, new_n14422_, new_n14423_,
    new_n14424_, new_n14425_, new_n14426_, new_n14427_, new_n14428_,
    new_n14429_, new_n14430_, new_n14431_, new_n14432_, new_n14433_,
    new_n14434_, new_n14435_, new_n14436_, new_n14437_, new_n14438_,
    new_n14439_, new_n14440_, new_n14441_, new_n14442_, new_n14443_,
    new_n14444_, new_n14445_, new_n14446_, new_n14447_, new_n14448_,
    new_n14449_, new_n14450_, new_n14451_, new_n14452_, new_n14453_,
    new_n14454_, new_n14455_, new_n14456_, new_n14457_, new_n14458_,
    new_n14459_, new_n14460_, new_n14461_, new_n14462_, new_n14463_,
    new_n14464_, new_n14465_, new_n14466_, new_n14467_, new_n14468_,
    new_n14469_, new_n14470_, new_n14471_, new_n14472_, new_n14473_,
    new_n14474_, new_n14475_, new_n14476_, new_n14477_, new_n14478_,
    new_n14479_, new_n14480_, new_n14481_, new_n14482_, new_n14483_,
    new_n14484_, new_n14485_, new_n14486_, new_n14487_, new_n14488_,
    new_n14489_, new_n14490_, new_n14491_, new_n14492_, new_n14493_,
    new_n14494_, new_n14495_, new_n14496_, new_n14497_, new_n14498_,
    new_n14499_, new_n14500_, new_n14501_, new_n14502_, new_n14503_,
    new_n14504_, new_n14505_, new_n14506_, new_n14507_, new_n14508_,
    new_n14509_, new_n14510_, new_n14511_, new_n14512_, new_n14513_,
    new_n14514_, new_n14515_, new_n14516_, new_n14517_, new_n14518_,
    new_n14519_, new_n14520_, new_n14521_, new_n14522_, new_n14523_,
    new_n14524_, new_n14525_, new_n14526_, new_n14527_, new_n14528_,
    new_n14529_, new_n14530_, new_n14531_, new_n14532_, new_n14533_,
    new_n14534_, new_n14535_, new_n14536_, new_n14537_, new_n14538_,
    new_n14539_, new_n14540_, new_n14541_, new_n14542_, new_n14543_,
    new_n14544_, new_n14545_, new_n14546_, new_n14547_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14589_, new_n14590_, new_n14591_, new_n14592_, new_n14593_,
    new_n14594_, new_n14595_, new_n14596_, new_n14597_, new_n14598_,
    new_n14599_, new_n14600_, new_n14601_, new_n14602_, new_n14603_,
    new_n14604_, new_n14605_, new_n14606_, new_n14607_, new_n14608_,
    new_n14609_, new_n14610_, new_n14611_, new_n14612_, new_n14613_,
    new_n14614_, new_n14615_, new_n14616_, new_n14617_, new_n14618_,
    new_n14619_, new_n14620_, new_n14621_, new_n14622_, new_n14623_,
    new_n14624_, new_n14625_, new_n14626_, new_n14627_, new_n14628_,
    new_n14629_, new_n14630_, new_n14631_, new_n14632_, new_n14633_,
    new_n14634_, new_n14635_, new_n14636_, new_n14637_, new_n14638_,
    new_n14639_, new_n14640_, new_n14641_, new_n14642_, new_n14643_,
    new_n14644_, new_n14645_, new_n14646_, new_n14647_, new_n14648_,
    new_n14649_, new_n14650_, new_n14651_, new_n14652_, new_n14653_,
    new_n14654_, new_n14655_, new_n14656_, new_n14657_, new_n14658_,
    new_n14659_, new_n14660_, new_n14661_, new_n14662_, new_n14663_,
    new_n14664_, new_n14665_, new_n14666_, new_n14667_, new_n14668_,
    new_n14669_, new_n14670_, new_n14671_, new_n14672_, new_n14673_,
    new_n14674_, new_n14675_, new_n14676_, new_n14677_, new_n14678_,
    new_n14679_, new_n14680_, new_n14681_, new_n14682_, new_n14683_,
    new_n14684_, new_n14685_, new_n14686_, new_n14687_, new_n14688_,
    new_n14689_, new_n14690_, new_n14691_, new_n14692_, new_n14693_,
    new_n14694_, new_n14695_, new_n14696_, new_n14697_, new_n14698_,
    new_n14699_, new_n14700_, new_n14701_, new_n14702_, new_n14703_,
    new_n14704_, new_n14705_, new_n14706_, new_n14707_, new_n14708_,
    new_n14709_, new_n14710_, new_n14711_, new_n14712_, new_n14713_,
    new_n14714_, new_n14715_, new_n14716_, new_n14717_, new_n14718_,
    new_n14719_, new_n14720_, new_n14721_, new_n14722_, new_n14723_,
    new_n14724_, new_n14725_, new_n14726_, new_n14727_, new_n14728_,
    new_n14729_, new_n14730_, new_n14731_, new_n14732_, new_n14733_,
    new_n14734_, new_n14735_, new_n14736_, new_n14737_, new_n14738_,
    new_n14739_, new_n14740_, new_n14741_, new_n14742_, new_n14743_,
    new_n14744_, new_n14745_, new_n14746_, new_n14747_, new_n14748_,
    new_n14749_, new_n14750_, new_n14751_, new_n14752_, new_n14753_,
    new_n14754_, new_n14755_, new_n14756_, new_n14757_, new_n14758_,
    new_n14759_, new_n14760_, new_n14761_, new_n14762_, new_n14763_,
    new_n14764_, new_n14765_, new_n14766_, new_n14767_, new_n14768_,
    new_n14769_, new_n14770_, new_n14771_, new_n14772_, new_n14773_,
    new_n14774_, new_n14775_, new_n14776_, new_n14777_, new_n14778_,
    new_n14779_, new_n14780_, new_n14781_, new_n14782_, new_n14783_,
    new_n14784_, new_n14785_, new_n14786_, new_n14787_, new_n14788_,
    new_n14789_, new_n14790_, new_n14791_, new_n14792_, new_n14793_,
    new_n14794_, new_n14795_, new_n14796_, new_n14797_, new_n14798_,
    new_n14799_, new_n14800_, new_n14801_, new_n14802_, new_n14803_,
    new_n14804_, new_n14805_, new_n14806_, new_n14807_, new_n14808_,
    new_n14809_, new_n14810_, new_n14811_, new_n14812_, new_n14813_,
    new_n14814_, new_n14815_, new_n14816_, new_n14817_, new_n14818_,
    new_n14819_, new_n14820_, new_n14821_, new_n14822_, new_n14823_,
    new_n14824_, new_n14825_, new_n14826_, new_n14827_, new_n14828_,
    new_n14829_, new_n14830_, new_n14831_, new_n14832_, new_n14833_,
    new_n14834_, new_n14835_, new_n14836_, new_n14837_, new_n14838_,
    new_n14839_, new_n14840_, new_n14841_, new_n14842_, new_n14843_,
    new_n14844_, new_n14845_, new_n14846_, new_n14847_, new_n14848_,
    new_n14849_, new_n14850_, new_n14851_, new_n14852_, new_n14853_,
    new_n14854_, new_n14855_, new_n14856_, new_n14857_, new_n14858_,
    new_n14859_, new_n14860_, new_n14861_, new_n14862_, new_n14863_,
    new_n14864_, new_n14865_, new_n14866_, new_n14867_, new_n14868_,
    new_n14869_, new_n14870_, new_n14871_, new_n14872_, new_n14873_,
    new_n14874_, new_n14875_, new_n14876_, new_n14877_, new_n14878_,
    new_n14879_, new_n14880_, new_n14881_, new_n14882_, new_n14883_,
    new_n14884_, new_n14885_, new_n14886_, new_n14887_, new_n14888_,
    new_n14889_, new_n14890_, new_n14891_, new_n14892_, new_n14893_,
    new_n14894_, new_n14895_, new_n14896_, new_n14897_, new_n14898_,
    new_n14899_, new_n14900_, new_n14901_, new_n14902_, new_n14903_,
    new_n14904_, new_n14905_, new_n14906_, new_n14907_, new_n14908_,
    new_n14909_, new_n14910_, new_n14911_, new_n14912_, new_n14913_,
    new_n14914_, new_n14915_, new_n14916_, new_n14917_, new_n14918_,
    new_n14919_, new_n14920_, new_n14921_, new_n14922_, new_n14923_,
    new_n14924_, new_n14925_, new_n14926_, new_n14927_, new_n14928_,
    new_n14929_, new_n14930_, new_n14931_, new_n14932_, new_n14933_,
    new_n14934_, new_n14935_, new_n14936_, new_n14937_, new_n14938_,
    new_n14939_, new_n14940_, new_n14941_, new_n14942_, new_n14943_,
    new_n14944_, new_n14945_, new_n14946_, new_n14947_, new_n14948_,
    new_n14949_, new_n14950_, new_n14951_, new_n14952_, new_n14953_,
    new_n14954_, new_n14955_, new_n14956_, new_n14957_, new_n14958_,
    new_n14959_, new_n14960_, new_n14961_, new_n14962_, new_n14963_,
    new_n14964_, new_n14965_, new_n14966_, new_n14967_, new_n14968_,
    new_n14969_, new_n14970_, new_n14971_, new_n14972_, new_n14973_,
    new_n14974_, new_n14975_, new_n14976_, new_n14977_, new_n14978_,
    new_n14979_, new_n14980_, new_n14981_, new_n14982_, new_n14983_,
    new_n14984_, new_n14985_, new_n14986_, new_n14987_, new_n14988_,
    new_n14989_, new_n14990_, new_n14991_, new_n14992_, new_n14993_,
    new_n14994_, new_n14995_, new_n14996_, new_n14997_, new_n14998_,
    new_n14999_, new_n15000_, new_n15001_, new_n15002_, new_n15003_,
    new_n15004_, new_n15005_, new_n15006_, new_n15007_, new_n15008_,
    new_n15009_, new_n15010_, new_n15011_, new_n15012_, new_n15013_,
    new_n15014_, new_n15015_, new_n15016_, new_n15017_, new_n15018_,
    new_n15019_, new_n15020_, new_n15021_, new_n15022_, new_n15023_,
    new_n15024_, new_n15025_, new_n15027_, new_n15028_, new_n15029_,
    new_n15030_, new_n15031_, new_n15032_, new_n15033_, new_n15034_,
    new_n15035_, new_n15036_, new_n15037_, new_n15038_, new_n15039_,
    new_n15040_, new_n15041_, new_n15042_, new_n15043_, new_n15044_,
    new_n15045_, new_n15046_, new_n15047_, new_n15048_, new_n15049_,
    new_n15050_, new_n15051_, new_n15052_, new_n15053_, new_n15054_,
    new_n15055_, new_n15056_, new_n15057_, new_n15061_, new_n15062_,
    new_n15063_, new_n15064_, new_n15065_, new_n15066_, new_n15067_,
    new_n15068_, new_n15069_, new_n15070_, new_n15072_, new_n15074_,
    new_n15075_, new_n15076_, new_n15079_, new_n15081_, new_n15084_,
    new_n15085_, new_n15088_, new_n15092_, new_n15093_, new_n15094_,
    new_n15095_, new_n15096_, new_n15098_, new_n15100_, new_n15101_,
    new_n15103_, new_n15104_, new_n15105_, new_n15106_, new_n15108_,
    new_n15109_, new_n15110_, new_n15111_, new_n15115_, new_n15116_,
    new_n15117_, new_n15118_, new_n15119_, new_n15120_, new_n15121_,
    new_n15122_, new_n15123_, new_n15124_, new_n15125_, new_n15126_,
    new_n15133_, new_n15134_, new_n15135_, new_n15136_, new_n15137_,
    new_n15138_, new_n15140_, new_n15146_, new_n15147_, new_n15148_,
    new_n15149_, new_n15150_, new_n15151_, new_n15152_, new_n15153_,
    new_n15154_, new_n15155_, new_n15156_, new_n15158_, new_n15159_,
    new_n15160_, new_n15161_, new_n15162_, new_n15163_, new_n15164_,
    new_n15165_, new_n15166_, new_n15167_, new_n15168_, new_n15169_,
    new_n15170_, new_n15171_, new_n15172_, new_n15173_, new_n15174_,
    new_n15175_, new_n15176_, new_n15177_, new_n15178_, new_n15179_,
    new_n15180_, new_n15181_, new_n15182_, new_n15183_, new_n15184_,
    new_n15185_, new_n15186_, new_n15187_, new_n15188_, new_n15189_,
    new_n15190_, new_n15191_, new_n15192_, new_n15193_, new_n15194_,
    new_n15195_, new_n15196_, new_n15197_, new_n15198_, new_n15199_,
    new_n15200_, new_n15201_, new_n15202_, new_n15203_, new_n15204_,
    new_n15205_, new_n15206_, new_n15207_, new_n15208_, new_n15209_,
    new_n15210_, new_n15211_, new_n15212_, new_n15213_, new_n15214_,
    new_n15215_, new_n15216_, new_n15217_, new_n15218_, new_n15219_,
    new_n15220_, new_n15221_, new_n15222_, new_n15223_, new_n15224_,
    new_n15225_, new_n15226_, new_n15227_, new_n15228_, new_n15229_,
    new_n15230_, new_n15231_, new_n15232_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15369_,
    new_n15370_, new_n15371_, new_n15372_, new_n15373_, new_n15374_,
    new_n15375_, new_n15376_, new_n15377_, new_n15378_, new_n15379_,
    new_n15380_, new_n15381_, new_n15382_, new_n15383_, new_n15384_,
    new_n15385_, new_n15386_, new_n15387_, new_n15388_, new_n15389_,
    new_n15390_, new_n15391_, new_n15392_, new_n15393_, new_n15394_,
    new_n15395_, new_n15396_, new_n15397_, new_n15398_, new_n15399_,
    new_n15400_, new_n15401_, new_n15402_, new_n15403_, new_n15404_,
    new_n15405_, new_n15406_, new_n15407_, new_n15408_, new_n15409_,
    new_n15410_, new_n15411_, new_n15412_, new_n15413_, new_n15414_,
    new_n15415_, new_n15416_, new_n15417_, new_n15418_, new_n15419_,
    new_n15420_, new_n15421_, new_n15422_, new_n15423_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15428_, new_n15429_,
    new_n15430_, new_n15431_, new_n15432_, new_n15433_, new_n15434_,
    new_n15435_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15469_,
    new_n15470_, new_n15471_, new_n15472_, new_n15473_, new_n15474_,
    new_n15475_, new_n15476_, new_n15477_, new_n15478_, new_n15479_,
    new_n15480_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15488_, new_n15489_,
    new_n15490_, new_n15491_, new_n15492_, new_n15493_, new_n15494_,
    new_n15495_, new_n15496_, new_n15497_, new_n15498_, new_n15499_,
    new_n15500_, new_n15501_, new_n15502_, new_n15503_, new_n15504_,
    new_n15505_, new_n15506_, new_n15507_, new_n15508_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15575_, new_n15576_, new_n15577_, new_n15578_, new_n15579_,
    new_n15580_, new_n15581_, new_n15582_, new_n15583_, new_n15584_,
    new_n15585_, new_n15586_, new_n15587_, new_n15588_, new_n15589_,
    new_n15590_, new_n15591_, new_n15592_, new_n15593_, new_n15594_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15601_, new_n15602_, new_n15603_, new_n15604_,
    new_n15605_, new_n15606_, new_n15607_, new_n15608_, new_n15609_,
    new_n15610_, new_n15611_, new_n15612_, new_n15613_, new_n15614_,
    new_n15615_, new_n15616_, new_n15617_, new_n15618_, new_n15619_,
    new_n15620_, new_n15621_, new_n15622_, new_n15623_, new_n15624_,
    new_n15625_, new_n15626_, new_n15627_, new_n15628_, new_n15629_,
    new_n15630_, new_n15631_, new_n15632_, new_n15633_, new_n15634_,
    new_n15635_, new_n15636_, new_n15637_, new_n15638_, new_n15639_,
    new_n15640_, new_n15641_, new_n15642_, new_n15643_, new_n15644_,
    new_n15645_, new_n15646_, new_n15647_, new_n15648_, new_n15649_,
    new_n15650_, new_n15651_, new_n15652_, new_n15653_, new_n15654_,
    new_n15655_, new_n15656_, new_n15657_, new_n15658_, new_n15659_,
    new_n15660_, new_n15661_, new_n15662_, new_n15663_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15674_,
    new_n15675_, new_n15676_, new_n15677_, new_n15678_, new_n15679_,
    new_n15680_, new_n15681_, new_n15682_, new_n15683_, new_n15684_,
    new_n15685_, new_n15686_, new_n15687_, new_n15688_, new_n15689_,
    new_n15690_, new_n15691_, new_n15692_, new_n15693_, new_n15694_,
    new_n15695_, new_n15696_, new_n15697_, new_n15698_, new_n15699_,
    new_n15700_, new_n15701_, new_n15702_, new_n15703_, new_n15704_,
    new_n15705_, new_n15706_, new_n15707_, new_n15708_, new_n15709_,
    new_n15710_, new_n15711_, new_n15712_, new_n15713_, new_n15714_,
    new_n15715_, new_n15716_, new_n15717_, new_n15718_, new_n15719_,
    new_n15720_, new_n15721_, new_n15722_, new_n15723_, new_n15724_,
    new_n15725_, new_n15726_, new_n15727_, new_n15728_, new_n15729_,
    new_n15730_, new_n15731_, new_n15732_, new_n15733_, new_n15734_,
    new_n15735_, new_n15736_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15755_, new_n15756_, new_n15757_, new_n15758_, new_n15759_,
    new_n15760_, new_n15761_, new_n15762_, new_n15763_, new_n15764_,
    new_n15765_, new_n15766_, new_n15767_, new_n15768_, new_n15769_,
    new_n15770_, new_n15771_, new_n15772_, new_n15773_, new_n15774_,
    new_n15775_, new_n15776_, new_n15777_, new_n15778_, new_n15779_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15786_, new_n15787_, new_n15788_, new_n15789_,
    new_n15790_, new_n15791_, new_n15792_, new_n15793_, new_n15794_,
    new_n15795_, new_n15796_, new_n15797_, new_n15798_, new_n15799_,
    new_n15800_, new_n15801_, new_n15802_, new_n15803_, new_n15804_,
    new_n15805_, new_n15806_, new_n15807_, new_n15808_, new_n15809_,
    new_n15810_, new_n15811_, new_n15812_, new_n15813_, new_n15814_,
    new_n15815_, new_n15816_, new_n15817_, new_n15818_, new_n15819_,
    new_n15820_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15865_, new_n15866_, new_n15867_, new_n15868_, new_n15869_,
    new_n15870_, new_n15871_, new_n15872_, new_n15873_, new_n15874_,
    new_n15875_, new_n15876_, new_n15877_, new_n15878_, new_n15879_,
    new_n15880_, new_n15881_, new_n15882_, new_n15883_, new_n15884_,
    new_n15885_, new_n15886_, new_n15887_, new_n15888_, new_n15889_,
    new_n15890_, new_n15891_, new_n15892_, new_n15893_, new_n15894_,
    new_n15895_, new_n15896_, new_n15897_, new_n15898_, new_n15899_,
    new_n15900_, new_n15901_, new_n15902_, new_n15903_, new_n15904_,
    new_n15905_, new_n15906_, new_n15907_, new_n15908_, new_n15909_,
    new_n15910_, new_n15911_, new_n15912_, new_n15913_, new_n15914_,
    new_n15915_, new_n15916_, new_n15917_, new_n15918_, new_n15919_,
    new_n15920_, new_n15921_, new_n15922_, new_n15923_, new_n15924_,
    new_n15925_, new_n15926_, new_n15927_, new_n15928_, new_n15929_,
    new_n15930_, new_n15931_, new_n15932_, new_n15933_, new_n15934_,
    new_n15935_, new_n15936_, new_n15937_, new_n15938_, new_n15939_,
    new_n15940_, new_n15941_, new_n15942_, new_n15943_, new_n15944_,
    new_n15945_, new_n15946_, new_n15947_, new_n15948_, new_n15949_,
    new_n15950_, new_n15951_, new_n15952_, new_n15953_, new_n15954_,
    new_n15955_, new_n15956_, new_n15957_, new_n15958_, new_n15959_,
    new_n15960_, new_n15961_, new_n15962_, new_n15963_, new_n15964_,
    new_n15965_, new_n15966_, new_n15967_, new_n15968_, new_n15969_,
    new_n15970_, new_n15971_, new_n15972_, new_n15973_, new_n15974_,
    new_n15975_, new_n15976_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15987_, new_n15988_, new_n15989_,
    new_n15990_, new_n15991_, new_n15992_, new_n15993_, new_n15994_,
    new_n15995_, new_n15996_, new_n15997_, new_n15998_, new_n15999_,
    new_n16000_, new_n16001_, new_n16002_, new_n16003_, new_n16004_,
    new_n16005_, new_n16006_, new_n16007_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16012_, new_n16013_, new_n16014_,
    new_n16015_, new_n16016_, new_n16017_, new_n16018_, new_n16019_,
    new_n16020_, new_n16021_, new_n16022_, new_n16023_, new_n16024_,
    new_n16025_, new_n16026_, new_n16027_, new_n16028_, new_n16029_,
    new_n16030_, new_n16031_, new_n16032_, new_n16033_, new_n16034_,
    new_n16035_, new_n16036_, new_n16037_, new_n16038_, new_n16039_,
    new_n16040_, new_n16041_, new_n16042_, new_n16043_, new_n16044_,
    new_n16045_, new_n16046_, new_n16047_, new_n16048_, new_n16049_,
    new_n16050_, new_n16051_, new_n16052_, new_n16053_, new_n16054_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16060_, new_n16061_, new_n16062_, new_n16063_, new_n16064_,
    new_n16065_, new_n16066_, new_n16067_, new_n16068_, new_n16069_,
    new_n16070_, new_n16071_, new_n16072_, new_n16073_, new_n16074_,
    new_n16075_, new_n16076_, new_n16077_, new_n16078_, new_n16079_,
    new_n16080_, new_n16081_, new_n16082_, new_n16083_, new_n16084_,
    new_n16085_, new_n16086_, new_n16087_, new_n16088_, new_n16089_,
    new_n16090_, new_n16091_, new_n16092_, new_n16093_, new_n16094_,
    new_n16095_, new_n16096_, new_n16097_, new_n16098_, new_n16099_,
    new_n16100_, new_n16101_, new_n16102_, new_n16103_, new_n16104_,
    new_n16105_, new_n16106_, new_n16107_, new_n16108_, new_n16109_,
    new_n16110_, new_n16111_, new_n16112_, new_n16113_, new_n16114_,
    new_n16115_, new_n16116_, new_n16117_, new_n16118_, new_n16119_,
    new_n16120_, new_n16121_, new_n16122_, new_n16123_, new_n16124_,
    new_n16125_, new_n16126_, new_n16127_, new_n16128_, new_n16129_,
    new_n16130_, new_n16131_, new_n16132_, new_n16133_, new_n16134_,
    new_n16135_, new_n16136_, new_n16137_, new_n16138_, new_n16139_,
    new_n16140_, new_n16141_, new_n16142_, new_n16143_, new_n16144_,
    new_n16145_, new_n16146_, new_n16147_, new_n16148_, new_n16149_,
    new_n16150_, new_n16151_, new_n16152_, new_n16153_, new_n16154_,
    new_n16155_, new_n16156_, new_n16157_, new_n16158_, new_n16159_,
    new_n16160_, new_n16161_, new_n16162_, new_n16163_, new_n16164_,
    new_n16165_, new_n16166_, new_n16167_, new_n16168_, new_n16169_,
    new_n16170_, new_n16171_, new_n16172_, new_n16173_, new_n16174_,
    new_n16175_, new_n16176_, new_n16177_, new_n16178_, new_n16179_,
    new_n16180_, new_n16181_, new_n16182_, new_n16183_, new_n16184_,
    new_n16185_, new_n16186_, new_n16187_, new_n16188_, new_n16189_,
    new_n16190_, new_n16191_, new_n16192_, new_n16193_, new_n16194_,
    new_n16195_, new_n16196_, new_n16197_, new_n16198_, new_n16199_,
    new_n16200_, new_n16201_, new_n16202_, new_n16203_, new_n16204_,
    new_n16205_, new_n16206_, new_n16207_, new_n16208_, new_n16209_,
    new_n16210_, new_n16211_, new_n16212_, new_n16213_, new_n16214_,
    new_n16215_, new_n16216_, new_n16217_, new_n16218_, new_n16219_,
    new_n16220_, new_n16221_, new_n16222_, new_n16223_, new_n16224_,
    new_n16225_, new_n16226_, new_n16227_, new_n16228_, new_n16229_,
    new_n16230_, new_n16231_, new_n16232_, new_n16233_, new_n16234_,
    new_n16235_, new_n16236_, new_n16237_, new_n16238_, new_n16239_,
    new_n16240_, new_n16241_, new_n16242_, new_n16243_, new_n16244_,
    new_n16245_, new_n16246_, new_n16247_, new_n16248_, new_n16249_,
    new_n16250_, new_n16251_, new_n16252_, new_n16253_, new_n16254_,
    new_n16255_, new_n16256_, new_n16257_, new_n16258_, new_n16259_,
    new_n16260_, new_n16261_, new_n16262_, new_n16263_, new_n16264_,
    new_n16265_, new_n16266_, new_n16267_, new_n16268_, new_n16269_,
    new_n16270_, new_n16271_, new_n16272_, new_n16273_, new_n16274_,
    new_n16275_, new_n16276_, new_n16277_, new_n16278_, new_n16279_,
    new_n16280_, new_n16281_, new_n16282_, new_n16283_, new_n16284_,
    new_n16285_, new_n16286_, new_n16287_, new_n16288_, new_n16289_,
    new_n16290_, new_n16291_, new_n16292_, new_n16293_, new_n16294_,
    new_n16295_, new_n16296_, new_n16297_, new_n16298_, new_n16299_,
    new_n16300_, new_n16301_, new_n16302_, new_n16303_, new_n16304_,
    new_n16305_, new_n16306_, new_n16307_, new_n16308_, new_n16309_,
    new_n16310_, new_n16311_, new_n16312_, new_n16313_, new_n16314_,
    new_n16315_, new_n16316_, new_n16317_, new_n16318_, new_n16319_,
    new_n16320_, new_n16321_, new_n16322_, new_n16323_, new_n16324_,
    new_n16325_, new_n16326_, new_n16327_, new_n16328_, new_n16329_,
    new_n16330_, new_n16331_, new_n16332_, new_n16333_, new_n16334_,
    new_n16335_, new_n16336_, new_n16337_, new_n16338_, new_n16339_,
    new_n16340_, new_n16341_, new_n16342_, new_n16343_, new_n16344_,
    new_n16345_, new_n16346_, new_n16347_, new_n16348_, new_n16349_,
    new_n16350_, new_n16351_, new_n16352_, new_n16353_, new_n16354_,
    new_n16355_, new_n16356_, new_n16357_, new_n16358_, new_n16359_,
    new_n16360_, new_n16361_, new_n16362_, new_n16363_, new_n16364_,
    new_n16365_, new_n16366_, new_n16367_, new_n16368_, new_n16369_,
    new_n16370_, new_n16371_, new_n16372_, new_n16373_, new_n16374_,
    new_n16375_, new_n16376_, new_n16377_, new_n16378_, new_n16379_,
    new_n16380_, new_n16381_, new_n16382_, new_n16383_, new_n16384_,
    new_n16385_, new_n16386_, new_n16387_, new_n16388_, new_n16389_,
    new_n16390_, new_n16391_, new_n16392_, new_n16393_, new_n16394_,
    new_n16395_, new_n16396_, new_n16397_, new_n16398_, new_n16399_,
    new_n16400_, new_n16401_, new_n16402_, new_n16403_, new_n16404_,
    new_n16405_, new_n16406_, new_n16407_, new_n16408_, new_n16409_,
    new_n16410_, new_n16411_, new_n16412_, new_n16413_, new_n16414_,
    new_n16415_, new_n16416_, new_n16417_, new_n16418_, new_n16419_,
    new_n16420_, new_n16421_, new_n16422_, new_n16423_, new_n16424_,
    new_n16425_, new_n16426_, new_n16427_, new_n16428_, new_n16429_,
    new_n16430_, new_n16431_, new_n16432_, new_n16433_, new_n16434_,
    new_n16435_, new_n16436_, new_n16437_, new_n16438_, new_n16439_,
    new_n16440_, new_n16441_, new_n16442_, new_n16443_, new_n16444_,
    new_n16445_, new_n16446_, new_n16447_, new_n16448_, new_n16449_,
    new_n16450_, new_n16451_, new_n16452_, new_n16453_, new_n16454_,
    new_n16455_, new_n16456_, new_n16457_, new_n16458_, new_n16459_,
    new_n16460_, new_n16461_, new_n16462_, new_n16463_, new_n16464_,
    new_n16465_, new_n16466_, new_n16467_, new_n16468_, new_n16469_,
    new_n16470_, new_n16471_, new_n16472_, new_n16473_, new_n16474_,
    new_n16475_, new_n16476_, new_n16477_, new_n16478_, new_n16479_,
    new_n16480_, new_n16481_, new_n16482_, new_n16483_, new_n16484_,
    new_n16485_, new_n16486_, new_n16487_, new_n16488_, new_n16489_,
    new_n16490_, new_n16491_, new_n16492_, new_n16493_, new_n16494_,
    new_n16495_, new_n16496_, new_n16497_, new_n16498_, new_n16499_,
    new_n16500_, new_n16501_, new_n16502_, new_n16503_, new_n16504_,
    new_n16505_, new_n16506_, new_n16507_, new_n16508_, new_n16509_,
    new_n16510_, new_n16511_, new_n16512_, new_n16513_, new_n16514_,
    new_n16515_, new_n16516_, new_n16517_, new_n16518_, new_n16519_,
    new_n16520_, new_n16521_, new_n16522_, new_n16523_, new_n16524_,
    new_n16525_, new_n16526_, new_n16527_, new_n16528_, new_n16529_,
    new_n16530_, new_n16531_, new_n16532_, new_n16533_, new_n16534_,
    new_n16535_, new_n16536_, new_n16537_, new_n16538_, new_n16539_,
    new_n16540_, new_n16541_, new_n16542_, new_n16543_, new_n16544_,
    new_n16545_, new_n16546_, new_n16547_, new_n16548_, new_n16549_,
    new_n16550_, new_n16551_, new_n16552_, new_n16553_, new_n16554_,
    new_n16555_, new_n16556_, new_n16557_, new_n16558_, new_n16559_,
    new_n16560_, new_n16561_, new_n16562_, new_n16563_, new_n16564_,
    new_n16565_, new_n16566_, new_n16567_, new_n16568_, new_n16569_,
    new_n16570_, new_n16571_, new_n16572_, new_n16573_, new_n16574_,
    new_n16575_, new_n16576_, new_n16577_, new_n16578_, new_n16579_,
    new_n16580_, new_n16581_, new_n16582_, new_n16583_, new_n16584_,
    new_n16585_, new_n16586_, new_n16587_, new_n16588_, new_n16589_,
    new_n16590_, new_n16591_, new_n16592_, new_n16593_, new_n16594_,
    new_n16595_, new_n16596_, new_n16597_, new_n16598_, new_n16599_,
    new_n16600_, new_n16601_, new_n16602_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16610_, new_n16611_, new_n16612_, new_n16613_, new_n16614_,
    new_n16615_, new_n16616_, new_n16617_, new_n16618_, new_n16619_,
    new_n16620_, new_n16621_, new_n16622_, new_n16623_, new_n16624_,
    new_n16625_, new_n16626_, new_n16627_, new_n16628_, new_n16629_,
    new_n16630_, new_n16631_, new_n16632_, new_n16633_, new_n16634_,
    new_n16635_, new_n16636_, new_n16637_, new_n16638_, new_n16639_,
    new_n16640_, new_n16641_, new_n16642_, new_n16643_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16650_, new_n16651_, new_n16652_, new_n16653_, new_n16654_,
    new_n16655_, new_n16656_, new_n16657_, new_n16658_, new_n16659_,
    new_n16660_, new_n16661_, new_n16662_, new_n16663_, new_n16664_,
    new_n16665_, new_n16666_, new_n16667_, new_n16668_, new_n16669_,
    new_n16670_, new_n16671_, new_n16672_, new_n16673_, new_n16674_,
    new_n16675_, new_n16676_, new_n16677_, new_n16678_, new_n16679_,
    new_n16680_, new_n16681_, new_n16682_, new_n16683_, new_n16684_,
    new_n16685_, new_n16686_, new_n16687_, new_n16688_, new_n16689_,
    new_n16690_, new_n16691_, new_n16692_, new_n16693_, new_n16694_,
    new_n16695_, new_n16696_, new_n16697_, new_n16698_, new_n16699_,
    new_n16700_, new_n16701_, new_n16702_, new_n16703_, new_n16704_,
    new_n16705_, new_n16706_, new_n16707_, new_n16708_, new_n16709_,
    new_n16710_, new_n16711_, new_n16712_, new_n16713_, new_n16714_,
    new_n16715_, new_n16716_, new_n16717_, new_n16718_, new_n16719_,
    new_n16720_, new_n16721_, new_n16722_, new_n16723_, new_n16724_,
    new_n16725_, new_n16726_, new_n16727_, new_n16728_, new_n16729_,
    new_n16730_, new_n16731_, new_n16732_, new_n16733_, new_n16734_,
    new_n16735_, new_n16736_, new_n16737_, new_n16738_, new_n16739_,
    new_n16740_, new_n16741_, new_n16742_, new_n16743_, new_n16744_,
    new_n16745_, new_n16746_, new_n16747_, new_n16748_, new_n16749_,
    new_n16750_, new_n16751_, new_n16752_, new_n16753_, new_n16754_,
    new_n16755_, new_n16756_, new_n16757_, new_n16758_, new_n16759_,
    new_n16760_, new_n16761_, new_n16762_, new_n16763_, new_n16764_,
    new_n16765_, new_n16766_, new_n16767_, new_n16768_, new_n16769_,
    new_n16770_, new_n16771_, new_n16772_, new_n16773_, new_n16774_,
    new_n16775_, new_n16776_, new_n16777_, new_n16778_, new_n16779_,
    new_n16780_, new_n16781_, new_n16782_, new_n16783_, new_n16784_,
    new_n16785_, new_n16786_, new_n16787_, new_n16788_, new_n16789_,
    new_n16790_, new_n16791_, new_n16792_, new_n16793_, new_n16794_,
    new_n16795_, new_n16796_, new_n16797_, new_n16798_, new_n16799_,
    new_n16800_, new_n16801_, new_n16802_, new_n16803_, new_n16804_,
    new_n16805_, new_n16806_, new_n16807_, new_n16808_, new_n16809_,
    new_n16810_, new_n16811_, new_n16812_, new_n16813_, new_n16814_,
    new_n16815_, new_n16816_, new_n16817_, new_n16818_, new_n16819_,
    new_n16820_, new_n16821_, new_n16822_, new_n16823_, new_n16824_,
    new_n16825_, new_n16826_, new_n16827_, new_n16828_, new_n16829_,
    new_n16830_, new_n16831_, new_n16832_, new_n16833_, new_n16834_,
    new_n16835_, new_n16836_, new_n16837_, new_n16838_, new_n16839_,
    new_n16840_, new_n16841_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16848_, new_n16849_,
    new_n16850_, new_n16851_, new_n16852_, new_n16853_, new_n16854_,
    new_n16855_, new_n16856_, new_n16857_, new_n16858_, new_n16859_,
    new_n16860_, new_n16861_, new_n16862_, new_n16863_, new_n16864_,
    new_n16865_, new_n16866_, new_n16867_, new_n16868_, new_n16869_,
    new_n16870_, new_n16871_, new_n16872_, new_n16873_, new_n16874_,
    new_n16875_, new_n16876_, new_n16877_, new_n16878_, new_n16879_,
    new_n16880_, new_n16881_, new_n16882_, new_n16883_, new_n16884_,
    new_n16885_, new_n16886_, new_n16887_, new_n16888_, new_n16889_,
    new_n16890_, new_n16891_, new_n16892_, new_n16893_, new_n16894_,
    new_n16895_, new_n16896_, new_n16897_, new_n16898_, new_n16899_,
    new_n16900_, new_n16901_, new_n16902_, new_n16903_, new_n16904_,
    new_n16905_, new_n16906_, new_n16907_, new_n16908_, new_n16909_,
    new_n16910_, new_n16911_, new_n16912_, new_n16913_, new_n16914_,
    new_n16915_, new_n16916_, new_n16917_, new_n16918_, new_n16919_,
    new_n16920_, new_n16921_, new_n16922_, new_n16923_, new_n16924_,
    new_n16925_, new_n16926_, new_n16927_, new_n16928_, new_n16929_,
    new_n16930_, new_n16931_, new_n16932_, new_n16933_, new_n16934_,
    new_n16935_, new_n16936_, new_n16937_, new_n16938_, new_n16939_,
    new_n16940_, new_n16941_, new_n16942_, new_n16943_, new_n16944_,
    new_n16945_, new_n16946_, new_n16947_, new_n16948_, new_n16949_,
    new_n16950_, new_n16951_, new_n16952_, new_n16953_, new_n16954_,
    new_n16955_, new_n16956_, new_n16957_, new_n16958_, new_n16959_,
    new_n16960_, new_n16961_, new_n16962_, new_n16963_, new_n16964_,
    new_n16965_, new_n16966_, new_n16967_, new_n16968_, new_n16969_,
    new_n16970_, new_n16971_, new_n16972_, new_n16973_, new_n16974_,
    new_n16975_, new_n16976_, new_n16977_, new_n16978_, new_n16979_,
    new_n16981_, new_n16982_, new_n16983_, new_n16984_, new_n16986_,
    new_n16987_, new_n16988_, new_n16989_, new_n16990_, new_n16991_,
    new_n16993_, new_n16995_, new_n16996_, new_n16997_, new_n16998_,
    new_n16999_, new_n17001_, new_n17002_, new_n17003_, new_n17004_,
    new_n17006_, new_n17007_, new_n17008_, new_n17009_, new_n17011_,
    new_n17012_, new_n17013_, new_n17014_, new_n17015_, new_n17016_,
    new_n17018_, new_n17020_, new_n17021_, new_n17022_, new_n17023_,
    new_n17024_, new_n17026_, new_n17027_, new_n17028_, new_n17029_,
    new_n17031_, new_n17032_, new_n17034_, new_n17035_, new_n17036_,
    new_n17037_, new_n17038_, new_n17039_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17090_, new_n17091_, new_n17092_, new_n17093_, new_n17094_,
    new_n17095_, new_n17096_, new_n17097_, new_n17098_, new_n17099_,
    new_n17100_, new_n17101_, new_n17102_, new_n17103_, new_n17104_,
    new_n17105_, new_n17106_, new_n17107_, new_n17108_, new_n17109_,
    new_n17110_, new_n17111_, new_n17112_, new_n17114_, new_n17115_,
    new_n17116_, new_n17117_, new_n17118_, new_n17119_, new_n17120_,
    new_n17121_, new_n17122_, new_n17123_, new_n17124_, new_n17125_,
    new_n17126_, new_n17127_, new_n17128_, new_n17129_, new_n17131_,
    new_n17132_, new_n17133_, new_n17134_, new_n17135_, new_n17136_,
    new_n17137_, new_n17138_, new_n17139_, new_n17140_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17166_, new_n17167_,
    new_n17168_, new_n17169_, new_n17170_, new_n17171_, new_n17172_,
    new_n17173_, new_n17174_, new_n17175_, new_n17176_, new_n17177_,
    new_n17178_, new_n17179_, new_n17180_, new_n17181_, new_n17182_,
    new_n17183_, new_n17184_, new_n17185_, new_n17186_, new_n17187_,
    new_n17188_, new_n17189_, new_n17190_, new_n17191_, new_n17192_,
    new_n17193_, new_n17194_, new_n17195_, new_n17196_, new_n17197_,
    new_n17198_, new_n17199_, new_n17200_, new_n17201_, new_n17202_,
    new_n17203_, new_n17204_, new_n17205_, new_n17206_, new_n17207_,
    new_n17208_, new_n17209_, new_n17210_, new_n17211_, new_n17212_,
    new_n17213_, new_n17214_, new_n17215_, new_n17216_, new_n17217_,
    new_n17218_, new_n17219_, new_n17220_, new_n17221_, new_n17222_,
    new_n17223_, new_n17224_, new_n17225_, new_n17226_, new_n17227_,
    new_n17228_, new_n17229_, new_n17230_, new_n17231_, new_n17232_,
    new_n17233_, new_n17234_, new_n17235_, new_n17236_, new_n17237_,
    new_n17238_, new_n17239_, new_n17240_, new_n17241_, new_n17242_,
    new_n17243_, new_n17244_, new_n17245_, new_n17246_, new_n17247_,
    new_n17248_, new_n17249_, new_n17250_, new_n17251_, new_n17252_,
    new_n17253_, new_n17254_, new_n17255_, new_n17256_, new_n17257_,
    new_n17258_, new_n17259_, new_n17260_, new_n17261_, new_n17262_,
    new_n17263_, new_n17264_, new_n17265_, new_n17266_, new_n17267_,
    new_n17268_, new_n17269_, new_n17270_, new_n17271_, new_n17272_,
    new_n17273_, new_n17274_, new_n17275_, new_n17276_, new_n17277_,
    new_n17278_, new_n17279_, new_n17280_, new_n17281_, new_n17282_,
    new_n17283_, new_n17284_, new_n17285_, new_n17286_, new_n17287_,
    new_n17288_, new_n17289_, new_n17290_, new_n17291_, new_n17292_,
    new_n17293_, new_n17294_, new_n17295_, new_n17296_, new_n17297_,
    new_n17298_, new_n17299_, new_n17300_, new_n17301_, new_n17302_,
    new_n17303_, new_n17304_, new_n17305_, new_n17306_, new_n17307_,
    new_n17308_, new_n17309_, new_n17310_, new_n17311_, new_n17312_,
    new_n17313_, new_n17314_, new_n17315_, new_n17316_, new_n17317_,
    new_n17318_, new_n17319_, new_n17320_, new_n17321_, new_n17322_,
    new_n17323_, new_n17324_, new_n17325_, new_n17326_, new_n17327_,
    new_n17328_, new_n17329_, new_n17330_, new_n17331_, new_n17332_,
    new_n17333_, new_n17334_, new_n17335_, new_n17336_, new_n17337_,
    new_n17338_, new_n17339_, new_n17340_, new_n17341_, new_n17342_,
    new_n17343_, new_n17344_, new_n17345_, new_n17346_, new_n17347_,
    new_n17348_, new_n17349_, new_n17350_, new_n17351_, new_n17352_,
    new_n17353_, new_n17354_, new_n17355_, new_n17356_, new_n17357_,
    new_n17359_, new_n17360_, new_n17361_, new_n17364_, new_n17365_,
    new_n17368_, new_n17369_, new_n17370_, new_n17372_, new_n17373_,
    new_n17374_, new_n17375_, new_n17377_, new_n17378_, new_n17379_,
    new_n17380_, new_n17381_, new_n17382_, new_n17384_, new_n17385_,
    new_n17386_, new_n17387_, new_n17388_, new_n17390_, new_n17391_,
    new_n17392_, new_n17393_, new_n17394_, new_n17395_, new_n17397_,
    new_n17398_, new_n17399_, new_n17401_, new_n17402_, new_n17405_,
    new_n17406_, new_n17407_, new_n17409_, new_n17410_, new_n17411_,
    new_n17412_, new_n17413_, new_n17415_, new_n17416_, new_n17417_,
    new_n17418_, new_n17419_, new_n17421_, new_n17422_, new_n17423_,
    new_n17424_, new_n17425_, new_n17427_, new_n17428_, new_n17429_,
    new_n17430_, new_n17431_, new_n17433_, new_n17434_, new_n17435_,
    new_n17436_, new_n17437_, new_n17439_, new_n17440_, new_n17441_,
    new_n17442_, new_n17443_, new_n17445_, new_n17446_, new_n17447_,
    new_n17448_, new_n17449_, new_n17451_, new_n17452_, new_n17453_,
    new_n17454_, new_n17455_, new_n17457_, new_n17458_, new_n17459_,
    new_n17460_, new_n17461_, new_n17463_, new_n17464_, new_n17465_,
    new_n17466_, new_n17467_, new_n17469_, new_n17470_, new_n17471_,
    new_n17472_, new_n17473_, new_n17475_, new_n17476_, new_n17477_,
    new_n17478_, new_n17479_, new_n17481_, new_n17482_, new_n17483_,
    new_n17484_, new_n17485_, new_n17487_, new_n17488_, new_n17489_,
    new_n17490_, new_n17491_, new_n17493_, new_n17494_, new_n17495_,
    new_n17496_, new_n17497_, new_n17499_, new_n17500_, new_n17501_,
    new_n17502_, new_n17503_, new_n17505_, new_n17506_, new_n17507_,
    new_n17508_, new_n17509_, new_n17511_, new_n17512_, new_n17513_,
    new_n17514_, new_n17515_, new_n17517_, new_n17518_, new_n17519_,
    new_n17520_, new_n17521_, new_n17523_, new_n17524_, new_n17525_,
    new_n17526_, new_n17527_, new_n17529_, new_n17530_, new_n17531_,
    new_n17532_, new_n17533_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17541_, new_n17542_, new_n17543_,
    new_n17544_, new_n17545_, new_n17547_, new_n17548_, new_n17549_,
    new_n17550_, new_n17551_, new_n17553_, new_n17554_, new_n17555_,
    new_n17556_, new_n17557_, new_n17559_, new_n17560_, new_n17561_,
    new_n17562_, new_n17563_, new_n17565_, new_n17566_, new_n17567_,
    new_n17568_, new_n17569_, new_n17571_, new_n17572_, new_n17573_,
    new_n17574_, new_n17575_, new_n17577_, new_n17578_, new_n17579_,
    new_n17580_, new_n17582_, new_n17583_, new_n17584_, new_n17585_,
    new_n17587_, new_n17588_, new_n17589_, new_n17590_, new_n17592_,
    new_n17594_, new_n17595_, new_n17597_, new_n17598_, new_n17600_,
    new_n17602_, new_n17603_, new_n17605_, new_n17606_, new_n17608_,
    new_n17610_, new_n17611_, new_n17613_, new_n17614_, new_n17616_,
    new_n17617_, new_n17618_, new_n17619_, new_n17620_, new_n17622_,
    new_n17624_, new_n17625_, new_n17626_, new_n17627_, new_n17628_,
    new_n17630_, new_n17631_, new_n17632_, new_n17633_, new_n17634_,
    new_n17636_, new_n17637_, new_n17639_, new_n17640_, new_n17641_,
    new_n17642_, new_n17643_, new_n17644_, new_n17645_, new_n17646_,
    new_n17647_, new_n17648_, new_n17650_, new_n17651_, new_n17652_,
    new_n17654_, new_n17655_, new_n17656_, new_n17657_, new_n17658_,
    new_n17659_, new_n17660_, new_n17661_, new_n17662_, new_n17664_,
    new_n17665_, new_n17666_, new_n17667_, new_n17668_, new_n17669_,
    new_n17672_, new_n17673_, new_n17674_, new_n17675_, new_n17676_,
    new_n17680_, new_n17681_, new_n17682_, new_n17684_, new_n17685_,
    new_n17686_, new_n17688_, new_n17689_, new_n17690_, new_n17691_,
    new_n17692_, new_n17693_, new_n17694_, new_n17695_, new_n17696_,
    new_n17697_, new_n17698_, new_n17699_, new_n17700_, new_n17702_,
    new_n17703_, new_n17704_, new_n17705_, new_n17706_, new_n17707_,
    new_n17708_, new_n17709_, new_n17710_, new_n17711_, new_n17712_,
    new_n17713_, new_n17714_, new_n17715_, new_n17716_, new_n17717_,
    new_n17718_, new_n17719_, new_n17720_, new_n17721_, new_n17722_,
    new_n17723_, new_n17724_, new_n17725_, new_n17726_, new_n17727_,
    new_n17728_, new_n17729_, new_n17730_, new_n17731_, new_n17732_,
    new_n17733_, new_n17735_, new_n17736_, new_n17737_, new_n17738_,
    new_n17739_, new_n17740_, new_n17742_, new_n17743_, new_n17744_,
    new_n17745_, new_n17746_, new_n17747_, new_n17748_, new_n17749_,
    new_n17750_, new_n17751_, new_n17752_, new_n17753_, new_n17754_,
    new_n17755_, new_n17756_, new_n17757_, new_n17758_, new_n17759_,
    new_n17760_, new_n17761_, new_n17763_, new_n17764_, new_n17765_,
    new_n17766_, new_n17767_, new_n17768_, new_n17771_, new_n17772_,
    new_n17773_, new_n17775_, new_n17776_, new_n17777_, new_n17778_,
    new_n17779_, new_n17780_, new_n17781_, new_n17782_, new_n17783_,
    new_n17784_, new_n17785_, new_n17786_, new_n17787_, new_n17788_,
    new_n17789_, new_n17790_, new_n17791_, new_n17792_, new_n17793_,
    new_n17794_, new_n17795_, new_n17796_, new_n17797_, new_n17798_,
    new_n17799_, new_n17800_, new_n17801_, new_n17802_, new_n17803_,
    new_n17804_, new_n17805_, new_n17806_, new_n17807_, new_n17808_,
    new_n17809_, new_n17810_, new_n17811_, new_n17812_, new_n17813_,
    new_n17814_, new_n17815_, new_n17816_, new_n17817_, new_n17818_,
    new_n17819_, new_n17820_, new_n17821_, new_n17822_, new_n17823_,
    new_n17824_, new_n17825_, new_n17826_, new_n17827_, new_n17828_,
    new_n17829_, new_n17830_, new_n17831_, new_n17832_, new_n17833_,
    new_n17834_, new_n17835_, new_n17836_, new_n17837_, new_n17839_,
    new_n17840_, new_n17841_, new_n17844_, new_n17845_, new_n17846_,
    new_n17847_, new_n17848_, new_n17849_, new_n17851_, new_n17852_,
    new_n17853_, new_n17855_, new_n17856_, new_n17857_, new_n17858_,
    new_n17860_, new_n17861_, new_n17862_, new_n17865_, new_n17866_,
    new_n17867_, new_n17868_, new_n17869_, new_n17870_, new_n17871_,
    new_n17872_, new_n17873_, new_n17874_, new_n17875_, new_n17876_,
    new_n17877_, new_n17878_, new_n17879_, new_n17880_, new_n17881_,
    new_n17882_, new_n17883_, new_n17884_, new_n17885_, new_n17886_,
    new_n17887_, new_n17888_, new_n17889_, new_n17890_, new_n17891_,
    new_n17892_, new_n17893_, new_n17894_, new_n17895_, new_n17896_,
    new_n17897_, new_n17898_, new_n17899_, new_n17900_, new_n17901_,
    new_n17902_, new_n17903_, new_n17904_, new_n17905_, new_n17906_,
    new_n17907_, new_n17908_, new_n17909_, new_n17910_, new_n17911_,
    new_n17912_, new_n17913_, new_n17914_, new_n17915_, new_n17916_,
    new_n17917_, new_n17918_, new_n17919_, new_n17920_, new_n17921_,
    new_n17922_, new_n17923_, new_n17924_, new_n17925_, new_n17926_,
    new_n17927_, new_n17928_, new_n17929_, new_n17930_, new_n17931_,
    new_n17932_, new_n17933_, new_n17934_, new_n17935_, new_n17936_,
    new_n17937_, new_n17938_, new_n17939_, new_n17940_, new_n17941_,
    new_n17942_, new_n17943_, new_n17944_, new_n17945_, new_n17946_,
    new_n17947_, new_n17948_, new_n17949_, new_n17950_, new_n17951_,
    new_n17952_, new_n17953_, new_n17954_, new_n17955_, new_n17956_,
    new_n17957_, new_n17958_, new_n17959_, new_n17960_, new_n17961_,
    new_n17962_, new_n17963_, new_n17964_, new_n17965_, new_n17966_,
    new_n17967_, new_n17968_, new_n17969_, new_n17970_, new_n17971_,
    new_n17972_, new_n17973_, new_n17974_, new_n17975_, new_n17976_,
    new_n17978_, new_n17979_, new_n17980_, new_n17981_, new_n17982_,
    new_n17983_, new_n17984_, new_n17985_, new_n17986_, new_n17987_,
    new_n17990_, new_n17991_, new_n17992_, new_n17993_, new_n17994_,
    new_n17995_, new_n17996_, new_n17999_, new_n18000_, new_n18001_,
    new_n18003_, new_n18004_, new_n18005_, new_n18006_, new_n18007_,
    new_n18008_, new_n18009_, new_n18010_, new_n18011_, new_n18012_,
    new_n18013_, new_n18014_, new_n18016_, new_n18017_, new_n18019_,
    new_n18020_, new_n18022_, new_n18023_, new_n18024_, new_n18025_,
    new_n18026_, new_n18027_, new_n18028_, new_n18029_, new_n18030_,
    new_n18031_, new_n18033_, new_n18034_, new_n18035_, new_n18037_,
    new_n18038_, new_n18039_, new_n18040_, new_n18041_, new_n18042_,
    new_n18043_, new_n18044_, new_n18045_, new_n18046_, new_n18048_,
    new_n18049_, new_n18050_, new_n18052_, new_n18055_, new_n18056_,
    new_n18057_, new_n18058_, new_n18059_, new_n18061_, new_n18062_,
    new_n18063_, new_n18064_, new_n18065_, new_n18066_, new_n18068_,
    new_n18069_, new_n18071_, new_n18072_, new_n18073_, new_n18075_,
    new_n18076_, new_n18077_, new_n18079_, new_n18080_, new_n18081_,
    new_n18083_, new_n18084_, new_n18085_, new_n18087_, new_n18088_,
    new_n18089_, new_n18091_, new_n18092_, new_n18093_, new_n18095_,
    new_n18096_, new_n18097_, new_n18099_, new_n18100_, new_n18101_,
    new_n18103_, new_n18104_, new_n18105_, new_n18107_, new_n18108_,
    new_n18109_, new_n18111_, new_n18112_, new_n18113_, new_n18115_,
    new_n18116_, new_n18117_, new_n18119_, new_n18120_, new_n18121_,
    new_n18123_, new_n18124_, new_n18125_, new_n18127_, new_n18128_,
    new_n18129_, new_n18130_, new_n18131_, new_n18132_, new_n18133_,
    new_n18134_, new_n18135_, new_n18136_, new_n18137_, new_n18138_,
    new_n18139_, new_n18140_, new_n18141_, new_n18142_, new_n18143_,
    new_n18144_, new_n18145_, new_n18147_, new_n18149_, new_n18150_,
    new_n18151_, new_n18152_, new_n18153_, new_n18154_, new_n18155_,
    new_n18156_, new_n18157_, new_n18158_, new_n18159_, new_n18161_,
    new_n18163_, new_n18164_, new_n18165_, new_n18167_, new_n18168_,
    new_n18169_, new_n18170_, new_n18171_, new_n18173_, new_n18175_,
    new_n18176_, new_n18177_, new_n18178_, new_n18179_, new_n18180_,
    new_n18181_, new_n18183_, new_n18185_, new_n18186_, new_n18187_,
    new_n18189_, new_n18190_, new_n18191_, new_n18192_, new_n18193_,
    new_n18194_, new_n18195_, new_n18197_, new_n18199_, new_n18200_,
    new_n18201_, new_n18203_, new_n18204_, new_n18205_, new_n18206_,
    new_n18207_, new_n18208_, new_n18209_, new_n18211_, new_n18212_,
    new_n18213_, new_n18214_, new_n18215_, new_n18216_, new_n18217_,
    new_n18218_, new_n18219_, new_n18220_, new_n18221_, new_n18222_,
    new_n18223_, new_n18224_, new_n18226_, new_n18227_, new_n18229_,
    new_n18230_, new_n18231_, new_n18233_, new_n18234_, new_n18235_,
    new_n18236_, new_n18238_, new_n18239_, new_n18240_, new_n18241_,
    new_n18242_, new_n18243_, new_n18244_, new_n18246_, new_n18248_,
    new_n18249_, new_n18250_, new_n18252_, new_n18253_, new_n18254_,
    new_n18255_, new_n18257_, new_n18258_, new_n18260_, new_n18261_,
    new_n18262_, new_n18263_, new_n18265_, new_n18266_, new_n18267_,
    new_n18268_, new_n18269_, new_n18270_, new_n18271_, new_n18273_,
    new_n18275_, new_n18276_, new_n18277_, new_n18279_, new_n18280_,
    new_n18281_, new_n18282_, new_n18284_, new_n18285_, new_n18287_,
    new_n18288_, new_n18289_, new_n18290_, new_n18292_, new_n18293_,
    new_n18294_, new_n18295_, new_n18296_, new_n18297_, new_n18298_,
    new_n18299_, new_n18301_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18311_,
    new_n18312_, new_n18313_, new_n18314_, new_n18316_, new_n18317_,
    new_n18319_, new_n18320_, new_n18321_, new_n18322_, new_n18324_,
    new_n18325_, new_n18326_, new_n18327_, new_n18328_, new_n18329_,
    new_n18330_, new_n18332_, new_n18334_, new_n18335_, new_n18336_,
    new_n18337_, new_n18338_, new_n18339_, new_n18341_, new_n18342_,
    new_n18343_, new_n18344_, new_n18346_, new_n18347_, new_n18349_,
    new_n18350_, new_n18351_, new_n18352_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18361_,
    new_n18363_, new_n18364_, new_n18365_, new_n18366_, new_n18367_,
    new_n18369_, new_n18370_, new_n18371_, new_n18372_, new_n18374_,
    new_n18375_, new_n18377_, new_n18378_, new_n18379_, new_n18380_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18389_, new_n18391_, new_n18392_, new_n18393_,
    new_n18394_, new_n18395_, new_n18397_, new_n18398_, new_n18399_,
    new_n18400_, new_n18402_, new_n18403_, new_n18405_, new_n18406_,
    new_n18407_, new_n18408_, new_n18410_, new_n18411_, new_n18412_,
    new_n18413_, new_n18414_, new_n18415_, new_n18417_, new_n18419_,
    new_n18420_, new_n18421_, new_n18422_, new_n18423_, new_n18425_,
    new_n18426_, new_n18427_, new_n18428_, new_n18430_, new_n18431_,
    new_n18433_, new_n18434_, new_n18435_, new_n18436_, new_n18438_,
    new_n18439_, new_n18440_, new_n18441_, new_n18442_, new_n18443_,
    new_n18445_, new_n18447_, new_n18448_, new_n18449_, new_n18450_,
    new_n18451_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18458_, new_n18459_, new_n18461_, new_n18462_, new_n18463_,
    new_n18464_, new_n18466_, new_n18467_, new_n18468_, new_n18469_,
    new_n18470_, new_n18471_, new_n18473_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18481_, new_n18482_,
    new_n18483_, new_n18484_, new_n18486_, new_n18487_, new_n18489_,
    new_n18490_, new_n18491_, new_n18492_, new_n18494_, new_n18495_,
    new_n18496_, new_n18497_, new_n18498_, new_n18499_, new_n18501_,
    new_n18503_, new_n18504_, new_n18505_, new_n18506_, new_n18507_,
    new_n18509_, new_n18510_, new_n18511_, new_n18512_, new_n18514_,
    new_n18515_, new_n18517_, new_n18518_, new_n18519_, new_n18520_,
    new_n18522_, new_n18523_, new_n18524_, new_n18525_, new_n18526_,
    new_n18527_, new_n18529_, new_n18531_, new_n18532_, new_n18533_,
    new_n18534_, new_n18535_, new_n18537_, new_n18538_, new_n18539_,
    new_n18540_, new_n18542_, new_n18543_, new_n18545_, new_n18546_,
    new_n18547_, new_n18548_, new_n18550_, new_n18551_, new_n18552_,
    new_n18553_, new_n18554_, new_n18555_, new_n18557_, new_n18559_,
    new_n18560_, new_n18561_, new_n18562_, new_n18563_, new_n18565_,
    new_n18566_, new_n18567_, new_n18568_, new_n18570_, new_n18571_,
    new_n18573_, new_n18574_, new_n18575_, new_n18576_, new_n18578_,
    new_n18579_, new_n18580_, new_n18581_, new_n18582_, new_n18583_,
    new_n18585_, new_n18587_, new_n18588_, new_n18589_, new_n18590_,
    new_n18591_, new_n18593_, new_n18594_, new_n18595_, new_n18596_,
    new_n18598_, new_n18599_, new_n18601_, new_n18602_, new_n18603_,
    new_n18604_, new_n18606_, new_n18607_, new_n18608_, new_n18609_,
    new_n18610_, new_n18611_, new_n18613_, new_n18615_, new_n18616_,
    new_n18617_, new_n18618_, new_n18619_, new_n18621_, new_n18622_,
    new_n18623_, new_n18624_, new_n18626_, new_n18627_, new_n18629_,
    new_n18630_, new_n18631_, new_n18632_, new_n18634_, new_n18635_,
    new_n18636_, new_n18637_, new_n18638_, new_n18639_, new_n18641_,
    new_n18643_, new_n18644_, new_n18645_, new_n18646_, new_n18647_,
    new_n18649_, new_n18650_, new_n18651_, new_n18652_, new_n18654_,
    new_n18655_, new_n18657_, new_n18658_, new_n18659_, new_n18660_,
    new_n18662_, new_n18663_, new_n18664_, new_n18665_, new_n18666_,
    new_n18667_, new_n18669_, new_n18671_, new_n18672_, new_n18673_,
    new_n18674_, new_n18675_, new_n18677_, new_n18678_, new_n18679_,
    new_n18680_, new_n18682_, new_n18683_, new_n18685_, new_n18686_,
    new_n18687_, new_n18688_, new_n18690_, new_n18691_, new_n18692_,
    new_n18693_, new_n18694_, new_n18695_, new_n18697_, new_n18699_,
    new_n18700_, new_n18701_, new_n18702_, new_n18703_, new_n18705_,
    new_n18706_, new_n18707_, new_n18708_, new_n18710_, new_n18711_,
    new_n18713_, new_n18714_, new_n18715_, new_n18716_, new_n18718_,
    new_n18719_, new_n18720_, new_n18721_, new_n18722_, new_n18723_,
    new_n18725_, new_n18727_, new_n18728_, new_n18729_, new_n18730_,
    new_n18731_, new_n18733_, new_n18734_, new_n18735_, new_n18736_,
    new_n18738_, new_n18739_, new_n18741_, new_n18742_, new_n18743_,
    new_n18744_, new_n18746_, new_n18747_, new_n18748_, new_n18749_,
    new_n18750_, new_n18751_, new_n18753_, new_n18755_, new_n18756_,
    new_n18757_, new_n18758_, new_n18759_, new_n18761_, new_n18762_,
    new_n18763_, new_n18764_, new_n18766_, new_n18767_, new_n18769_,
    new_n18770_, new_n18771_, new_n18772_, new_n18774_, new_n18775_,
    new_n18776_, new_n18777_, new_n18778_, new_n18779_, new_n18781_,
    new_n18783_, new_n18784_, new_n18785_, new_n18786_, new_n18787_,
    new_n18789_, new_n18790_, new_n18791_, new_n18792_, new_n18794_,
    new_n18795_, new_n18797_, new_n18798_, new_n18799_, new_n18800_,
    new_n18802_, new_n18803_, new_n18804_, new_n18805_, new_n18806_,
    new_n18807_, new_n18809_, new_n18811_, new_n18812_, new_n18813_,
    new_n18814_, new_n18815_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18822_, new_n18823_, new_n18825_, new_n18826_,
    new_n18828_, new_n18829_, new_n18831_, new_n18832_, new_n18834_,
    new_n18835_, new_n18837_, new_n18838_, new_n18840_, new_n18841_,
    new_n18843_, new_n18844_, new_n18846_, new_n18847_, new_n18849_,
    new_n18850_, new_n18852_, new_n18853_, new_n18855_, new_n18856_,
    new_n18858_, new_n18859_, new_n18860_, new_n18861_, new_n18862_,
    new_n18864_, new_n18865_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18873_, new_n18874_, new_n18876_,
    new_n18877_, new_n18878_, new_n18879_, new_n18880_, new_n18882_,
    new_n18883_, new_n18885_, new_n18886_, new_n18887_, new_n18888_,
    new_n18889_, new_n18891_, new_n18892_, new_n18894_, new_n18895_,
    new_n18896_, new_n18897_, new_n18898_, new_n18900_, new_n18901_,
    new_n18903_, new_n18904_, new_n18905_, new_n18906_, new_n18907_,
    new_n18909_, new_n18910_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18918_, new_n18919_, new_n18921_,
    new_n18922_, new_n18923_, new_n18924_, new_n18925_, new_n18927_,
    new_n18928_, new_n18930_, new_n18931_, new_n18932_, new_n18933_,
    new_n18934_, new_n18936_, new_n18937_, new_n18939_, new_n18940_,
    new_n18941_, new_n18942_, new_n18943_, new_n18945_, new_n18946_,
    new_n18948_, new_n18949_, new_n18950_, new_n18951_, new_n18952_,
    new_n18954_, new_n18955_, new_n18957_, new_n18958_, new_n18959_,
    new_n18960_, new_n18961_, new_n18963_, new_n18964_, new_n18966_,
    new_n18967_, new_n18968_, new_n18969_, new_n18970_, new_n18972_,
    new_n18973_, new_n18975_, new_n18976_, new_n18977_, new_n18978_,
    new_n18979_, new_n18981_, new_n18982_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18990_, new_n18991_,
    new_n18993_, new_n18994_, new_n18995_, new_n18996_, new_n18997_,
    new_n18999_, new_n19000_, new_n19002_, new_n19003_, new_n19004_,
    new_n19005_, new_n19006_, new_n19008_, new_n19009_, new_n19011_,
    new_n19012_, new_n19013_, new_n19014_, new_n19015_, new_n19017_,
    new_n19018_, new_n19020_, new_n19021_, new_n19022_, new_n19023_,
    new_n19024_, new_n19026_, new_n19027_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19035_, new_n19036_,
    new_n19038_, new_n19039_, new_n19040_, new_n19041_, new_n19042_,
    new_n19044_, new_n19045_, new_n19047_, new_n19048_, new_n19049_,
    new_n19050_, new_n19051_, new_n19053_, new_n19054_, new_n19056_,
    new_n19057_, new_n19058_, new_n19059_, new_n19060_, new_n19062_,
    new_n19063_, new_n19065_, new_n19066_, new_n19067_, new_n19068_,
    new_n19069_, new_n19071_, new_n19072_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19080_, new_n19081_,
    new_n19083_, new_n19084_, new_n19085_, new_n19086_, new_n19087_,
    new_n19089_, new_n19090_, new_n19092_, new_n19093_, new_n19094_,
    new_n19095_, new_n19096_, new_n19098_, new_n19099_, new_n19101_,
    new_n19102_, new_n19103_, new_n19104_, new_n19105_, new_n19107_,
    new_n19108_, new_n19110_, new_n19111_, new_n19112_, new_n19113_,
    new_n19114_, new_n19116_, new_n19117_, new_n19119_, new_n19120_,
    new_n19121_, new_n19122_, new_n19123_, new_n19125_, new_n19126_,
    new_n19128_, new_n19129_, new_n19130_, new_n19131_, new_n19132_,
    new_n19134_, new_n19135_, new_n19137_, new_n19138_, new_n19139_,
    new_n19140_, new_n19141_, new_n19143_, new_n19144_, new_n19146_,
    new_n19148_, new_n19149_, new_n19151_, new_n19152_, new_n19153_,
    new_n19154_, new_n19156_, new_n19157_, new_n19158_, new_n19159_,
    new_n19160_, new_n19162_, new_n19163_, new_n19166_, new_n19167_,
    new_n19168_, new_n19169_, new_n19170_, new_n19171_, new_n19172_,
    new_n19173_, new_n19174_, new_n19175_, new_n19176_, new_n19177_,
    new_n19178_, new_n19180_, new_n19181_, new_n19183_, new_n19184_,
    new_n19186_, new_n19187_, new_n19189_, new_n19190_, new_n19191_,
    new_n19193_, new_n19194_, new_n19195_, new_n19196_, new_n19197_,
    new_n19198_, new_n19199_, new_n19200_, new_n19201_, new_n19202_,
    new_n19203_, new_n19205_, new_n19206_, new_n19208_, new_n19209_,
    new_n19210_, new_n19212_, new_n19213_, new_n19214_, new_n19216_,
    new_n19217_, new_n19218_, new_n19220_, new_n19221_, new_n19222_,
    new_n19224_, new_n19225_, new_n19226_, new_n19228_, new_n19229_,
    new_n19230_, new_n19231_, new_n19232_, new_n19234_, new_n19235_,
    new_n19236_, new_n19238_, new_n19240_, new_n19241_, new_n19242_,
    new_n19243_, new_n19244_, new_n19246_, new_n19247_, new_n19248_,
    new_n19250_, new_n19251_, new_n19252_, new_n19253_, new_n19254_,
    new_n19255_, new_n19256_, new_n19257_, new_n19258_, new_n19259_,
    new_n19260_, new_n19261_, new_n19262_, new_n19263_, new_n19264_,
    new_n19265_, new_n19266_, new_n19267_, new_n19268_, new_n19269_,
    new_n19270_, new_n19271_, new_n19272_, new_n19273_, new_n19274_,
    new_n19275_, new_n19276_, new_n19277_, new_n19278_, new_n19279_,
    new_n19280_, new_n19281_, new_n19282_, new_n19283_, new_n19284_,
    new_n19285_, new_n19286_, new_n19287_, new_n19288_, new_n19289_,
    new_n19290_, new_n19291_, new_n19292_, new_n19293_, new_n19294_,
    new_n19295_, new_n19296_, new_n19297_, new_n19298_, new_n19299_,
    new_n19300_, new_n19301_, new_n19302_, new_n19303_, new_n19304_,
    new_n19305_, new_n19306_, new_n19307_, new_n19308_, new_n19309_,
    new_n19310_, new_n19311_, new_n19312_, new_n19313_, new_n19314_,
    new_n19315_, new_n19316_, new_n19317_, new_n19318_, new_n19319_,
    new_n19320_, new_n19321_, new_n19322_, new_n19323_, new_n19324_,
    new_n19325_, new_n19326_, new_n19327_, new_n19328_, new_n19329_,
    new_n19330_, new_n19331_, new_n19332_, new_n19333_, new_n19334_,
    new_n19335_, new_n19336_, new_n19337_, new_n19338_, new_n19339_,
    new_n19340_, new_n19341_, new_n19342_, new_n19343_, new_n19344_,
    new_n19345_, new_n19346_, new_n19347_, new_n19348_, new_n19349_,
    new_n19350_, new_n19351_, new_n19352_, new_n19353_, new_n19354_,
    new_n19355_, new_n19356_, new_n19357_, new_n19358_, new_n19359_,
    new_n19360_, new_n19361_, new_n19362_, new_n19363_, new_n19364_,
    new_n19365_, new_n19366_, new_n19367_, new_n19368_, new_n19369_,
    new_n19370_, new_n19371_, new_n19372_, new_n19373_, new_n19374_,
    new_n19375_, new_n19376_, new_n19377_, new_n19378_, new_n19379_,
    new_n19380_, new_n19381_, new_n19382_, new_n19383_, new_n19384_,
    new_n19385_, new_n19386_, new_n19387_, new_n19388_, new_n19389_,
    new_n19390_, new_n19391_, new_n19392_, new_n19393_, new_n19394_,
    new_n19395_, new_n19396_, new_n19397_, new_n19398_, new_n19399_,
    new_n19400_, new_n19401_, new_n19402_, new_n19403_, new_n19404_,
    new_n19405_, new_n19406_, new_n19407_, new_n19408_, new_n19409_,
    new_n19410_, new_n19411_, new_n19412_, new_n19413_, new_n19414_,
    new_n19415_, new_n19416_, new_n19417_, new_n19418_, new_n19419_,
    new_n19420_, new_n19421_, new_n19422_, new_n19423_, new_n19424_,
    new_n19425_, new_n19426_, new_n19427_, new_n19428_, new_n19429_,
    new_n19430_, new_n19431_, new_n19432_, new_n19433_, new_n19434_,
    new_n19435_, new_n19436_, new_n19437_, new_n19438_, new_n19439_,
    new_n19440_, new_n19441_, new_n19442_, new_n19443_, new_n19444_,
    new_n19445_, new_n19446_, new_n19447_, new_n19448_, new_n19449_,
    new_n19450_, new_n19451_, new_n19452_, new_n19453_, new_n19454_,
    new_n19455_, new_n19456_, new_n19457_, new_n19458_, new_n19459_,
    new_n19460_, new_n19461_, new_n19462_, new_n19463_, new_n19464_,
    new_n19465_, new_n19466_, new_n19467_, new_n19468_, new_n19469_,
    new_n19470_, new_n19471_, new_n19472_, new_n19473_, new_n19474_,
    new_n19475_, new_n19476_, new_n19477_, new_n19478_, new_n19479_,
    new_n19480_, new_n19481_, new_n19482_, new_n19483_, new_n19484_,
    new_n19485_, new_n19486_, new_n19487_, new_n19488_, new_n19489_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19514_,
    new_n19515_, new_n19516_, new_n19517_, new_n19518_, new_n19519_,
    new_n19520_, new_n19521_, new_n19522_, new_n19523_, new_n19524_,
    new_n19525_, new_n19526_, new_n19527_, new_n19528_, new_n19529_,
    new_n19530_, new_n19531_, new_n19532_, new_n19533_, new_n19534_,
    new_n19535_, new_n19536_, new_n19537_, new_n19538_, new_n19539_,
    new_n19540_, new_n19541_, new_n19542_, new_n19543_, new_n19544_,
    new_n19545_, new_n19546_, new_n19547_, new_n19548_, new_n19549_,
    new_n19550_, new_n19551_, new_n19552_, new_n19553_, new_n19554_,
    new_n19555_, new_n19556_, new_n19557_, new_n19558_, new_n19559_,
    new_n19560_, new_n19561_, new_n19562_, new_n19563_, new_n19564_,
    new_n19565_, new_n19566_, new_n19567_, new_n19568_, new_n19569_,
    new_n19570_, new_n19571_, new_n19572_, new_n19573_, new_n19574_,
    new_n19575_, new_n19576_, new_n19577_, new_n19578_, new_n19579_,
    new_n19580_, new_n19581_, new_n19582_, new_n19583_, new_n19584_,
    new_n19585_, new_n19586_, new_n19587_, new_n19588_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19735_,
    new_n19736_, new_n19737_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19804_, new_n19805_, new_n19806_,
    new_n19807_, new_n19808_, new_n19809_, new_n19810_, new_n19811_,
    new_n19812_, new_n19813_, new_n19814_, new_n19815_, new_n19816_,
    new_n19817_, new_n19818_, new_n19819_, new_n19820_, new_n19821_,
    new_n19822_, new_n19823_, new_n19824_, new_n19825_, new_n19826_,
    new_n19827_, new_n19828_, new_n19829_, new_n19830_, new_n19831_,
    new_n19832_, new_n19833_, new_n19834_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19840_, new_n19841_,
    new_n19843_, new_n19844_, new_n19845_, new_n19846_, new_n19847_,
    new_n19848_, new_n19849_, new_n19850_, new_n19851_, new_n19852_,
    new_n19853_, new_n19854_, new_n19855_, new_n19856_, new_n19857_,
    new_n19858_, new_n19859_, new_n19860_, new_n19861_, new_n19862_,
    new_n19863_, new_n19864_, new_n19865_, new_n19866_, new_n19867_,
    new_n19868_, new_n19869_, new_n19870_, new_n19871_, new_n19872_,
    new_n19873_, new_n19874_, new_n19875_, new_n19876_, new_n19877_,
    new_n19878_, new_n19879_, new_n19880_, new_n19881_, new_n19882_,
    new_n19883_, new_n19884_, new_n19885_, new_n19886_, new_n19887_,
    new_n19888_, new_n19889_, new_n19890_, new_n19891_, new_n19892_,
    new_n19893_, new_n19894_, new_n19895_, new_n19896_, new_n19897_,
    new_n19898_, new_n19899_, new_n19900_, new_n19901_, new_n19902_,
    new_n19903_, new_n19904_, new_n19905_, new_n19906_, new_n19907_,
    new_n19908_, new_n19909_, new_n19910_, new_n19911_, new_n19912_,
    new_n19913_, new_n19914_, new_n19915_, new_n19916_, new_n19917_,
    new_n19918_, new_n19919_, new_n19920_, new_n19921_, new_n19922_,
    new_n19923_, new_n19924_, new_n19925_, new_n19926_, new_n19927_,
    new_n19928_, new_n19929_, new_n19930_, new_n19931_, new_n19932_,
    new_n19933_, new_n19934_, new_n19935_, new_n19936_, new_n19937_,
    new_n19938_, new_n19939_, new_n19940_, new_n19941_, new_n19942_,
    new_n19943_, new_n19944_, new_n19945_, new_n19946_, new_n19947_,
    new_n19948_, new_n19950_, new_n19951_, new_n19952_, new_n19953_,
    new_n19954_, new_n19955_, new_n19956_, new_n19957_, new_n19958_,
    new_n19959_, new_n19960_, new_n19961_, new_n19962_, new_n19963_,
    new_n19964_, new_n19965_, new_n19966_, new_n19967_, new_n19968_,
    new_n19969_, new_n19970_, new_n19971_, new_n19972_, new_n19973_,
    new_n19974_, new_n19975_, new_n19976_, new_n19977_, new_n19978_,
    new_n19979_, new_n19980_, new_n19981_, new_n19982_, new_n19983_,
    new_n19984_, new_n19985_, new_n19986_, new_n19987_, new_n19988_,
    new_n19989_, new_n19990_, new_n19991_, new_n19992_, new_n19993_,
    new_n19994_, new_n19995_, new_n19996_, new_n19997_, new_n19998_,
    new_n19999_, new_n20000_, new_n20001_, new_n20002_, new_n20003_,
    new_n20004_, new_n20005_, new_n20006_, new_n20007_, new_n20008_,
    new_n20009_, new_n20010_, new_n20011_, new_n20012_, new_n20013_,
    new_n20014_, new_n20015_, new_n20016_, new_n20017_, new_n20018_,
    new_n20019_, new_n20020_, new_n20021_, new_n20022_, new_n20023_,
    new_n20024_, new_n20025_, new_n20026_, new_n20027_, new_n20028_,
    new_n20030_, new_n20031_, new_n20032_, new_n20033_, new_n20034_,
    new_n20035_, new_n20036_, new_n20037_, new_n20038_, new_n20039_,
    new_n20040_, new_n20041_, new_n20042_, new_n20043_, new_n20044_,
    new_n20045_, new_n20046_, new_n20047_, new_n20048_, new_n20049_,
    new_n20050_, new_n20051_, new_n20052_, new_n20053_, new_n20054_,
    new_n20055_, new_n20056_, new_n20057_, new_n20058_, new_n20059_,
    new_n20060_, new_n20061_, new_n20062_, new_n20063_, new_n20064_,
    new_n20065_, new_n20066_, new_n20067_, new_n20068_, new_n20069_,
    new_n20070_, new_n20071_, new_n20072_, new_n20073_, new_n20074_,
    new_n20075_, new_n20076_, new_n20077_, new_n20078_, new_n20079_,
    new_n20080_, new_n20081_, new_n20082_, new_n20083_, new_n20084_,
    new_n20085_, new_n20086_, new_n20087_, new_n20088_, new_n20089_,
    new_n20090_, new_n20091_, new_n20092_, new_n20093_, new_n20094_,
    new_n20095_, new_n20096_, new_n20097_, new_n20098_, new_n20099_,
    new_n20100_, new_n20101_, new_n20102_, new_n20103_, new_n20104_,
    new_n20105_, new_n20106_, new_n20107_, new_n20108_, new_n20109_,
    new_n20110_, new_n20111_, new_n20112_, new_n20113_, new_n20115_,
    new_n20116_, new_n20117_, new_n20118_, new_n20119_, new_n20120_,
    new_n20121_, new_n20122_, new_n20123_, new_n20124_, new_n20125_,
    new_n20126_, new_n20127_, new_n20128_, new_n20129_, new_n20130_,
    new_n20131_, new_n20132_, new_n20133_, new_n20134_, new_n20135_,
    new_n20136_, new_n20137_, new_n20138_, new_n20139_, new_n20140_,
    new_n20141_, new_n20142_, new_n20143_, new_n20144_, new_n20145_,
    new_n20146_, new_n20147_, new_n20148_, new_n20149_, new_n20150_,
    new_n20151_, new_n20152_, new_n20153_, new_n20154_, new_n20155_,
    new_n20156_, new_n20157_, new_n20158_, new_n20159_, new_n20160_,
    new_n20161_, new_n20162_, new_n20163_, new_n20164_, new_n20165_,
    new_n20166_, new_n20167_, new_n20168_, new_n20169_, new_n20170_,
    new_n20171_, new_n20172_, new_n20173_, new_n20174_, new_n20175_,
    new_n20176_, new_n20177_, new_n20178_, new_n20179_, new_n20180_,
    new_n20181_, new_n20182_, new_n20183_, new_n20184_, new_n20185_,
    new_n20186_, new_n20187_, new_n20188_, new_n20189_, new_n20190_,
    new_n20191_, new_n20192_, new_n20193_, new_n20194_, new_n20195_,
    new_n20196_, new_n20197_, new_n20198_, new_n20200_, new_n20201_,
    new_n20202_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20210_, new_n20211_,
    new_n20212_, new_n20213_, new_n20214_, new_n20215_, new_n20216_,
    new_n20217_, new_n20218_, new_n20219_, new_n20220_, new_n20221_,
    new_n20222_, new_n20223_, new_n20224_, new_n20225_, new_n20226_,
    new_n20227_, new_n20228_, new_n20229_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20283_, new_n20284_, new_n20285_, new_n20286_, new_n20287_,
    new_n20288_, new_n20289_, new_n20290_, new_n20291_, new_n20292_,
    new_n20293_, new_n20294_, new_n20295_, new_n20296_, new_n20297_,
    new_n20298_, new_n20299_, new_n20300_, new_n20301_, new_n20302_,
    new_n20303_, new_n20304_, new_n20305_, new_n20306_, new_n20307_,
    new_n20308_, new_n20309_, new_n20310_, new_n20311_, new_n20312_,
    new_n20313_, new_n20314_, new_n20315_, new_n20316_, new_n20317_,
    new_n20318_, new_n20319_, new_n20320_, new_n20321_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20351_, new_n20352_, new_n20353_,
    new_n20354_, new_n20355_, new_n20356_, new_n20357_, new_n20358_,
    new_n20359_, new_n20360_, new_n20361_, new_n20362_, new_n20363_,
    new_n20364_, new_n20365_, new_n20366_, new_n20367_, new_n20368_,
    new_n20369_, new_n20370_, new_n20371_, new_n20372_, new_n20373_,
    new_n20374_, new_n20375_, new_n20376_, new_n20377_, new_n20378_,
    new_n20379_, new_n20380_, new_n20381_, new_n20382_, new_n20383_,
    new_n20384_, new_n20385_, new_n20386_, new_n20387_, new_n20388_,
    new_n20389_, new_n20390_, new_n20391_, new_n20392_, new_n20393_,
    new_n20394_, new_n20395_, new_n20396_, new_n20397_, new_n20398_,
    new_n20399_, new_n20400_, new_n20401_, new_n20402_, new_n20403_,
    new_n20404_, new_n20405_, new_n20406_, new_n20407_, new_n20408_,
    new_n20409_, new_n20410_, new_n20411_, new_n20412_, new_n20413_,
    new_n20414_, new_n20415_, new_n20416_, new_n20417_, new_n20418_,
    new_n20419_, new_n20420_, new_n20421_, new_n20422_, new_n20424_,
    new_n20425_, new_n20426_, new_n20427_, new_n20428_, new_n20429_,
    new_n20430_, new_n20431_, new_n20432_, new_n20433_, new_n20434_,
    new_n20435_, new_n20436_, new_n20437_, new_n20438_, new_n20439_,
    new_n20440_, new_n20441_, new_n20442_, new_n20443_, new_n20444_,
    new_n20445_, new_n20446_, new_n20447_, new_n20448_, new_n20449_,
    new_n20450_, new_n20451_, new_n20452_, new_n20453_, new_n20454_,
    new_n20455_, new_n20456_, new_n20457_, new_n20458_, new_n20459_,
    new_n20460_, new_n20461_, new_n20462_, new_n20463_, new_n20464_,
    new_n20465_, new_n20466_, new_n20467_, new_n20468_, new_n20469_,
    new_n20470_, new_n20471_, new_n20472_, new_n20473_, new_n20474_,
    new_n20475_, new_n20476_, new_n20477_, new_n20478_, new_n20479_,
    new_n20480_, new_n20481_, new_n20482_, new_n20483_, new_n20484_,
    new_n20485_, new_n20486_, new_n20487_, new_n20488_, new_n20489_,
    new_n20490_, new_n20491_, new_n20492_, new_n20493_, new_n20494_,
    new_n20495_, new_n20497_, new_n20498_, new_n20499_, new_n20500_,
    new_n20501_, new_n20502_, new_n20503_, new_n20504_, new_n20505_,
    new_n20506_, new_n20507_, new_n20508_, new_n20509_, new_n20510_,
    new_n20511_, new_n20512_, new_n20513_, new_n20514_, new_n20515_,
    new_n20516_, new_n20517_, new_n20518_, new_n20519_, new_n20520_,
    new_n20521_, new_n20522_, new_n20523_, new_n20524_, new_n20525_,
    new_n20526_, new_n20527_, new_n20528_, new_n20529_, new_n20530_,
    new_n20531_, new_n20532_, new_n20533_, new_n20534_, new_n20535_,
    new_n20536_, new_n20537_, new_n20538_, new_n20539_, new_n20540_,
    new_n20541_, new_n20542_, new_n20543_, new_n20544_, new_n20545_,
    new_n20546_, new_n20547_, new_n20548_, new_n20549_, new_n20550_,
    new_n20551_, new_n20552_, new_n20553_, new_n20554_, new_n20555_,
    new_n20556_, new_n20557_, new_n20558_, new_n20559_, new_n20560_,
    new_n20561_, new_n20562_, new_n20563_, new_n20564_, new_n20565_,
    new_n20566_, new_n20567_, new_n20568_, new_n20570_, new_n20571_,
    new_n20572_, new_n20573_, new_n20574_, new_n20575_, new_n20576_,
    new_n20577_, new_n20578_, new_n20579_, new_n20580_, new_n20581_,
    new_n20582_, new_n20583_, new_n20584_, new_n20585_, new_n20586_,
    new_n20587_, new_n20588_, new_n20589_, new_n20590_, new_n20591_,
    new_n20592_, new_n20593_, new_n20594_, new_n20595_, new_n20596_,
    new_n20597_, new_n20598_, new_n20599_, new_n20600_, new_n20601_,
    new_n20602_, new_n20603_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20643_, new_n20644_, new_n20645_, new_n20646_, new_n20647_,
    new_n20648_, new_n20649_, new_n20650_, new_n20651_, new_n20652_,
    new_n20653_, new_n20654_, new_n20655_, new_n20656_, new_n20657_,
    new_n20658_, new_n20659_, new_n20660_, new_n20661_, new_n20662_,
    new_n20663_, new_n20664_, new_n20665_, new_n20666_, new_n20667_,
    new_n20668_, new_n20669_, new_n20670_, new_n20671_, new_n20672_,
    new_n20673_, new_n20674_, new_n20675_, new_n20676_, new_n20677_,
    new_n20678_, new_n20679_, new_n20680_, new_n20681_, new_n20682_,
    new_n20683_, new_n20684_, new_n20685_, new_n20686_, new_n20687_,
    new_n20688_, new_n20689_, new_n20690_, new_n20691_, new_n20692_,
    new_n20693_, new_n20694_, new_n20695_, new_n20696_, new_n20697_,
    new_n20698_, new_n20699_, new_n20700_, new_n20701_, new_n20702_,
    new_n20703_, new_n20704_, new_n20705_, new_n20706_, new_n20707_,
    new_n20708_, new_n20709_, new_n20710_, new_n20711_, new_n20712_,
    new_n20713_, new_n20714_, new_n20716_, new_n20717_, new_n20718_,
    new_n20719_, new_n20720_, new_n20721_, new_n20722_, new_n20723_,
    new_n20724_, new_n20725_, new_n20726_, new_n20727_, new_n20728_,
    new_n20729_, new_n20730_, new_n20731_, new_n20732_, new_n20733_,
    new_n20734_, new_n20735_, new_n20736_, new_n20737_, new_n20738_,
    new_n20739_, new_n20740_, new_n20741_, new_n20742_, new_n20743_,
    new_n20744_, new_n20745_, new_n20746_, new_n20747_, new_n20748_,
    new_n20749_, new_n20750_, new_n20751_, new_n20752_, new_n20753_,
    new_n20754_, new_n20755_, new_n20756_, new_n20757_, new_n20758_,
    new_n20759_, new_n20760_, new_n20761_, new_n20762_, new_n20763_,
    new_n20764_, new_n20765_, new_n20766_, new_n20767_, new_n20768_,
    new_n20769_, new_n20770_, new_n20771_, new_n20772_, new_n20773_,
    new_n20774_, new_n20775_, new_n20776_, new_n20777_, new_n20778_,
    new_n20779_, new_n20780_, new_n20781_, new_n20782_, new_n20783_,
    new_n20784_, new_n20785_, new_n20786_, new_n20787_, new_n20789_,
    new_n20790_, new_n20791_, new_n20792_, new_n20793_, new_n20794_,
    new_n20795_, new_n20796_, new_n20797_, new_n20798_, new_n20799_,
    new_n20800_, new_n20801_, new_n20802_, new_n20803_, new_n20804_,
    new_n20805_, new_n20806_, new_n20807_, new_n20808_, new_n20809_,
    new_n20810_, new_n20811_, new_n20812_, new_n20813_, new_n20814_,
    new_n20815_, new_n20816_, new_n20817_, new_n20818_, new_n20819_,
    new_n20820_, new_n20821_, new_n20822_, new_n20823_, new_n20824_,
    new_n20825_, new_n20826_, new_n20827_, new_n20828_, new_n20829_,
    new_n20830_, new_n20831_, new_n20832_, new_n20833_, new_n20834_,
    new_n20835_, new_n20836_, new_n20837_, new_n20838_, new_n20839_,
    new_n20840_, new_n20841_, new_n20842_, new_n20843_, new_n20844_,
    new_n20845_, new_n20846_, new_n20847_, new_n20848_, new_n20849_,
    new_n20850_, new_n20851_, new_n20852_, new_n20853_, new_n20854_,
    new_n20855_, new_n20856_, new_n20857_, new_n20858_, new_n20860_,
    new_n20861_, new_n20862_, new_n20863_, new_n20864_, new_n20865_,
    new_n20866_, new_n20867_, new_n20868_, new_n20869_, new_n20870_,
    new_n20871_, new_n20872_, new_n20873_, new_n20874_, new_n20875_,
    new_n20876_, new_n20877_, new_n20878_, new_n20879_, new_n20880_,
    new_n20881_, new_n20882_, new_n20883_, new_n20884_, new_n20885_,
    new_n20886_, new_n20887_, new_n20888_, new_n20889_, new_n20890_,
    new_n20891_, new_n20892_, new_n20893_, new_n20894_, new_n20895_,
    new_n20896_, new_n20897_, new_n20898_, new_n20899_, new_n20900_,
    new_n20901_, new_n20902_, new_n20903_, new_n20904_, new_n20905_,
    new_n20906_, new_n20907_, new_n20908_, new_n20909_, new_n20910_,
    new_n20911_, new_n20912_, new_n20913_, new_n20914_, new_n20915_,
    new_n20916_, new_n20917_, new_n20918_, new_n20919_, new_n20920_,
    new_n20921_, new_n20922_, new_n20924_, new_n20925_, new_n20926_,
    new_n20927_, new_n20928_, new_n20929_, new_n20930_, new_n20931_,
    new_n20932_, new_n20933_, new_n20934_, new_n20935_, new_n20936_,
    new_n20937_, new_n20938_, new_n20939_, new_n20940_, new_n20941_,
    new_n20942_, new_n20943_, new_n20944_, new_n20945_, new_n20946_,
    new_n20947_, new_n20948_, new_n20949_, new_n20950_, new_n20951_,
    new_n20952_, new_n20953_, new_n20954_, new_n20955_, new_n20956_,
    new_n20957_, new_n20958_, new_n20959_, new_n20960_, new_n20961_,
    new_n20962_, new_n20963_, new_n20964_, new_n20965_, new_n20966_,
    new_n20967_, new_n20968_, new_n20969_, new_n20970_, new_n20971_,
    new_n20972_, new_n20973_, new_n20974_, new_n20975_, new_n20976_,
    new_n20977_, new_n20978_, new_n20979_, new_n20980_, new_n20981_,
    new_n20982_, new_n20983_, new_n20984_, new_n20985_, new_n20986_,
    new_n20987_, new_n20988_, new_n20989_, new_n20990_, new_n20991_,
    new_n20993_, new_n20994_, new_n20995_, new_n20996_, new_n20997_,
    new_n20998_, new_n20999_, new_n21000_, new_n21001_, new_n21002_,
    new_n21003_, new_n21004_, new_n21005_, new_n21006_, new_n21007_,
    new_n21008_, new_n21009_, new_n21010_, new_n21011_, new_n21012_,
    new_n21013_, new_n21014_, new_n21015_, new_n21016_, new_n21017_,
    new_n21018_, new_n21019_, new_n21020_, new_n21021_, new_n21022_,
    new_n21023_, new_n21024_, new_n21025_, new_n21026_, new_n21027_,
    new_n21028_, new_n21029_, new_n21030_, new_n21031_, new_n21032_,
    new_n21033_, new_n21034_, new_n21035_, new_n21036_, new_n21037_,
    new_n21038_, new_n21039_, new_n21040_, new_n21041_, new_n21042_,
    new_n21043_, new_n21044_, new_n21045_, new_n21046_, new_n21047_,
    new_n21048_, new_n21049_, new_n21050_, new_n21051_, new_n21052_,
    new_n21053_, new_n21054_, new_n21055_, new_n21056_, new_n21057_,
    new_n21058_, new_n21059_, new_n21061_, new_n21062_, new_n21063_,
    new_n21064_, new_n21065_, new_n21066_, new_n21067_, new_n21068_,
    new_n21069_, new_n21070_, new_n21071_, new_n21072_, new_n21073_,
    new_n21074_, new_n21075_, new_n21076_, new_n21077_, new_n21078_,
    new_n21079_, new_n21080_, new_n21081_, new_n21082_, new_n21083_,
    new_n21084_, new_n21085_, new_n21086_, new_n21087_, new_n21088_,
    new_n21089_, new_n21090_, new_n21091_, new_n21092_, new_n21093_,
    new_n21094_, new_n21095_, new_n21096_, new_n21097_, new_n21098_,
    new_n21099_, new_n21100_, new_n21101_, new_n21102_, new_n21103_,
    new_n21104_, new_n21105_, new_n21106_, new_n21107_, new_n21108_,
    new_n21109_, new_n21110_, new_n21111_, new_n21112_, new_n21113_,
    new_n21114_, new_n21115_, new_n21116_, new_n21117_, new_n21118_,
    new_n21119_, new_n21120_, new_n21121_, new_n21122_, new_n21123_,
    new_n21124_, new_n21125_, new_n21126_, new_n21127_, new_n21129_,
    new_n21130_, new_n21131_, new_n21132_, new_n21133_, new_n21134_,
    new_n21135_, new_n21136_, new_n21137_, new_n21138_, new_n21139_,
    new_n21140_, new_n21141_, new_n21142_, new_n21143_, new_n21144_,
    new_n21145_, new_n21146_, new_n21147_, new_n21148_, new_n21149_,
    new_n21150_, new_n21151_, new_n21152_, new_n21153_, new_n21154_,
    new_n21155_, new_n21156_, new_n21157_, new_n21158_, new_n21159_,
    new_n21160_, new_n21161_, new_n21162_, new_n21163_, new_n21164_,
    new_n21165_, new_n21166_, new_n21167_, new_n21168_, new_n21169_,
    new_n21170_, new_n21171_, new_n21172_, new_n21173_, new_n21174_,
    new_n21175_, new_n21176_, new_n21177_, new_n21178_, new_n21179_,
    new_n21180_, new_n21181_, new_n21182_, new_n21183_, new_n21184_,
    new_n21185_, new_n21186_, new_n21187_, new_n21188_, new_n21189_,
    new_n21190_, new_n21191_, new_n21192_, new_n21193_, new_n21194_,
    new_n21195_, new_n21197_, new_n21198_, new_n21199_, new_n21200_,
    new_n21201_, new_n21202_, new_n21203_, new_n21204_, new_n21205_,
    new_n21206_, new_n21207_, new_n21208_, new_n21209_, new_n21210_,
    new_n21211_, new_n21212_, new_n21213_, new_n21214_, new_n21215_,
    new_n21216_, new_n21217_, new_n21218_, new_n21219_, new_n21220_,
    new_n21221_, new_n21222_, new_n21223_, new_n21224_, new_n21225_,
    new_n21226_, new_n21227_, new_n21228_, new_n21229_, new_n21230_,
    new_n21231_, new_n21232_, new_n21233_, new_n21234_, new_n21235_,
    new_n21236_, new_n21237_, new_n21238_, new_n21239_, new_n21240_,
    new_n21241_, new_n21242_, new_n21243_, new_n21244_, new_n21245_,
    new_n21246_, new_n21247_, new_n21248_, new_n21249_, new_n21250_,
    new_n21251_, new_n21252_, new_n21253_, new_n21254_, new_n21255_,
    new_n21256_, new_n21257_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21265_, new_n21266_,
    new_n21267_, new_n21268_, new_n21269_, new_n21270_, new_n21271_,
    new_n21272_, new_n21273_, new_n21274_, new_n21275_, new_n21276_,
    new_n21277_, new_n21278_, new_n21279_, new_n21280_, new_n21281_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21297_, new_n21298_, new_n21299_, new_n21300_, new_n21301_,
    new_n21302_, new_n21303_, new_n21304_, new_n21305_, new_n21306_,
    new_n21307_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21333_, new_n21334_, new_n21335_, new_n21336_, new_n21337_,
    new_n21338_, new_n21339_, new_n21340_, new_n21341_, new_n21342_,
    new_n21343_, new_n21344_, new_n21345_, new_n21346_, new_n21347_,
    new_n21348_, new_n21349_, new_n21350_, new_n21351_, new_n21352_,
    new_n21353_, new_n21354_, new_n21355_, new_n21356_, new_n21357_,
    new_n21358_, new_n21359_, new_n21360_, new_n21361_, new_n21362_,
    new_n21363_, new_n21364_, new_n21365_, new_n21366_, new_n21367_,
    new_n21368_, new_n21369_, new_n21370_, new_n21371_, new_n21372_,
    new_n21373_, new_n21374_, new_n21375_, new_n21376_, new_n21377_,
    new_n21378_, new_n21379_, new_n21380_, new_n21381_, new_n21382_,
    new_n21383_, new_n21384_, new_n21385_, new_n21386_, new_n21387_,
    new_n21388_, new_n21389_, new_n21390_, new_n21391_, new_n21392_,
    new_n21393_, new_n21394_, new_n21395_, new_n21396_, new_n21397_,
    new_n21398_, new_n21399_, new_n21401_, new_n21402_, new_n21403_,
    new_n21404_, new_n21405_, new_n21406_, new_n21407_, new_n21408_,
    new_n21409_, new_n21410_, new_n21411_, new_n21412_, new_n21413_,
    new_n21414_, new_n21415_, new_n21416_, new_n21417_, new_n21418_,
    new_n21419_, new_n21420_, new_n21421_, new_n21422_, new_n21423_,
    new_n21424_, new_n21425_, new_n21426_, new_n21427_, new_n21428_,
    new_n21429_, new_n21430_, new_n21431_, new_n21432_, new_n21433_,
    new_n21434_, new_n21435_, new_n21436_, new_n21437_, new_n21438_,
    new_n21439_, new_n21440_, new_n21441_, new_n21442_, new_n21443_,
    new_n21444_, new_n21445_, new_n21446_, new_n21447_, new_n21448_,
    new_n21449_, new_n21450_, new_n21451_, new_n21452_, new_n21453_,
    new_n21454_, new_n21455_, new_n21456_, new_n21457_, new_n21458_,
    new_n21459_, new_n21460_, new_n21461_, new_n21462_, new_n21463_,
    new_n21464_, new_n21465_, new_n21467_, new_n21468_, new_n21469_,
    new_n21470_, new_n21471_, new_n21472_, new_n21473_, new_n21474_,
    new_n21475_, new_n21476_, new_n21477_, new_n21478_, new_n21479_,
    new_n21480_, new_n21481_, new_n21482_, new_n21483_, new_n21484_,
    new_n21485_, new_n21486_, new_n21487_, new_n21488_, new_n21489_,
    new_n21490_, new_n21491_, new_n21492_, new_n21493_, new_n21494_,
    new_n21495_, new_n21496_, new_n21497_, new_n21498_, new_n21499_,
    new_n21500_, new_n21501_, new_n21502_, new_n21503_, new_n21504_,
    new_n21505_, new_n21506_, new_n21507_, new_n21508_, new_n21509_,
    new_n21510_, new_n21511_, new_n21512_, new_n21513_, new_n21514_,
    new_n21515_, new_n21516_, new_n21517_, new_n21518_, new_n21519_,
    new_n21520_, new_n21521_, new_n21522_, new_n21523_, new_n21524_,
    new_n21525_, new_n21526_, new_n21527_, new_n21528_, new_n21529_,
    new_n21530_, new_n21531_, new_n21532_, new_n21533_, new_n21535_,
    new_n21536_, new_n21537_, new_n21538_, new_n21539_, new_n21540_,
    new_n21541_, new_n21542_, new_n21543_, new_n21544_, new_n21545_,
    new_n21546_, new_n21547_, new_n21548_, new_n21549_, new_n21550_,
    new_n21551_, new_n21552_, new_n21553_, new_n21554_, new_n21555_,
    new_n21556_, new_n21557_, new_n21558_, new_n21559_, new_n21560_,
    new_n21561_, new_n21562_, new_n21563_, new_n21564_, new_n21565_,
    new_n21566_, new_n21567_, new_n21568_, new_n21569_, new_n21570_,
    new_n21571_, new_n21572_, new_n21573_, new_n21574_, new_n21575_,
    new_n21576_, new_n21577_, new_n21578_, new_n21579_, new_n21580_,
    new_n21581_, new_n21582_, new_n21583_, new_n21584_, new_n21585_,
    new_n21586_, new_n21587_, new_n21588_, new_n21589_, new_n21590_,
    new_n21591_, new_n21592_, new_n21593_, new_n21594_, new_n21595_,
    new_n21596_, new_n21597_, new_n21598_, new_n21599_, new_n21600_,
    new_n21601_, new_n21603_, new_n21604_, new_n21605_, new_n21606_,
    new_n21607_, new_n21608_, new_n21609_, new_n21610_, new_n21611_,
    new_n21612_, new_n21613_, new_n21614_, new_n21615_, new_n21616_,
    new_n21617_, new_n21618_, new_n21619_, new_n21620_, new_n21621_,
    new_n21622_, new_n21623_, new_n21624_, new_n21625_, new_n21626_,
    new_n21627_, new_n21628_, new_n21629_, new_n21630_, new_n21631_,
    new_n21632_, new_n21633_, new_n21634_, new_n21635_, new_n21636_,
    new_n21637_, new_n21638_, new_n21639_, new_n21640_, new_n21641_,
    new_n21642_, new_n21643_, new_n21644_, new_n21645_, new_n21646_,
    new_n21647_, new_n21648_, new_n21649_, new_n21650_, new_n21651_,
    new_n21652_, new_n21653_, new_n21654_, new_n21655_, new_n21656_,
    new_n21657_, new_n21658_, new_n21659_, new_n21660_, new_n21661_,
    new_n21662_, new_n21663_, new_n21664_, new_n21665_, new_n21666_,
    new_n21667_, new_n21668_, new_n21669_, new_n21671_, new_n21672_,
    new_n21673_, new_n21674_, new_n21675_, new_n21676_, new_n21677_,
    new_n21678_, new_n21679_, new_n21680_, new_n21681_, new_n21682_,
    new_n21683_, new_n21684_, new_n21685_, new_n21686_, new_n21687_,
    new_n21688_, new_n21689_, new_n21690_, new_n21691_, new_n21692_,
    new_n21693_, new_n21694_, new_n21695_, new_n21696_, new_n21697_,
    new_n21698_, new_n21699_, new_n21700_, new_n21701_, new_n21702_,
    new_n21703_, new_n21704_, new_n21705_, new_n21706_, new_n21707_,
    new_n21708_, new_n21709_, new_n21710_, new_n21711_, new_n21712_,
    new_n21713_, new_n21714_, new_n21715_, new_n21716_, new_n21717_,
    new_n21718_, new_n21719_, new_n21720_, new_n21721_, new_n21722_,
    new_n21723_, new_n21724_, new_n21725_, new_n21726_, new_n21727_,
    new_n21728_, new_n21729_, new_n21730_, new_n21731_, new_n21732_,
    new_n21733_, new_n21734_, new_n21735_, new_n21737_, new_n21738_,
    new_n21739_, new_n21740_, new_n21741_, new_n21742_, new_n21743_,
    new_n21744_, new_n21745_, new_n21746_, new_n21747_, new_n21748_,
    new_n21749_, new_n21750_, new_n21751_, new_n21752_, new_n21753_,
    new_n21754_, new_n21755_, new_n21756_, new_n21757_, new_n21758_,
    new_n21759_, new_n21760_, new_n21761_, new_n21762_, new_n21763_,
    new_n21764_, new_n21765_, new_n21766_, new_n21767_, new_n21768_,
    new_n21769_, new_n21770_, new_n21771_, new_n21772_, new_n21773_,
    new_n21774_, new_n21775_, new_n21776_, new_n21777_, new_n21778_,
    new_n21779_, new_n21780_, new_n21781_, new_n21782_, new_n21783_,
    new_n21784_, new_n21785_, new_n21786_, new_n21787_, new_n21788_,
    new_n21789_, new_n21790_, new_n21791_, new_n21792_, new_n21793_,
    new_n21794_, new_n21795_, new_n21796_, new_n21797_, new_n21798_,
    new_n21800_, new_n21801_, new_n21802_, new_n21803_, new_n21804_,
    new_n21805_, new_n21806_, new_n21807_, new_n21808_, new_n21809_,
    new_n21810_, new_n21811_, new_n21812_, new_n21813_, new_n21814_,
    new_n21815_, new_n21816_, new_n21817_, new_n21818_, new_n21819_,
    new_n21820_, new_n21821_, new_n21822_, new_n21823_, new_n21824_,
    new_n21825_, new_n21826_, new_n21827_, new_n21828_, new_n21829_,
    new_n21830_, new_n21831_, new_n21832_, new_n21833_, new_n21834_,
    new_n21835_, new_n21836_, new_n21837_, new_n21838_, new_n21839_,
    new_n21840_, new_n21841_, new_n21842_, new_n21843_, new_n21844_,
    new_n21845_, new_n21846_, new_n21847_, new_n21848_, new_n21849_,
    new_n21850_, new_n21851_, new_n21852_, new_n21853_, new_n21854_,
    new_n21855_, new_n21856_, new_n21857_, new_n21858_, new_n21859_,
    new_n21860_, new_n21861_, new_n21863_, new_n21864_, new_n21865_,
    new_n21866_, new_n21867_, new_n21868_, new_n21869_, new_n21870_,
    new_n21871_, new_n21872_, new_n21873_, new_n21874_, new_n21875_,
    new_n21876_, new_n21877_, new_n21878_, new_n21879_, new_n21880_,
    new_n21881_, new_n21882_, new_n21883_, new_n21884_, new_n21885_,
    new_n21886_, new_n21887_, new_n21888_, new_n21889_, new_n21890_,
    new_n21891_, new_n21892_, new_n21893_, new_n21894_, new_n21895_,
    new_n21896_, new_n21897_, new_n21898_, new_n21899_, new_n21900_,
    new_n21901_, new_n21902_, new_n21903_, new_n21904_, new_n21905_,
    new_n21906_, new_n21907_, new_n21908_, new_n21909_, new_n21910_,
    new_n21911_, new_n21912_, new_n21913_, new_n21914_, new_n21915_,
    new_n21916_, new_n21917_, new_n21918_, new_n21919_, new_n21920_,
    new_n21921_, new_n21922_, new_n21924_, new_n21926_, new_n21928_,
    new_n21930_, new_n21932_, new_n21934_, new_n21936_, new_n21938_,
    new_n21940_, new_n21942_, new_n21944_, new_n21946_, new_n21948_,
    new_n21950_, new_n21952_, new_n21954_, new_n21956_, new_n21958_,
    new_n21960_, new_n21962_, new_n21964_, new_n21966_, new_n21968_,
    new_n21970_, new_n21972_, new_n21974_, new_n21976_, new_n21978_,
    new_n21980_, new_n21982_, new_n21983_, new_n21985_, new_n21986_,
    new_n21988_, new_n21989_, new_n21990_, new_n21991_, new_n21992_,
    new_n21993_, new_n21994_, new_n21995_, new_n21996_, new_n21997_,
    new_n21999_, new_n22000_, new_n22001_, new_n22002_, new_n22003_,
    new_n22004_, new_n22005_, new_n22006_, new_n22007_, new_n22009_,
    new_n22010_, new_n22011_, new_n22012_, new_n22013_, new_n22014_,
    new_n22015_, new_n22016_, new_n22018_, new_n22019_, new_n22020_,
    new_n22021_, new_n22022_, new_n22023_, new_n22024_, new_n22025_,
    new_n22027_, new_n22028_, new_n22029_, new_n22030_, new_n22031_,
    new_n22032_, new_n22033_, new_n22034_, new_n22036_, new_n22037_,
    new_n22038_, new_n22039_, new_n22040_, new_n22041_, new_n22042_,
    new_n22043_, new_n22045_, new_n22046_, new_n22047_, new_n22048_,
    new_n22049_, new_n22050_, new_n22051_, new_n22052_, new_n22054_,
    new_n22055_, new_n22056_, new_n22057_, new_n22058_, new_n22059_,
    new_n22060_, new_n22061_, new_n22063_, new_n22064_, new_n22065_,
    new_n22066_, new_n22067_, new_n22068_, new_n22069_, new_n22070_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22080_, new_n22081_, new_n22082_,
    new_n22083_, new_n22084_, new_n22085_, new_n22086_, new_n22088_,
    new_n22089_, new_n22090_, new_n22091_, new_n22092_, new_n22093_,
    new_n22094_, new_n22096_, new_n22097_, new_n22098_, new_n22099_,
    new_n22100_, new_n22101_, new_n22102_, new_n22104_, new_n22105_,
    new_n22106_, new_n22107_, new_n22108_, new_n22109_, new_n22110_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22120_, new_n22121_, new_n22122_,
    new_n22123_, new_n22124_, new_n22125_, new_n22126_, new_n22128_,
    new_n22129_, new_n22130_, new_n22131_, new_n22132_, new_n22133_,
    new_n22134_, new_n22136_, new_n22137_, new_n22138_, new_n22139_,
    new_n22140_, new_n22141_, new_n22143_, new_n22144_, new_n22145_,
    new_n22146_, new_n22147_, new_n22148_, new_n22150_, new_n22151_,
    new_n22152_, new_n22153_, new_n22154_, new_n22155_, new_n22157_,
    new_n22158_, new_n22159_, new_n22160_, new_n22161_, new_n22162_,
    new_n22164_, new_n22165_, new_n22166_, new_n22167_, new_n22168_,
    new_n22169_, new_n22171_, new_n22172_, new_n22173_, new_n22174_,
    new_n22175_, new_n22176_, new_n22178_, new_n22179_, new_n22180_,
    new_n22181_, new_n22182_, new_n22183_, new_n22185_, new_n22186_,
    new_n22187_, new_n22188_, new_n22189_, new_n22190_, new_n22192_,
    new_n22193_, new_n22194_, new_n22195_, new_n22196_, new_n22197_,
    new_n22199_, new_n22200_, new_n22201_, new_n22202_, new_n22203_,
    new_n22204_, new_n22206_, new_n22207_, new_n22208_, new_n22209_,
    new_n22210_, new_n22211_, new_n22213_, new_n22214_, new_n22215_,
    new_n22216_, new_n22217_, new_n22218_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22227_,
    new_n22228_, new_n22229_, new_n22230_, new_n22231_, new_n22232_,
    new_n22234_, new_n22235_, new_n22236_, new_n22237_, new_n22238_,
    new_n22239_, new_n22241_, new_n22242_, new_n22243_, new_n22244_,
    new_n22245_, new_n22246_, new_n22248_, new_n22249_, new_n22250_,
    new_n22251_, new_n22252_, new_n22253_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22262_,
    new_n22263_, new_n22264_, new_n22265_, new_n22266_, new_n22267_,
    new_n22269_, new_n22270_, new_n22271_, new_n22272_, new_n22273_,
    new_n22274_, new_n22276_, new_n22277_, new_n22278_, new_n22279_,
    new_n22280_, new_n22281_, new_n22283_, new_n22284_, new_n22285_,
    new_n22286_, new_n22287_, new_n22288_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22297_,
    new_n22298_, new_n22299_, new_n22300_, new_n22301_, new_n22302_,
    new_n22304_, new_n22305_, new_n22306_, new_n22307_, new_n22308_,
    new_n22309_, new_n22311_, new_n22312_, new_n22313_, new_n22314_,
    new_n22315_, new_n22316_, new_n22318_, new_n22319_, new_n22320_,
    new_n22321_, new_n22322_, new_n22323_, new_n22325_, new_n22326_,
    new_n22327_, new_n22328_, new_n22329_, new_n22330_, new_n22332_,
    new_n22333_, new_n22334_, new_n22335_, new_n22336_, new_n22337_,
    new_n22339_, new_n22340_, new_n22341_, new_n22342_, new_n22343_,
    new_n22344_, new_n22346_, new_n22347_, new_n22348_, new_n22349_,
    new_n22350_, new_n22351_, new_n22353_, new_n22354_, new_n22355_,
    new_n22356_, new_n22357_, new_n22358_, new_n22360_, new_n22361_,
    new_n22362_, new_n22363_, new_n22364_, new_n22365_, new_n22367_,
    new_n22368_, new_n22369_, new_n22370_, new_n22371_, new_n22372_,
    new_n22374_, new_n22375_, new_n22376_, new_n22377_, new_n22378_,
    new_n22379_, new_n22381_, new_n22382_, new_n22383_, new_n22384_,
    new_n22385_, new_n22386_, new_n22388_, new_n22389_, new_n22390_,
    new_n22391_, new_n22392_, new_n22393_, new_n22395_, new_n22396_,
    new_n22397_, new_n22398_, new_n22399_, new_n22400_, new_n22402_,
    new_n22403_, new_n22404_, new_n22405_, new_n22406_, new_n22407_,
    new_n22409_, new_n22410_, new_n22411_, new_n22412_, new_n22413_,
    new_n22414_, new_n22416_, new_n22417_, new_n22418_, new_n22419_,
    new_n22420_, new_n22421_, new_n22423_, new_n22424_, new_n22425_,
    new_n22426_, new_n22427_, new_n22428_, new_n22430_, new_n22431_,
    new_n22432_, new_n22433_, new_n22434_, new_n22435_, new_n22437_,
    new_n22438_, new_n22439_, new_n22440_, new_n22441_, new_n22442_,
    new_n22444_, new_n22445_, new_n22446_, new_n22447_, new_n22448_,
    new_n22449_, new_n22451_, new_n22452_, new_n22453_, new_n22454_,
    new_n22455_, new_n22456_, new_n22458_, new_n22459_, new_n22460_,
    new_n22461_, new_n22462_, new_n22463_, new_n22465_, new_n22466_,
    new_n22467_, new_n22468_, new_n22469_, new_n22470_, new_n22472_,
    new_n22473_, new_n22474_, new_n22475_, new_n22476_, new_n22477_,
    new_n22478_, new_n22479_, new_n22480_, new_n22481_, new_n22482_,
    new_n22484_, new_n22485_, new_n22487_, new_n22488_, new_n22490_,
    new_n22491_, new_n22493_, new_n22494_, new_n22495_, new_n22496_,
    new_n22498_, new_n22499_, new_n22501_, new_n22502_, new_n22503_,
    new_n22505_, new_n22506_, new_n22507_, new_n22509_, new_n22510_,
    new_n22511_, new_n22513_, new_n22514_, new_n22516_, new_n22517_,
    new_n22518_, new_n22520_, new_n22521_, new_n22522_, new_n22524_,
    new_n22525_, new_n22526_, new_n22528_, new_n22529_, new_n22530_,
    new_n22532_, new_n22533_, new_n22534_, new_n22536_, new_n22537_,
    new_n22538_, new_n22540_, new_n22541_, new_n22542_, new_n22544_,
    new_n22545_, new_n22547_, new_n22548_, new_n22549_, new_n22550_,
    new_n22551_, new_n22553_, new_n22554_, new_n22555_, new_n22556_,
    new_n22557_, new_n22559_, new_n22560_, new_n22561_, new_n22562_,
    new_n22563_, new_n22564_, new_n22566_, new_n22567_, new_n22568_,
    new_n22569_, new_n22570_, new_n22572_, new_n22573_, new_n22574_,
    new_n22575_, new_n22576_, new_n22577_, new_n22579_, new_n22580_,
    new_n22581_, new_n22582_, new_n22583_, new_n22584_, new_n22586_,
    new_n22587_, new_n22588_, new_n22589_, new_n22590_, new_n22591_,
    new_n22593_, new_n22594_, new_n22595_, new_n22596_, new_n22597_,
    new_n22599_, new_n22600_, new_n22601_, new_n22602_, new_n22603_,
    new_n22604_, new_n22606_, new_n22607_, new_n22608_, new_n22609_,
    new_n22610_, new_n22611_, new_n22613_, new_n22614_, new_n22615_,
    new_n22616_, new_n22617_, new_n22618_, new_n22620_, new_n22621_,
    new_n22622_, new_n22623_, new_n22624_, new_n22626_, new_n22627_,
    new_n22628_, new_n22629_, new_n22630_, new_n22631_, new_n22632_,
    new_n22633_, new_n22634_, new_n22635_, new_n22636_, new_n22637_,
    new_n22638_, new_n22639_, new_n22640_, new_n22641_, new_n22643_,
    new_n22644_, new_n22645_, new_n22646_, new_n22647_, new_n22649_,
    new_n22650_, new_n22651_, new_n22652_, new_n22653_, new_n22654_,
    new_n22655_, new_n22656_, new_n22657_, new_n22658_, new_n22659_,
    new_n22660_, new_n22661_, new_n22662_, new_n22663_, new_n22664_,
    new_n22665_, new_n22666_, new_n22667_, new_n22668_, new_n22669_,
    new_n22670_, new_n22671_, new_n22672_, new_n22673_, new_n22674_,
    new_n22675_, new_n22676_, new_n22677_, new_n22678_, new_n22679_,
    new_n22680_, new_n22681_, new_n22682_, new_n22683_, new_n22684_,
    new_n22685_, new_n22686_, new_n22687_, new_n22688_, new_n22689_,
    new_n22690_, new_n22691_, new_n22692_, new_n22693_, new_n22694_,
    new_n22695_, new_n22696_, new_n22697_, new_n22698_, new_n22699_,
    new_n22700_, new_n22701_, new_n22702_, new_n22703_, new_n22704_,
    new_n22705_, new_n22706_, new_n22707_, new_n22708_, new_n22709_,
    new_n22710_, new_n22711_, new_n22712_, new_n22713_, new_n22714_,
    new_n22715_, new_n22716_, new_n22717_, new_n22718_, new_n22719_,
    new_n22720_, new_n22721_, new_n22722_, new_n22723_, new_n22724_,
    new_n22725_, new_n22726_, new_n22727_, new_n22728_, new_n22730_,
    new_n22731_, new_n22732_, new_n22733_, new_n22734_, new_n22735_,
    new_n22736_, new_n22737_, new_n22738_, new_n22739_, new_n22740_,
    new_n22741_, new_n22742_, new_n22743_, new_n22745_, new_n22746_,
    new_n22747_, new_n22748_, new_n22749_, new_n22750_, new_n22751_,
    new_n22752_, new_n22753_, new_n22754_, new_n22755_, new_n22756_,
    new_n22757_, new_n22758_, new_n22760_, new_n22761_, new_n22762_,
    new_n22763_, new_n22764_, new_n22765_, new_n22766_, new_n22767_,
    new_n22768_, new_n22769_, new_n22770_, new_n22771_, new_n22772_,
    new_n22773_, new_n22775_, new_n22776_, new_n22777_, new_n22778_,
    new_n22779_, new_n22780_, new_n22781_, new_n22782_, new_n22783_,
    new_n22784_, new_n22785_, new_n22786_, new_n22787_, new_n22788_,
    new_n22790_, new_n22791_, new_n22792_, new_n22793_, new_n22794_,
    new_n22796_, new_n22797_, new_n22798_, new_n22799_, new_n22800_,
    new_n22801_, new_n22802_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22877_, new_n22878_, new_n22879_, new_n22880_, new_n22881_,
    new_n22882_, new_n22883_, new_n22884_, new_n22885_, new_n22886_,
    new_n22887_, new_n22888_, new_n22889_, new_n22890_, new_n22892_,
    new_n22893_, new_n22894_, new_n22895_, new_n22896_, new_n22897_,
    new_n22898_, new_n22899_, new_n22900_, new_n22901_, new_n22902_,
    new_n22903_, new_n22904_, new_n22905_, new_n22907_, new_n22908_,
    new_n22909_, new_n22910_, new_n22911_, new_n22912_, new_n22913_,
    new_n22914_, new_n22915_, new_n22916_, new_n22917_, new_n22918_,
    new_n22919_, new_n22920_, new_n22922_, new_n22923_, new_n22924_,
    new_n22925_, new_n22926_, new_n22927_, new_n22928_, new_n22929_,
    new_n22930_, new_n22931_, new_n22932_, new_n22933_, new_n22934_,
    new_n22935_, new_n22937_, new_n22938_, new_n22939_, new_n22940_,
    new_n22941_, new_n22943_, new_n22944_, new_n22945_, new_n22946_,
    new_n22947_, new_n22948_, new_n22949_, new_n22950_, new_n22951_,
    new_n22952_, new_n22953_, new_n22954_, new_n22955_, new_n22956_,
    new_n22957_, new_n22958_, new_n22959_, new_n22960_, new_n22961_,
    new_n22962_, new_n22963_, new_n22964_, new_n22965_, new_n22966_,
    new_n22967_, new_n22968_, new_n22969_, new_n22970_, new_n22971_,
    new_n22972_, new_n22973_, new_n22974_, new_n22975_, new_n22976_,
    new_n22977_, new_n22978_, new_n22979_, new_n22980_, new_n22981_,
    new_n22982_, new_n22983_, new_n22984_, new_n22985_, new_n22986_,
    new_n22987_, new_n22988_, new_n22989_, new_n22990_, new_n22991_,
    new_n22992_, new_n22993_, new_n22994_, new_n22995_, new_n22996_,
    new_n22997_, new_n22998_, new_n22999_, new_n23000_, new_n23001_,
    new_n23002_, new_n23003_, new_n23004_, new_n23005_, new_n23006_,
    new_n23007_, new_n23008_, new_n23009_, new_n23010_, new_n23011_,
    new_n23012_, new_n23013_, new_n23014_, new_n23015_, new_n23016_,
    new_n23017_, new_n23018_, new_n23019_, new_n23020_, new_n23021_,
    new_n23022_, new_n23024_, new_n23025_, new_n23026_, new_n23027_,
    new_n23028_, new_n23029_, new_n23030_, new_n23031_, new_n23032_,
    new_n23033_, new_n23034_, new_n23035_, new_n23036_, new_n23037_,
    new_n23039_, new_n23040_, new_n23041_, new_n23042_, new_n23043_,
    new_n23044_, new_n23045_, new_n23046_, new_n23047_, new_n23048_,
    new_n23049_, new_n23050_, new_n23051_, new_n23052_, new_n23054_,
    new_n23055_, new_n23056_, new_n23057_, new_n23058_, new_n23059_,
    new_n23060_, new_n23061_, new_n23062_, new_n23063_, new_n23064_,
    new_n23065_, new_n23066_, new_n23067_, new_n23069_, new_n23070_,
    new_n23071_, new_n23072_, new_n23073_, new_n23074_, new_n23075_,
    new_n23076_, new_n23077_, new_n23078_, new_n23079_, new_n23080_,
    new_n23081_, new_n23082_, new_n23084_, new_n23085_, new_n23086_,
    new_n23087_, new_n23088_, new_n23091_, new_n23092_, new_n23093_,
    new_n23094_, new_n23095_, new_n23096_, new_n23097_, new_n23098_,
    new_n23099_, new_n23102_, new_n23103_, new_n23105_, new_n23106_,
    new_n23107_, new_n23108_, new_n23109_, new_n23110_, new_n23111_,
    new_n23112_, new_n23113_, new_n23114_, new_n23115_, new_n23117_,
    new_n23118_, new_n23119_, new_n23120_, new_n23121_, new_n23122_,
    new_n23123_, new_n23124_, new_n23125_, new_n23126_, new_n23127_,
    new_n23128_, new_n23129_, new_n23130_, new_n23131_, new_n23132_,
    new_n23133_, new_n23134_, new_n23135_, new_n23136_, new_n23137_,
    new_n23138_, new_n23139_, new_n23140_, new_n23141_, new_n23142_,
    new_n23144_, new_n23145_, new_n23146_, new_n23147_, new_n23148_,
    new_n23149_, new_n23150_, new_n23151_, new_n23153_, new_n23154_,
    new_n23155_, new_n23156_, new_n23157_, new_n23158_, new_n23160_,
    new_n23161_, new_n23163_, new_n23164_, new_n23165_, new_n23167_,
    new_n23168_, new_n23169_, new_n23170_, new_n23171_, new_n23172_,
    new_n23173_, new_n23174_, new_n23175_, new_n23176_, new_n23177_,
    new_n23178_, new_n23179_, new_n23180_, new_n23181_, new_n23182_,
    new_n23184_, new_n23185_, new_n23186_, new_n23187_, new_n23188_,
    new_n23189_, new_n23190_, new_n23192_, new_n23193_, new_n23194_,
    new_n23195_, new_n23196_, new_n23197_, new_n23198_, new_n23199_,
    new_n23200_, new_n23201_, new_n23202_, new_n23203_, new_n23204_,
    new_n23206_, new_n23207_, new_n23208_, new_n23209_, new_n23210_,
    new_n23211_, new_n23214_, new_n23215_, new_n23216_, new_n23217_,
    new_n23219_, new_n23220_, new_n23221_, new_n23222_, new_n23223_,
    new_n23224_, new_n23225_, new_n23226_, new_n23227_, new_n23228_,
    new_n23229_, new_n23230_, new_n23231_, new_n23232_, new_n23233_,
    new_n23234_, new_n23235_, new_n23236_, new_n23237_, new_n23238_,
    new_n23239_, new_n23240_, new_n23241_, new_n23244_, new_n23245_,
    new_n23246_, new_n23247_, new_n23248_, new_n23249_, new_n23250_,
    new_n23251_, new_n23252_, new_n23255_, new_n23256_, new_n23258_,
    new_n23259_, new_n23260_, new_n23261_, new_n23262_, new_n23263_,
    new_n23264_, new_n23265_, new_n23266_, new_n23267_, new_n23268_,
    new_n23270_, new_n23271_, new_n23272_, new_n23273_, new_n23274_,
    new_n23275_, new_n23277_, new_n23278_, new_n23279_, new_n23280_,
    new_n23281_, new_n23282_, new_n23283_, new_n23284_, new_n23285_,
    new_n23286_, new_n23287_, new_n23288_, new_n23289_, new_n23290_,
    new_n23291_, new_n23292_, new_n23293_, new_n23294_, new_n23295_,
    new_n23296_, new_n23297_, new_n23298_, new_n23299_, new_n23300_,
    new_n23301_, new_n23302_, new_n23304_, new_n23305_, new_n23306_,
    new_n23307_, new_n23308_, new_n23309_, new_n23310_, new_n23311_,
    new_n23312_, new_n23314_, new_n23315_, new_n23316_, new_n23317_,
    new_n23318_, new_n23319_, new_n23320_, new_n23321_, new_n23322_,
    new_n23323_, new_n23324_, new_n23325_, new_n23326_, new_n23327_,
    new_n23328_, new_n23329_, new_n23330_, new_n23331_, new_n23332_,
    new_n23333_, new_n23334_, new_n23335_, new_n23336_, new_n23337_,
    new_n23338_, new_n23339_, new_n23340_, new_n23341_, new_n23343_,
    new_n23344_, new_n23345_, new_n23346_, new_n23347_, new_n23348_,
    new_n23349_, new_n23350_, new_n23352_, new_n23353_, new_n23354_,
    new_n23355_, new_n23356_, new_n23357_, new_n23358_, new_n23359_,
    new_n23360_, new_n23361_, new_n23362_, new_n23363_, new_n23364_,
    new_n23365_, new_n23366_, new_n23367_, new_n23368_, new_n23369_,
    new_n23370_, new_n23371_, new_n23372_, new_n23373_, new_n23374_,
    new_n23375_, new_n23376_, new_n23377_, new_n23378_, new_n23379_,
    new_n23381_, new_n23382_, new_n23383_, new_n23384_, new_n23385_,
    new_n23386_, new_n23387_, new_n23388_, new_n23390_, new_n23391_,
    new_n23392_, new_n23393_, new_n23394_, new_n23395_, new_n23396_,
    new_n23397_, new_n23398_, new_n23399_, new_n23400_, new_n23401_,
    new_n23402_, new_n23403_, new_n23404_, new_n23405_, new_n23406_,
    new_n23407_, new_n23408_, new_n23409_, new_n23410_, new_n23411_,
    new_n23412_, new_n23413_, new_n23414_, new_n23415_, new_n23416_,
    new_n23417_, new_n23418_, new_n23419_, new_n23420_, new_n23422_,
    new_n23423_, new_n23424_, new_n23425_, new_n23426_, new_n23427_,
    new_n23428_, new_n23429_, new_n23431_, new_n23432_, new_n23433_,
    new_n23434_, new_n23435_, new_n23436_, new_n23437_, new_n23438_,
    new_n23439_, new_n23440_, new_n23441_, new_n23442_, new_n23443_,
    new_n23444_, new_n23445_, new_n23446_, new_n23447_, new_n23448_,
    new_n23449_, new_n23450_, new_n23451_, new_n23452_, new_n23453_,
    new_n23454_, new_n23455_, new_n23456_, new_n23457_, new_n23458_,
    new_n23459_, new_n23461_, new_n23462_, new_n23463_, new_n23464_,
    new_n23465_, new_n23466_, new_n23467_, new_n23468_, new_n23470_,
    new_n23471_, new_n23472_, new_n23473_, new_n23474_, new_n23475_,
    new_n23476_, new_n23477_, new_n23478_, new_n23479_, new_n23480_,
    new_n23481_, new_n23482_, new_n23483_, new_n23484_, new_n23485_,
    new_n23486_, new_n23487_, new_n23488_, new_n23489_, new_n23490_,
    new_n23491_, new_n23492_, new_n23493_, new_n23494_, new_n23495_,
    new_n23496_, new_n23497_, new_n23498_, new_n23499_, new_n23500_,
    new_n23502_, new_n23503_, new_n23504_, new_n23505_, new_n23506_,
    new_n23507_, new_n23508_, new_n23509_, new_n23510_, new_n23511_,
    new_n23512_, new_n23514_, new_n23515_, new_n23516_, new_n23517_,
    new_n23518_, new_n23519_, new_n23520_, new_n23521_, new_n23522_,
    new_n23523_, new_n23524_, new_n23525_, new_n23526_, new_n23528_,
    new_n23529_, new_n23530_, new_n23532_, new_n23533_, new_n23534_,
    new_n23536_, new_n23537_, new_n23538_, new_n23539_, new_n23540_,
    new_n23541_, new_n23542_, new_n23543_, new_n23544_, new_n23545_,
    new_n23548_, new_n23549_, new_n23550_, new_n23551_, new_n23553_,
    new_n23554_, new_n23555_, new_n23556_, new_n23557_, new_n23559_,
    new_n23560_, new_n23562_, new_n23563_, new_n23564_, new_n23565_,
    new_n23566_, new_n23567_, new_n23568_, new_n23569_, new_n23570_,
    new_n23571_, new_n23572_, new_n23573_, new_n23574_, new_n23575_,
    new_n23576_, new_n23577_, new_n23578_, new_n23579_, new_n23580_,
    new_n23581_, new_n23582_, new_n23583_, new_n23584_, new_n23585_,
    new_n23586_, new_n23587_, new_n23588_, new_n23589_, new_n23590_,
    new_n23591_, new_n23592_, new_n23593_, new_n23594_, new_n23595_,
    new_n23596_, new_n23597_, new_n23598_, new_n23599_, new_n23600_,
    new_n23601_, new_n23602_, new_n23603_, new_n23604_, new_n23605_,
    new_n23606_, new_n23607_, new_n23608_, new_n23609_, new_n23610_,
    new_n23611_, new_n23612_, new_n23614_, new_n23615_, new_n23616_,
    new_n23617_, new_n23618_, new_n23619_, new_n23620_, new_n23621_,
    new_n23622_, new_n23623_, new_n23625_, new_n23626_, new_n23627_,
    new_n23628_, new_n23630_, new_n23632_, new_n23635_, new_n23636_,
    new_n23637_, new_n23639_, new_n23640_, new_n23641_, new_n23642_,
    new_n23643_, new_n23645_, new_n23646_, new_n23647_, new_n23648_,
    new_n23649_, new_n23650_, new_n23651_, new_n23652_, new_n23653_,
    new_n23654_, new_n23656_, new_n23657_, new_n23658_, new_n23659_,
    new_n23661_, new_n23662_, new_n23663_, new_n23664_, new_n23665_,
    new_n23668_, new_n23669_, new_n23670_, new_n23672_, new_n23673_,
    new_n23674_, new_n23675_, new_n23676_, new_n23679_, new_n23680_,
    new_n23681_, new_n23682_, new_n23683_, new_n23684_, new_n23685_,
    new_n23686_, new_n23687_, new_n23690_, new_n23691_, new_n23693_,
    new_n23694_, new_n23695_, new_n23696_, new_n23697_, new_n23698_,
    new_n23699_, new_n23700_, new_n23701_, new_n23702_, new_n23703_,
    new_n23705_, new_n23706_, new_n23707_, new_n23708_, new_n23709_,
    new_n23710_, new_n23711_, new_n23712_, new_n23713_, new_n23714_,
    new_n23715_, new_n23716_, new_n23717_, new_n23718_, new_n23719_,
    new_n23720_, new_n23721_, new_n23722_, new_n23723_, new_n23724_,
    new_n23725_, new_n23726_, new_n23727_, new_n23728_, new_n23729_,
    new_n23730_, new_n23731_, new_n23732_, new_n23733_, new_n23734_,
    new_n23735_, new_n23736_, new_n23737_, new_n23738_, new_n23739_,
    new_n23740_, new_n23741_, new_n23742_, new_n23743_, new_n23744_,
    new_n23745_, new_n23746_, new_n23747_, new_n23748_, new_n23749_,
    new_n23750_, new_n23751_, new_n23752_, new_n23753_, new_n23754_,
    new_n23755_, new_n23756_, new_n23757_, new_n23758_, new_n23759_,
    new_n23760_, new_n23761_, new_n23762_, new_n23763_, new_n23764_,
    new_n23765_, new_n23767_, new_n23768_, new_n23769_, new_n23770_,
    new_n23771_, new_n23772_, new_n23773_, new_n23774_, new_n23775_,
    new_n23776_, new_n23777_, new_n23778_, new_n23779_, new_n23780_,
    new_n23782_, new_n23783_, new_n23784_, new_n23785_, new_n23786_,
    new_n23787_, new_n23788_, new_n23789_, new_n23790_, new_n23791_,
    new_n23792_, new_n23793_, new_n23794_, new_n23795_, new_n23797_,
    new_n23798_, new_n23799_, new_n23800_, new_n23801_, new_n23802_,
    new_n23803_, new_n23804_, new_n23805_, new_n23806_, new_n23807_,
    new_n23808_, new_n23809_, new_n23810_, new_n23812_, new_n23813_,
    new_n23814_, new_n23815_, new_n23816_, new_n23817_, new_n23818_,
    new_n23819_, new_n23820_, new_n23821_, new_n23822_, new_n23823_,
    new_n23824_, new_n23825_, new_n23827_, new_n23828_, new_n23829_,
    new_n23830_, new_n23831_, new_n23832_, new_n23833_, new_n23834_,
    new_n23835_, new_n23836_, new_n23837_, new_n23838_, new_n23839_,
    new_n23840_, new_n23842_, new_n23843_, new_n23844_, new_n23845_,
    new_n23846_, new_n23847_, new_n23848_, new_n23849_, new_n23850_,
    new_n23851_, new_n23852_, new_n23853_, new_n23854_, new_n23855_,
    new_n23857_, new_n23858_, new_n23859_, new_n23860_, new_n23861_,
    new_n23862_, new_n23863_, new_n23864_, new_n23865_, new_n23866_,
    new_n23867_, new_n23868_, new_n23869_, new_n23870_, new_n23872_,
    new_n23873_, new_n23874_, new_n23875_, new_n23876_, new_n23877_,
    new_n23879_, new_n23880_, new_n23882_, new_n23883_, new_n23885_,
    new_n23886_, new_n23888_, new_n23889_, new_n23891_, new_n23892_,
    new_n23894_, new_n23895_, new_n23897_, new_n23898_, new_n23900_,
    new_n23901_, new_n23902_, new_n23903_, new_n23904_, new_n23905_,
    new_n23906_, new_n23907_, new_n23908_, new_n23909_, new_n23910_,
    new_n23911_, new_n23912_, new_n23913_, new_n23915_, new_n23916_,
    new_n23917_, new_n23918_, new_n23919_, new_n23920_, new_n23921_,
    new_n23922_, new_n23923_, new_n23924_, new_n23925_, new_n23926_,
    new_n23927_, new_n23928_, new_n23930_, new_n23931_, new_n23932_,
    new_n23933_, new_n23934_, new_n23935_, new_n23936_, new_n23937_,
    new_n23938_, new_n23939_, new_n23940_, new_n23941_, new_n23942_,
    new_n23943_, new_n23945_, new_n23946_, new_n23947_, new_n23948_,
    new_n23949_, new_n23950_, new_n23951_, new_n23952_, new_n23953_,
    new_n23954_, new_n23955_, new_n23956_, new_n23957_, new_n23958_,
    new_n23960_, new_n23961_, new_n23962_, new_n23963_, new_n23964_,
    new_n23965_, new_n23966_, new_n23967_, new_n23968_, new_n23969_,
    new_n23970_, new_n23971_, new_n23972_, new_n23973_, new_n23975_,
    new_n23976_, new_n23977_, new_n23978_, new_n23979_, new_n23980_,
    new_n23981_, new_n23982_, new_n23983_, new_n23984_, new_n23985_,
    new_n23986_, new_n23987_, new_n23988_, new_n23990_, new_n23991_,
    new_n23992_, new_n23993_, new_n23994_, new_n23995_, new_n23996_,
    new_n23997_, new_n23998_, new_n23999_, new_n24000_, new_n24001_,
    new_n24002_, new_n24003_, new_n24005_, new_n24006_, new_n24007_,
    new_n24008_, new_n24009_, new_n24010_, new_n24011_, new_n24012_,
    new_n24013_, new_n24014_, new_n24015_, new_n24016_, new_n24017_,
    new_n24018_, new_n24020_, new_n24021_, new_n24022_, new_n24023_,
    new_n24024_, new_n24025_, new_n24027_, new_n24028_, new_n24030_,
    new_n24031_, new_n24033_, new_n24034_, new_n24036_, new_n24037_,
    new_n24039_, new_n24040_, new_n24042_, new_n24043_, new_n24045_,
    new_n24046_, new_n24048_, new_n24049_, new_n24050_, new_n24051_,
    new_n24052_, new_n24053_, new_n24054_, new_n24055_, new_n24056_,
    new_n24057_, new_n24058_, new_n24059_, new_n24060_, new_n24061_,
    new_n24062_, new_n24063_, new_n24064_, new_n24065_, new_n24066_,
    new_n24067_, new_n24068_, new_n24069_, new_n24070_, new_n24071_,
    new_n24072_, new_n24073_, new_n24075_, new_n24076_, new_n24077_,
    new_n24078_, new_n24079_, new_n24080_, new_n24081_, new_n24082_,
    new_n24083_, new_n24084_, new_n24085_, new_n24086_, new_n24087_,
    new_n24088_, new_n24089_, new_n24090_, new_n24091_, new_n24093_,
    new_n24094_, new_n24095_, new_n24096_, new_n24097_, new_n24098_,
    new_n24099_, new_n24100_, new_n24101_, new_n24102_, new_n24103_,
    new_n24104_, new_n24105_, new_n24106_, new_n24107_, new_n24108_,
    new_n24109_, new_n24111_, new_n24112_, new_n24113_, new_n24114_,
    new_n24115_, new_n24116_, new_n24117_, new_n24118_, new_n24119_,
    new_n24120_, new_n24121_, new_n24122_, new_n24123_, new_n24124_,
    new_n24125_, new_n24126_, new_n24127_, new_n24129_, new_n24130_,
    new_n24131_, new_n24132_, new_n24133_, new_n24134_, new_n24135_,
    new_n24136_, new_n24137_, new_n24138_, new_n24139_, new_n24140_,
    new_n24141_, new_n24142_, new_n24143_, new_n24144_, new_n24145_,
    new_n24147_, new_n24148_, new_n24149_, new_n24150_, new_n24151_,
    new_n24152_, new_n24153_, new_n24154_, new_n24155_, new_n24156_,
    new_n24157_, new_n24158_, new_n24159_, new_n24160_, new_n24161_,
    new_n24162_, new_n24163_, new_n24165_, new_n24166_, new_n24167_,
    new_n24168_, new_n24169_, new_n24170_, new_n24171_, new_n24172_,
    new_n24173_, new_n24174_, new_n24175_, new_n24176_, new_n24177_,
    new_n24178_, new_n24179_, new_n24180_, new_n24181_, new_n24183_,
    new_n24184_, new_n24185_, new_n24186_, new_n24187_, new_n24188_,
    new_n24189_, new_n24190_, new_n24191_, new_n24192_, new_n24193_,
    new_n24194_, new_n24195_, new_n24196_, new_n24197_, new_n24198_,
    new_n24199_, new_n24201_, new_n24202_, new_n24203_, new_n24204_,
    new_n24205_, new_n24206_, new_n24208_, new_n24209_, new_n24211_,
    new_n24212_, new_n24214_, new_n24215_, new_n24217_, new_n24218_,
    new_n24220_, new_n24221_, new_n24223_, new_n24224_, new_n24226_,
    new_n24227_, new_n24229_, new_n24230_, new_n24231_, new_n24232_,
    new_n24233_, new_n24234_, new_n24235_, new_n24236_, new_n24237_,
    new_n24238_, new_n24239_, new_n24240_, new_n24241_, new_n24242_,
    new_n24243_, new_n24244_, new_n24245_, new_n24246_, new_n24247_,
    new_n24248_, new_n24249_, new_n24250_, new_n24251_, new_n24252_,
    new_n24253_, new_n24254_, new_n24255_, new_n24256_, new_n24257_,
    new_n24258_, new_n24259_, new_n24261_, new_n24262_, new_n24263_,
    new_n24264_, new_n24265_, new_n24266_, new_n24267_, new_n24268_,
    new_n24269_, new_n24270_, new_n24271_, new_n24272_, new_n24273_,
    new_n24274_, new_n24275_, new_n24276_, new_n24277_, new_n24278_,
    new_n24280_, new_n24281_, new_n24282_, new_n24283_, new_n24284_,
    new_n24285_, new_n24286_, new_n24287_, new_n24288_, new_n24289_,
    new_n24290_, new_n24291_, new_n24292_, new_n24293_, new_n24294_,
    new_n24295_, new_n24296_, new_n24297_, new_n24299_, new_n24300_,
    new_n24301_, new_n24302_, new_n24303_, new_n24304_, new_n24305_,
    new_n24306_, new_n24307_, new_n24308_, new_n24309_, new_n24310_,
    new_n24311_, new_n24312_, new_n24313_, new_n24314_, new_n24315_,
    new_n24316_, new_n24318_, new_n24319_, new_n24320_, new_n24321_,
    new_n24322_, new_n24323_, new_n24324_, new_n24325_, new_n24326_,
    new_n24327_, new_n24328_, new_n24329_, new_n24330_, new_n24331_,
    new_n24332_, new_n24333_, new_n24334_, new_n24335_, new_n24337_,
    new_n24338_, new_n24339_, new_n24340_, new_n24341_, new_n24342_,
    new_n24343_, new_n24344_, new_n24345_, new_n24346_, new_n24347_,
    new_n24348_, new_n24349_, new_n24350_, new_n24351_, new_n24352_,
    new_n24353_, new_n24354_, new_n24356_, new_n24357_, new_n24358_,
    new_n24359_, new_n24360_, new_n24361_, new_n24362_, new_n24363_,
    new_n24364_, new_n24365_, new_n24366_, new_n24367_, new_n24368_,
    new_n24369_, new_n24370_, new_n24371_, new_n24372_, new_n24373_,
    new_n24375_, new_n24376_, new_n24377_, new_n24378_, new_n24379_,
    new_n24380_, new_n24381_, new_n24382_, new_n24383_, new_n24384_,
    new_n24385_, new_n24386_, new_n24387_, new_n24388_, new_n24389_,
    new_n24390_, new_n24391_, new_n24392_, new_n24394_, new_n24395_,
    new_n24396_, new_n24397_, new_n24398_, new_n24399_, new_n24400_,
    new_n24401_, new_n24403_, new_n24404_, new_n24405_, new_n24407_,
    new_n24408_, new_n24410_, new_n24411_, new_n24413_, new_n24414_,
    new_n24416_, new_n24417_, new_n24419_, new_n24420_, new_n24422_,
    new_n24423_, new_n24425_, new_n24426_, new_n24427_, new_n24428_,
    new_n24429_, new_n24430_, new_n24431_, new_n24432_, new_n24433_,
    new_n24434_, new_n24435_, new_n24436_, new_n24437_, new_n24438_,
    new_n24440_, new_n24441_, new_n24442_, new_n24443_, new_n24444_,
    new_n24445_, new_n24447_, new_n24448_, new_n24450_, new_n24452_,
    new_n24453_, new_n24454_, new_n24455_, new_n24456_, new_n24458_,
    new_n24459_, new_n24460_, new_n24462_, new_n24463_, new_n24464_,
    new_n24465_, new_n24466_, new_n24467_, new_n24468_, new_n24469_,
    new_n24470_, new_n24471_, new_n24472_, new_n24473_, new_n24474_,
    new_n24475_, new_n24476_, new_n24478_, new_n24479_, new_n24480_,
    new_n24481_, new_n24482_, new_n24483_, new_n24484_, new_n24485_,
    new_n24486_, new_n24487_, new_n24488_, new_n24489_, new_n24490_,
    new_n24492_, new_n24493_, new_n24494_, new_n24495_, new_n24496_,
    new_n24497_, new_n24498_, new_n24499_, new_n24500_, new_n24501_,
    new_n24502_, new_n24503_, new_n24505_, new_n24506_, new_n24507_,
    new_n24508_, new_n24509_, new_n24510_, new_n24512_, new_n24513_,
    new_n24514_, new_n24515_, new_n24517_, new_n24518_, new_n24520_,
    new_n24521_, new_n24522_, new_n24523_, new_n24524_, new_n24527_,
    new_n24528_, new_n24529_, new_n24530_, new_n24531_, new_n24532_,
    new_n24533_, new_n24534_, new_n24535_, new_n24536_, new_n24537_,
    new_n24538_, new_n24539_, new_n24541_, new_n24542_, new_n24543_,
    new_n24545_, new_n24546_, new_n24547_, new_n24549_, new_n24550_,
    new_n24551_, new_n24552_, new_n24553_, new_n24554_, new_n24555_,
    new_n24556_, new_n24557_, new_n24558_, new_n24559_, new_n24560_,
    new_n24561_, new_n24562_, new_n24563_, new_n24564_, new_n24565_,
    new_n24566_, new_n24567_, new_n24568_, new_n24569_, new_n24570_,
    new_n24571_, new_n24572_, new_n24573_, new_n24574_, new_n24575_,
    new_n24576_, new_n24577_, new_n24578_, new_n24579_, new_n24580_,
    new_n24581_, new_n24582_, new_n24583_, new_n24585_, new_n24586_,
    new_n24587_, new_n24588_, new_n24589_, new_n24590_, new_n24591_,
    new_n24592_, new_n24593_, new_n24595_, new_n24597_, new_n24599_,
    new_n24600_, new_n24601_, new_n24603_, new_n24604_, new_n24605_,
    new_n24606_, new_n24610_, new_n24611_, new_n24612_, new_n24613_,
    new_n24614_, new_n24615_, new_n24616_, new_n24617_, new_n24618_,
    new_n24619_, new_n24620_, new_n24621_, new_n24622_, new_n24623_,
    new_n24624_, new_n24625_, new_n24626_, new_n24627_, new_n24628_,
    new_n24629_, new_n24630_, new_n24631_, new_n24632_, new_n24633_,
    new_n24634_, new_n24635_, new_n24636_, new_n24637_, new_n24638_,
    new_n24639_, new_n24640_, new_n24641_, new_n24642_, new_n24643_,
    new_n24644_, new_n24645_, new_n24646_, new_n24647_, new_n24648_,
    new_n24649_, new_n24650_, new_n24651_, new_n24652_, new_n24653_,
    new_n24654_, new_n24655_, new_n24656_, new_n24657_, new_n24658_,
    new_n24659_, new_n24660_, new_n24661_, new_n24662_, new_n24663_,
    new_n24664_, new_n24665_, new_n24666_, new_n24667_, new_n24668_,
    new_n24669_, new_n24670_, new_n24671_, new_n24672_, new_n24673_,
    new_n24674_, new_n24675_, new_n24676_, new_n24677_, new_n24678_,
    new_n24679_, new_n24680_, new_n24681_, new_n24682_, new_n24683_,
    new_n24684_, new_n24685_, new_n24686_, new_n24687_, new_n24688_,
    new_n24689_, new_n24690_, new_n24691_, new_n24692_, new_n24693_,
    new_n24694_, new_n24695_, new_n24696_, new_n24697_, new_n24698_,
    new_n24699_, new_n24700_, new_n24701_, new_n24702_, new_n24703_,
    new_n24704_, new_n24705_, new_n24706_, new_n24707_, new_n24708_,
    new_n24709_, new_n24710_, new_n24711_, new_n24712_, new_n24713_,
    new_n24714_, new_n24715_, new_n24716_, new_n24717_, new_n24718_,
    new_n24719_, new_n24720_, new_n24721_, new_n24722_, new_n24723_,
    new_n24724_, new_n24725_, new_n24726_, new_n24727_, new_n24728_,
    new_n24729_, new_n24730_, new_n24731_, new_n24732_, new_n24733_,
    new_n24734_, new_n24735_, new_n24736_, new_n24737_, new_n24738_,
    new_n24739_, new_n24740_, new_n24741_, new_n24742_, new_n24743_,
    new_n24744_, new_n24745_, new_n24746_, new_n24747_, new_n24748_,
    new_n24749_, new_n24750_, new_n24751_, new_n24752_, new_n24753_,
    new_n24754_, new_n24755_, new_n24756_, new_n24757_, new_n24758_,
    new_n24759_, new_n24760_, new_n24761_, new_n24762_, new_n24763_,
    new_n24764_, new_n24765_, new_n24766_, new_n24767_, new_n24768_,
    new_n24769_, new_n24770_, new_n24771_, new_n24772_, new_n24773_,
    new_n24774_, new_n24775_, new_n24776_, new_n24777_, new_n24778_,
    new_n24779_, new_n24780_, new_n24781_, new_n24782_, new_n24783_,
    new_n24784_, new_n24785_, new_n24786_, new_n24787_, new_n24788_,
    new_n24789_, new_n24790_, new_n24791_, new_n24792_, new_n24793_,
    new_n24794_, new_n24795_, new_n24796_, new_n24797_, new_n24798_,
    new_n24799_, new_n24800_, new_n24801_, new_n24802_, new_n24803_,
    new_n24804_, new_n24805_, new_n24806_, new_n24807_, new_n24808_,
    new_n24809_, new_n24810_, new_n24811_, new_n24812_, new_n24813_,
    new_n24814_, new_n24815_, new_n24816_, new_n24817_, new_n24818_,
    new_n24819_, new_n24820_, new_n24821_, new_n24822_, new_n24823_,
    new_n24824_, new_n24825_, new_n24826_, new_n24827_, new_n24828_,
    new_n24829_, new_n24830_, new_n24831_, new_n24832_, new_n24833_,
    new_n24834_, new_n24835_, new_n24836_, new_n24837_, new_n24838_,
    new_n24839_, new_n24840_, new_n24841_, new_n24842_, new_n24843_,
    new_n24844_, new_n24845_, new_n24846_, new_n24847_, new_n24848_,
    new_n24849_, new_n24850_, new_n24851_, new_n24852_, new_n24853_,
    new_n24854_, new_n24855_, new_n24856_, new_n24857_, new_n24858_,
    new_n24859_, new_n24860_, new_n24861_, new_n24862_, new_n24863_,
    new_n24864_, new_n24865_, new_n24866_, new_n24867_, new_n24868_,
    new_n24869_, new_n24870_, new_n24871_, new_n24872_, new_n24873_,
    new_n24874_, new_n24875_, new_n24876_, new_n24877_, new_n24878_,
    new_n24879_, new_n24880_, new_n24881_, new_n24882_, new_n24883_,
    new_n24884_, new_n24885_, new_n24886_, new_n24887_, new_n24888_,
    new_n24889_, new_n24890_, new_n24891_, new_n24892_, new_n24893_,
    new_n24894_, new_n24895_, new_n24896_, new_n24897_, new_n24898_,
    new_n24899_, new_n24900_, new_n24901_, new_n24902_, new_n24903_,
    new_n24904_, new_n24905_, new_n24906_, new_n24907_, new_n24908_,
    new_n24909_, new_n24910_, new_n24911_, new_n24912_, new_n24913_,
    new_n24914_, new_n24915_, new_n24916_, new_n24917_, new_n24918_,
    new_n24919_, new_n24920_, new_n24921_, new_n24922_, new_n24923_,
    new_n24924_, new_n24925_, new_n24926_, new_n24927_, new_n24928_,
    new_n24929_, new_n24930_, new_n24931_, new_n24932_, new_n24933_,
    new_n24934_, new_n24935_, new_n24936_, new_n24937_, new_n24938_,
    new_n24939_, new_n24940_, new_n24941_, new_n24942_, new_n24943_,
    new_n24944_, new_n24945_, new_n24946_, new_n24947_, new_n24948_,
    new_n24949_, new_n24950_, new_n24951_, new_n24952_, new_n24953_,
    new_n24954_, new_n24955_, new_n24956_, new_n24957_, new_n24958_,
    new_n24959_, new_n24960_, new_n24961_, new_n24962_, new_n24963_,
    new_n24964_, new_n24965_, new_n24966_, new_n24967_, new_n24968_,
    new_n24969_, new_n24970_, new_n24971_, new_n24972_, new_n24973_,
    new_n24974_, new_n24975_, new_n24976_, new_n24977_, new_n24978_,
    new_n24979_, new_n24980_, new_n24981_, new_n24982_, new_n24983_,
    new_n24984_, new_n24985_, new_n24986_, new_n24987_, new_n24988_,
    new_n24989_, new_n24990_, new_n24991_, new_n24992_, new_n24993_,
    new_n24994_, new_n24995_, new_n24996_, new_n24997_, new_n24998_,
    new_n24999_, new_n25000_, new_n25001_, new_n25002_, new_n25003_,
    new_n25004_, new_n25005_, new_n25006_, new_n25007_, new_n25008_,
    new_n25009_, new_n25010_, new_n25011_, new_n25012_, new_n25013_,
    new_n25014_, new_n25015_, new_n25016_, new_n25017_, new_n25018_,
    new_n25019_, new_n25020_, new_n25021_, new_n25022_, new_n25023_,
    new_n25024_, new_n25025_, new_n25026_, new_n25027_, new_n25028_,
    new_n25029_, new_n25030_, new_n25031_, new_n25032_, new_n25033_,
    new_n25034_, new_n25035_, new_n25036_, new_n25037_, new_n25038_,
    new_n25039_, new_n25040_, new_n25041_, new_n25042_, new_n25043_,
    new_n25044_, new_n25045_, new_n25046_, new_n25047_, new_n25048_,
    new_n25049_, new_n25050_, new_n25051_, new_n25052_, new_n25053_,
    new_n25054_, new_n25055_, new_n25056_, new_n25057_, new_n25058_,
    new_n25059_, new_n25060_, new_n25061_, new_n25062_, new_n25063_,
    new_n25064_, new_n25065_, new_n25066_, new_n25067_, new_n25068_,
    new_n25069_, new_n25070_, new_n25071_, new_n25072_, new_n25073_,
    new_n25074_, new_n25075_, new_n25076_, new_n25077_, new_n25078_,
    new_n25079_, new_n25080_, new_n25081_, new_n25082_, new_n25083_,
    new_n25084_, new_n25085_, new_n25086_, new_n25087_, new_n25088_,
    new_n25089_, new_n25090_, new_n25091_, new_n25092_, new_n25093_,
    new_n25094_, new_n25095_, new_n25096_, new_n25097_, new_n25098_,
    new_n25099_, new_n25100_, new_n25101_, new_n25102_, new_n25103_,
    new_n25104_, new_n25105_, new_n25106_, new_n25107_, new_n25108_,
    new_n25109_, new_n25110_, new_n25111_, new_n25112_, new_n25113_,
    new_n25114_, new_n25115_, new_n25116_, new_n25117_, new_n25118_,
    new_n25119_, new_n25120_, new_n25121_, new_n25122_, new_n25123_,
    new_n25124_, new_n25125_, new_n25126_, new_n25127_, new_n25128_,
    new_n25129_, new_n25130_, new_n25131_, new_n25132_, new_n25133_,
    new_n25134_, new_n25135_, new_n25136_, new_n25137_, new_n25138_,
    new_n25139_, new_n25140_, new_n25141_, new_n25142_, new_n25143_,
    new_n25144_, new_n25145_, new_n25146_, new_n25147_, new_n25148_,
    new_n25149_, new_n25150_, new_n25151_, new_n25152_, new_n25153_,
    new_n25154_, new_n25155_, new_n25156_, new_n25157_, new_n25158_,
    new_n25159_, new_n25160_, new_n25161_, new_n25162_, new_n25163_,
    new_n25164_, new_n25165_, new_n25166_, new_n25167_, new_n25168_,
    new_n25169_, new_n25170_, new_n25171_, new_n25172_, new_n25173_,
    new_n25174_, new_n25175_, new_n25176_, new_n25177_, new_n25178_,
    new_n25179_, new_n25180_, new_n25181_, new_n25182_, new_n25183_,
    new_n25184_, new_n25185_, new_n25186_, new_n25187_, new_n25188_,
    new_n25189_, new_n25190_, new_n25191_, new_n25192_, new_n25193_,
    new_n25194_, new_n25195_, new_n25196_, new_n25197_, new_n25198_,
    new_n25199_, new_n25200_, new_n25201_, new_n25202_, new_n25203_,
    new_n25204_, new_n25205_, new_n25206_, new_n25207_, new_n25208_,
    new_n25209_, new_n25210_, new_n25211_, new_n25212_, new_n25213_,
    new_n25214_, new_n25215_, new_n25216_, new_n25217_, new_n25218_,
    new_n25219_, new_n25220_, new_n25221_, new_n25222_, new_n25223_,
    new_n25224_, new_n25225_, new_n25226_, new_n25227_, new_n25228_,
    new_n25229_, new_n25230_, new_n25231_, new_n25232_, new_n25233_,
    new_n25234_, new_n25235_, new_n25236_, new_n25237_, new_n25238_,
    new_n25239_, new_n25240_, new_n25241_, new_n25242_, new_n25243_,
    new_n25244_, new_n25245_, new_n25246_, new_n25247_, new_n25248_,
    new_n25249_, new_n25250_, new_n25251_, new_n25252_, new_n25253_,
    new_n25254_, new_n25255_, new_n25256_, new_n25257_, new_n25258_,
    new_n25259_, new_n25260_, new_n25261_, new_n25262_, new_n25263_,
    new_n25264_, new_n25265_, new_n25266_, new_n25267_, new_n25268_,
    new_n25269_, new_n25270_, new_n25271_, new_n25272_, new_n25273_,
    new_n25274_, new_n25275_, new_n25276_, new_n25277_, new_n25278_,
    new_n25279_, new_n25280_, new_n25281_, new_n25282_, new_n25283_,
    new_n25284_, new_n25285_, new_n25286_, new_n25287_, new_n25288_,
    new_n25289_, new_n25290_, new_n25291_, new_n25292_, new_n25293_,
    new_n25294_, new_n25295_, new_n25296_, new_n25297_, new_n25298_,
    new_n25299_, new_n25300_, new_n25301_, new_n25302_, new_n25303_,
    new_n25304_, new_n25305_, new_n25306_, new_n25307_, new_n25308_,
    new_n25309_, new_n25310_, new_n25311_, new_n25312_, new_n25313_,
    new_n25314_, new_n25315_, new_n25316_, new_n25317_, new_n25318_,
    new_n25319_, new_n25320_, new_n25321_, new_n25322_, new_n25323_,
    new_n25324_, new_n25325_, new_n25326_, new_n25327_, new_n25328_,
    new_n25329_, new_n25330_, new_n25331_, new_n25332_, new_n25333_,
    new_n25334_, new_n25335_, new_n25336_, new_n25337_, new_n25338_,
    new_n25339_, new_n25340_, new_n25341_, new_n25342_, new_n25343_,
    new_n25344_, new_n25345_, new_n25346_, new_n25347_, new_n25348_,
    new_n25349_, new_n25350_, new_n25351_, new_n25352_, new_n25353_,
    new_n25354_, new_n25355_, new_n25356_, new_n25357_, new_n25358_,
    new_n25359_, new_n25360_, new_n25361_, new_n25362_, new_n25363_,
    new_n25364_, new_n25365_, new_n25366_, new_n25367_, new_n25368_,
    new_n25369_, new_n25370_, new_n25371_, new_n25372_, new_n25373_,
    new_n25374_, new_n25375_, new_n25376_, new_n25377_, new_n25378_,
    new_n25379_, new_n25380_, new_n25381_, new_n25382_, new_n25383_,
    new_n25384_, new_n25385_, new_n25386_, new_n25387_, new_n25388_,
    new_n25389_, new_n25390_, new_n25391_, new_n25392_, new_n25393_,
    new_n25394_, new_n25395_, new_n25396_, new_n25397_, new_n25398_,
    new_n25399_, new_n25400_, new_n25401_, new_n25402_, new_n25403_,
    new_n25404_, new_n25405_, new_n25406_, new_n25408_, new_n25409_,
    new_n25410_, new_n25411_, new_n25412_, new_n25413_, new_n25414_,
    new_n25415_, new_n25416_, new_n25417_, new_n25418_, new_n25419_,
    new_n25420_, new_n25421_, new_n25422_, new_n25423_, new_n25424_,
    new_n25425_, new_n25426_, new_n25427_, new_n25428_, new_n25429_,
    new_n25430_, new_n25431_, new_n25432_, new_n25433_, new_n25434_,
    new_n25435_, new_n25436_, new_n25437_, new_n25438_, new_n25439_,
    new_n25440_, new_n25441_, new_n25442_, new_n25443_, new_n25444_,
    new_n25445_, new_n25446_, new_n25447_, new_n25448_, new_n25449_,
    new_n25450_, new_n25451_, new_n25452_, new_n25453_, new_n25454_,
    new_n25455_, new_n25456_, new_n25457_, new_n25458_, new_n25459_,
    new_n25460_, new_n25461_, new_n25462_, new_n25463_, new_n25464_,
    new_n25465_, new_n25466_, new_n25467_, new_n25468_, new_n25469_,
    new_n25470_, new_n25471_, new_n25472_, new_n25474_, new_n25475_,
    new_n25476_, new_n25477_, new_n25478_, new_n25479_, new_n25480_,
    new_n25481_, new_n25482_, new_n25483_, new_n25484_, new_n25485_,
    new_n25486_, new_n25487_, new_n25488_, new_n25489_, new_n25490_,
    new_n25491_, new_n25492_, new_n25493_, new_n25494_, new_n25495_,
    new_n25496_, new_n25497_, new_n25498_, new_n25499_, new_n25500_,
    new_n25501_, new_n25502_, new_n25503_, new_n25504_, new_n25505_,
    new_n25506_, new_n25507_, new_n25508_, new_n25509_, new_n25510_,
    new_n25511_, new_n25512_, new_n25513_, new_n25514_, new_n25515_,
    new_n25516_, new_n25517_, new_n25518_, new_n25519_, new_n25520_,
    new_n25521_, new_n25522_, new_n25523_, new_n25524_, new_n25525_,
    new_n25526_, new_n25527_, new_n25528_, new_n25529_, new_n25530_,
    new_n25531_, new_n25532_, new_n25533_, new_n25534_, new_n25535_,
    new_n25536_, new_n25537_, new_n25538_, new_n25539_, new_n25540_,
    new_n25541_, new_n25542_, new_n25543_, new_n25544_, new_n25546_,
    new_n25547_, new_n25548_, new_n25549_, new_n25550_, new_n25551_,
    new_n25552_, new_n25553_, new_n25554_, new_n25555_, new_n25556_,
    new_n25557_, new_n25558_, new_n25559_, new_n25560_, new_n25561_,
    new_n25562_, new_n25563_, new_n25564_, new_n25565_, new_n25566_,
    new_n25567_, new_n25568_, new_n25569_, new_n25570_, new_n25571_,
    new_n25572_, new_n25573_, new_n25574_, new_n25575_, new_n25576_,
    new_n25577_, new_n25578_, new_n25579_, new_n25580_, new_n25581_,
    new_n25582_, new_n25583_, new_n25584_, new_n25585_, new_n25586_,
    new_n25587_, new_n25588_, new_n25589_, new_n25590_, new_n25591_,
    new_n25592_, new_n25593_, new_n25594_, new_n25595_, new_n25596_,
    new_n25597_, new_n25598_, new_n25599_, new_n25600_, new_n25601_,
    new_n25602_, new_n25603_, new_n25604_, new_n25605_, new_n25606_,
    new_n25607_, new_n25608_, new_n25609_, new_n25610_, new_n25611_,
    new_n25612_, new_n25613_, new_n25614_, new_n25615_, new_n25616_,
    new_n25617_, new_n25618_, new_n25619_, new_n25621_, new_n25622_,
    new_n25623_, new_n25624_, new_n25625_, new_n25626_, new_n25627_,
    new_n25628_, new_n25629_, new_n25630_, new_n25631_, new_n25632_,
    new_n25633_, new_n25634_, new_n25635_, new_n25636_, new_n25637_,
    new_n25638_, new_n25639_, new_n25640_, new_n25641_, new_n25642_,
    new_n25643_, new_n25644_, new_n25645_, new_n25646_, new_n25647_,
    new_n25648_, new_n25649_, new_n25650_, new_n25651_, new_n25652_,
    new_n25653_, new_n25654_, new_n25655_, new_n25656_, new_n25657_,
    new_n25658_, new_n25659_, new_n25660_, new_n25661_, new_n25662_,
    new_n25663_, new_n25664_, new_n25665_, new_n25666_, new_n25667_,
    new_n25668_, new_n25669_, new_n25670_, new_n25671_, new_n25672_,
    new_n25673_, new_n25674_, new_n25675_, new_n25676_, new_n25677_,
    new_n25678_, new_n25679_, new_n25680_, new_n25681_, new_n25682_,
    new_n25683_, new_n25684_, new_n25685_, new_n25686_, new_n25687_,
    new_n25688_, new_n25689_, new_n25690_, new_n25691_, new_n25692_,
    new_n25693_, new_n25694_, new_n25695_, new_n25696_, new_n25698_,
    new_n25699_, new_n25700_, new_n25701_, new_n25702_, new_n25703_,
    new_n25704_, new_n25705_, new_n25706_, new_n25707_, new_n25708_,
    new_n25709_, new_n25710_, new_n25711_, new_n25712_, new_n25713_,
    new_n25714_, new_n25715_, new_n25716_, new_n25717_, new_n25718_,
    new_n25719_, new_n25720_, new_n25721_, new_n25722_, new_n25723_,
    new_n25724_, new_n25725_, new_n25726_, new_n25727_, new_n25728_,
    new_n25729_, new_n25730_, new_n25731_, new_n25732_, new_n25733_,
    new_n25734_, new_n25735_, new_n25736_, new_n25737_, new_n25738_,
    new_n25739_, new_n25740_, new_n25741_, new_n25742_, new_n25743_,
    new_n25744_, new_n25745_, new_n25746_, new_n25747_, new_n25748_,
    new_n25749_, new_n25750_, new_n25751_, new_n25752_, new_n25753_,
    new_n25754_, new_n25755_, new_n25756_, new_n25757_, new_n25758_,
    new_n25759_, new_n25760_, new_n25761_, new_n25762_, new_n25763_,
    new_n25764_, new_n25765_, new_n25766_, new_n25767_, new_n25768_,
    new_n25769_, new_n25770_, new_n25771_, new_n25772_, new_n25774_,
    new_n25775_, new_n25776_, new_n25777_, new_n25778_, new_n25779_,
    new_n25780_, new_n25781_, new_n25782_, new_n25783_, new_n25784_,
    new_n25785_, new_n25786_, new_n25787_, new_n25788_, new_n25789_,
    new_n25790_, new_n25791_, new_n25792_, new_n25793_, new_n25794_,
    new_n25795_, new_n25796_, new_n25797_, new_n25798_, new_n25799_,
    new_n25800_, new_n25801_, new_n25802_, new_n25803_, new_n25804_,
    new_n25805_, new_n25806_, new_n25807_, new_n25808_, new_n25809_,
    new_n25810_, new_n25811_, new_n25812_, new_n25813_, new_n25814_,
    new_n25815_, new_n25816_, new_n25817_, new_n25818_, new_n25819_,
    new_n25820_, new_n25821_, new_n25822_, new_n25823_, new_n25824_,
    new_n25825_, new_n25826_, new_n25827_, new_n25828_, new_n25829_,
    new_n25830_, new_n25831_, new_n25832_, new_n25833_, new_n25834_,
    new_n25835_, new_n25836_, new_n25837_, new_n25838_, new_n25839_,
    new_n25840_, new_n25841_, new_n25842_, new_n25843_, new_n25844_,
    new_n25845_, new_n25846_, new_n25847_, new_n25848_, new_n25849_,
    new_n25850_, new_n25851_, new_n25852_, new_n25854_, new_n25855_,
    new_n25856_, new_n25857_, new_n25858_, new_n25859_, new_n25860_,
    new_n25861_, new_n25862_, new_n25863_, new_n25864_, new_n25865_,
    new_n25866_, new_n25867_, new_n25868_, new_n25869_, new_n25870_,
    new_n25871_, new_n25872_, new_n25873_, new_n25874_, new_n25875_,
    new_n25876_, new_n25877_, new_n25878_, new_n25879_, new_n25880_,
    new_n25881_, new_n25882_, new_n25883_, new_n25884_, new_n25885_,
    new_n25886_, new_n25887_, new_n25888_, new_n25889_, new_n25890_,
    new_n25891_, new_n25892_, new_n25893_, new_n25894_, new_n25895_,
    new_n25896_, new_n25897_, new_n25898_, new_n25899_, new_n25900_,
    new_n25901_, new_n25902_, new_n25903_, new_n25904_, new_n25905_,
    new_n25906_, new_n25907_, new_n25908_, new_n25909_, new_n25910_,
    new_n25911_, new_n25912_, new_n25913_, new_n25914_, new_n25915_,
    new_n25916_, new_n25917_, new_n25918_, new_n25919_, new_n25920_,
    new_n25921_, new_n25922_, new_n25923_, new_n25924_, new_n25925_,
    new_n25926_, new_n25927_, new_n25928_, new_n25930_, new_n25931_,
    new_n25932_, new_n25933_, new_n25934_, new_n25935_, new_n25936_,
    new_n25937_, new_n25938_, new_n25939_, new_n25940_, new_n25941_,
    new_n25942_, new_n25943_, new_n25944_, new_n25945_, new_n25946_,
    new_n25947_, new_n25948_, new_n25949_, new_n25950_, new_n25951_,
    new_n25952_, new_n25953_, new_n25954_, new_n25955_, new_n25956_,
    new_n25957_, new_n25958_, new_n25959_, new_n25960_, new_n25961_,
    new_n25962_, new_n25963_, new_n25964_, new_n25965_, new_n25966_,
    new_n25967_, new_n25968_, new_n25969_, new_n25970_, new_n25971_,
    new_n25972_, new_n25973_, new_n25974_, new_n25975_, new_n25976_,
    new_n25977_, new_n25978_, new_n25979_, new_n25980_, new_n25981_,
    new_n25982_, new_n25983_, new_n25984_, new_n25985_, new_n25986_,
    new_n25987_, new_n25988_, new_n25989_, new_n25990_, new_n25991_,
    new_n25992_, new_n25993_, new_n25994_, new_n25995_, new_n25996_,
    new_n25997_, new_n25998_, new_n25999_, new_n26000_, new_n26001_,
    new_n26002_, new_n26003_, new_n26004_, new_n26005_, new_n26006_,
    new_n26007_, new_n26008_, new_n26009_, new_n26011_, new_n26012_,
    new_n26013_, new_n26014_, new_n26015_, new_n26016_, new_n26017_,
    new_n26018_, new_n26019_, new_n26020_, new_n26021_, new_n26022_,
    new_n26023_, new_n26024_, new_n26025_, new_n26026_, new_n26027_,
    new_n26028_, new_n26029_, new_n26030_, new_n26031_, new_n26032_,
    new_n26033_, new_n26034_, new_n26035_, new_n26036_, new_n26037_,
    new_n26038_, new_n26039_, new_n26040_, new_n26041_, new_n26042_,
    new_n26043_, new_n26044_, new_n26045_, new_n26046_, new_n26047_,
    new_n26048_, new_n26049_, new_n26050_, new_n26051_, new_n26052_,
    new_n26053_, new_n26054_, new_n26055_, new_n26056_, new_n26057_,
    new_n26058_, new_n26059_, new_n26060_, new_n26061_, new_n26062_,
    new_n26063_, new_n26064_, new_n26065_, new_n26066_, new_n26067_,
    new_n26068_, new_n26069_, new_n26070_, new_n26071_, new_n26072_,
    new_n26073_, new_n26074_, new_n26075_, new_n26076_, new_n26077_,
    new_n26078_, new_n26079_, new_n26080_, new_n26081_, new_n26082_,
    new_n26083_, new_n26084_, new_n26085_, new_n26087_, new_n26088_,
    new_n26089_, new_n26090_, new_n26091_, new_n26092_, new_n26093_,
    new_n26094_, new_n26095_, new_n26096_, new_n26097_, new_n26098_,
    new_n26099_, new_n26100_, new_n26101_, new_n26102_, new_n26103_,
    new_n26104_, new_n26105_, new_n26106_, new_n26107_, new_n26108_,
    new_n26109_, new_n26110_, new_n26111_, new_n26112_, new_n26113_,
    new_n26114_, new_n26115_, new_n26116_, new_n26117_, new_n26118_,
    new_n26119_, new_n26120_, new_n26121_, new_n26122_, new_n26123_,
    new_n26124_, new_n26125_, new_n26126_, new_n26127_, new_n26128_,
    new_n26129_, new_n26130_, new_n26131_, new_n26132_, new_n26133_,
    new_n26134_, new_n26135_, new_n26136_, new_n26137_, new_n26138_,
    new_n26139_, new_n26140_, new_n26141_, new_n26142_, new_n26143_,
    new_n26144_, new_n26145_, new_n26146_, new_n26147_, new_n26148_,
    new_n26149_, new_n26150_, new_n26151_, new_n26152_, new_n26153_,
    new_n26154_, new_n26155_, new_n26156_, new_n26157_, new_n26158_,
    new_n26159_, new_n26160_, new_n26161_, new_n26162_, new_n26163_,
    new_n26164_, new_n26165_, new_n26167_, new_n26168_, new_n26169_,
    new_n26170_, new_n26171_, new_n26172_, new_n26173_, new_n26174_,
    new_n26175_, new_n26176_, new_n26177_, new_n26178_, new_n26179_,
    new_n26180_, new_n26181_, new_n26182_, new_n26183_, new_n26184_,
    new_n26185_, new_n26186_, new_n26187_, new_n26188_, new_n26189_,
    new_n26190_, new_n26191_, new_n26192_, new_n26193_, new_n26194_,
    new_n26195_, new_n26196_, new_n26197_, new_n26198_, new_n26199_,
    new_n26200_, new_n26201_, new_n26202_, new_n26203_, new_n26204_,
    new_n26205_, new_n26206_, new_n26207_, new_n26208_, new_n26209_,
    new_n26210_, new_n26211_, new_n26212_, new_n26213_, new_n26214_,
    new_n26215_, new_n26216_, new_n26217_, new_n26218_, new_n26219_,
    new_n26220_, new_n26221_, new_n26222_, new_n26223_, new_n26224_,
    new_n26225_, new_n26226_, new_n26227_, new_n26228_, new_n26229_,
    new_n26230_, new_n26231_, new_n26232_, new_n26233_, new_n26234_,
    new_n26235_, new_n26236_, new_n26237_, new_n26238_, new_n26239_,
    new_n26240_, new_n26241_, new_n26243_, new_n26244_, new_n26245_,
    new_n26246_, new_n26247_, new_n26248_, new_n26249_, new_n26250_,
    new_n26251_, new_n26252_, new_n26253_, new_n26254_, new_n26255_,
    new_n26256_, new_n26257_, new_n26258_, new_n26259_, new_n26260_,
    new_n26261_, new_n26262_, new_n26263_, new_n26264_, new_n26265_,
    new_n26266_, new_n26267_, new_n26268_, new_n26269_, new_n26270_,
    new_n26271_, new_n26272_, new_n26273_, new_n26274_, new_n26275_,
    new_n26276_, new_n26277_, new_n26278_, new_n26279_, new_n26280_,
    new_n26281_, new_n26282_, new_n26283_, new_n26284_, new_n26285_,
    new_n26286_, new_n26287_, new_n26288_, new_n26289_, new_n26290_,
    new_n26291_, new_n26292_, new_n26293_, new_n26294_, new_n26295_,
    new_n26296_, new_n26297_, new_n26298_, new_n26299_, new_n26300_,
    new_n26301_, new_n26302_, new_n26303_, new_n26304_, new_n26305_,
    new_n26306_, new_n26307_, new_n26308_, new_n26309_, new_n26310_,
    new_n26311_, new_n26312_, new_n26313_, new_n26314_, new_n26315_,
    new_n26316_, new_n26317_, new_n26318_, new_n26319_, new_n26320_,
    new_n26321_, new_n26322_, new_n26323_, new_n26324_, new_n26325_,
    new_n26327_, new_n26328_, new_n26329_, new_n26330_, new_n26331_,
    new_n26332_, new_n26333_, new_n26334_, new_n26335_, new_n26336_,
    new_n26337_, new_n26338_, new_n26339_, new_n26340_, new_n26341_,
    new_n26342_, new_n26343_, new_n26344_, new_n26345_, new_n26346_,
    new_n26347_, new_n26348_, new_n26349_, new_n26350_, new_n26351_,
    new_n26352_, new_n26353_, new_n26354_, new_n26355_, new_n26356_,
    new_n26357_, new_n26358_, new_n26359_, new_n26360_, new_n26361_,
    new_n26362_, new_n26363_, new_n26364_, new_n26365_, new_n26366_,
    new_n26367_, new_n26368_, new_n26369_, new_n26370_, new_n26371_,
    new_n26372_, new_n26373_, new_n26374_, new_n26375_, new_n26376_,
    new_n26377_, new_n26378_, new_n26379_, new_n26380_, new_n26381_,
    new_n26382_, new_n26383_, new_n26384_, new_n26385_, new_n26386_,
    new_n26387_, new_n26388_, new_n26389_, new_n26390_, new_n26391_,
    new_n26392_, new_n26393_, new_n26394_, new_n26395_, new_n26396_,
    new_n26397_, new_n26398_, new_n26399_, new_n26400_, new_n26401_,
    new_n26403_, new_n26404_, new_n26405_, new_n26406_, new_n26407_,
    new_n26408_, new_n26409_, new_n26410_, new_n26411_, new_n26412_,
    new_n26413_, new_n26414_, new_n26415_, new_n26416_, new_n26417_,
    new_n26418_, new_n26419_, new_n26420_, new_n26421_, new_n26422_,
    new_n26423_, new_n26424_, new_n26425_, new_n26426_, new_n26427_,
    new_n26428_, new_n26429_, new_n26430_, new_n26431_, new_n26432_,
    new_n26433_, new_n26434_, new_n26435_, new_n26436_, new_n26437_,
    new_n26438_, new_n26439_, new_n26440_, new_n26441_, new_n26442_,
    new_n26443_, new_n26444_, new_n26445_, new_n26446_, new_n26447_,
    new_n26448_, new_n26449_, new_n26450_, new_n26451_, new_n26452_,
    new_n26453_, new_n26454_, new_n26455_, new_n26456_, new_n26457_,
    new_n26458_, new_n26459_, new_n26460_, new_n26461_, new_n26462_,
    new_n26463_, new_n26464_, new_n26465_, new_n26466_, new_n26467_,
    new_n26468_, new_n26469_, new_n26470_, new_n26471_, new_n26472_,
    new_n26473_, new_n26474_, new_n26475_, new_n26476_, new_n26477_,
    new_n26478_, new_n26479_, new_n26480_, new_n26481_, new_n26483_,
    new_n26484_, new_n26485_, new_n26486_, new_n26487_, new_n26488_,
    new_n26489_, new_n26490_, new_n26491_, new_n26492_, new_n26493_,
    new_n26494_, new_n26495_, new_n26496_, new_n26497_, new_n26498_,
    new_n26499_, new_n26500_, new_n26501_, new_n26502_, new_n26503_,
    new_n26504_, new_n26505_, new_n26506_, new_n26507_, new_n26508_,
    new_n26509_, new_n26510_, new_n26511_, new_n26512_, new_n26513_,
    new_n26514_, new_n26515_, new_n26516_, new_n26517_, new_n26518_,
    new_n26519_, new_n26520_, new_n26521_, new_n26522_, new_n26523_,
    new_n26524_, new_n26525_, new_n26526_, new_n26527_, new_n26528_,
    new_n26529_, new_n26530_, new_n26531_, new_n26532_, new_n26533_,
    new_n26534_, new_n26535_, new_n26536_, new_n26537_, new_n26538_,
    new_n26539_, new_n26540_, new_n26541_, new_n26542_, new_n26543_,
    new_n26544_, new_n26545_, new_n26546_, new_n26547_, new_n26548_,
    new_n26549_, new_n26550_, new_n26551_, new_n26552_, new_n26553_,
    new_n26554_, new_n26555_, new_n26557_, new_n26558_, new_n26559_,
    new_n26560_, new_n26561_, new_n26562_, new_n26563_, new_n26564_,
    new_n26565_, new_n26566_, new_n26567_, new_n26568_, new_n26569_,
    new_n26570_, new_n26571_, new_n26572_, new_n26573_, new_n26574_,
    new_n26575_, new_n26576_, new_n26577_, new_n26578_, new_n26579_,
    new_n26580_, new_n26581_, new_n26582_, new_n26583_, new_n26584_,
    new_n26585_, new_n26586_, new_n26587_, new_n26588_, new_n26589_,
    new_n26590_, new_n26591_, new_n26592_, new_n26593_, new_n26594_,
    new_n26595_, new_n26596_, new_n26597_, new_n26598_, new_n26599_,
    new_n26600_, new_n26601_, new_n26602_, new_n26603_, new_n26604_,
    new_n26605_, new_n26606_, new_n26607_, new_n26608_, new_n26609_,
    new_n26610_, new_n26611_, new_n26612_, new_n26613_, new_n26614_,
    new_n26615_, new_n26616_, new_n26617_, new_n26618_, new_n26619_,
    new_n26620_, new_n26621_, new_n26622_, new_n26623_, new_n26624_,
    new_n26625_, new_n26626_, new_n26627_, new_n26628_, new_n26629_,
    new_n26630_, new_n26631_, new_n26632_, new_n26633_, new_n26634_,
    new_n26635_, new_n26636_, new_n26637_, new_n26638_, new_n26639_,
    new_n26640_, new_n26641_, new_n26642_, new_n26643_, new_n26644_,
    new_n26645_, new_n26646_, new_n26648_, new_n26649_, new_n26650_,
    new_n26651_, new_n26652_, new_n26653_, new_n26654_, new_n26655_,
    new_n26656_, new_n26657_, new_n26658_, new_n26659_, new_n26660_,
    new_n26661_, new_n26662_, new_n26663_, new_n26664_, new_n26665_,
    new_n26666_, new_n26667_, new_n26668_, new_n26669_, new_n26670_,
    new_n26671_, new_n26673_, new_n26674_, new_n26675_, new_n26676_,
    new_n26677_, new_n26678_, new_n26679_, new_n26680_, new_n26681_,
    new_n26682_, new_n26683_, new_n26684_, new_n26685_, new_n26686_,
    new_n26687_, new_n26688_, new_n26689_, new_n26690_, new_n26691_,
    new_n26692_, new_n26693_, new_n26694_, new_n26695_, new_n26696_,
    new_n26697_, new_n26698_, new_n26700_, new_n26701_, new_n26702_,
    new_n26703_, new_n26704_, new_n26705_, new_n26706_, new_n26707_,
    new_n26708_, new_n26709_, new_n26710_, new_n26711_, new_n26712_,
    new_n26713_, new_n26714_, new_n26715_, new_n26716_, new_n26717_,
    new_n26718_, new_n26719_, new_n26720_, new_n26721_, new_n26722_,
    new_n26723_, new_n26724_, new_n26725_, new_n26727_, new_n26728_,
    new_n26729_, new_n26730_, new_n26731_, new_n26732_, new_n26733_,
    new_n26734_, new_n26735_, new_n26736_, new_n26737_, new_n26738_,
    new_n26739_, new_n26740_, new_n26741_, new_n26742_, new_n26743_,
    new_n26744_, new_n26745_, new_n26746_, new_n26747_, new_n26748_,
    new_n26749_, new_n26750_, new_n26751_, new_n26752_, new_n26753_,
    new_n26754_, new_n26755_, new_n26757_, new_n26758_, new_n26759_,
    new_n26760_, new_n26761_, new_n26762_, new_n26763_, new_n26764_,
    new_n26765_, new_n26766_, new_n26767_, new_n26768_, new_n26769_,
    new_n26770_, new_n26771_, new_n26772_, new_n26773_, new_n26774_,
    new_n26775_, new_n26776_, new_n26777_, new_n26778_, new_n26779_,
    new_n26780_, new_n26781_, new_n26782_, new_n26784_, new_n26785_,
    new_n26786_, new_n26787_, new_n26788_, new_n26789_, new_n26790_,
    new_n26791_, new_n26792_, new_n26793_, new_n26794_, new_n26795_,
    new_n26796_, new_n26797_, new_n26798_, new_n26799_, new_n26800_,
    new_n26801_, new_n26802_, new_n26803_, new_n26804_, new_n26805_,
    new_n26806_, new_n26807_, new_n26808_, new_n26809_, new_n26810_,
    new_n26811_, new_n26812_, new_n26814_, new_n26815_, new_n26816_,
    new_n26817_, new_n26818_, new_n26819_, new_n26820_, new_n26821_,
    new_n26822_, new_n26823_, new_n26824_, new_n26825_, new_n26826_,
    new_n26827_, new_n26828_, new_n26829_, new_n26830_, new_n26831_,
    new_n26832_, new_n26833_, new_n26834_, new_n26835_, new_n26836_,
    new_n26837_, new_n26838_, new_n26839_, new_n26841_, new_n26842_,
    new_n26843_, new_n26844_, new_n26845_, new_n26846_, new_n26847_,
    new_n26848_, new_n26849_, new_n26850_, new_n26851_, new_n26852_,
    new_n26853_, new_n26854_, new_n26855_, new_n26856_, new_n26857_,
    new_n26858_, new_n26859_, new_n26860_, new_n26861_, new_n26862_,
    new_n26863_, new_n26864_, new_n26865_, new_n26866_, new_n26867_,
    new_n26868_, new_n26869_, new_n26870_, new_n26871_, new_n26872_,
    new_n26874_, new_n26875_, new_n26876_, new_n26877_, new_n26878_,
    new_n26879_, new_n26880_, new_n26881_, new_n26882_, new_n26883_,
    new_n26884_, new_n26885_, new_n26886_, new_n26887_, new_n26888_,
    new_n26889_, new_n26890_, new_n26891_, new_n26892_, new_n26893_,
    new_n26894_, new_n26895_, new_n26896_, new_n26897_, new_n26898_,
    new_n26899_, new_n26901_, new_n26902_, new_n26903_, new_n26904_,
    new_n26905_, new_n26906_, new_n26907_, new_n26908_, new_n26909_,
    new_n26910_, new_n26911_, new_n26912_, new_n26913_, new_n26914_,
    new_n26915_, new_n26916_, new_n26917_, new_n26918_, new_n26919_,
    new_n26920_, new_n26921_, new_n26922_, new_n26923_, new_n26924_,
    new_n26925_, new_n26926_, new_n26927_, new_n26928_, new_n26929_,
    new_n26931_, new_n26932_, new_n26933_, new_n26934_, new_n26935_,
    new_n26936_, new_n26937_, new_n26938_, new_n26939_, new_n26940_,
    new_n26941_, new_n26942_, new_n26943_, new_n26944_, new_n26945_,
    new_n26946_, new_n26947_, new_n26948_, new_n26949_, new_n26950_,
    new_n26951_, new_n26952_, new_n26953_, new_n26954_, new_n26955_,
    new_n26956_, new_n26958_, new_n26959_, new_n26960_, new_n26961_,
    new_n26962_, new_n26963_, new_n26964_, new_n26965_, new_n26966_,
    new_n26967_, new_n26968_, new_n26969_, new_n26970_, new_n26971_,
    new_n26972_, new_n26973_, new_n26974_, new_n26975_, new_n26976_,
    new_n26977_, new_n26978_, new_n26979_, new_n26980_, new_n26981_,
    new_n26982_, new_n26983_, new_n26984_, new_n26985_, new_n26986_,
    new_n26987_, new_n26988_, new_n26989_, new_n26991_, new_n26992_,
    new_n26993_, new_n26994_, new_n26995_, new_n26996_, new_n26997_,
    new_n26998_, new_n26999_, new_n27000_, new_n27001_, new_n27002_,
    new_n27003_, new_n27004_, new_n27005_, new_n27006_, new_n27007_,
    new_n27008_, new_n27009_, new_n27010_, new_n27011_, new_n27012_,
    new_n27013_, new_n27014_, new_n27015_, new_n27016_, new_n27018_,
    new_n27019_, new_n27020_, new_n27021_, new_n27022_, new_n27023_,
    new_n27024_, new_n27025_, new_n27026_, new_n27027_, new_n27028_,
    new_n27029_, new_n27030_, new_n27031_, new_n27032_, new_n27033_,
    new_n27034_, new_n27035_, new_n27036_, new_n27037_, new_n27038_,
    new_n27039_, new_n27040_, new_n27041_, new_n27042_, new_n27043_,
    new_n27044_, new_n27045_, new_n27046_, new_n27048_, new_n27049_,
    new_n27050_, new_n27051_, new_n27052_, new_n27053_, new_n27054_,
    new_n27055_, new_n27056_, new_n27057_, new_n27058_, new_n27059_,
    new_n27060_, new_n27061_, new_n27062_, new_n27063_, new_n27064_,
    new_n27065_, new_n27066_, new_n27067_, new_n27068_, new_n27069_,
    new_n27070_, new_n27071_, new_n27072_, new_n27073_, new_n27075_,
    new_n27076_, new_n27077_, new_n27078_, new_n27079_, new_n27080_,
    new_n27081_, new_n27082_, new_n27083_, new_n27084_, new_n27085_,
    new_n27086_, new_n27087_, new_n27088_, new_n27089_, new_n27090_,
    new_n27091_, new_n27092_, new_n27093_, new_n27094_, new_n27095_,
    new_n27096_, new_n27097_, new_n27098_, new_n27100_, new_n27101_,
    new_n27102_, new_n27103_, new_n27104_, new_n27105_, new_n27106_,
    new_n27107_, new_n27108_, new_n27110_, new_n27111_, new_n27112_,
    new_n27114_, new_n27115_, new_n27116_, new_n27117_, new_n27118_,
    new_n27119_, new_n27120_, new_n27121_, new_n27122_, new_n27124_,
    new_n27125_, new_n27126_, new_n27127_, new_n27128_, new_n27129_,
    new_n27130_, new_n27131_, new_n27132_, new_n27134_, new_n27135_,
    new_n27136_, new_n27137_, new_n27138_, new_n27139_, new_n27140_,
    new_n27141_, new_n27142_, new_n27144_, new_n27145_, new_n27146_,
    new_n27147_, new_n27148_, new_n27149_, new_n27150_, new_n27151_,
    new_n27152_, new_n27154_, new_n27155_, new_n27156_, new_n27157_,
    new_n27158_, new_n27159_, new_n27160_, new_n27161_, new_n27162_,
    new_n27164_, new_n27165_, new_n27166_, new_n27167_, new_n27168_,
    new_n27169_, new_n27170_, new_n27171_, new_n27172_, new_n27174_,
    new_n27175_, new_n27176_, new_n27177_, new_n27178_, new_n27179_,
    new_n27180_, new_n27181_, new_n27182_, new_n27184_, new_n27185_,
    new_n27186_, new_n27187_, new_n27188_, new_n27189_, new_n27190_,
    new_n27191_, new_n27192_, new_n27194_, new_n27195_, new_n27196_,
    new_n27197_, new_n27198_, new_n27199_, new_n27200_, new_n27201_,
    new_n27202_, new_n27204_, new_n27205_, new_n27206_, new_n27207_,
    new_n27208_, new_n27209_, new_n27210_, new_n27211_, new_n27212_,
    new_n27214_, new_n27215_, new_n27216_, new_n27217_, new_n27218_,
    new_n27219_, new_n27220_, new_n27221_, new_n27222_, new_n27224_,
    new_n27225_, new_n27226_, new_n27227_, new_n27228_, new_n27229_,
    new_n27230_, new_n27231_, new_n27232_, new_n27234_, new_n27235_,
    new_n27236_, new_n27237_, new_n27238_, new_n27239_, new_n27240_,
    new_n27241_, new_n27242_, new_n27244_, new_n27245_, new_n27246_,
    new_n27247_, new_n27248_, new_n27249_, new_n27250_, new_n27251_,
    new_n27252_, new_n27254_, new_n27255_, new_n27256_, new_n27257_,
    new_n27258_, new_n27259_, new_n27260_, new_n27261_, new_n27262_,
    new_n27264_, new_n27265_, new_n27266_, new_n27267_, new_n27268_,
    new_n27269_, new_n27270_, new_n27271_, new_n27272_, new_n27274_,
    new_n27275_, new_n27276_, new_n27278_, new_n27279_, new_n27280_,
    new_n27281_, new_n27282_, new_n27283_, new_n27284_, new_n27285_,
    new_n27286_, new_n27288_, new_n27289_, new_n27291_, new_n27292_,
    new_n27294_, new_n27295_, new_n27297_, new_n27298_, new_n27300_,
    new_n27301_, new_n27302_, new_n27303_, new_n27304_, new_n27305_,
    new_n27306_, new_n27307_, new_n27308_, new_n27309_, new_n27311_,
    new_n27312_, new_n27313_, new_n27314_, new_n27315_, new_n27316_,
    new_n27317_, new_n27318_, new_n27319_, new_n27320_, new_n27322_,
    new_n27323_, new_n27324_, new_n27325_, new_n27326_, new_n27327_,
    new_n27328_, new_n27329_, new_n27330_, new_n27331_, new_n27333_,
    new_n27334_, new_n27335_, new_n27336_, new_n27337_, new_n27338_,
    new_n27339_, new_n27340_, new_n27341_, new_n27342_, new_n27343_,
    new_n27345_, new_n27346_, new_n27347_, new_n27348_, new_n27350_,
    new_n27351_, new_n27352_, new_n27353_, new_n27354_, new_n27356_,
    new_n27357_, new_n27359_, new_n27360_, new_n27361_, new_n27362_,
    new_n27363_, new_n27364_, new_n27365_, new_n27366_, new_n27367_,
    new_n27368_, new_n27369_, new_n27370_, new_n27371_, new_n27373_,
    new_n27374_, new_n27376_, new_n27377_, new_n27378_, new_n27379_,
    new_n27380_, new_n27381_, new_n27382_, new_n27383_, new_n27384_,
    new_n27386_, new_n27387_, new_n27388_, new_n27389_, new_n27390_,
    new_n27391_, new_n27392_, new_n27394_, new_n27395_, new_n27396_,
    new_n27397_, new_n27399_, new_n27405_, new_n27406_, new_n27407_,
    new_n27408_, new_n27409_, new_n27410_, new_n27411_, new_n27412_,
    new_n27414_, new_n27415_, new_n27416_, new_n27417_, new_n27419_,
    new_n27420_, new_n27421_, new_n27422_, new_n27423_, new_n27425_,
    new_n27426_, new_n27427_, new_n27428_, new_n27429_, new_n27430_,
    new_n27431_, new_n27432_, new_n27433_, new_n27434_, new_n27435_,
    new_n27436_, new_n27438_, new_n27440_, new_n27441_, new_n27442_,
    new_n27444_, new_n27445_, new_n27446_, new_n27447_, new_n27448_,
    new_n27449_, new_n27450_, new_n27451_, new_n27452_, new_n27453_,
    new_n27454_, new_n27455_, new_n27457_, new_n27458_, new_n27459_,
    new_n27460_, new_n27462_, new_n27463_, new_n27464_, new_n27465_,
    new_n27466_, new_n27467_, new_n27468_, new_n27469_, new_n27470_,
    new_n27471_, new_n27472_, new_n27473_, new_n27474_, new_n27476_,
    new_n27477_, new_n27478_, new_n27479_, new_n27480_, new_n27481_,
    new_n27482_, new_n27483_, new_n27484_, new_n27486_, new_n27487_,
    new_n27488_, new_n27489_, new_n27490_, new_n27491_, new_n27492_,
    new_n27493_, new_n27494_, new_n27495_, new_n27497_, new_n27498_,
    new_n27499_, new_n27500_, new_n27501_, new_n27502_, new_n27503_,
    new_n27504_, new_n27505_, new_n27506_, new_n27508_, new_n27509_,
    new_n27510_, new_n27511_, new_n27512_, new_n27513_, new_n27514_,
    new_n27515_, new_n27516_, new_n27518_, new_n27519_, new_n27520_,
    new_n27521_, new_n27522_, new_n27523_, new_n27524_, new_n27525_,
    new_n27526_, new_n27528_, new_n27529_, new_n27530_, new_n27531_,
    new_n27532_, new_n27533_, new_n27534_, new_n27535_, new_n27536_,
    new_n27538_, new_n27539_, new_n27540_, new_n27541_, new_n27542_,
    new_n27543_, new_n27544_, new_n27545_, new_n27546_, new_n27548_,
    new_n27549_, new_n27550_, new_n27551_, new_n27552_, new_n27553_,
    new_n27554_, new_n27555_, new_n27556_, new_n27558_, new_n27559_,
    new_n27560_, new_n27561_, new_n27562_, new_n27563_, new_n27564_,
    new_n27565_, new_n27566_, new_n27568_, new_n27569_, new_n27570_,
    new_n27571_, new_n27572_, new_n27573_, new_n27574_, new_n27575_,
    new_n27576_, new_n27578_, new_n27579_, new_n27580_, new_n27581_,
    new_n27582_, new_n27583_, new_n27584_, new_n27585_, new_n27586_,
    new_n27588_, new_n27589_, new_n27590_, new_n27591_, new_n27592_,
    new_n27593_, new_n27594_, new_n27595_, new_n27596_, new_n27598_,
    new_n27599_, new_n27600_, new_n27601_, new_n27602_, new_n27603_,
    new_n27604_, new_n27605_, new_n27606_, new_n27608_, new_n27609_,
    new_n27610_, new_n27611_, new_n27612_, new_n27613_, new_n27614_,
    new_n27615_, new_n27616_, new_n27618_, new_n27619_, new_n27620_,
    new_n27621_, new_n27622_, new_n27623_, new_n27624_, new_n27625_,
    new_n27626_, new_n27628_, new_n27629_, new_n27630_, new_n27631_,
    new_n27632_, new_n27633_, new_n27634_, new_n27635_, new_n27636_,
    new_n27638_, new_n27639_, new_n27640_, new_n27641_, new_n27642_,
    new_n27643_, new_n27644_, new_n27645_, new_n27646_, new_n27648_,
    new_n27649_, new_n27650_, new_n27651_, new_n27652_, new_n27653_,
    new_n27654_, new_n27655_, new_n27656_, new_n27658_, new_n27659_,
    new_n27660_, new_n27661_, new_n27662_, new_n27663_, new_n27664_,
    new_n27665_, new_n27666_, new_n27667_, new_n27669_, new_n27670_,
    new_n27671_, new_n27672_, new_n27673_, new_n27674_, new_n27675_,
    new_n27676_, new_n27677_, new_n27678_, new_n27680_, new_n27681_,
    new_n27682_, new_n27683_, new_n27684_, new_n27685_, new_n27686_,
    new_n27687_, new_n27688_, new_n27690_, new_n27691_, new_n27692_,
    new_n27693_, new_n27694_, new_n27695_, new_n27696_, new_n27697_,
    new_n27698_, new_n27700_, new_n27701_, new_n27702_, new_n27703_,
    new_n27704_, new_n27705_, new_n27706_, new_n27707_, new_n27708_,
    new_n27710_, new_n27711_, new_n27712_, new_n27713_, new_n27714_,
    new_n27715_, new_n27716_, new_n27717_, new_n27718_, new_n27720_,
    new_n27721_, new_n27722_, new_n27723_, new_n27724_, new_n27725_,
    new_n27726_, new_n27727_, new_n27728_, new_n27730_, new_n27731_,
    new_n27732_, new_n27733_, new_n27734_, new_n27735_, new_n27736_,
    new_n27737_, new_n27738_, new_n27739_, new_n27741_, new_n27742_,
    new_n27743_, new_n27744_, new_n27745_, new_n27746_, new_n27747_,
    new_n27748_, new_n27749_, new_n27751_, new_n27752_, new_n27753_,
    new_n27754_, new_n27755_, new_n27756_, new_n27757_, new_n27758_,
    new_n27759_, new_n27761_, new_n27762_, new_n27763_, new_n27764_,
    new_n27765_, new_n27766_, new_n27767_, new_n27768_, new_n27769_,
    new_n27770_, new_n27772_, new_n27773_, new_n27774_, new_n27775_,
    new_n27776_, new_n27777_, new_n27778_, new_n27779_, new_n27780_,
    new_n27782_, new_n27783_, new_n27784_, new_n27785_, new_n27786_,
    new_n27787_, new_n27788_, new_n27789_, new_n27790_, new_n27792_,
    new_n27793_, new_n27794_, new_n27795_, new_n27796_, new_n27797_,
    new_n27798_, new_n27799_, new_n27800_, new_n27801_, new_n27802_,
    new_n27803_, new_n27804_, new_n27805_, new_n27806_, new_n27807_,
    new_n27808_, new_n27809_, new_n27810_, new_n27811_, new_n27812_,
    new_n27813_, new_n27814_, new_n27815_, new_n27816_, new_n27817_,
    new_n27818_, new_n27819_, new_n27820_, new_n27821_, new_n27822_,
    new_n27823_, new_n27824_, new_n27825_, new_n27826_, new_n27827_,
    new_n27828_, new_n27830_, new_n27831_, new_n27832_, new_n27833_,
    new_n27834_, new_n27835_, new_n27836_, new_n27837_, new_n27838_,
    new_n27839_, new_n27840_, new_n27841_, new_n27843_, new_n27844_,
    new_n27845_, new_n27846_, new_n27847_, new_n27848_, new_n27850_,
    new_n27851_, new_n27852_, new_n27853_, new_n27854_, new_n27855_,
    new_n27857_, new_n27858_, new_n27859_, new_n27860_, new_n27861_,
    new_n27862_, new_n27868_, new_n27869_, new_n27870_, new_n27871_,
    new_n27872_, new_n27873_, new_n27874_, new_n27875_, new_n27876_,
    new_n27877_, new_n27879_, new_n27880_, new_n27881_, new_n27882_,
    new_n27883_, new_n27885_, new_n27886_, new_n27887_, new_n27888_,
    new_n27889_, new_n27891_, new_n27892_, new_n27893_, new_n27894_,
    new_n27895_, new_n27897_, new_n27898_, new_n27899_, new_n27900_,
    new_n27901_, new_n27902_, new_n27903_, new_n27904_, new_n27905_,
    new_n27906_, new_n27907_, new_n27908_, new_n27909_, new_n27910_,
    new_n27911_, new_n27912_, new_n27913_, new_n27914_, new_n27915_,
    new_n27916_, new_n27917_, new_n27918_, new_n27919_, new_n27920_,
    new_n27921_, new_n27922_, new_n27923_, new_n27924_, new_n27925_,
    new_n27926_, new_n27927_, new_n27928_, new_n27929_, new_n27930_,
    new_n27931_, new_n27932_, new_n27933_, new_n27934_, new_n27935_,
    new_n27936_, new_n27937_, new_n27938_, new_n27939_, new_n27940_,
    new_n27941_, new_n27942_, new_n27943_, new_n27944_, new_n27945_,
    new_n27946_, new_n27947_, new_n27948_, new_n27949_, new_n27950_,
    new_n27951_, new_n27952_, new_n27953_, new_n27954_, new_n27955_,
    new_n27956_, new_n27957_, new_n27958_, new_n27959_, new_n27960_,
    new_n27961_, new_n27962_, new_n27963_, new_n27964_, new_n27965_,
    new_n27966_, new_n27967_, new_n27968_, new_n27969_, new_n27970_,
    new_n27971_, new_n27972_, new_n27973_, new_n27974_, new_n27975_,
    new_n27976_, new_n27977_, new_n27978_, new_n27979_, new_n27980_,
    new_n27981_, new_n27982_, new_n27983_, new_n27984_, new_n27985_,
    new_n27986_, new_n27987_, new_n27988_, new_n27989_, new_n27990_,
    new_n27991_, new_n27992_, new_n27993_, new_n27994_, new_n27995_,
    new_n27996_, new_n27997_, new_n27998_, new_n27999_, new_n28000_,
    new_n28001_, new_n28002_, new_n28003_, new_n28004_, new_n28005_,
    new_n28006_, new_n28007_, new_n28008_, new_n28009_, new_n28010_,
    new_n28011_, new_n28012_, new_n28013_, new_n28014_, new_n28015_,
    new_n28016_, new_n28017_, new_n28018_, new_n28020_, new_n28021_,
    new_n28022_, new_n28023_, new_n28024_, new_n28025_, new_n28026_,
    new_n28027_, new_n28028_, new_n28029_, new_n28030_, new_n28031_,
    new_n28032_, new_n28033_, new_n28034_, new_n28035_, new_n28036_,
    new_n28037_, new_n28038_, new_n28039_, new_n28040_, new_n28041_,
    new_n28042_, new_n28043_, new_n28044_, new_n28045_, new_n28046_,
    new_n28047_, new_n28048_, new_n28049_, new_n28050_, new_n28051_,
    new_n28052_, new_n28053_, new_n28054_, new_n28055_, new_n28056_,
    new_n28057_, new_n28058_, new_n28059_, new_n28060_, new_n28061_,
    new_n28062_, new_n28063_, new_n28064_, new_n28065_, new_n28066_,
    new_n28067_, new_n28068_, new_n28069_, new_n28070_, new_n28071_,
    new_n28072_, new_n28073_, new_n28074_, new_n28075_, new_n28076_,
    new_n28077_, new_n28078_, new_n28079_, new_n28080_, new_n28081_,
    new_n28082_, new_n28083_, new_n28084_, new_n28085_, new_n28086_,
    new_n28087_, new_n28088_, new_n28089_, new_n28090_, new_n28091_,
    new_n28092_, new_n28093_, new_n28094_, new_n28095_, new_n28096_,
    new_n28097_, new_n28098_, new_n28099_, new_n28100_, new_n28101_,
    new_n28102_, new_n28103_, new_n28104_, new_n28105_, new_n28106_,
    new_n28108_, new_n28109_, new_n28110_, new_n28111_, new_n28112_,
    new_n28113_, new_n28114_, new_n28115_, new_n28116_, new_n28117_,
    new_n28118_, new_n28119_, new_n28120_, new_n28121_, new_n28122_,
    new_n28123_, new_n28124_, new_n28125_, new_n28126_, new_n28127_,
    new_n28128_, new_n28129_, new_n28130_, new_n28131_, new_n28132_,
    new_n28133_, new_n28134_, new_n28135_, new_n28136_, new_n28137_,
    new_n28138_, new_n28139_, new_n28140_, new_n28141_, new_n28142_,
    new_n28143_, new_n28144_, new_n28145_, new_n28146_, new_n28147_,
    new_n28148_, new_n28149_, new_n28150_, new_n28151_, new_n28152_,
    new_n28153_, new_n28154_, new_n28155_, new_n28156_, new_n28157_,
    new_n28158_, new_n28159_, new_n28160_, new_n28161_, new_n28162_,
    new_n28163_, new_n28164_, new_n28165_, new_n28166_, new_n28167_,
    new_n28168_, new_n28169_, new_n28170_, new_n28171_, new_n28172_,
    new_n28173_, new_n28174_, new_n28175_, new_n28176_, new_n28177_,
    new_n28178_, new_n28179_, new_n28180_, new_n28181_, new_n28182_,
    new_n28183_, new_n28184_, new_n28185_, new_n28186_, new_n28187_,
    new_n28188_, new_n28189_, new_n28190_, new_n28191_, new_n28192_,
    new_n28193_, new_n28194_, new_n28196_, new_n28197_, new_n28198_,
    new_n28199_, new_n28200_, new_n28201_, new_n28202_, new_n28203_,
    new_n28204_, new_n28205_, new_n28206_, new_n28207_, new_n28208_,
    new_n28209_, new_n28210_, new_n28211_, new_n28212_, new_n28213_,
    new_n28214_, new_n28215_, new_n28216_, new_n28217_, new_n28218_,
    new_n28219_, new_n28220_, new_n28221_, new_n28222_, new_n28223_,
    new_n28224_, new_n28225_, new_n28226_, new_n28227_, new_n28228_,
    new_n28229_, new_n28230_, new_n28231_, new_n28232_, new_n28233_,
    new_n28234_, new_n28235_, new_n28236_, new_n28237_, new_n28238_,
    new_n28239_, new_n28240_, new_n28241_, new_n28242_, new_n28243_,
    new_n28244_, new_n28245_, new_n28246_, new_n28247_, new_n28248_,
    new_n28249_, new_n28250_, new_n28251_, new_n28252_, new_n28253_,
    new_n28254_, new_n28255_, new_n28256_, new_n28257_, new_n28258_,
    new_n28259_, new_n28260_, new_n28261_, new_n28262_, new_n28263_,
    new_n28264_, new_n28265_, new_n28266_, new_n28267_, new_n28268_,
    new_n28269_, new_n28270_, new_n28271_, new_n28272_, new_n28273_,
    new_n28274_, new_n28275_, new_n28276_, new_n28277_, new_n28278_,
    new_n28279_, new_n28280_, new_n28281_, new_n28282_, new_n28284_,
    new_n28285_, new_n28286_, new_n28287_, new_n28288_, new_n28289_,
    new_n28290_, new_n28291_, new_n28292_, new_n28293_, new_n28294_,
    new_n28295_, new_n28296_, new_n28297_, new_n28298_, new_n28299_,
    new_n28300_, new_n28301_, new_n28302_, new_n28303_, new_n28304_,
    new_n28305_, new_n28306_, new_n28307_, new_n28308_, new_n28309_,
    new_n28310_, new_n28311_, new_n28312_, new_n28313_, new_n28314_,
    new_n28315_, new_n28316_, new_n28317_, new_n28318_, new_n28319_,
    new_n28320_, new_n28321_, new_n28322_, new_n28323_, new_n28324_,
    new_n28325_, new_n28326_, new_n28327_, new_n28328_, new_n28329_,
    new_n28330_, new_n28331_, new_n28332_, new_n28333_, new_n28334_,
    new_n28335_, new_n28336_, new_n28337_, new_n28338_, new_n28339_,
    new_n28340_, new_n28341_, new_n28342_, new_n28343_, new_n28344_,
    new_n28345_, new_n28346_, new_n28347_, new_n28348_, new_n28349_,
    new_n28350_, new_n28351_, new_n28352_, new_n28353_, new_n28354_,
    new_n28355_, new_n28356_, new_n28357_, new_n28358_, new_n28359_,
    new_n28360_, new_n28361_, new_n28362_, new_n28363_, new_n28364_,
    new_n28365_, new_n28366_, new_n28367_, new_n28368_, new_n28369_,
    new_n28370_, new_n28372_, new_n28373_, new_n28374_, new_n28375_,
    new_n28376_, new_n28377_, new_n28378_, new_n28379_, new_n28380_,
    new_n28381_, new_n28382_, new_n28383_, new_n28384_, new_n28385_,
    new_n28386_, new_n28387_, new_n28388_, new_n28389_, new_n28390_,
    new_n28391_, new_n28392_, new_n28393_, new_n28394_, new_n28395_,
    new_n28396_, new_n28397_, new_n28398_, new_n28399_, new_n28400_,
    new_n28401_, new_n28402_, new_n28403_, new_n28404_, new_n28405_,
    new_n28406_, new_n28407_, new_n28408_, new_n28409_, new_n28410_,
    new_n28411_, new_n28412_, new_n28413_, new_n28414_, new_n28415_,
    new_n28416_, new_n28417_, new_n28418_, new_n28419_, new_n28420_,
    new_n28421_, new_n28422_, new_n28423_, new_n28424_, new_n28425_,
    new_n28426_, new_n28427_, new_n28428_, new_n28429_, new_n28430_,
    new_n28431_, new_n28432_, new_n28433_, new_n28434_, new_n28435_,
    new_n28436_, new_n28437_, new_n28438_, new_n28439_, new_n28440_,
    new_n28441_, new_n28442_, new_n28443_, new_n28444_, new_n28445_,
    new_n28446_, new_n28447_, new_n28448_, new_n28449_, new_n28450_,
    new_n28451_, new_n28452_, new_n28453_, new_n28454_, new_n28455_,
    new_n28456_, new_n28457_, new_n28458_, new_n28460_, new_n28461_,
    new_n28462_, new_n28463_, new_n28464_, new_n28465_, new_n28466_,
    new_n28467_, new_n28468_, new_n28469_, new_n28470_, new_n28471_,
    new_n28472_, new_n28473_, new_n28474_, new_n28475_, new_n28476_,
    new_n28477_, new_n28478_, new_n28479_, new_n28480_, new_n28481_,
    new_n28482_, new_n28483_, new_n28484_, new_n28485_, new_n28486_,
    new_n28487_, new_n28488_, new_n28489_, new_n28490_, new_n28491_,
    new_n28492_, new_n28493_, new_n28494_, new_n28495_, new_n28496_,
    new_n28497_, new_n28498_, new_n28499_, new_n28500_, new_n28501_,
    new_n28502_, new_n28503_, new_n28504_, new_n28505_, new_n28506_,
    new_n28507_, new_n28508_, new_n28509_, new_n28510_, new_n28511_,
    new_n28512_, new_n28513_, new_n28514_, new_n28515_, new_n28516_,
    new_n28517_, new_n28518_, new_n28519_, new_n28520_, new_n28521_,
    new_n28522_, new_n28523_, new_n28524_, new_n28525_, new_n28526_,
    new_n28527_, new_n28528_, new_n28529_, new_n28530_, new_n28531_,
    new_n28532_, new_n28533_, new_n28534_, new_n28535_, new_n28536_,
    new_n28537_, new_n28538_, new_n28539_, new_n28540_, new_n28541_,
    new_n28542_, new_n28543_, new_n28544_, new_n28545_, new_n28546_,
    new_n28548_, new_n28549_, new_n28550_, new_n28551_, new_n28552_,
    new_n28553_, new_n28554_, new_n28555_, new_n28556_, new_n28557_,
    new_n28558_, new_n28559_, new_n28560_, new_n28561_, new_n28562_,
    new_n28563_, new_n28564_, new_n28565_, new_n28566_, new_n28567_,
    new_n28568_, new_n28569_, new_n28570_, new_n28571_, new_n28572_,
    new_n28573_, new_n28574_, new_n28575_, new_n28576_, new_n28577_,
    new_n28578_, new_n28579_, new_n28580_, new_n28581_, new_n28582_,
    new_n28583_, new_n28584_, new_n28585_, new_n28586_, new_n28587_,
    new_n28588_, new_n28589_, new_n28590_, new_n28591_, new_n28592_,
    new_n28593_, new_n28594_, new_n28595_, new_n28596_, new_n28597_,
    new_n28598_, new_n28599_, new_n28600_, new_n28601_, new_n28602_,
    new_n28603_, new_n28604_, new_n28605_, new_n28606_, new_n28607_,
    new_n28608_, new_n28609_, new_n28610_, new_n28611_, new_n28612_,
    new_n28613_, new_n28614_, new_n28615_, new_n28616_, new_n28617_,
    new_n28618_, new_n28619_, new_n28620_, new_n28621_, new_n28622_,
    new_n28623_, new_n28624_, new_n28625_, new_n28626_, new_n28627_,
    new_n28628_, new_n28629_, new_n28630_, new_n28631_, new_n28632_,
    new_n28633_, new_n28634_, new_n28636_, new_n28637_, new_n28638_,
    new_n28639_, new_n28640_, new_n28641_, new_n28642_, new_n28643_,
    new_n28644_, new_n28645_, new_n28646_, new_n28647_, new_n28648_,
    new_n28649_, new_n28650_, new_n28651_, new_n28652_, new_n28653_,
    new_n28654_, new_n28655_, new_n28656_, new_n28657_, new_n28658_,
    new_n28659_, new_n28660_, new_n28661_, new_n28662_, new_n28663_,
    new_n28664_, new_n28665_, new_n28666_, new_n28667_, new_n28668_,
    new_n28669_, new_n28670_, new_n28671_, new_n28672_, new_n28673_,
    new_n28674_, new_n28675_, new_n28676_, new_n28677_, new_n28678_,
    new_n28679_, new_n28680_, new_n28681_, new_n28682_, new_n28683_,
    new_n28684_, new_n28685_, new_n28686_, new_n28687_, new_n28688_,
    new_n28689_, new_n28690_, new_n28691_, new_n28692_, new_n28693_,
    new_n28694_, new_n28695_, new_n28696_, new_n28697_, new_n28698_,
    new_n28699_, new_n28700_, new_n28701_, new_n28702_, new_n28703_,
    new_n28704_, new_n28705_, new_n28706_, new_n28707_, new_n28708_,
    new_n28709_, new_n28710_, new_n28711_, new_n28712_, new_n28713_,
    new_n28714_, new_n28715_, new_n28716_, new_n28717_, new_n28718_,
    new_n28719_, new_n28720_, new_n28721_, new_n28722_, new_n28724_,
    new_n28725_, new_n28726_, new_n28727_, new_n28728_, new_n28729_,
    new_n28730_, new_n28731_, new_n28732_, new_n28733_, new_n28734_,
    new_n28735_, new_n28736_, new_n28737_, new_n28738_, new_n28739_,
    new_n28740_, new_n28741_, new_n28742_, new_n28743_, new_n28744_,
    new_n28745_, new_n28746_, new_n28747_, new_n28748_, new_n28749_,
    new_n28750_, new_n28751_, new_n28752_, new_n28753_, new_n28754_,
    new_n28755_, new_n28756_, new_n28757_, new_n28758_, new_n28759_,
    new_n28760_, new_n28761_, new_n28762_, new_n28763_, new_n28764_,
    new_n28765_, new_n28766_, new_n28767_, new_n28768_, new_n28769_,
    new_n28770_, new_n28771_, new_n28772_, new_n28773_, new_n28774_,
    new_n28775_, new_n28776_, new_n28777_, new_n28778_, new_n28779_,
    new_n28780_, new_n28781_, new_n28782_, new_n28783_, new_n28784_,
    new_n28785_, new_n28786_, new_n28787_, new_n28788_, new_n28789_,
    new_n28790_, new_n28791_, new_n28792_, new_n28793_, new_n28794_,
    new_n28795_, new_n28796_, new_n28797_, new_n28798_, new_n28799_,
    new_n28800_, new_n28801_, new_n28802_, new_n28803_, new_n28804_,
    new_n28805_, new_n28806_, new_n28807_, new_n28808_, new_n28809_,
    new_n28810_, new_n28812_, new_n28813_, new_n28814_, new_n28815_,
    new_n28816_, new_n28817_, new_n28818_, new_n28819_, new_n28820_,
    new_n28821_, new_n28822_, new_n28823_, new_n28824_, new_n28825_,
    new_n28826_, new_n28827_, new_n28828_, new_n28829_, new_n28830_,
    new_n28831_, new_n28832_, new_n28833_, new_n28834_, new_n28835_,
    new_n28836_, new_n28837_, new_n28838_, new_n28839_, new_n28840_,
    new_n28841_, new_n28842_, new_n28843_, new_n28844_, new_n28845_,
    new_n28846_, new_n28847_, new_n28848_, new_n28849_, new_n28850_,
    new_n28851_, new_n28852_, new_n28853_, new_n28854_, new_n28855_,
    new_n28856_, new_n28857_, new_n28858_, new_n28859_, new_n28860_,
    new_n28861_, new_n28862_, new_n28863_, new_n28864_, new_n28865_,
    new_n28866_, new_n28867_, new_n28868_, new_n28869_, new_n28870_,
    new_n28871_, new_n28872_, new_n28873_, new_n28874_, new_n28875_,
    new_n28876_, new_n28877_, new_n28878_, new_n28879_, new_n28880_,
    new_n28881_, new_n28882_, new_n28883_, new_n28884_, new_n28885_,
    new_n28886_, new_n28887_, new_n28888_, new_n28889_, new_n28890_,
    new_n28891_, new_n28892_, new_n28893_, new_n28894_, new_n28895_,
    new_n28896_, new_n28897_, new_n28898_, new_n28900_, new_n28901_,
    new_n28902_, new_n28903_, new_n28904_, new_n28905_, new_n28906_,
    new_n28907_, new_n28908_, new_n28909_, new_n28910_, new_n28911_,
    new_n28912_, new_n28913_, new_n28914_, new_n28915_, new_n28916_,
    new_n28917_, new_n28918_, new_n28919_, new_n28920_, new_n28921_,
    new_n28922_, new_n28923_, new_n28924_, new_n28925_, new_n28926_,
    new_n28927_, new_n28928_, new_n28929_, new_n28930_, new_n28931_,
    new_n28932_, new_n28933_, new_n28934_, new_n28935_, new_n28936_,
    new_n28937_, new_n28938_, new_n28939_, new_n28940_, new_n28941_,
    new_n28942_, new_n28943_, new_n28944_, new_n28945_, new_n28946_,
    new_n28947_, new_n28948_, new_n28949_, new_n28950_, new_n28951_,
    new_n28952_, new_n28953_, new_n28954_, new_n28955_, new_n28956_,
    new_n28957_, new_n28958_, new_n28959_, new_n28960_, new_n28961_,
    new_n28962_, new_n28963_, new_n28964_, new_n28965_, new_n28966_,
    new_n28967_, new_n28968_, new_n28969_, new_n28970_, new_n28971_,
    new_n28972_, new_n28973_, new_n28974_, new_n28975_, new_n28976_,
    new_n28977_, new_n28978_, new_n28979_, new_n28980_, new_n28981_,
    new_n28982_, new_n28983_, new_n28984_, new_n28985_, new_n28986_,
    new_n28988_, new_n28989_, new_n28990_, new_n28991_, new_n28992_,
    new_n28993_, new_n28994_, new_n28995_, new_n28996_, new_n28997_,
    new_n28998_, new_n28999_, new_n29000_, new_n29001_, new_n29002_,
    new_n29003_, new_n29004_, new_n29005_, new_n29006_, new_n29007_,
    new_n29008_, new_n29009_, new_n29010_, new_n29011_, new_n29012_,
    new_n29013_, new_n29014_, new_n29015_, new_n29016_, new_n29017_,
    new_n29018_, new_n29019_, new_n29020_, new_n29021_, new_n29022_,
    new_n29023_, new_n29024_, new_n29025_, new_n29026_, new_n29027_,
    new_n29028_, new_n29029_, new_n29030_, new_n29031_, new_n29032_,
    new_n29033_, new_n29034_, new_n29035_, new_n29036_, new_n29037_,
    new_n29038_, new_n29039_, new_n29040_, new_n29041_, new_n29042_,
    new_n29043_, new_n29044_, new_n29045_, new_n29046_, new_n29047_,
    new_n29048_, new_n29049_, new_n29050_, new_n29051_, new_n29052_,
    new_n29053_, new_n29054_, new_n29055_, new_n29056_, new_n29057_,
    new_n29058_, new_n29059_, new_n29060_, new_n29061_, new_n29062_,
    new_n29063_, new_n29064_, new_n29065_, new_n29066_, new_n29067_,
    new_n29068_, new_n29069_, new_n29070_, new_n29071_, new_n29072_,
    new_n29073_, new_n29074_, new_n29076_, new_n29077_, new_n29078_,
    new_n29079_, new_n29080_, new_n29081_, new_n29082_, new_n29083_,
    new_n29084_, new_n29085_, new_n29086_, new_n29087_, new_n29088_,
    new_n29089_, new_n29090_, new_n29091_, new_n29092_, new_n29093_,
    new_n29094_, new_n29095_, new_n29096_, new_n29097_, new_n29098_,
    new_n29099_, new_n29100_, new_n29101_, new_n29102_, new_n29103_,
    new_n29104_, new_n29105_, new_n29106_, new_n29107_, new_n29108_,
    new_n29109_, new_n29110_, new_n29111_, new_n29112_, new_n29113_,
    new_n29114_, new_n29115_, new_n29116_, new_n29117_, new_n29118_,
    new_n29119_, new_n29120_, new_n29121_, new_n29122_, new_n29123_,
    new_n29124_, new_n29125_, new_n29126_, new_n29127_, new_n29128_,
    new_n29129_, new_n29130_, new_n29131_, new_n29132_, new_n29133_,
    new_n29134_, new_n29135_, new_n29136_, new_n29137_, new_n29138_,
    new_n29139_, new_n29140_, new_n29141_, new_n29142_, new_n29143_,
    new_n29144_, new_n29145_, new_n29146_, new_n29147_, new_n29148_,
    new_n29149_, new_n29150_, new_n29151_, new_n29152_, new_n29153_,
    new_n29154_, new_n29155_, new_n29156_, new_n29157_, new_n29158_,
    new_n29159_, new_n29160_, new_n29161_, new_n29162_, new_n29164_,
    new_n29165_, new_n29166_, new_n29167_, new_n29168_, new_n29169_,
    new_n29170_, new_n29171_, new_n29172_, new_n29173_, new_n29174_,
    new_n29175_, new_n29176_, new_n29177_, new_n29178_, new_n29179_,
    new_n29180_, new_n29181_, new_n29182_, new_n29183_, new_n29184_,
    new_n29185_, new_n29186_, new_n29187_, new_n29188_, new_n29189_,
    new_n29190_, new_n29191_, new_n29192_, new_n29193_, new_n29194_,
    new_n29195_, new_n29196_, new_n29197_, new_n29198_, new_n29199_,
    new_n29200_, new_n29201_, new_n29202_, new_n29203_, new_n29204_,
    new_n29205_, new_n29206_, new_n29207_, new_n29208_, new_n29209_,
    new_n29210_, new_n29211_, new_n29212_, new_n29213_, new_n29214_,
    new_n29215_, new_n29216_, new_n29217_, new_n29218_, new_n29219_,
    new_n29220_, new_n29221_, new_n29222_, new_n29223_, new_n29224_,
    new_n29225_, new_n29226_, new_n29227_, new_n29228_, new_n29229_,
    new_n29230_, new_n29231_, new_n29232_, new_n29233_, new_n29234_,
    new_n29235_, new_n29236_, new_n29237_, new_n29238_, new_n29239_,
    new_n29240_, new_n29241_, new_n29242_, new_n29243_, new_n29244_,
    new_n29245_, new_n29246_, new_n29247_, new_n29248_, new_n29249_,
    new_n29250_, new_n29252_, new_n29253_, new_n29254_, new_n29255_,
    new_n29256_, new_n29257_, new_n29258_, new_n29259_, new_n29260_,
    new_n29261_, new_n29262_, new_n29263_, new_n29264_, new_n29265_,
    new_n29266_, new_n29267_, new_n29268_, new_n29269_, new_n29270_,
    new_n29271_, new_n29272_, new_n29273_, new_n29274_, new_n29275_,
    new_n29276_, new_n29277_, new_n29278_, new_n29279_, new_n29280_,
    new_n29281_, new_n29282_, new_n29283_, new_n29284_, new_n29285_,
    new_n29286_, new_n29287_, new_n29288_, new_n29289_, new_n29290_,
    new_n29291_, new_n29292_, new_n29293_, new_n29294_, new_n29295_,
    new_n29296_, new_n29297_, new_n29298_, new_n29299_, new_n29300_,
    new_n29301_, new_n29302_, new_n29303_, new_n29304_, new_n29305_,
    new_n29306_, new_n29307_, new_n29308_, new_n29309_, new_n29310_,
    new_n29311_, new_n29312_, new_n29313_, new_n29314_, new_n29315_,
    new_n29316_, new_n29317_, new_n29318_, new_n29319_, new_n29320_,
    new_n29321_, new_n29322_, new_n29323_, new_n29324_, new_n29325_,
    new_n29326_, new_n29327_, new_n29328_, new_n29329_, new_n29330_,
    new_n29331_, new_n29332_, new_n29333_, new_n29334_, new_n29335_,
    new_n29336_, new_n29337_, new_n29338_, new_n29340_, new_n29341_,
    new_n29342_, new_n29343_, new_n29344_, new_n29345_, new_n29346_,
    new_n29347_, new_n29348_, new_n29349_, new_n29350_, new_n29351_,
    new_n29352_, new_n29353_, new_n29354_, new_n29355_, new_n29356_,
    new_n29357_, new_n29358_, new_n29359_, new_n29360_, new_n29361_,
    new_n29362_, new_n29363_, new_n29364_, new_n29365_, new_n29366_,
    new_n29367_, new_n29368_, new_n29369_, new_n29370_, new_n29371_,
    new_n29372_, new_n29373_, new_n29374_, new_n29375_, new_n29376_,
    new_n29377_, new_n29378_, new_n29379_, new_n29380_, new_n29381_,
    new_n29382_, new_n29383_, new_n29384_, new_n29385_, new_n29386_,
    new_n29387_, new_n29388_, new_n29389_, new_n29390_, new_n29391_,
    new_n29392_, new_n29393_, new_n29394_, new_n29395_, new_n29396_,
    new_n29397_, new_n29398_, new_n29399_, new_n29400_, new_n29401_,
    new_n29402_, new_n29403_, new_n29404_, new_n29405_, new_n29406_,
    new_n29407_, new_n29408_, new_n29409_, new_n29410_, new_n29411_,
    new_n29412_, new_n29413_, new_n29414_, new_n29415_, new_n29416_,
    new_n29417_, new_n29418_, new_n29419_, new_n29420_, new_n29421_,
    new_n29422_, new_n29423_, new_n29424_, new_n29425_, new_n29426_,
    new_n29428_, new_n29429_, new_n29430_, new_n29431_, new_n29432_,
    new_n29433_, new_n29434_, new_n29435_, new_n29436_, new_n29437_,
    new_n29438_, new_n29439_, new_n29440_, new_n29441_, new_n29442_,
    new_n29443_, new_n29444_, new_n29445_, new_n29446_, new_n29447_,
    new_n29448_, new_n29449_, new_n29450_, new_n29451_, new_n29452_,
    new_n29453_, new_n29454_, new_n29455_, new_n29456_, new_n29457_,
    new_n29458_, new_n29459_, new_n29460_, new_n29461_, new_n29462_,
    new_n29463_, new_n29464_, new_n29465_, new_n29466_, new_n29467_,
    new_n29468_, new_n29469_, new_n29470_, new_n29471_, new_n29472_,
    new_n29473_, new_n29474_, new_n29475_, new_n29476_, new_n29477_,
    new_n29478_, new_n29479_, new_n29480_, new_n29481_, new_n29482_,
    new_n29483_, new_n29484_, new_n29485_, new_n29486_, new_n29487_,
    new_n29488_, new_n29489_, new_n29490_, new_n29491_, new_n29492_,
    new_n29493_, new_n29494_, new_n29495_, new_n29496_, new_n29497_,
    new_n29498_, new_n29499_, new_n29500_, new_n29501_, new_n29502_,
    new_n29503_, new_n29504_, new_n29505_, new_n29506_, new_n29507_,
    new_n29508_, new_n29509_, new_n29510_, new_n29511_, new_n29512_,
    new_n29513_, new_n29514_, new_n29516_, new_n29517_, new_n29518_,
    new_n29519_, new_n29520_, new_n29521_, new_n29522_, new_n29523_,
    new_n29524_, new_n29525_, new_n29526_, new_n29527_, new_n29528_,
    new_n29529_, new_n29530_, new_n29531_, new_n29532_, new_n29533_,
    new_n29534_, new_n29535_, new_n29536_, new_n29537_, new_n29538_,
    new_n29539_, new_n29540_, new_n29541_, new_n29542_, new_n29543_,
    new_n29544_, new_n29545_, new_n29546_, new_n29547_, new_n29548_,
    new_n29549_, new_n29550_, new_n29551_, new_n29552_, new_n29553_,
    new_n29554_, new_n29555_, new_n29556_, new_n29557_, new_n29558_,
    new_n29559_, new_n29560_, new_n29561_, new_n29562_, new_n29563_,
    new_n29564_, new_n29565_, new_n29566_, new_n29567_, new_n29568_,
    new_n29569_, new_n29570_, new_n29571_, new_n29572_, new_n29573_,
    new_n29574_, new_n29575_, new_n29576_, new_n29577_, new_n29578_,
    new_n29579_, new_n29580_, new_n29581_, new_n29582_, new_n29583_,
    new_n29584_, new_n29585_, new_n29586_, new_n29587_, new_n29588_,
    new_n29589_, new_n29590_, new_n29591_, new_n29592_, new_n29593_,
    new_n29594_, new_n29595_, new_n29596_, new_n29597_, new_n29598_,
    new_n29599_, new_n29600_, new_n29601_, new_n29602_, new_n29604_,
    new_n29605_, new_n29606_, new_n29607_, new_n29608_, new_n29609_,
    new_n29610_, new_n29611_, new_n29612_, new_n29613_, new_n29614_,
    new_n29615_, new_n29616_, new_n29617_, new_n29618_, new_n29619_,
    new_n29620_, new_n29621_, new_n29622_, new_n29623_, new_n29624_,
    new_n29625_, new_n29626_, new_n29627_, new_n29628_, new_n29629_,
    new_n29630_, new_n29631_, new_n29632_, new_n29633_, new_n29634_,
    new_n29635_, new_n29636_, new_n29637_, new_n29638_, new_n29639_,
    new_n29640_, new_n29641_, new_n29642_, new_n29643_, new_n29644_,
    new_n29645_, new_n29646_, new_n29647_, new_n29648_, new_n29649_,
    new_n29650_, new_n29651_, new_n29652_, new_n29653_, new_n29654_,
    new_n29655_, new_n29656_, new_n29657_, new_n29658_, new_n29659_,
    new_n29660_, new_n29661_, new_n29662_, new_n29663_, new_n29664_,
    new_n29665_, new_n29666_, new_n29667_, new_n29668_, new_n29669_,
    new_n29670_, new_n29671_, new_n29672_, new_n29673_, new_n29674_,
    new_n29675_, new_n29676_, new_n29677_, new_n29678_, new_n29679_,
    new_n29680_, new_n29681_, new_n29682_, new_n29683_, new_n29684_,
    new_n29685_, new_n29686_, new_n29687_, new_n29688_, new_n29689_,
    new_n29690_, new_n29691_, new_n29692_, new_n29693_, new_n29694_,
    new_n29695_, new_n29697_, new_n29698_, new_n29699_, new_n29700_,
    new_n29701_, new_n29702_, new_n29703_, new_n29704_, new_n29705_,
    new_n29706_, new_n29707_, new_n29708_, new_n29709_, new_n29710_,
    new_n29711_, new_n29712_, new_n29713_, new_n29714_, new_n29715_,
    new_n29716_, new_n29717_, new_n29718_, new_n29719_, new_n29720_,
    new_n29721_, new_n29722_, new_n29723_, new_n29724_, new_n29725_,
    new_n29726_, new_n29727_, new_n29728_, new_n29729_, new_n29730_,
    new_n29731_, new_n29732_, new_n29733_, new_n29734_, new_n29735_,
    new_n29736_, new_n29737_, new_n29738_, new_n29739_, new_n29740_,
    new_n29741_, new_n29742_, new_n29743_, new_n29744_, new_n29745_,
    new_n29746_, new_n29747_, new_n29748_, new_n29749_, new_n29750_,
    new_n29751_, new_n29752_, new_n29753_, new_n29754_, new_n29755_,
    new_n29756_, new_n29757_, new_n29758_, new_n29759_, new_n29760_,
    new_n29761_, new_n29762_, new_n29763_, new_n29764_, new_n29765_,
    new_n29766_, new_n29767_, new_n29768_, new_n29769_, new_n29770_,
    new_n29771_, new_n29772_, new_n29773_, new_n29774_, new_n29775_,
    new_n29776_, new_n29777_, new_n29778_, new_n29779_, new_n29780_,
    new_n29781_, new_n29782_, new_n29783_, new_n29785_, new_n29786_,
    new_n29787_, new_n29788_, new_n29789_, new_n29790_, new_n29791_,
    new_n29792_, new_n29793_, new_n29794_, new_n29795_, new_n29796_,
    new_n29797_, new_n29798_, new_n29799_, new_n29800_, new_n29801_,
    new_n29802_, new_n29803_, new_n29804_, new_n29805_, new_n29806_,
    new_n29807_, new_n29808_, new_n29809_, new_n29810_, new_n29811_,
    new_n29812_, new_n29813_, new_n29814_, new_n29815_, new_n29816_,
    new_n29817_, new_n29818_, new_n29819_, new_n29820_, new_n29821_,
    new_n29822_, new_n29823_, new_n29824_, new_n29825_, new_n29826_,
    new_n29827_, new_n29828_, new_n29829_, new_n29830_, new_n29831_,
    new_n29832_, new_n29833_, new_n29834_, new_n29835_, new_n29836_,
    new_n29837_, new_n29838_, new_n29839_, new_n29840_, new_n29841_,
    new_n29842_, new_n29843_, new_n29844_, new_n29845_, new_n29846_,
    new_n29847_, new_n29848_, new_n29849_, new_n29850_, new_n29851_,
    new_n29852_, new_n29853_, new_n29854_, new_n29855_, new_n29856_,
    new_n29857_, new_n29858_, new_n29859_, new_n29860_, new_n29861_,
    new_n29862_, new_n29863_, new_n29864_, new_n29865_, new_n29866_,
    new_n29867_, new_n29868_, new_n29869_, new_n29870_, new_n29871_,
    new_n29873_, new_n29874_, new_n29875_, new_n29876_, new_n29877_,
    new_n29878_, new_n29879_, new_n29880_, new_n29881_, new_n29882_,
    new_n29883_, new_n29884_, new_n29885_, new_n29886_, new_n29887_,
    new_n29888_, new_n29889_, new_n29890_, new_n29891_, new_n29892_,
    new_n29893_, new_n29894_, new_n29895_, new_n29896_, new_n29897_,
    new_n29898_, new_n29899_, new_n29900_, new_n29901_, new_n29902_,
    new_n29903_, new_n29904_, new_n29905_, new_n29906_, new_n29907_,
    new_n29908_, new_n29909_, new_n29910_, new_n29911_, new_n29912_,
    new_n29913_, new_n29914_, new_n29915_, new_n29916_, new_n29917_,
    new_n29918_, new_n29919_, new_n29920_, new_n29921_, new_n29922_,
    new_n29923_, new_n29924_, new_n29925_, new_n29926_, new_n29927_,
    new_n29928_, new_n29929_, new_n29930_, new_n29931_, new_n29932_,
    new_n29933_, new_n29934_, new_n29935_, new_n29936_, new_n29937_,
    new_n29938_, new_n29939_, new_n29940_, new_n29941_, new_n29942_,
    new_n29943_, new_n29944_, new_n29945_, new_n29946_, new_n29947_,
    new_n29948_, new_n29949_, new_n29950_, new_n29951_, new_n29952_,
    new_n29953_, new_n29954_, new_n29955_, new_n29956_, new_n29957_,
    new_n29958_, new_n29959_, new_n29961_, new_n29962_, new_n29963_,
    new_n29964_, new_n29965_, new_n29966_, new_n29967_, new_n29968_,
    new_n29969_, new_n29970_, new_n29971_, new_n29972_, new_n29973_,
    new_n29974_, new_n29975_, new_n29976_, new_n29977_, new_n29978_,
    new_n29979_, new_n29980_, new_n29981_, new_n29982_, new_n29983_,
    new_n29984_, new_n29985_, new_n29986_, new_n29987_, new_n29988_,
    new_n29989_, new_n29990_, new_n29991_, new_n29992_, new_n29993_,
    new_n29994_, new_n29995_, new_n29996_, new_n29997_, new_n29998_,
    new_n29999_, new_n30000_, new_n30001_, new_n30002_, new_n30003_,
    new_n30004_, new_n30005_, new_n30006_, new_n30007_, new_n30008_,
    new_n30009_, new_n30010_, new_n30011_, new_n30012_, new_n30013_,
    new_n30014_, new_n30015_, new_n30016_, new_n30017_, new_n30018_,
    new_n30019_, new_n30020_, new_n30021_, new_n30022_, new_n30023_,
    new_n30024_, new_n30025_, new_n30026_, new_n30027_, new_n30028_,
    new_n30029_, new_n30030_, new_n30031_, new_n30032_, new_n30033_,
    new_n30034_, new_n30035_, new_n30037_, new_n30038_, new_n30039_,
    new_n30040_, new_n30041_, new_n30042_, new_n30043_, new_n30044_,
    new_n30045_, new_n30046_, new_n30047_, new_n30048_, new_n30049_,
    new_n30050_, new_n30051_, new_n30052_, new_n30053_, new_n30054_,
    new_n30055_, new_n30056_, new_n30057_, new_n30058_, new_n30059_,
    new_n30060_, new_n30061_, new_n30062_, new_n30063_, new_n30064_,
    new_n30065_, new_n30066_, new_n30067_, new_n30068_, new_n30069_,
    new_n30070_, new_n30071_, new_n30072_, new_n30073_, new_n30074_,
    new_n30075_, new_n30076_, new_n30077_, new_n30078_, new_n30079_,
    new_n30080_, new_n30081_, new_n30082_, new_n30083_, new_n30084_,
    new_n30085_, new_n30086_, new_n30087_, new_n30088_, new_n30089_,
    new_n30090_, new_n30091_, new_n30092_, new_n30093_, new_n30094_,
    new_n30095_, new_n30096_, new_n30097_, new_n30098_, new_n30099_,
    new_n30100_, new_n30101_, new_n30102_, new_n30103_, new_n30104_,
    new_n30105_, new_n30106_, new_n30107_, new_n30108_, new_n30109_,
    new_n30110_, new_n30111_, new_n30112_, new_n30113_, new_n30114_,
    new_n30115_, new_n30116_, new_n30117_, new_n30118_, new_n30119_,
    new_n30121_, new_n30122_, new_n30123_, new_n30124_, new_n30125_,
    new_n30126_, new_n30127_, new_n30128_, new_n30129_, new_n30130_,
    new_n30131_, new_n30132_, new_n30133_, new_n30134_, new_n30135_,
    new_n30136_, new_n30137_, new_n30138_, new_n30139_, new_n30140_,
    new_n30141_, new_n30142_, new_n30143_, new_n30144_, new_n30145_,
    new_n30146_, new_n30147_, new_n30148_, new_n30149_, new_n30150_,
    new_n30151_, new_n30152_, new_n30153_, new_n30154_, new_n30155_,
    new_n30156_, new_n30157_, new_n30158_, new_n30159_, new_n30160_,
    new_n30161_, new_n30162_, new_n30163_, new_n30164_, new_n30165_,
    new_n30166_, new_n30167_, new_n30168_, new_n30169_, new_n30170_,
    new_n30171_, new_n30172_, new_n30173_, new_n30174_, new_n30175_,
    new_n30176_, new_n30177_, new_n30178_, new_n30179_, new_n30180_,
    new_n30181_, new_n30182_, new_n30183_, new_n30184_, new_n30185_,
    new_n30186_, new_n30187_, new_n30188_, new_n30189_, new_n30190_,
    new_n30191_, new_n30192_, new_n30193_, new_n30194_, new_n30195_,
    new_n30196_, new_n30197_, new_n30198_, new_n30199_, new_n30200_,
    new_n30201_, new_n30202_, new_n30203_, new_n30204_, new_n30205_,
    new_n30206_, new_n30207_, new_n30208_, new_n30209_, new_n30210_,
    new_n30211_, new_n30212_, new_n30213_, new_n30214_, new_n30215_,
    new_n30216_, new_n30217_, new_n30218_, new_n30219_, new_n30220_,
    new_n30221_, new_n30222_, new_n30223_, new_n30224_, new_n30225_,
    new_n30226_, new_n30227_, new_n30228_, new_n30229_, new_n30230_,
    new_n30231_, new_n30232_, new_n30233_, new_n30234_, new_n30235_,
    new_n30236_, new_n30237_, new_n30238_, new_n30239_, new_n30241_,
    new_n30242_, new_n30243_, new_n30244_, new_n30245_, new_n30246_,
    new_n30247_, new_n30248_, new_n30249_, new_n30250_, new_n30251_,
    new_n30252_, new_n30253_, new_n30254_, new_n30255_, new_n30256_,
    new_n30257_, new_n30258_, new_n30259_, new_n30260_, new_n30261_,
    new_n30262_, new_n30263_, new_n30264_, new_n30265_, new_n30266_,
    new_n30267_, new_n30268_, new_n30269_, new_n30270_, new_n30271_,
    new_n30272_, new_n30273_, new_n30274_, new_n30275_, new_n30276_,
    new_n30277_, new_n30278_, new_n30279_, new_n30280_, new_n30281_,
    new_n30282_, new_n30283_, new_n30284_, new_n30285_, new_n30286_,
    new_n30287_, new_n30288_, new_n30289_, new_n30290_, new_n30291_,
    new_n30292_, new_n30293_, new_n30294_, new_n30295_, new_n30296_,
    new_n30297_, new_n30298_, new_n30299_, new_n30300_, new_n30301_,
    new_n30302_, new_n30303_, new_n30304_, new_n30305_, new_n30306_,
    new_n30307_, new_n30308_, new_n30309_, new_n30310_, new_n30311_,
    new_n30312_, new_n30313_, new_n30314_, new_n30315_, new_n30316_,
    new_n30317_, new_n30318_, new_n30319_, new_n30320_, new_n30321_,
    new_n30322_, new_n30323_, new_n30324_, new_n30325_, new_n30326_,
    new_n30327_, new_n30328_, new_n30329_, new_n30330_, new_n30331_,
    new_n30332_, new_n30333_, new_n30334_, new_n30335_, new_n30336_,
    new_n30337_, new_n30338_, new_n30340_, new_n30341_, new_n30342_,
    new_n30343_, new_n30344_, new_n30345_, new_n30346_, new_n30347_,
    new_n30348_, new_n30349_, new_n30350_, new_n30351_, new_n30352_,
    new_n30353_, new_n30354_, new_n30355_, new_n30356_, new_n30357_,
    new_n30358_, new_n30359_, new_n30360_, new_n30361_, new_n30362_,
    new_n30363_, new_n30364_, new_n30365_, new_n30366_, new_n30367_,
    new_n30368_, new_n30369_, new_n30370_, new_n30371_, new_n30372_,
    new_n30373_, new_n30374_, new_n30375_, new_n30376_, new_n30377_,
    new_n30378_, new_n30379_, new_n30380_, new_n30381_, new_n30382_,
    new_n30383_, new_n30384_, new_n30385_, new_n30386_, new_n30387_,
    new_n30388_, new_n30389_, new_n30390_, new_n30391_, new_n30392_,
    new_n30393_, new_n30394_, new_n30395_, new_n30396_, new_n30397_,
    new_n30398_, new_n30399_, new_n30400_, new_n30401_, new_n30402_,
    new_n30403_, new_n30404_, new_n30405_, new_n30406_, new_n30407_,
    new_n30408_, new_n30409_, new_n30410_, new_n30411_, new_n30412_,
    new_n30413_, new_n30414_, new_n30415_, new_n30416_, new_n30417_,
    new_n30418_, new_n30419_, new_n30420_, new_n30421_, new_n30422_,
    new_n30423_, new_n30424_, new_n30425_, new_n30426_, new_n30427_,
    new_n30428_, new_n30429_, new_n30430_, new_n30431_, new_n30432_,
    new_n30433_, new_n30434_, new_n30435_, new_n30436_, new_n30437_,
    new_n30438_, new_n30440_, new_n30441_, new_n30442_, new_n30443_,
    new_n30444_, new_n30445_, new_n30446_, new_n30447_, new_n30448_,
    new_n30449_, new_n30450_, new_n30451_, new_n30452_, new_n30453_,
    new_n30454_, new_n30455_, new_n30456_, new_n30457_, new_n30458_,
    new_n30459_, new_n30460_, new_n30461_, new_n30462_, new_n30463_,
    new_n30464_, new_n30465_, new_n30466_, new_n30467_, new_n30468_,
    new_n30469_, new_n30470_, new_n30471_, new_n30472_, new_n30473_,
    new_n30474_, new_n30475_, new_n30476_, new_n30477_, new_n30478_,
    new_n30479_, new_n30480_, new_n30481_, new_n30482_, new_n30483_,
    new_n30484_, new_n30485_, new_n30486_, new_n30487_, new_n30488_,
    new_n30489_, new_n30490_, new_n30491_, new_n30492_, new_n30493_,
    new_n30494_, new_n30495_, new_n30496_, new_n30497_, new_n30498_,
    new_n30499_, new_n30500_, new_n30501_, new_n30502_, new_n30503_,
    new_n30504_, new_n30505_, new_n30506_, new_n30507_, new_n30508_,
    new_n30509_, new_n30510_, new_n30511_, new_n30512_, new_n30513_,
    new_n30514_, new_n30515_, new_n30516_, new_n30517_, new_n30518_,
    new_n30519_, new_n30520_, new_n30521_, new_n30522_, new_n30523_,
    new_n30524_, new_n30525_, new_n30526_, new_n30527_, new_n30528_,
    new_n30529_, new_n30530_, new_n30531_, new_n30532_, new_n30533_,
    new_n30534_, new_n30535_, new_n30536_, new_n30537_, new_n30538_,
    new_n30540_, new_n30541_, new_n30542_, new_n30543_, new_n30544_,
    new_n30545_, new_n30546_, new_n30547_, new_n30548_, new_n30549_,
    new_n30550_, new_n30551_, new_n30552_, new_n30553_, new_n30554_,
    new_n30555_, new_n30556_, new_n30557_, new_n30558_, new_n30559_,
    new_n30560_, new_n30561_, new_n30562_, new_n30563_, new_n30564_,
    new_n30565_, new_n30566_, new_n30567_, new_n30568_, new_n30569_,
    new_n30570_, new_n30571_, new_n30572_, new_n30573_, new_n30574_,
    new_n30575_, new_n30576_, new_n30577_, new_n30578_, new_n30579_,
    new_n30580_, new_n30581_, new_n30582_, new_n30583_, new_n30584_,
    new_n30585_, new_n30586_, new_n30587_, new_n30588_, new_n30589_,
    new_n30590_, new_n30591_, new_n30592_, new_n30593_, new_n30594_,
    new_n30595_, new_n30596_, new_n30597_, new_n30598_, new_n30599_,
    new_n30600_, new_n30601_, new_n30602_, new_n30603_, new_n30604_,
    new_n30605_, new_n30606_, new_n30607_, new_n30608_, new_n30609_,
    new_n30610_, new_n30611_, new_n30612_, new_n30613_, new_n30614_,
    new_n30615_, new_n30616_, new_n30617_, new_n30618_, new_n30619_,
    new_n30620_, new_n30621_, new_n30622_, new_n30623_, new_n30624_,
    new_n30625_, new_n30626_, new_n30627_, new_n30628_, new_n30629_,
    new_n30630_, new_n30631_, new_n30632_, new_n30633_, new_n30634_,
    new_n30635_, new_n30636_, new_n30637_, new_n30638_, new_n30640_,
    new_n30641_, new_n30642_, new_n30643_, new_n30644_, new_n30645_,
    new_n30646_, new_n30647_, new_n30648_, new_n30649_, new_n30650_,
    new_n30651_, new_n30652_, new_n30653_, new_n30654_, new_n30655_,
    new_n30656_, new_n30657_, new_n30658_, new_n30659_, new_n30660_,
    new_n30661_, new_n30662_, new_n30663_, new_n30664_, new_n30665_,
    new_n30666_, new_n30667_, new_n30668_, new_n30669_, new_n30670_,
    new_n30671_, new_n30672_, new_n30673_, new_n30674_, new_n30675_,
    new_n30676_, new_n30677_, new_n30678_, new_n30679_, new_n30680_,
    new_n30681_, new_n30682_, new_n30683_, new_n30684_, new_n30685_,
    new_n30686_, new_n30687_, new_n30688_, new_n30689_, new_n30690_,
    new_n30691_, new_n30692_, new_n30693_, new_n30694_, new_n30695_,
    new_n30696_, new_n30697_, new_n30698_, new_n30699_, new_n30700_,
    new_n30701_, new_n30702_, new_n30703_, new_n30704_, new_n30705_,
    new_n30706_, new_n30707_, new_n30708_, new_n30709_, new_n30710_,
    new_n30711_, new_n30712_, new_n30713_, new_n30714_, new_n30715_,
    new_n30716_, new_n30717_, new_n30718_, new_n30719_, new_n30720_,
    new_n30721_, new_n30722_, new_n30723_, new_n30724_, new_n30725_,
    new_n30726_, new_n30727_, new_n30728_, new_n30729_, new_n30731_,
    new_n30732_, new_n30733_, new_n30734_, new_n30735_, new_n30736_,
    new_n30737_, new_n30738_, new_n30739_, new_n30740_, new_n30741_,
    new_n30742_, new_n30743_, new_n30744_, new_n30745_, new_n30746_,
    new_n30747_, new_n30748_, new_n30749_, new_n30750_, new_n30751_,
    new_n30752_, new_n30753_, new_n30754_, new_n30755_, new_n30756_,
    new_n30757_, new_n30758_, new_n30759_, new_n30760_, new_n30761_,
    new_n30762_, new_n30763_, new_n30764_, new_n30765_, new_n30766_,
    new_n30767_, new_n30768_, new_n30769_, new_n30770_, new_n30771_,
    new_n30772_, new_n30773_, new_n30774_, new_n30775_, new_n30776_,
    new_n30777_, new_n30778_, new_n30779_, new_n30780_, new_n30781_,
    new_n30782_, new_n30783_, new_n30784_, new_n30785_, new_n30786_,
    new_n30787_, new_n30788_, new_n30789_, new_n30790_, new_n30791_,
    new_n30792_, new_n30793_, new_n30794_, new_n30795_, new_n30796_,
    new_n30797_, new_n30798_, new_n30799_, new_n30800_, new_n30801_,
    new_n30802_, new_n30803_, new_n30804_, new_n30805_, new_n30806_,
    new_n30807_, new_n30808_, new_n30809_, new_n30810_, new_n30811_,
    new_n30812_, new_n30813_, new_n30814_, new_n30815_, new_n30816_,
    new_n30817_, new_n30818_, new_n30819_, new_n30820_, new_n30822_,
    new_n30823_, new_n30824_, new_n30825_, new_n30826_, new_n30827_,
    new_n30829_, new_n30830_, new_n30831_, new_n30832_, new_n30833_,
    new_n30834_, new_n30835_, new_n30836_, new_n30838_, new_n30839_,
    new_n30840_, new_n30841_, new_n30842_, new_n30843_, new_n30844_,
    new_n30845_, new_n30846_, new_n30848_, new_n30849_, new_n30850_,
    new_n30851_, new_n30852_, new_n30853_, new_n30854_, new_n30855_,
    new_n30856_, new_n30858_, new_n30859_, new_n30860_, new_n30861_,
    new_n30862_, new_n30863_, new_n30864_, new_n30865_, new_n30866_,
    new_n30867_, new_n30869_, new_n30870_, new_n30871_, new_n30872_,
    new_n30873_, new_n30874_, new_n30875_, new_n30876_, new_n30877_,
    new_n30879_, new_n30880_, new_n30881_, new_n30882_, new_n30883_,
    new_n30884_, new_n30885_, new_n30886_, new_n30887_, new_n30888_,
    new_n30889_, new_n30891_, new_n30892_, new_n30893_, new_n30894_,
    new_n30895_, new_n30896_, new_n30897_, new_n30898_, new_n30899_,
    new_n30901_, new_n30902_, new_n30903_, new_n30904_, new_n30905_,
    new_n30906_, new_n30907_, new_n30908_, new_n30909_, new_n30910_,
    new_n30912_, new_n30913_, new_n30914_, new_n30915_, new_n30916_,
    new_n30917_, new_n30918_, new_n30919_, new_n30920_, new_n30922_,
    new_n30923_, new_n30924_, new_n30925_, new_n30926_, new_n30927_,
    new_n30928_, new_n30929_, new_n30930_, new_n30931_, new_n30932_,
    new_n30934_, new_n30935_, new_n30936_, new_n30937_, new_n30938_,
    new_n30939_, new_n30940_, new_n30941_, new_n30942_, new_n30944_,
    new_n30945_, new_n30946_, new_n30947_, new_n30948_, new_n30949_,
    new_n30950_, new_n30951_, new_n30952_, new_n30953_, new_n30955_,
    new_n30956_, new_n30957_, new_n30958_, new_n30959_, new_n30960_,
    new_n30961_, new_n30962_, new_n30963_, new_n30965_, new_n30966_,
    new_n30967_, new_n30968_, new_n30969_, new_n30970_, new_n30971_,
    new_n30972_, new_n30973_, new_n30974_, new_n30975_, new_n30976_,
    new_n30978_, new_n30979_, new_n30980_, new_n30981_, new_n30982_,
    new_n30983_, new_n30984_, new_n30985_, new_n30986_, new_n30988_,
    new_n30989_, new_n30990_, new_n30991_, new_n30992_, new_n30993_,
    new_n30994_, new_n30995_, new_n30996_, new_n30997_, new_n30999_,
    new_n31000_, new_n31001_, new_n31002_, new_n31003_, new_n31004_,
    new_n31005_, new_n31006_, new_n31007_, new_n31009_, new_n31010_,
    new_n31011_, new_n31012_, new_n31013_, new_n31014_, new_n31015_,
    new_n31016_, new_n31017_, new_n31018_, new_n31019_, new_n31021_,
    new_n31022_, new_n31023_, new_n31024_, new_n31025_, new_n31026_,
    new_n31027_, new_n31028_, new_n31029_, new_n31031_, new_n31032_,
    new_n31033_, new_n31034_, new_n31035_, new_n31036_, new_n31037_,
    new_n31038_, new_n31039_, new_n31040_, new_n31042_, new_n31043_,
    new_n31044_, new_n31045_, new_n31046_, new_n31047_, new_n31048_,
    new_n31049_, new_n31050_, new_n31052_, new_n31053_, new_n31054_,
    new_n31055_, new_n31056_, new_n31057_, new_n31058_, new_n31059_,
    new_n31060_, new_n31061_, new_n31062_, new_n31063_, new_n31065_,
    new_n31066_, new_n31067_, new_n31068_, new_n31069_, new_n31070_,
    new_n31071_, new_n31072_, new_n31073_, new_n31075_, new_n31076_,
    new_n31077_, new_n31078_, new_n31079_, new_n31080_, new_n31081_,
    new_n31082_, new_n31083_, new_n31084_, new_n31086_, new_n31087_,
    new_n31088_, new_n31089_, new_n31090_, new_n31091_, new_n31092_,
    new_n31093_, new_n31094_, new_n31096_, new_n31097_, new_n31098_,
    new_n31099_, new_n31100_, new_n31101_, new_n31102_, new_n31103_,
    new_n31104_, new_n31105_, new_n31106_, new_n31108_, new_n31109_,
    new_n31110_, new_n31111_, new_n31112_, new_n31113_, new_n31114_,
    new_n31115_, new_n31116_, new_n31118_, new_n31119_, new_n31120_,
    new_n31121_, new_n31122_, new_n31123_, new_n31124_, new_n31125_,
    new_n31126_, new_n31127_, new_n31129_, new_n31130_, new_n31131_,
    new_n31132_, new_n31133_, new_n31134_, new_n31135_, new_n31136_,
    new_n31137_, new_n31139_, new_n31141_, new_n31144_, new_n31146_,
    new_n31148_, new_n31149_, new_n31150_, new_n31151_, new_n31152_,
    new_n31156_, new_n31157_, new_n31159_, new_n31160_, new_n31161_,
    new_n31162_, new_n31163_, new_n31164_, new_n31165_, new_n31166_,
    new_n31167_, new_n31168_, new_n31169_, new_n31170_, new_n31171_,
    new_n31172_, new_n31173_, new_n31174_, new_n31175_, new_n31176_,
    new_n31177_, new_n31178_, new_n31180_, new_n31181_, new_n31182_,
    new_n31183_, new_n31184_, new_n31185_, new_n31186_, new_n31187_,
    new_n31188_, new_n31189_, new_n31190_, new_n31191_, new_n31192_,
    new_n31193_, new_n31194_, new_n31195_, new_n31196_, new_n31197_,
    new_n31199_, new_n31200_, new_n31201_, new_n31202_, new_n31203_,
    new_n31204_, new_n31205_, new_n31206_, new_n31207_, new_n31208_,
    new_n31209_, new_n31210_, new_n31211_, new_n31212_, new_n31213_,
    new_n31214_, new_n31215_, new_n31216_, new_n31218_, new_n31219_,
    new_n31220_, new_n31221_, new_n31222_, new_n31223_, new_n31224_,
    new_n31225_, new_n31226_, new_n31227_, new_n31228_, new_n31229_,
    new_n31230_, new_n31231_, new_n31232_, new_n31233_, new_n31234_,
    new_n31235_, new_n31237_, new_n31238_, new_n31239_, new_n31240_,
    new_n31241_, new_n31242_, new_n31243_, new_n31244_, new_n31245_,
    new_n31246_, new_n31247_, new_n31248_, new_n31249_, new_n31250_,
    new_n31251_, new_n31252_, new_n31253_, new_n31254_, new_n31256_,
    new_n31257_, new_n31258_, new_n31259_, new_n31260_, new_n31261_,
    new_n31262_, new_n31263_, new_n31264_, new_n31265_, new_n31266_,
    new_n31267_, new_n31268_, new_n31269_, new_n31270_, new_n31271_,
    new_n31272_, new_n31273_, new_n31275_, new_n31276_, new_n31277_,
    new_n31278_, new_n31279_, new_n31280_, new_n31281_, new_n31282_,
    new_n31283_, new_n31284_, new_n31285_, new_n31286_, new_n31287_,
    new_n31288_, new_n31289_, new_n31290_, new_n31291_, new_n31292_,
    new_n31294_, new_n31295_, new_n31296_, new_n31297_, new_n31298_,
    new_n31299_, new_n31300_, new_n31301_, new_n31302_, new_n31303_,
    new_n31304_, new_n31305_, new_n31306_, new_n31307_, new_n31308_,
    new_n31309_, new_n31310_, new_n31311_, new_n31313_, new_n31314_,
    new_n31315_, new_n31316_, new_n31317_, new_n31318_, new_n31319_,
    new_n31320_, new_n31321_, new_n31322_, new_n31323_, new_n31324_,
    new_n31325_, new_n31326_, new_n31327_, new_n31328_, new_n31329_,
    new_n31330_, new_n31331_, new_n31332_, new_n31334_, new_n31335_,
    new_n31336_, new_n31337_, new_n31338_, new_n31339_, new_n31340_,
    new_n31341_, new_n31342_, new_n31343_, new_n31344_, new_n31345_,
    new_n31346_, new_n31347_, new_n31348_, new_n31349_, new_n31350_,
    new_n31351_, new_n31352_, new_n31353_, new_n31355_, new_n31356_,
    new_n31357_, new_n31358_, new_n31359_, new_n31360_, new_n31361_,
    new_n31362_, new_n31363_, new_n31364_, new_n31365_, new_n31366_,
    new_n31367_, new_n31368_, new_n31369_, new_n31370_, new_n31371_,
    new_n31372_, new_n31374_, new_n31375_, new_n31376_, new_n31377_,
    new_n31378_, new_n31379_, new_n31380_, new_n31381_, new_n31382_,
    new_n31383_, new_n31384_, new_n31385_, new_n31386_, new_n31387_,
    new_n31388_, new_n31389_, new_n31390_, new_n31391_, new_n31392_,
    new_n31393_, new_n31395_, new_n31396_, new_n31397_, new_n31398_,
    new_n31399_, new_n31400_, new_n31401_, new_n31402_, new_n31403_,
    new_n31404_, new_n31405_, new_n31406_, new_n31407_, new_n31408_,
    new_n31409_, new_n31410_, new_n31411_, new_n31412_, new_n31413_,
    new_n31414_, new_n31416_, new_n31417_, new_n31418_, new_n31419_,
    new_n31420_, new_n31421_, new_n31422_, new_n31423_, new_n31424_,
    new_n31425_, new_n31426_, new_n31427_, new_n31428_, new_n31429_,
    new_n31430_, new_n31431_, new_n31432_, new_n31433_, new_n31435_,
    new_n31436_, new_n31437_, new_n31438_, new_n31439_, new_n31440_,
    new_n31441_, new_n31442_, new_n31443_, new_n31444_, new_n31445_,
    new_n31446_, new_n31447_, new_n31448_, new_n31449_, new_n31450_,
    new_n31451_, new_n31452_, new_n31454_, new_n31455_, new_n31456_,
    new_n31457_, new_n31458_, new_n31459_, new_n31460_, new_n31461_,
    new_n31462_, new_n31463_, new_n31464_, new_n31465_, new_n31466_,
    new_n31467_, new_n31468_, new_n31469_, new_n31470_, new_n31471_,
    new_n31473_, new_n31474_, new_n31475_, new_n31476_, new_n31477_,
    new_n31478_, new_n31479_, new_n31480_, new_n31481_, new_n31482_,
    new_n31483_, new_n31484_, new_n31485_, new_n31486_, new_n31487_,
    new_n31488_, new_n31489_, new_n31490_, new_n31491_, new_n31493_,
    new_n31494_, new_n31495_, new_n31496_, new_n31497_, new_n31498_,
    new_n31499_, new_n31500_, new_n31501_, new_n31502_, new_n31503_,
    new_n31504_, new_n31505_, new_n31506_, new_n31507_, new_n31508_,
    new_n31509_, new_n31510_, new_n31512_, new_n31513_, new_n31514_,
    new_n31515_, new_n31516_, new_n31517_, new_n31518_, new_n31519_,
    new_n31520_, new_n31521_, new_n31522_, new_n31523_, new_n31524_,
    new_n31525_, new_n31526_, new_n31527_, new_n31528_, new_n31529_,
    new_n31531_, new_n31532_, new_n31533_, new_n31534_, new_n31535_,
    new_n31536_, new_n31537_, new_n31538_, new_n31539_, new_n31540_,
    new_n31541_, new_n31542_, new_n31543_, new_n31544_, new_n31545_,
    new_n31546_, new_n31547_, new_n31548_, new_n31550_, new_n31551_,
    new_n31552_, new_n31553_, new_n31554_, new_n31555_, new_n31556_,
    new_n31557_, new_n31558_, new_n31559_, new_n31560_, new_n31561_,
    new_n31562_, new_n31563_, new_n31564_, new_n31565_, new_n31566_,
    new_n31567_, new_n31569_, new_n31570_, new_n31571_, new_n31572_,
    new_n31573_, new_n31574_, new_n31575_, new_n31576_, new_n31577_,
    new_n31578_, new_n31579_, new_n31580_, new_n31581_, new_n31582_,
    new_n31583_, new_n31584_, new_n31585_, new_n31586_, new_n31588_,
    new_n31589_, new_n31590_, new_n31591_, new_n31592_, new_n31593_,
    new_n31594_, new_n31595_, new_n31596_, new_n31597_, new_n31598_,
    new_n31599_, new_n31600_, new_n31601_, new_n31602_, new_n31603_,
    new_n31604_, new_n31605_, new_n31607_, new_n31608_, new_n31609_,
    new_n31610_, new_n31611_, new_n31612_, new_n31613_, new_n31614_,
    new_n31615_, new_n31616_, new_n31617_, new_n31618_, new_n31619_,
    new_n31620_, new_n31621_, new_n31622_, new_n31623_, new_n31624_,
    new_n31625_, new_n31627_, new_n31628_, new_n31629_, new_n31630_,
    new_n31631_, new_n31632_, new_n31633_, new_n31634_, new_n31635_,
    new_n31636_, new_n31637_, new_n31638_, new_n31639_, new_n31640_,
    new_n31641_, new_n31642_, new_n31643_, new_n31644_, new_n31646_,
    new_n31647_, new_n31648_, new_n31649_, new_n31650_, new_n31651_,
    new_n31652_, new_n31653_, new_n31654_, new_n31655_, new_n31656_,
    new_n31657_, new_n31658_, new_n31659_, new_n31660_, new_n31661_,
    new_n31662_, new_n31663_, new_n31665_, new_n31666_, new_n31667_,
    new_n31668_, new_n31669_, new_n31670_, new_n31671_, new_n31672_,
    new_n31673_, new_n31674_, new_n31675_, new_n31676_, new_n31677_,
    new_n31678_, new_n31679_, new_n31680_, new_n31681_, new_n31682_,
    new_n31683_, new_n31684_, new_n31686_, new_n31687_, new_n31688_,
    new_n31689_, new_n31690_, new_n31691_, new_n31692_, new_n31693_,
    new_n31694_, new_n31695_, new_n31696_, new_n31697_, new_n31698_,
    new_n31699_, new_n31700_, new_n31701_, new_n31702_, new_n31703_,
    new_n31704_, new_n31705_, new_n31707_, new_n31708_, new_n31709_,
    new_n31710_, new_n31711_, new_n31712_, new_n31713_, new_n31714_,
    new_n31715_, new_n31716_, new_n31717_, new_n31718_, new_n31719_,
    new_n31720_, new_n31721_, new_n31722_, new_n31723_, new_n31724_,
    new_n31726_, new_n31727_, new_n31728_, new_n31729_, new_n31730_,
    new_n31731_, new_n31732_, new_n31733_, new_n31734_, new_n31735_,
    new_n31736_, new_n31737_, new_n31738_, new_n31739_, new_n31740_,
    new_n31741_, new_n31742_, new_n31743_, new_n31745_, new_n31746_,
    new_n31747_, new_n31748_, new_n31749_, new_n31750_, new_n31751_,
    new_n31752_, new_n31753_, new_n31754_, new_n31755_, new_n31756_,
    new_n31757_, new_n31758_, new_n31759_, new_n31760_, new_n31761_,
    new_n31762_, new_n31764_, new_n31765_, new_n31766_, new_n31767_,
    new_n31768_, new_n31769_, new_n31770_, new_n31771_, new_n31772_,
    new_n31773_, new_n31774_, new_n31775_, new_n31776_, new_n31777_,
    new_n31778_, new_n31779_, new_n31780_, new_n31781_, new_n31782_,
    new_n31783_, new_n31784_, new_n31785_, new_n31787_, new_n31788_,
    new_n31789_, new_n31790_, new_n31791_, new_n31792_, new_n31793_,
    new_n31794_, new_n31795_, new_n31796_, new_n31797_, new_n31798_,
    new_n31799_, new_n31800_, new_n31802_, new_n31803_, new_n31804_,
    new_n31805_, new_n31806_, new_n31807_, new_n31808_, new_n31809_,
    new_n31810_, new_n31811_, new_n31812_, new_n31813_, new_n31814_,
    new_n31815_, new_n31817_, new_n31818_, new_n31819_, new_n31820_,
    new_n31821_, new_n31822_, new_n31823_, new_n31824_, new_n31825_,
    new_n31826_, new_n31827_, new_n31828_, new_n31829_, new_n31830_,
    new_n31832_, new_n31833_, new_n31834_, new_n31835_, new_n31836_,
    new_n31837_, new_n31838_, new_n31839_, new_n31840_, new_n31841_,
    new_n31842_, new_n31843_, new_n31844_, new_n31845_, new_n31847_,
    new_n31848_, new_n31849_, new_n31850_, new_n31851_, new_n31852_,
    new_n31853_, new_n31854_, new_n31855_, new_n31856_, new_n31857_,
    new_n31858_, new_n31859_, new_n31860_, new_n31862_, new_n31863_,
    new_n31864_, new_n31865_, new_n31866_, new_n31867_, new_n31868_,
    new_n31869_, new_n31870_, new_n31871_, new_n31872_, new_n31873_,
    new_n31874_, new_n31875_, new_n31877_, new_n31878_, new_n31879_,
    new_n31880_, new_n31881_, new_n31882_, new_n31883_, new_n31884_,
    new_n31885_, new_n31886_, new_n31887_, new_n31888_, new_n31890_,
    new_n31891_, new_n31892_, new_n31893_, new_n31894_, new_n31895_,
    new_n31896_, new_n31897_, new_n31898_, new_n31899_, new_n31900_,
    new_n31901_, new_n31902_, new_n31903_, new_n31905_, new_n31906_,
    new_n31907_, new_n31908_, new_n31909_, new_n31910_, new_n31911_,
    new_n31912_, new_n31913_, new_n31914_, new_n31915_, new_n31916_,
    new_n31917_, new_n31918_, new_n31920_, new_n31921_, new_n31922_,
    new_n31923_, new_n31924_, new_n31925_, new_n31926_, new_n31927_,
    new_n31928_, new_n31929_, new_n31930_, new_n31931_, new_n31932_,
    new_n31933_, new_n31935_, new_n31936_, new_n31937_, new_n31938_,
    new_n31939_, new_n31940_, new_n31941_, new_n31942_, new_n31943_,
    new_n31944_, new_n31945_, new_n31946_, new_n31948_, new_n31949_,
    new_n31950_, new_n31951_, new_n31952_, new_n31953_, new_n31954_,
    new_n31955_, new_n31956_, new_n31957_, new_n31958_, new_n31959_,
    new_n31960_, new_n31961_, new_n31963_, new_n31964_, new_n31965_,
    new_n31966_, new_n31967_, new_n31968_, new_n31969_, new_n31970_,
    new_n31971_, new_n31972_, new_n31973_, new_n31974_, new_n31975_,
    new_n31976_, new_n31978_, new_n31979_, new_n31980_, new_n31981_,
    new_n31982_, new_n31983_, new_n31984_, new_n31985_, new_n31986_,
    new_n31987_, new_n31988_, new_n31989_, new_n31991_, new_n31992_,
    new_n31993_, new_n31994_, new_n31995_, new_n31996_, new_n31997_,
    new_n31998_, new_n31999_, new_n32000_, new_n32001_, new_n32002_,
    new_n32003_, new_n32004_, new_n32006_, new_n32007_, new_n32008_,
    new_n32009_, new_n32010_, new_n32011_, new_n32012_, new_n32013_,
    new_n32014_, new_n32015_, new_n32016_, new_n32017_, new_n32018_,
    new_n32019_, new_n32021_, new_n32022_, new_n32023_, new_n32024_,
    new_n32025_, new_n32026_, new_n32027_, new_n32028_, new_n32029_,
    new_n32030_, new_n32031_, new_n32032_, new_n32033_, new_n32034_,
    new_n32036_, new_n32037_, new_n32038_, new_n32039_, new_n32040_,
    new_n32041_, new_n32042_, new_n32043_, new_n32044_, new_n32045_,
    new_n32046_, new_n32047_, new_n32048_, new_n32049_, new_n32051_,
    new_n32052_, new_n32053_, new_n32054_, new_n32055_, new_n32056_,
    new_n32057_, new_n32058_, new_n32059_, new_n32060_, new_n32061_,
    new_n32062_, new_n32063_, new_n32064_, new_n32066_, new_n32067_,
    new_n32068_, new_n32069_, new_n32070_, new_n32071_, new_n32072_,
    new_n32073_, new_n32074_, new_n32075_, new_n32076_, new_n32077_,
    new_n32078_, new_n32079_, new_n32081_, new_n32082_, new_n32083_,
    new_n32084_, new_n32085_, new_n32086_, new_n32087_, new_n32088_,
    new_n32089_, new_n32090_, new_n32091_, new_n32092_, new_n32093_,
    new_n32094_, new_n32096_, new_n32097_, new_n32098_, new_n32099_,
    new_n32100_, new_n32101_, new_n32102_, new_n32103_, new_n32104_,
    new_n32105_, new_n32106_, new_n32107_, new_n32108_, new_n32110_,
    new_n32111_, new_n32112_, new_n32113_, new_n32114_, new_n32115_,
    new_n32116_, new_n32117_, new_n32118_, new_n32119_, new_n32120_,
    new_n32121_, new_n32122_, new_n32123_, new_n32125_, new_n32126_,
    new_n32127_, new_n32128_, new_n32129_, new_n32130_, new_n32131_,
    new_n32132_, new_n32133_, new_n32134_, new_n32135_, new_n32136_,
    new_n32137_, new_n32138_, new_n32140_, new_n32141_, new_n32142_,
    new_n32143_, new_n32144_, new_n32145_, new_n32146_, new_n32147_,
    new_n32148_, new_n32149_, new_n32150_, new_n32151_, new_n32152_,
    new_n32153_, new_n32155_, new_n32156_, new_n32157_, new_n32158_,
    new_n32159_, new_n32160_, new_n32161_, new_n32162_, new_n32163_,
    new_n32164_, new_n32165_, new_n32166_, new_n32167_, new_n32168_,
    new_n32170_, new_n32171_, new_n32172_, new_n32173_, new_n32174_,
    new_n32175_, new_n32176_, new_n32177_, new_n32178_, new_n32179_,
    new_n32180_, new_n32181_, new_n32183_, new_n32184_, new_n32185_,
    new_n32186_, new_n32187_, new_n32188_, new_n32189_, new_n32190_,
    new_n32191_, new_n32192_, new_n32193_, new_n32194_, new_n32196_,
    new_n32197_, new_n32198_, new_n32199_, new_n32200_, new_n32201_,
    new_n32202_, new_n32203_, new_n32204_, new_n32205_, new_n32206_,
    new_n32207_, new_n32209_, new_n32210_, new_n32211_, new_n32212_,
    new_n32213_, new_n32214_, new_n32215_, new_n32216_, new_n32217_,
    new_n32218_, new_n32219_, new_n32220_, new_n32222_, new_n32223_,
    new_n32224_, new_n32225_, new_n32226_, new_n32227_, new_n32228_,
    new_n32229_, new_n32230_, new_n32231_, new_n32232_, new_n32233_,
    new_n32235_, new_n32236_, new_n32237_, new_n32238_, new_n32239_,
    new_n32240_, new_n32241_, new_n32242_, new_n32243_, new_n32244_,
    new_n32245_, new_n32246_, new_n32247_, new_n32248_, new_n32250_,
    new_n32251_, new_n32252_, new_n32253_, new_n32254_, new_n32255_,
    new_n32256_, new_n32257_, new_n32258_, new_n32259_, new_n32260_,
    new_n32261_, new_n32262_, new_n32263_, new_n32265_, new_n32266_,
    new_n32267_, new_n32268_, new_n32269_, new_n32270_, new_n32271_,
    new_n32272_, new_n32273_, new_n32274_, new_n32275_, new_n32276_,
    new_n32277_, new_n32278_, new_n32280_, new_n32281_, new_n32282_,
    new_n32283_, new_n32284_, new_n32285_, new_n32286_, new_n32287_,
    new_n32288_, new_n32289_, new_n32290_, new_n32291_, new_n32292_,
    new_n32293_, new_n32295_, new_n32296_, new_n32297_, new_n32298_,
    new_n32299_, new_n32300_, new_n32301_, new_n32302_, new_n32303_,
    new_n32304_, new_n32305_, new_n32306_, new_n32307_, new_n32308_,
    new_n32310_, new_n32311_, new_n32312_, new_n32313_, new_n32314_,
    new_n32315_, new_n32316_, new_n32317_, new_n32318_, new_n32319_,
    new_n32320_, new_n32321_, new_n32322_, new_n32323_, new_n32325_,
    new_n32326_, new_n32327_, new_n32328_, new_n32329_, new_n32330_,
    new_n32331_, new_n32332_, new_n32333_, new_n32334_, new_n32335_,
    new_n32336_, new_n32337_, new_n32338_, new_n32340_, new_n32341_,
    new_n32342_, new_n32343_, new_n32344_, new_n32345_, new_n32346_,
    new_n32347_, new_n32348_, new_n32349_, new_n32350_, new_n32351_,
    new_n32352_, new_n32353_, new_n32355_, new_n32356_, new_n32357_,
    new_n32358_, new_n32359_, new_n32360_, new_n32361_, new_n32362_,
    new_n32363_, new_n32364_, new_n32365_, new_n32366_, new_n32367_,
    new_n32368_, new_n32370_, new_n32371_, new_n32372_, new_n32373_,
    new_n32374_, new_n32375_, new_n32376_, new_n32377_, new_n32378_,
    new_n32379_, new_n32380_, new_n32381_, new_n32382_, new_n32383_,
    new_n32385_, new_n32386_, new_n32387_, new_n32388_, new_n32389_,
    new_n32390_, new_n32391_, new_n32392_, new_n32393_, new_n32394_,
    new_n32395_, new_n32396_, new_n32397_, new_n32398_, new_n32400_,
    new_n32401_, new_n32402_, new_n32403_, new_n32404_, new_n32405_,
    new_n32406_, new_n32407_, new_n32408_, new_n32409_, new_n32410_,
    new_n32411_, new_n32412_, new_n32413_, new_n32415_, new_n32416_,
    new_n32417_, new_n32418_, new_n32419_, new_n32420_, new_n32421_,
    new_n32422_, new_n32423_, new_n32424_, new_n32425_, new_n32426_,
    new_n32427_, new_n32428_, new_n32430_, new_n32431_, new_n32432_,
    new_n32433_, new_n32434_, new_n32435_, new_n32436_, new_n32437_,
    new_n32438_, new_n32439_, new_n32440_, new_n32441_, new_n32442_,
    new_n32443_, new_n32445_, new_n32446_, new_n32447_, new_n32448_,
    new_n32449_, new_n32450_, new_n32451_, new_n32452_, new_n32453_,
    new_n32454_, new_n32455_, new_n32456_, new_n32457_, new_n32458_,
    new_n32460_, new_n32461_, new_n32462_, new_n32463_, new_n32464_,
    new_n32465_, new_n32466_, new_n32467_, new_n32468_, new_n32469_,
    new_n32470_, new_n32471_, new_n32472_, new_n32473_, new_n32475_,
    new_n32476_, new_n32477_, new_n32478_, new_n32479_, new_n32480_,
    new_n32481_, new_n32482_, new_n32483_, new_n32484_, new_n32485_,
    new_n32486_, new_n32487_, new_n32488_, new_n32490_, new_n32491_,
    new_n32492_, new_n32493_, new_n32494_, new_n32495_, new_n32496_,
    new_n32497_, new_n32498_, new_n32499_, new_n32500_, new_n32501_,
    new_n32502_, new_n32503_, new_n32505_, new_n32506_, new_n32507_,
    new_n32508_, new_n32509_, new_n32510_, new_n32511_, new_n32512_,
    new_n32513_, new_n32514_, new_n32515_, new_n32516_, new_n32517_,
    new_n32518_, new_n32520_, new_n32521_, new_n32522_, new_n32523_,
    new_n32524_, new_n32525_, new_n32526_, new_n32527_, new_n32528_,
    new_n32529_, new_n32530_, new_n32531_, new_n32532_, new_n32533_,
    new_n32535_, new_n32536_, new_n32537_, new_n32538_, new_n32539_,
    new_n32540_, new_n32541_, new_n32542_, new_n32543_, new_n32544_,
    new_n32545_, new_n32546_, new_n32547_, new_n32548_, new_n32550_,
    new_n32551_, new_n32552_, new_n32553_, new_n32554_, new_n32555_,
    new_n32556_, new_n32557_, new_n32558_, new_n32559_, new_n32560_,
    new_n32561_, new_n32562_, new_n32563_, new_n32565_, new_n32566_,
    new_n32567_, new_n32568_, new_n32569_, new_n32570_, new_n32571_,
    new_n32572_, new_n32573_, new_n32574_, new_n32575_, new_n32576_,
    new_n32577_, new_n32578_, new_n32580_, new_n32581_, new_n32582_,
    new_n32583_, new_n32584_, new_n32585_, new_n32586_, new_n32587_,
    new_n32588_, new_n32589_, new_n32590_, new_n32591_, new_n32592_,
    new_n32593_, new_n32595_, new_n32596_, new_n32597_, new_n32598_,
    new_n32599_, new_n32600_, new_n32601_, new_n32602_, new_n32603_,
    new_n32604_, new_n32605_, new_n32606_, new_n32607_, new_n32608_,
    new_n32610_, new_n32611_, new_n32612_, new_n32613_, new_n32614_,
    new_n32615_, new_n32616_, new_n32617_, new_n32618_, new_n32619_,
    new_n32620_, new_n32621_, new_n32622_, new_n32623_, new_n32625_,
    new_n32626_, new_n32627_, new_n32628_, new_n32629_, new_n32630_,
    new_n32631_, new_n32632_, new_n32633_, new_n32634_, new_n32635_,
    new_n32636_, new_n32637_, new_n32638_, new_n32640_, new_n32641_,
    new_n32642_, new_n32643_, new_n32644_, new_n32645_, new_n32646_,
    new_n32647_, new_n32648_, new_n32649_, new_n32650_, new_n32651_,
    new_n32652_, new_n32653_, new_n32655_, new_n32656_, new_n32657_,
    new_n32658_, new_n32659_, new_n32660_, new_n32661_, new_n32662_,
    new_n32663_, new_n32664_, new_n32665_, new_n32666_, new_n32667_,
    new_n32668_, new_n32670_, new_n32671_, new_n32672_, new_n32673_,
    new_n32674_, new_n32675_, new_n32676_, new_n32677_, new_n32678_,
    new_n32679_, new_n32680_, new_n32681_, new_n32682_, new_n32683_,
    new_n32685_, new_n32686_, new_n32687_, new_n32688_, new_n32689_,
    new_n32690_, new_n32691_, new_n32692_, new_n32693_, new_n32694_,
    new_n32695_, new_n32696_, new_n32697_, new_n32698_, new_n32700_,
    new_n32701_, new_n32702_, new_n32703_, new_n32704_, new_n32705_,
    new_n32706_, new_n32707_, new_n32708_, new_n32709_, new_n32710_,
    new_n32711_, new_n32712_, new_n32713_, new_n32715_, new_n32716_,
    new_n32717_, new_n32718_, new_n32719_, new_n32720_, new_n32721_,
    new_n32722_, new_n32723_, new_n32724_, new_n32725_, new_n32726_,
    new_n32727_, new_n32728_, new_n33366_, new_n33367_, new_n33368_,
    new_n33369_, new_n33370_, new_n33371_, new_n33372_, new_n33373_,
    new_n33374_, new_n33375_, new_n33376_, new_n33377_, new_n33378_,
    new_n33379_, new_n33380_, new_n33381_, new_n33382_, new_n33383_,
    new_n33384_, new_n33385_, new_n33386_, new_n33387_, new_n33388_,
    new_n33389_, new_n33390_, new_n33391_, new_n33392_, new_n33393_,
    new_n33394_, new_n33395_, new_n33396_, new_n33397_, new_n33398_,
    new_n33399_, new_n33400_, new_n33401_, new_n33402_, new_n33403_,
    new_n33404_, new_n33405_, new_n33406_, new_n33407_, new_n33408_,
    new_n33409_, new_n33410_, new_n33411_, new_n33412_, new_n33413_,
    new_n33414_, new_n33415_, new_n33416_, new_n33417_, new_n33418_,
    new_n33419_, new_n33420_, new_n33421_, new_n33422_, new_n33423_,
    new_n33424_, new_n33425_, new_n33426_, new_n33427_, new_n33428_,
    new_n33429_, new_n33430_, new_n33431_, new_n33432_, new_n33433_,
    new_n33434_, new_n33435_, new_n33436_, new_n33437_, new_n33438_,
    new_n33439_, new_n33440_, new_n33441_, new_n33442_, new_n33443_,
    new_n33444_, new_n33445_, new_n33446_, new_n33447_, new_n33448_,
    new_n33449_, new_n33450_, new_n33451_, new_n33452_, new_n33453_,
    new_n33454_, new_n33455_, new_n33456_, new_n33457_, new_n33458_,
    new_n33459_, new_n33460_, new_n33461_, new_n33462_, new_n33463_,
    new_n33464_, new_n33465_, new_n33466_, new_n33467_, new_n33468_,
    new_n33469_, new_n33470_, new_n33471_, new_n33472_, new_n33473_,
    new_n33474_, new_n33475_, new_n33476_, new_n33477_, new_n33478_,
    new_n33479_, new_n33480_, new_n33481_, new_n33482_, new_n33483_,
    new_n33484_, new_n33485_, new_n33486_, new_n33487_, new_n33488_,
    new_n33489_, new_n33490_, new_n33491_, new_n33492_, new_n33493_,
    new_n33494_, new_n33495_, new_n33496_, new_n33497_, new_n33498_,
    new_n33499_, new_n33500_, new_n33501_, new_n33502_, new_n33503_,
    new_n33504_, new_n33505_, new_n33506_, new_n33507_, new_n33508_,
    new_n33509_, new_n33510_, new_n33511_, new_n33512_, new_n33513_,
    new_n33514_, new_n33515_, new_n33516_, new_n33517_, new_n33518_,
    new_n33519_, new_n33520_, new_n33521_, new_n33522_, new_n33523_,
    new_n33524_, new_n33525_, new_n33526_, new_n33527_, new_n33528_,
    new_n33529_, new_n33530_, new_n33531_, new_n33532_, new_n33533_,
    new_n33534_, new_n33535_, new_n33536_, new_n33537_, new_n33538_,
    new_n33539_, new_n33540_, new_n33541_, new_n33542_, new_n33543_,
    new_n33544_, new_n33545_, new_n33546_, new_n33547_, new_n33548_,
    new_n33549_, new_n33550_, new_n33551_, new_n33552_, new_n33553_,
    new_n33554_, new_n33555_, new_n33556_, new_n33557_, new_n33558_,
    new_n33559_, new_n33560_, new_n33561_, new_n33562_, new_n33563_,
    new_n33564_, new_n33565_, new_n33566_, new_n33567_, new_n33568_,
    new_n33569_, new_n33570_, new_n33571_, new_n33572_, new_n33573_,
    new_n33574_, new_n33575_, new_n33576_, new_n33577_, new_n33578_,
    new_n33579_, new_n33580_, new_n33581_, new_n33582_, new_n33583_,
    new_n33584_, new_n33585_, new_n33586_, new_n33587_, new_n33588_,
    new_n33589_, new_n33590_, new_n33591_, new_n33592_, new_n33593_,
    new_n33594_, new_n33595_, new_n33596_, new_n33597_, new_n33598_,
    new_n33599_, new_n33600_, new_n33601_, new_n33602_, new_n33603_,
    new_n33604_, new_n33605_, new_n33606_, new_n33607_, new_n33608_,
    new_n33609_, new_n33610_, new_n33611_, new_n33612_, new_n33613_,
    new_n33614_, new_n33615_, new_n33616_, new_n33617_, new_n33618_,
    new_n33619_, new_n33620_, new_n33621_, new_n33622_, new_n33623_,
    new_n33624_, new_n33625_, new_n33626_, new_n33627_, new_n33628_,
    new_n33629_, new_n33630_, new_n33631_, new_n33632_, new_n33633_,
    new_n33634_, new_n33635_, new_n33636_, new_n33637_, new_n33638_,
    new_n33639_, new_n33640_, new_n33641_, new_n33642_, new_n33643_,
    new_n33644_, new_n33645_, new_n33646_, new_n33647_, new_n33648_,
    new_n33649_, new_n33650_, new_n33651_, new_n33652_, new_n33653_,
    new_n33654_, new_n33655_, new_n33656_, new_n33657_, new_n33658_,
    new_n33659_, new_n33660_, new_n33661_, new_n33662_, new_n33663_,
    new_n33664_, new_n33665_, new_n33666_, new_n33667_, new_n33668_,
    new_n33669_, new_n33670_, new_n33671_, new_n33672_, new_n33673_,
    new_n33674_, new_n33675_, new_n33676_, new_n33677_, new_n33678_,
    new_n33679_, new_n33680_, new_n33681_, new_n33682_, new_n33683_,
    new_n33684_, new_n33685_, new_n33686_, new_n33687_, new_n33688_,
    new_n33689_, new_n33690_, new_n33691_, new_n33692_, new_n33693_,
    new_n33694_, new_n33695_, new_n33696_, new_n33697_, new_n33698_,
    new_n33699_, new_n33700_, new_n33702_, new_n33703_, new_n33704_,
    new_n33705_, new_n33706_, new_n33707_, new_n33708_, new_n33709_,
    new_n33710_, new_n33711_, new_n33712_, new_n33713_, new_n33714_,
    new_n33715_, new_n33716_, new_n33717_, new_n33718_, new_n33719_,
    new_n33720_, new_n33721_, new_n33722_, new_n33723_, new_n33724_,
    new_n33725_, new_n33726_, new_n33727_, new_n33728_, new_n33729_,
    new_n33730_, new_n33731_, new_n33732_, new_n33733_, new_n33734_,
    new_n33735_, new_n33736_, new_n33737_, new_n33738_, new_n33739_,
    new_n33740_, new_n33741_, new_n33742_, new_n33743_, new_n33744_,
    new_n33745_, new_n33746_, new_n33747_, new_n33748_, new_n33749_,
    new_n33750_, new_n33751_, new_n33752_, new_n33753_, new_n33754_,
    new_n33755_, new_n33756_, new_n33757_, new_n33758_, new_n33759_,
    new_n33760_, new_n33761_, new_n33762_, new_n33763_, new_n33764_,
    new_n33765_, new_n33766_, new_n33767_, new_n33768_, new_n33769_,
    new_n33770_, new_n33771_, new_n33772_, new_n33773_, new_n33774_,
    new_n33775_, new_n33776_, new_n33777_, new_n33778_, new_n33779_,
    new_n33780_, new_n33781_, new_n33782_, new_n33783_, new_n33784_,
    new_n33785_, new_n33786_, new_n33787_, new_n33788_, new_n33789_,
    new_n33790_, new_n33791_, new_n33792_, new_n33793_, new_n33794_,
    new_n33795_, new_n33796_, new_n33797_, new_n33798_, new_n33799_,
    new_n33800_, new_n33801_, new_n33802_, new_n33803_, new_n33804_,
    new_n33805_, new_n33806_, new_n33807_, new_n33808_, new_n33809_,
    new_n33810_, new_n33811_, new_n33812_, new_n33813_, new_n33814_,
    new_n33815_, new_n33816_, new_n33817_, new_n33818_, new_n33819_,
    new_n33820_, new_n33821_, new_n33822_, new_n33823_, new_n33824_,
    new_n33825_, new_n33826_, new_n33827_, new_n33828_, new_n33829_,
    new_n33830_, new_n33831_, new_n33832_, new_n33833_, new_n33834_,
    new_n33835_, new_n33836_, new_n33837_, new_n33838_, new_n33839_,
    new_n33840_, new_n33841_, new_n33842_, new_n33843_, new_n33844_,
    new_n33845_, new_n33846_, new_n33847_, new_n33848_, new_n33849_,
    new_n33850_, new_n33851_, new_n33852_, new_n33853_, new_n33854_,
    new_n33855_, new_n33856_, new_n33857_, new_n33858_, new_n33859_,
    new_n33860_, new_n33861_, new_n33862_, new_n33863_, new_n33864_,
    new_n33865_, new_n33866_, new_n33867_, new_n33868_, new_n33869_,
    new_n33870_, new_n33871_, new_n33872_, new_n33873_, new_n33874_,
    new_n33875_, new_n33876_, new_n33877_, new_n33878_, new_n33879_,
    new_n33880_, new_n33881_, new_n33882_, new_n33883_, new_n33884_,
    new_n33885_, new_n33886_, new_n33887_, new_n33888_, new_n33889_,
    new_n33890_, new_n33891_, new_n33892_, new_n33893_, new_n33894_,
    new_n33895_, new_n33896_, new_n33897_, new_n33898_, new_n33899_,
    new_n33900_, new_n33901_, new_n33902_, new_n33903_, new_n33904_,
    new_n33905_, new_n33906_, new_n33907_, new_n33908_, new_n33909_,
    new_n33910_, new_n33911_, new_n33912_, new_n33913_, new_n33914_,
    new_n33915_, new_n33916_, new_n33917_, new_n33918_, new_n33919_,
    new_n33920_, new_n33921_, new_n33922_, new_n33923_, new_n33924_,
    new_n33925_, new_n33926_, new_n33927_, new_n33928_, new_n33929_,
    new_n33930_, new_n33931_, new_n33932_, new_n33933_, new_n33934_,
    new_n33935_, new_n33936_, new_n33937_, new_n33938_, new_n33939_,
    new_n33940_, new_n33941_, new_n33942_, new_n33943_, new_n33944_,
    new_n33945_, new_n33946_, new_n33947_, new_n33948_, new_n33949_,
    new_n33950_, new_n33951_, new_n33952_, new_n33953_, new_n33954_,
    new_n33955_, new_n33956_, new_n33957_, new_n33958_, new_n33959_,
    new_n33960_, new_n33961_, new_n33962_, new_n33963_, new_n33964_,
    new_n33965_, new_n33966_, new_n33967_, new_n33968_, new_n33969_,
    new_n33970_, new_n33971_, new_n33972_, new_n33973_, new_n33974_,
    new_n33975_, new_n33976_, new_n33977_, new_n33978_, new_n33979_,
    new_n33980_, new_n33981_, new_n33982_, new_n33983_, new_n33984_,
    new_n33985_, new_n33986_, new_n33987_, new_n33988_, new_n33989_,
    new_n33990_, new_n33991_, new_n33992_, new_n33993_, new_n33994_,
    new_n33995_, new_n33996_, new_n33997_, new_n33998_, new_n33999_,
    new_n34000_, new_n34001_, new_n34002_, new_n34003_, new_n34004_,
    new_n34005_, new_n34006_, new_n34007_, new_n34008_, new_n34009_,
    new_n34010_, new_n34011_, new_n34012_, new_n34013_, new_n34014_,
    new_n34015_, new_n34016_, new_n34017_, new_n34018_, new_n34019_,
    new_n34020_, new_n34021_, new_n34022_, new_n34023_, new_n34024_,
    new_n34025_, new_n34026_, new_n34027_, new_n34029_, new_n34030_,
    new_n34031_, new_n34032_, new_n34033_, new_n34034_, new_n34035_,
    new_n34036_, new_n34037_, new_n34038_, new_n34039_, new_n34040_,
    new_n34041_, new_n34042_, new_n34043_, new_n34044_, new_n34045_,
    new_n34046_, new_n34047_, new_n34048_, new_n34049_, new_n34050_,
    new_n34051_, new_n34052_, new_n34053_, new_n34054_, new_n34055_,
    new_n34056_, new_n34057_, new_n34058_, new_n34059_, new_n34060_,
    new_n34061_, new_n34062_, new_n34063_, new_n34064_, new_n34065_,
    new_n34066_, new_n34067_, new_n34068_, new_n34069_, new_n34070_,
    new_n34071_, new_n34072_, new_n34073_, new_n34074_, new_n34075_,
    new_n34076_, new_n34077_, new_n34078_, new_n34079_, new_n34080_,
    new_n34081_, new_n34082_, new_n34083_, new_n34084_, new_n34085_,
    new_n34086_, new_n34087_, new_n34088_, new_n34089_, new_n34090_,
    new_n34091_, new_n34092_, new_n34093_, new_n34094_, new_n34095_,
    new_n34096_, new_n34097_, new_n34098_, new_n34099_, new_n34100_,
    new_n34101_, new_n34102_, new_n34103_, new_n34104_, new_n34105_,
    new_n34106_, new_n34107_, new_n34108_, new_n34109_, new_n34110_,
    new_n34111_, new_n34112_, new_n34113_, new_n34114_, new_n34115_,
    new_n34116_, new_n34117_, new_n34118_, new_n34119_, new_n34120_,
    new_n34121_, new_n34122_, new_n34123_, new_n34124_, new_n34125_,
    new_n34126_, new_n34127_, new_n34128_, new_n34129_, new_n34130_,
    new_n34131_, new_n34132_, new_n34133_, new_n34134_, new_n34135_,
    new_n34136_, new_n34137_, new_n34138_, new_n34139_, new_n34140_,
    new_n34141_, new_n34142_, new_n34143_, new_n34144_, new_n34145_,
    new_n34146_, new_n34147_, new_n34148_, new_n34149_, new_n34150_,
    new_n34151_, new_n34152_, new_n34153_, new_n34154_, new_n34155_,
    new_n34156_, new_n34157_, new_n34158_, new_n34159_, new_n34160_,
    new_n34161_, new_n34162_, new_n34163_, new_n34164_, new_n34165_,
    new_n34166_, new_n34167_, new_n34168_, new_n34169_, new_n34170_,
    new_n34171_, new_n34172_, new_n34173_, new_n34174_, new_n34175_,
    new_n34176_, new_n34177_, new_n34178_, new_n34179_, new_n34180_,
    new_n34181_, new_n34182_, new_n34183_, new_n34184_, new_n34185_,
    new_n34186_, new_n34187_, new_n34188_, new_n34189_, new_n34190_,
    new_n34191_, new_n34192_, new_n34193_, new_n34194_, new_n34195_,
    new_n34196_, new_n34197_, new_n34198_, new_n34199_, new_n34200_,
    new_n34201_, new_n34202_, new_n34203_, new_n34204_, new_n34205_,
    new_n34206_, new_n34207_, new_n34208_, new_n34209_, new_n34210_,
    new_n34211_, new_n34212_, new_n34213_, new_n34214_, new_n34215_,
    new_n34216_, new_n34217_, new_n34218_, new_n34219_, new_n34220_,
    new_n34221_, new_n34222_, new_n34223_, new_n34224_, new_n34225_,
    new_n34226_, new_n34227_, new_n34228_, new_n34229_, new_n34230_,
    new_n34231_, new_n34232_, new_n34233_, new_n34234_, new_n34235_,
    new_n34236_, new_n34237_, new_n34238_, new_n34239_, new_n34240_,
    new_n34241_, new_n34242_, new_n34243_, new_n34244_, new_n34245_,
    new_n34246_, new_n34247_, new_n34248_, new_n34249_, new_n34250_,
    new_n34251_, new_n34252_, new_n34253_, new_n34254_, new_n34255_,
    new_n34256_, new_n34257_, new_n34258_, new_n34259_, new_n34260_,
    new_n34261_, new_n34262_, new_n34263_, new_n34264_, new_n34265_,
    new_n34266_, new_n34267_, new_n34268_, new_n34269_, new_n34270_,
    new_n34271_, new_n34272_, new_n34273_, new_n34274_, new_n34275_,
    new_n34276_, new_n34277_, new_n34278_, new_n34279_, new_n34280_,
    new_n34281_, new_n34282_, new_n34283_, new_n34284_, new_n34285_,
    new_n34286_, new_n34287_, new_n34288_, new_n34289_, new_n34290_,
    new_n34291_, new_n34292_, new_n34293_, new_n34294_, new_n34295_,
    new_n34296_, new_n34297_, new_n34298_, new_n34299_, new_n34300_,
    new_n34301_, new_n34302_, new_n34303_, new_n34304_, new_n34305_,
    new_n34306_, new_n34307_, new_n34308_, new_n34309_, new_n34310_,
    new_n34311_, new_n34312_, new_n34313_, new_n34314_, new_n34315_,
    new_n34316_, new_n34317_, new_n34318_, new_n34319_, new_n34320_,
    new_n34321_, new_n34322_, new_n34323_, new_n34324_, new_n34325_,
    new_n34326_, new_n34327_, new_n34328_, new_n34329_, new_n34330_,
    new_n34331_, new_n34332_, new_n34333_, new_n34334_, new_n34335_,
    new_n34336_, new_n34337_, new_n34338_, new_n34339_, new_n34340_,
    new_n34341_, new_n34342_, new_n34343_, new_n34344_, new_n34345_,
    new_n34346_, new_n34347_, new_n34348_, new_n34349_, new_n34350_,
    new_n34351_, new_n34352_, new_n34353_, new_n34354_, new_n34356_,
    new_n34357_, new_n34358_, new_n34359_, new_n34360_, new_n34361_,
    new_n34362_, new_n34363_, new_n34364_, new_n34365_, new_n34366_,
    new_n34367_, new_n34368_, new_n34369_, new_n34370_, new_n34371_,
    new_n34372_, new_n34373_, new_n34374_, new_n34375_, new_n34376_,
    new_n34377_, new_n34378_, new_n34379_, new_n34380_, new_n34381_,
    new_n34382_, new_n34383_, new_n34384_, new_n34385_, new_n34386_,
    new_n34387_, new_n34388_, new_n34389_, new_n34390_, new_n34391_,
    new_n34392_, new_n34393_, new_n34394_, new_n34395_, new_n34396_,
    new_n34397_, new_n34398_, new_n34399_, new_n34400_, new_n34401_,
    new_n34402_, new_n34403_, new_n34404_, new_n34405_, new_n34406_,
    new_n34407_, new_n34408_, new_n34409_, new_n34410_, new_n34411_,
    new_n34412_, new_n34413_, new_n34414_, new_n34415_, new_n34416_,
    new_n34417_, new_n34418_, new_n34419_, new_n34420_, new_n34421_,
    new_n34422_, new_n34423_, new_n34424_, new_n34425_, new_n34426_,
    new_n34427_, new_n34428_, new_n34429_, new_n34430_, new_n34431_,
    new_n34432_, new_n34433_, new_n34434_, new_n34435_, new_n34436_,
    new_n34437_, new_n34438_, new_n34439_, new_n34440_, new_n34441_,
    new_n34442_, new_n34443_, new_n34444_, new_n34445_, new_n34446_,
    new_n34447_, new_n34448_, new_n34449_, new_n34450_, new_n34451_,
    new_n34452_, new_n34453_, new_n34454_, new_n34455_, new_n34456_,
    new_n34457_, new_n34458_, new_n34459_, new_n34460_, new_n34461_,
    new_n34462_, new_n34463_, new_n34464_, new_n34465_, new_n34466_,
    new_n34467_, new_n34468_, new_n34469_, new_n34470_, new_n34471_,
    new_n34472_, new_n34473_, new_n34474_, new_n34475_, new_n34476_,
    new_n34477_, new_n34478_, new_n34479_, new_n34480_, new_n34481_,
    new_n34482_, new_n34483_, new_n34484_, new_n34485_, new_n34486_,
    new_n34487_, new_n34488_, new_n34489_, new_n34490_, new_n34491_,
    new_n34492_, new_n34493_, new_n34494_, new_n34495_, new_n34496_,
    new_n34497_, new_n34498_, new_n34499_, new_n34500_, new_n34501_,
    new_n34502_, new_n34503_, new_n34504_, new_n34505_, new_n34506_,
    new_n34507_, new_n34508_, new_n34509_, new_n34510_, new_n34511_,
    new_n34512_, new_n34513_, new_n34514_, new_n34515_, new_n34516_,
    new_n34517_, new_n34518_, new_n34519_, new_n34520_, new_n34521_,
    new_n34522_, new_n34523_, new_n34524_, new_n34525_, new_n34526_,
    new_n34527_, new_n34528_, new_n34529_, new_n34530_, new_n34531_,
    new_n34532_, new_n34533_, new_n34534_, new_n34535_, new_n34536_,
    new_n34537_, new_n34538_, new_n34539_, new_n34540_, new_n34541_,
    new_n34542_, new_n34543_, new_n34544_, new_n34545_, new_n34546_,
    new_n34547_, new_n34548_, new_n34549_, new_n34550_, new_n34551_,
    new_n34552_, new_n34553_, new_n34554_, new_n34555_, new_n34556_,
    new_n34557_, new_n34558_, new_n34559_, new_n34560_, new_n34561_,
    new_n34562_, new_n34563_, new_n34564_, new_n34565_, new_n34566_,
    new_n34567_, new_n34568_, new_n34569_, new_n34570_, new_n34571_,
    new_n34572_, new_n34573_, new_n34574_, new_n34575_, new_n34576_,
    new_n34577_, new_n34578_, new_n34579_, new_n34580_, new_n34581_,
    new_n34582_, new_n34583_, new_n34584_, new_n34585_, new_n34586_,
    new_n34587_, new_n34588_, new_n34589_, new_n34590_, new_n34591_,
    new_n34592_, new_n34593_, new_n34594_, new_n34595_, new_n34596_,
    new_n34597_, new_n34598_, new_n34599_, new_n34600_, new_n34601_,
    new_n34602_, new_n34603_, new_n34604_, new_n34605_, new_n34606_,
    new_n34607_, new_n34608_, new_n34609_, new_n34610_, new_n34611_,
    new_n34612_, new_n34613_, new_n34614_, new_n34615_, new_n34616_,
    new_n34617_, new_n34618_, new_n34619_, new_n34620_, new_n34621_,
    new_n34622_, new_n34623_, new_n34624_, new_n34625_, new_n34626_,
    new_n34627_, new_n34628_, new_n34629_, new_n34630_, new_n34631_,
    new_n34632_, new_n34633_, new_n34634_, new_n34635_, new_n34636_,
    new_n34637_, new_n34638_, new_n34639_, new_n34640_, new_n34641_,
    new_n34642_, new_n34643_, new_n34644_, new_n34645_, new_n34646_,
    new_n34647_, new_n34648_, new_n34649_, new_n34650_, new_n34651_,
    new_n34652_, new_n34653_, new_n34654_, new_n34655_, new_n34656_,
    new_n34657_, new_n34658_, new_n34659_, new_n34660_, new_n34661_,
    new_n34662_, new_n34663_, new_n34664_, new_n34665_, new_n34666_,
    new_n34667_, new_n34668_, new_n34669_, new_n34670_, new_n34671_,
    new_n34672_, new_n34673_, new_n34674_, new_n34675_, new_n34676_,
    new_n34677_, new_n34678_, new_n34679_, new_n34680_, new_n34681_,
    new_n34682_, new_n34683_, new_n34684_, new_n34685_, new_n34687_,
    new_n34688_, new_n34689_, new_n34690_, new_n34691_, new_n34692_,
    new_n34693_, new_n34694_, new_n34695_, new_n34696_, new_n34697_,
    new_n34699_, new_n34700_, new_n34701_, new_n34702_, new_n34703_,
    new_n34704_, new_n34705_, new_n34706_, new_n34707_, new_n34708_,
    new_n34709_, new_n34710_, new_n34711_, new_n34712_, new_n34713_,
    new_n34715_, new_n34716_, new_n34717_, new_n34718_, new_n34719_,
    new_n34721_, new_n34722_, new_n34724_, new_n34725_, new_n34727_,
    new_n34728_, new_n34729_, new_n34730_, new_n34731_, new_n34732_,
    new_n34734_, new_n34735_, new_n34737_, new_n34738_, new_n34740_,
    new_n34741_, new_n34743_, new_n34744_, new_n34746_, new_n34747_,
    new_n34749_, new_n34750_, new_n34752_, new_n34753_, new_n34755_,
    new_n34756_, new_n34758_, new_n34759_, new_n34761_, new_n34762_,
    new_n34764_, new_n34765_, new_n34767_, new_n34768_, new_n34770_,
    new_n34771_, new_n34773_, new_n34774_, new_n34776_, new_n34777_,
    new_n34779_, new_n34780_, new_n34782_, new_n34783_, new_n34785_,
    new_n34786_, new_n34788_, new_n34789_, new_n34791_, new_n34792_,
    new_n34794_, new_n34795_, new_n34797_, new_n34798_, new_n34800_,
    new_n34801_, new_n34803_, new_n34804_, new_n34806_, new_n34807_,
    new_n34809_, new_n34810_, new_n34812_, new_n34813_, new_n34815_,
    new_n34816_, new_n34818_, new_n34819_, new_n34821_, new_n34822_,
    new_n34824_, new_n34825_, new_n34827_, new_n34828_, new_n34829_,
    new_n34831_, new_n34832_, new_n34834_, new_n34835_, new_n34837_,
    new_n34838_, new_n34840_, new_n34841_, new_n34843_, new_n34844_,
    new_n34846_, new_n34847_, new_n34849_, new_n34850_, new_n34852_,
    new_n34853_, new_n34855_, new_n34856_, new_n34858_, new_n34859_,
    new_n34861_, new_n34862_, new_n34864_, new_n34865_, new_n34867_,
    new_n34868_, new_n34870_, new_n34871_, new_n34873_, new_n34874_,
    new_n34876_, new_n34877_, new_n34879_, new_n34880_, new_n34882_,
    new_n34883_, new_n34885_, new_n34886_, new_n34888_, new_n34889_,
    new_n34891_, new_n34892_, new_n34894_, new_n34895_, new_n34897_,
    new_n34898_, new_n34900_, new_n34901_, new_n34903_, new_n34904_,
    new_n34906_, new_n34907_, new_n34909_, new_n34910_, new_n34912_,
    new_n34913_, new_n34915_, new_n34916_, new_n34918_, new_n34919_,
    new_n34921_, new_n34922_, new_n34925_, new_n34926_, new_n34930_,
    new_n34931_, new_n34933_, new_n34934_, new_n34936_, new_n34937_,
    new_n34939_, new_n34940_, new_n34941_, new_n34943_, new_n34944_,
    new_n34945_, new_n34946_, new_n34947_, new_n34949_, new_n34950_,
    new_n34951_, new_n34953_, new_n34954_, new_n34955_, new_n34957_,
    new_n34958_, new_n34959_, new_n34960_, new_n34962_, new_n34963_,
    new_n34965_, new_n34966_, new_n34968_, new_n34969_, new_n34971_,
    new_n34972_, new_n34973_, new_n34975_, new_n34976_, new_n34978_,
    new_n34979_, new_n34981_, new_n34982_, new_n34984_, new_n34985_,
    new_n34986_, new_n34988_, new_n34989_, new_n34991_, new_n34992_,
    new_n34994_, new_n34995_, new_n34997_, new_n34998_, new_n34999_,
    new_n35001_, new_n35003_, new_n35005_, new_n35007_, new_n35009_,
    new_n35011_, new_n35013_, new_n35015_, new_n35017_, new_n35019_,
    new_n35021_, new_n35023_, new_n35025_, new_n35027_, new_n35029_,
    new_n35031_, new_n35032_, new_n35034_, new_n35035_, new_n35036_,
    new_n35037_, new_n35038_, new_n35040_, new_n35041_, new_n35042_,
    new_n35043_, new_n35044_, new_n35045_, new_n35046_, new_n35047_,
    new_n35048_, new_n35049_, new_n35050_, new_n35051_, new_n35052_,
    new_n35053_, new_n35055_, new_n35056_, new_n35057_, new_n35058_,
    new_n35059_, new_n35060_, new_n35061_, new_n35062_, new_n35063_,
    new_n35064_, new_n35065_, new_n35066_, new_n35067_, new_n35068_,
    new_n35069_, new_n35070_, new_n35071_, new_n35072_, new_n35073_,
    new_n35074_, new_n35075_, new_n35076_, new_n35078_, new_n35079_,
    new_n35080_, new_n35081_, new_n35082_, new_n35084_, new_n35085_,
    new_n35086_, new_n35087_, new_n35088_, new_n35089_, new_n35090_,
    new_n35091_, new_n35092_, new_n35093_, new_n35094_, new_n35095_,
    new_n35096_, new_n35097_, new_n35098_, new_n35099_, new_n35100_,
    new_n35101_, new_n35102_, new_n35104_, new_n35105_, new_n35106_,
    new_n35107_, new_n35108_, new_n35109_, new_n35110_, new_n35112_,
    new_n35113_, new_n35114_, new_n35115_, new_n35116_, new_n35117_,
    new_n35118_, new_n35119_, new_n35120_, new_n35121_, new_n35122_,
    new_n35123_, new_n35124_, new_n35125_, new_n35126_, new_n35127_,
    new_n35128_, new_n35129_, new_n35130_, new_n35131_, new_n35133_,
    new_n35134_, new_n35135_, new_n35136_, new_n35137_, new_n35138_,
    new_n35139_, new_n35141_, new_n35142_, new_n35143_, new_n35144_,
    new_n35145_, new_n35146_, new_n35147_, new_n35148_, new_n35149_,
    new_n35150_, new_n35151_, new_n35152_, new_n35153_, new_n35154_,
    new_n35155_, new_n35156_, new_n35157_, new_n35158_, new_n35159_,
    new_n35160_, new_n35161_, new_n35162_, new_n35164_, new_n35165_,
    new_n35166_, new_n35167_, new_n35168_, new_n35169_, new_n35171_,
    new_n35172_, new_n35173_, new_n35174_, new_n35175_, new_n35176_,
    new_n35177_, new_n35178_, new_n35179_, new_n35180_, new_n35181_,
    new_n35182_, new_n35183_, new_n35184_, new_n35185_, new_n35186_,
    new_n35187_, new_n35188_, new_n35189_, new_n35190_, new_n35192_,
    new_n35193_, new_n35194_, new_n35195_, new_n35196_, new_n35197_,
    new_n35199_, new_n35200_, new_n35201_, new_n35202_, new_n35203_,
    new_n35204_, new_n35205_, new_n35206_, new_n35207_, new_n35208_,
    new_n35209_, new_n35210_, new_n35211_, new_n35212_, new_n35213_,
    new_n35214_, new_n35215_, new_n35216_, new_n35217_, new_n35218_,
    new_n35220_, new_n35221_, new_n35222_, new_n35223_, new_n35224_,
    new_n35225_, new_n35226_, new_n35227_, new_n35228_, new_n35229_,
    new_n35230_, new_n35231_, new_n35232_, new_n35234_, new_n35235_,
    new_n35236_, new_n35237_, new_n35238_, new_n35239_, new_n35240_,
    new_n35241_, new_n35242_, new_n35243_, new_n35244_, new_n35245_,
    new_n35246_, new_n35247_, new_n35248_, new_n35249_, new_n35250_,
    new_n35252_, new_n35253_, new_n35254_, new_n35255_, new_n35256_,
    new_n35257_, new_n35258_, new_n35259_, new_n35260_, new_n35261_,
    new_n35262_, new_n35263_, new_n35264_, new_n35265_, new_n35266_,
    new_n35267_, new_n35268_, new_n35269_, new_n35270_, new_n35271_,
    new_n35272_, new_n35273_, new_n35275_, new_n35276_, new_n35277_,
    new_n35278_, new_n35279_, new_n35280_, new_n35281_, new_n35282_,
    new_n35283_, new_n35284_, new_n35285_, new_n35286_, new_n35287_,
    new_n35288_, new_n35290_, new_n35291_, new_n35292_, new_n35293_,
    new_n35294_, new_n35295_, new_n35296_, new_n35297_, new_n35298_,
    new_n35299_, new_n35300_, new_n35301_, new_n35302_, new_n35303_,
    new_n35305_, new_n35306_, new_n35307_, new_n35308_, new_n35309_,
    new_n35310_, new_n35311_, new_n35312_, new_n35313_, new_n35314_,
    new_n35315_, new_n35316_, new_n35317_, new_n35318_, new_n35320_,
    new_n35321_, new_n35322_, new_n35323_, new_n35324_, new_n35325_,
    new_n35326_, new_n35327_, new_n35328_, new_n35329_, new_n35330_,
    new_n35331_, new_n35332_, new_n35333_, new_n35334_, new_n35335_,
    new_n35336_, new_n35338_, new_n35339_, new_n35340_, new_n35341_,
    new_n35342_, new_n35343_, new_n35344_, new_n35345_, new_n35346_,
    new_n35347_, new_n35348_, new_n35349_, new_n35350_, new_n35351_,
    new_n35353_, new_n35354_, new_n35355_, new_n35356_, new_n35357_,
    new_n35358_, new_n35359_, new_n35360_, new_n35361_, new_n35362_,
    new_n35363_, new_n35364_, new_n35365_, new_n35366_, new_n35367_,
    new_n35368_, new_n35370_, new_n35371_, new_n35372_, new_n35373_,
    new_n35374_, new_n35375_, new_n35376_, new_n35377_, new_n35378_,
    new_n35379_, new_n35380_, new_n35381_, new_n35382_, new_n35383_,
    new_n35384_, new_n35385_, new_n35387_, new_n35388_, new_n35389_,
    new_n35390_, new_n35391_, new_n35392_, new_n35393_, new_n35394_,
    new_n35395_, new_n35396_, new_n35397_, new_n35398_, new_n35400_,
    new_n35401_, new_n35402_, new_n35403_, new_n35404_, new_n35405_,
    new_n35406_, new_n35407_, new_n35408_, new_n35410_, new_n35411_,
    new_n35412_, new_n35413_, new_n35414_, new_n35415_, new_n35416_,
    new_n35417_, new_n35418_, new_n35419_, new_n35420_, new_n35422_,
    new_n35423_, new_n35424_, new_n35425_, new_n35426_, new_n35427_,
    new_n35428_, new_n35429_, new_n35430_, new_n35431_, new_n35432_,
    new_n35434_, new_n35435_, new_n35436_, new_n35437_, new_n35438_,
    new_n35439_, new_n35440_, new_n35441_, new_n35442_, new_n35444_,
    new_n35445_, new_n35446_, new_n35447_, new_n35448_, new_n35449_,
    new_n35450_, new_n35451_, new_n35452_, new_n35454_, new_n35455_,
    new_n35456_, new_n35457_, new_n35458_, new_n35459_, new_n35460_,
    new_n35461_, new_n35462_, new_n35463_, new_n35464_, new_n35465_,
    new_n35466_, new_n35468_, new_n35469_, new_n35470_, new_n35471_,
    new_n35472_, new_n35473_, new_n35474_, new_n35475_, new_n35476_,
    new_n35478_, new_n35479_, new_n35480_, new_n35481_, new_n35482_,
    new_n35483_, new_n35484_, new_n35485_, new_n35486_, new_n35488_,
    new_n35489_, new_n35490_, new_n35491_, new_n35492_, new_n35493_,
    new_n35494_, new_n35495_, new_n35496_, new_n35498_, new_n35499_,
    new_n35500_, new_n35501_, new_n35502_, new_n35503_, new_n35504_,
    new_n35505_, new_n35506_, new_n35508_, new_n35509_, new_n35510_,
    new_n35511_, new_n35512_, new_n35513_, new_n35514_, new_n35515_,
    new_n35516_, new_n35518_, new_n35519_, new_n35520_, new_n35521_,
    new_n35522_, new_n35523_, new_n35524_, new_n35525_, new_n35526_,
    new_n35527_, new_n35528_, new_n35529_, new_n35530_, new_n35531_,
    new_n35533_, new_n35534_, new_n35535_, new_n35536_, new_n35537_,
    new_n35538_, new_n35539_, new_n35540_, new_n35541_, new_n35542_,
    new_n35543_, new_n35544_, new_n35545_, new_n35546_, new_n35547_,
    new_n35548_, new_n35550_, new_n35551_, new_n35552_, new_n35553_,
    new_n35554_, new_n35555_, new_n35556_, new_n35557_, new_n35558_,
    new_n35559_, new_n35560_, new_n35561_, new_n35562_, new_n35563_,
    new_n35565_, new_n35566_, new_n35567_, new_n35568_, new_n35569_,
    new_n35570_, new_n35571_, new_n35572_, new_n35573_, new_n35574_,
    new_n35575_, new_n35576_, new_n35577_, new_n35578_, new_n35579_,
    new_n35580_, new_n35581_, new_n35583_, new_n35584_, new_n35585_,
    new_n35586_, new_n35587_, new_n35588_, new_n35589_, new_n35591_,
    new_n35592_, new_n35594_, new_n35595_, new_n35597_, new_n35598_,
    new_n35600_, new_n35601_, new_n35603_, new_n35604_, new_n35606_,
    new_n35607_, new_n35609_, new_n35610_, new_n35612_, new_n35613_,
    new_n35615_, new_n35616_, new_n35618_, new_n35619_, new_n35621_,
    new_n35622_, new_n35624_, new_n35625_, new_n35627_, new_n35628_,
    new_n35630_, new_n35631_, new_n35633_, new_n35634_, new_n35636_,
    new_n35637_, new_n35639_, new_n35640_, new_n35642_, new_n35643_,
    new_n35645_, new_n35646_, new_n35648_, new_n35649_, new_n35651_,
    new_n35652_, new_n35654_, new_n35655_, new_n35657_, new_n35658_,
    new_n35660_, new_n35661_, new_n35663_, new_n35664_, new_n35666_,
    new_n35667_, new_n35669_, new_n35670_, new_n35672_, new_n35673_,
    new_n35675_, new_n35676_, new_n35678_, new_n35679_, new_n35681_,
    new_n35682_, new_n35684_, new_n35685_, new_n35686_, new_n35687_,
    new_n35688_, new_n35689_, new_n35690_, new_n35691_, new_n35692_,
    new_n35693_, new_n35694_, new_n35695_, new_n35696_, new_n35697_,
    new_n35698_, new_n35699_, new_n35700_, new_n35701_, new_n35702_,
    new_n35703_, new_n35705_, new_n35706_, new_n35707_, new_n35708_,
    new_n35709_, new_n35710_, new_n35711_, new_n35712_, new_n35713_,
    new_n35714_, new_n35715_, new_n35716_, new_n35717_, new_n35718_,
    new_n35719_, new_n35720_, new_n35721_, new_n35722_, new_n35723_,
    new_n35724_, new_n35725_, new_n35726_, new_n35727_, new_n35729_,
    new_n35730_, new_n35731_, new_n35732_, new_n35733_, new_n35734_,
    new_n35735_, new_n35736_, new_n35737_, new_n35738_, new_n35739_,
    new_n35740_, new_n35741_, new_n35742_, new_n35743_, new_n35744_,
    new_n35745_, new_n35746_, new_n35747_, new_n35748_, new_n35749_,
    new_n35750_, new_n35751_, new_n35752_, new_n35753_, new_n35754_,
    new_n35755_, new_n35756_, new_n35758_, new_n35759_, new_n35760_,
    new_n35761_, new_n35762_, new_n35763_, new_n35764_, new_n35765_,
    new_n35766_, new_n35767_, new_n35768_, new_n35769_, new_n35770_,
    new_n35771_, new_n35772_, new_n35773_, new_n35774_, new_n35775_,
    new_n35776_, new_n35777_, new_n35778_, new_n35779_, new_n35780_,
    new_n35781_, new_n35782_, new_n35783_, new_n35784_, new_n35785_,
    new_n35787_, new_n35788_, new_n35789_, new_n35790_, new_n35791_,
    new_n35792_, new_n35793_, new_n35794_, new_n35795_, new_n35796_,
    new_n35797_, new_n35798_, new_n35799_, new_n35800_, new_n35801_,
    new_n35802_, new_n35803_, new_n35804_, new_n35805_, new_n35806_,
    new_n35807_, new_n35808_, new_n35809_, new_n35810_, new_n35811_,
    new_n35812_, new_n35813_, new_n35814_, new_n35816_, new_n35817_,
    new_n35818_, new_n35819_, new_n35820_, new_n35821_, new_n35822_,
    new_n35823_, new_n35824_, new_n35825_, new_n35826_, new_n35827_,
    new_n35828_, new_n35829_, new_n35830_, new_n35831_, new_n35832_,
    new_n35833_, new_n35834_, new_n35835_, new_n35836_, new_n35837_,
    new_n35838_, new_n35839_, new_n35840_, new_n35841_, new_n35842_,
    new_n35843_, new_n35845_, new_n35846_, new_n35847_, new_n35848_,
    new_n35849_, new_n35850_, new_n35851_, new_n35852_, new_n35853_,
    new_n35854_, new_n35855_, new_n35856_, new_n35857_, new_n35858_,
    new_n35859_, new_n35860_, new_n35861_, new_n35862_, new_n35863_,
    new_n35864_, new_n35865_, new_n35866_, new_n35867_, new_n35868_,
    new_n35869_, new_n35870_, new_n35871_, new_n35872_, new_n35874_,
    new_n35875_, new_n35876_, new_n35877_, new_n35878_, new_n35879_,
    new_n35880_, new_n35881_, new_n35882_, new_n35883_, new_n35884_,
    new_n35885_, new_n35886_, new_n35887_, new_n35888_, new_n35889_,
    new_n35890_, new_n35891_, new_n35892_, new_n35893_, new_n35894_,
    new_n35895_, new_n35896_, new_n35897_, new_n35898_, new_n35899_,
    new_n35900_, new_n35901_, new_n35903_, new_n35904_, new_n35905_,
    new_n35906_, new_n35907_, new_n35908_, new_n35909_, new_n35910_,
    new_n35911_, new_n35912_, new_n35913_, new_n35914_, new_n35915_,
    new_n35916_, new_n35917_, new_n35918_, new_n35919_, new_n35920_,
    new_n35921_, new_n35922_, new_n35923_, new_n35924_, new_n35925_,
    new_n35926_, new_n35927_, new_n35928_, new_n35929_, new_n35930_,
    new_n35932_, new_n35933_, new_n35934_, new_n35935_, new_n35936_,
    new_n35937_, new_n35938_, new_n35939_, new_n35940_, new_n35941_,
    new_n35942_, new_n35943_, new_n35944_, new_n35945_, new_n35946_,
    new_n35947_, new_n35948_, new_n35949_, new_n35950_, new_n35951_,
    new_n35952_, new_n35953_, new_n35954_, new_n35955_, new_n35956_,
    new_n35957_, new_n35959_, new_n35960_, new_n35961_, new_n35962_,
    new_n35963_, new_n35964_, new_n35965_, new_n35966_, new_n35967_,
    new_n35968_, new_n35969_, new_n35970_, new_n35971_, new_n35972_,
    new_n35973_, new_n35974_, new_n35975_, new_n35976_, new_n35977_,
    new_n35978_, new_n35979_, new_n35980_, new_n35981_, new_n35982_,
    new_n35983_, new_n35984_, new_n35985_, new_n35986_, new_n35988_,
    new_n35989_, new_n35990_, new_n35991_, new_n35992_, new_n35993_,
    new_n35994_, new_n35995_, new_n35996_, new_n35997_, new_n35998_,
    new_n35999_, new_n36000_, new_n36001_, new_n36002_, new_n36003_,
    new_n36004_, new_n36005_, new_n36006_, new_n36007_, new_n36008_,
    new_n36009_, new_n36010_, new_n36011_, new_n36012_, new_n36013_,
    new_n36014_, new_n36015_, new_n36016_, new_n36017_, new_n36018_,
    new_n36019_, new_n36020_, new_n36021_, new_n36022_, new_n36024_,
    new_n36025_, new_n36026_, new_n36027_, new_n36028_, new_n36029_,
    new_n36030_, new_n36031_, new_n36032_, new_n36033_, new_n36034_,
    new_n36035_, new_n36036_, new_n36037_, new_n36038_, new_n36039_,
    new_n36040_, new_n36041_, new_n36042_, new_n36043_, new_n36044_,
    new_n36045_, new_n36046_, new_n36047_, new_n36048_, new_n36049_,
    new_n36050_, new_n36051_, new_n36052_, new_n36053_, new_n36054_,
    new_n36055_, new_n36056_, new_n36057_, new_n36058_, new_n36059_,
    new_n36060_, new_n36062_, new_n36063_, new_n36064_, new_n36065_,
    new_n36066_, new_n36067_, new_n36068_, new_n36069_, new_n36070_,
    new_n36071_, new_n36072_, new_n36073_, new_n36074_, new_n36075_,
    new_n36076_, new_n36077_, new_n36078_, new_n36079_, new_n36080_,
    new_n36081_, new_n36082_, new_n36083_, new_n36084_, new_n36085_,
    new_n36086_, new_n36087_, new_n36088_, new_n36089_, new_n36090_,
    new_n36091_, new_n36092_, new_n36093_, new_n36094_, new_n36095_,
    new_n36096_, new_n36097_, new_n36098_, new_n36099_, new_n36100_,
    new_n36101_, new_n36103_, new_n36104_, new_n36105_, new_n36106_,
    new_n36107_, new_n36108_, new_n36109_, new_n36110_, new_n36111_,
    new_n36112_, new_n36113_, new_n36114_, new_n36115_, new_n36116_,
    new_n36117_, new_n36118_, new_n36119_, new_n36120_, new_n36121_,
    new_n36122_, new_n36123_, new_n36124_, new_n36125_, new_n36126_,
    new_n36127_, new_n36128_, new_n36129_, new_n36130_, new_n36131_,
    new_n36132_, new_n36133_, new_n36134_, new_n36135_, new_n36136_,
    new_n36137_, new_n36138_, new_n36139_, new_n36140_, new_n36141_,
    new_n36142_, new_n36144_, new_n36145_, new_n36146_, new_n36147_,
    new_n36148_, new_n36149_, new_n36150_, new_n36151_, new_n36152_,
    new_n36153_, new_n36154_, new_n36155_, new_n36156_, new_n36157_,
    new_n36158_, new_n36159_, new_n36160_, new_n36161_, new_n36162_,
    new_n36163_, new_n36164_, new_n36165_, new_n36166_, new_n36167_,
    new_n36168_, new_n36169_, new_n36170_, new_n36171_, new_n36172_,
    new_n36173_, new_n36174_, new_n36175_, new_n36176_, new_n36177_,
    new_n36178_, new_n36179_, new_n36180_, new_n36181_, new_n36182_,
    new_n36183_, new_n36184_, new_n36185_, new_n36186_, new_n36187_,
    new_n36188_, new_n36189_, new_n36190_, new_n36191_, new_n36193_,
    new_n36194_, new_n36195_, new_n36196_, new_n36197_, new_n36198_,
    new_n36199_, new_n36200_, new_n36201_, new_n36202_, new_n36203_,
    new_n36204_, new_n36205_, new_n36206_, new_n36207_, new_n36208_,
    new_n36209_, new_n36210_, new_n36211_, new_n36212_, new_n36213_,
    new_n36214_, new_n36215_, new_n36216_, new_n36217_, new_n36218_,
    new_n36219_, new_n36220_, new_n36221_, new_n36222_, new_n36223_,
    new_n36224_, new_n36225_, new_n36226_, new_n36227_, new_n36228_,
    new_n36229_, new_n36230_, new_n36231_, new_n36232_, new_n36233_,
    new_n36234_, new_n36235_, new_n36237_, new_n36238_, new_n36239_,
    new_n36240_, new_n36241_, new_n36242_, new_n36243_, new_n36244_,
    new_n36245_, new_n36246_, new_n36247_, new_n36248_, new_n36249_,
    new_n36250_, new_n36251_, new_n36252_, new_n36253_, new_n36254_,
    new_n36255_, new_n36256_, new_n36257_, new_n36258_, new_n36259_,
    new_n36260_, new_n36261_, new_n36262_, new_n36263_, new_n36264_,
    new_n36265_, new_n36266_, new_n36267_, new_n36268_, new_n36269_,
    new_n36270_, new_n36271_, new_n36272_, new_n36273_, new_n36274_,
    new_n36275_, new_n36276_, new_n36277_, new_n36278_, new_n36279_,
    new_n36281_, new_n36282_, new_n36283_, new_n36284_, new_n36285_,
    new_n36286_, new_n36287_, new_n36288_, new_n36289_, new_n36290_,
    new_n36291_, new_n36292_, new_n36293_, new_n36294_, new_n36295_,
    new_n36296_, new_n36297_, new_n36298_, new_n36299_, new_n36300_,
    new_n36301_, new_n36302_, new_n36303_, new_n36304_, new_n36305_,
    new_n36306_, new_n36307_, new_n36308_, new_n36309_, new_n36310_,
    new_n36311_, new_n36312_, new_n36313_, new_n36314_, new_n36315_,
    new_n36316_, new_n36317_, new_n36318_, new_n36319_, new_n36320_,
    new_n36322_, new_n36323_, new_n36324_, new_n36325_, new_n36326_,
    new_n36327_, new_n36328_, new_n36329_, new_n36330_, new_n36331_,
    new_n36332_, new_n36333_, new_n36334_, new_n36335_, new_n36336_,
    new_n36337_, new_n36338_, new_n36339_, new_n36340_, new_n36341_,
    new_n36342_, new_n36343_, new_n36344_, new_n36345_, new_n36346_,
    new_n36347_, new_n36348_, new_n36349_, new_n36350_, new_n36351_,
    new_n36352_, new_n36353_, new_n36354_, new_n36355_, new_n36356_,
    new_n36357_, new_n36358_, new_n36359_, new_n36360_, new_n36361_,
    new_n36362_, new_n36363_, new_n36364_, new_n36366_, new_n36367_,
    new_n36368_, new_n36369_, new_n36370_, new_n36371_, new_n36372_,
    new_n36373_, new_n36374_, new_n36375_, new_n36376_, new_n36377_,
    new_n36378_, new_n36379_, new_n36380_, new_n36381_, new_n36382_,
    new_n36383_, new_n36384_, new_n36385_, new_n36386_, new_n36387_,
    new_n36388_, new_n36389_, new_n36390_, new_n36391_, new_n36392_,
    new_n36393_, new_n36394_, new_n36395_, new_n36396_, new_n36397_,
    new_n36398_, new_n36399_, new_n36400_, new_n36401_, new_n36402_,
    new_n36403_, new_n36404_, new_n36405_, new_n36406_, new_n36407_,
    new_n36408_, new_n36410_, new_n36411_, new_n36412_, new_n36413_,
    new_n36414_, new_n36415_, new_n36416_, new_n36417_, new_n36418_,
    new_n36419_, new_n36420_, new_n36421_, new_n36422_, new_n36423_,
    new_n36424_, new_n36425_, new_n36426_, new_n36427_, new_n36428_,
    new_n36429_, new_n36430_, new_n36431_, new_n36432_, new_n36433_,
    new_n36434_, new_n36435_, new_n36436_, new_n36437_, new_n36438_,
    new_n36439_, new_n36440_, new_n36441_, new_n36442_, new_n36443_,
    new_n36444_, new_n36445_, new_n36446_, new_n36447_, new_n36448_,
    new_n36449_, new_n36453_, new_n36454_, new_n36455_, new_n36456_,
    new_n36457_, new_n36458_, new_n36459_, new_n36460_, new_n36461_,
    new_n36462_, new_n36463_, new_n36464_, new_n36465_, new_n36466_,
    new_n36467_, new_n36468_, new_n36469_, new_n36470_, new_n36471_,
    new_n36472_, new_n36473_, new_n36474_, new_n36475_, new_n36476_,
    new_n36477_, new_n36478_, new_n36479_, new_n36480_, new_n36481_,
    new_n36482_, new_n36483_, new_n36484_, new_n36485_, new_n36486_,
    new_n36487_, new_n36488_, new_n36489_, new_n36490_, new_n36491_,
    new_n36492_, new_n36493_, new_n36494_, new_n36495_, new_n36496_,
    new_n36497_, new_n36498_, new_n36499_, new_n36500_, new_n36501_,
    new_n36502_, new_n36503_, new_n36504_, new_n36505_, new_n36506_,
    new_n36507_, new_n36508_, new_n36509_, new_n36510_, new_n36511_,
    new_n36512_, new_n36513_, new_n36514_, new_n36515_, new_n36516_,
    new_n36517_, new_n36518_, new_n36519_, new_n36520_, new_n36521_,
    new_n36522_, new_n36523_, new_n36524_, new_n36525_, new_n36526_,
    new_n36527_, new_n36528_, new_n36529_, new_n36530_, new_n36531_,
    new_n36532_, new_n36533_, new_n36534_, new_n36535_, new_n36536_,
    new_n36537_, new_n36538_, new_n36539_, new_n36540_, new_n36541_,
    new_n36542_, new_n36543_, new_n36544_, new_n36545_, new_n36546_,
    new_n36547_, new_n36548_, new_n36549_, new_n36550_, new_n36551_,
    new_n36552_, new_n36553_, new_n36554_, new_n36555_, new_n36556_,
    new_n36557_, new_n36558_, new_n36559_, new_n36560_, new_n36561_,
    new_n36562_, new_n36563_, new_n36564_, new_n36565_, new_n36566_,
    new_n36568_, new_n36569_, new_n36570_, new_n36571_, new_n36572_,
    new_n36573_, new_n36574_, new_n36575_, new_n36576_, new_n36577_,
    new_n36578_, new_n36579_, new_n36580_, new_n36581_, new_n36582_,
    new_n36583_, new_n36584_, new_n36585_, new_n36586_, new_n36587_,
    new_n36588_, new_n36589_, new_n36590_, new_n36591_, new_n36592_,
    new_n36594_, new_n36595_, new_n36596_, new_n36597_, new_n36598_,
    new_n36599_, new_n36600_, new_n36601_, new_n36602_, new_n36603_,
    new_n36604_, new_n36605_, new_n36606_, new_n36607_, new_n36608_,
    new_n36609_, new_n36610_, new_n36611_, new_n36612_, new_n36613_,
    new_n36614_, new_n36615_, new_n36616_, new_n36617_, new_n36618_,
    new_n36619_, new_n36620_, new_n36621_, new_n36622_, new_n36623_,
    new_n36625_, new_n36626_, new_n36627_, new_n36628_, new_n36629_,
    new_n36630_, new_n36631_, new_n36632_, new_n36633_, new_n36634_,
    new_n36635_, new_n36636_, new_n36637_, new_n36638_, new_n36639_,
    new_n36640_, new_n36641_, new_n36642_, new_n36643_, new_n36644_,
    new_n36645_, new_n36646_, new_n36647_, new_n36648_, new_n36649_,
    new_n36650_, new_n36651_, new_n36652_, new_n36653_, new_n36654_,
    new_n36655_, new_n36656_, new_n36657_, new_n36658_, new_n36659_,
    new_n36660_, new_n36662_, new_n36663_, new_n36664_, new_n36665_,
    new_n36666_, new_n36667_, new_n36668_, new_n36669_, new_n36670_,
    new_n36671_, new_n36672_, new_n36673_, new_n36674_, new_n36675_,
    new_n36676_, new_n36677_, new_n36678_, new_n36679_, new_n36680_,
    new_n36681_, new_n36682_, new_n36683_, new_n36684_, new_n36685_,
    new_n36686_, new_n36687_, new_n36688_, new_n36689_, new_n36690_,
    new_n36691_, new_n36692_, new_n36693_, new_n36694_, new_n36695_,
    new_n36696_, new_n36697_, new_n36698_, new_n36699_, new_n36700_,
    new_n36701_, new_n36703_, new_n36704_, new_n36705_, new_n36706_,
    new_n36707_, new_n36708_, new_n36709_, new_n36710_, new_n36711_,
    new_n36712_, new_n36713_, new_n36714_, new_n36715_, new_n36716_,
    new_n36717_, new_n36718_, new_n36719_, new_n36720_, new_n36721_,
    new_n36722_, new_n36723_, new_n36724_, new_n36725_, new_n36726_,
    new_n36727_, new_n36728_, new_n36729_, new_n36730_, new_n36731_,
    new_n36732_, new_n36733_, new_n36734_, new_n36735_, new_n36736_,
    new_n36737_, new_n36738_, new_n36739_, new_n36740_, new_n36741_,
    new_n36742_, new_n36743_, new_n36744_, new_n36746_, new_n36747_,
    new_n36748_, new_n36749_, new_n36750_, new_n36751_, new_n36752_,
    new_n36753_, new_n36754_, new_n36755_, new_n36756_, new_n36757_,
    new_n36758_, new_n36759_, new_n36760_, new_n36761_, new_n36762_,
    new_n36763_, new_n36764_, new_n36765_, new_n36766_, new_n36767_,
    new_n36768_, new_n36769_, new_n36770_, new_n36771_, new_n36772_,
    new_n36773_, new_n36774_, new_n36775_, new_n36776_, new_n36777_,
    new_n36778_, new_n36779_, new_n36780_, new_n36781_, new_n36782_,
    new_n36783_, new_n36784_, new_n36785_, new_n36786_, new_n36787_,
    new_n36789_, new_n36790_, new_n36791_, new_n36792_, new_n36793_,
    new_n36794_, new_n36795_, new_n36796_, new_n36797_, new_n36798_,
    new_n36799_, new_n36800_, new_n36801_, new_n36802_, new_n36803_,
    new_n36804_, new_n36805_, new_n36806_, new_n36807_, new_n36808_,
    new_n36809_, new_n36810_, new_n36811_, new_n36812_, new_n36813_,
    new_n36814_, new_n36815_, new_n36816_, new_n36817_, new_n36818_,
    new_n36819_, new_n36821_, new_n36822_, new_n36823_, new_n36824_,
    new_n36825_, new_n36826_, new_n36827_, new_n36828_, new_n36829_,
    new_n36830_, new_n36831_, new_n36832_, new_n36833_, new_n36834_,
    new_n36835_, new_n36836_, new_n36837_, new_n36838_, new_n36839_,
    new_n36840_, new_n36841_, new_n36842_, new_n36843_, new_n36844_,
    new_n36845_, new_n36846_, new_n36847_, new_n36848_, new_n36849_,
    new_n36850_, new_n36851_, new_n36853_, new_n36854_, new_n36855_,
    new_n36856_, new_n36857_, new_n36858_, new_n36859_, new_n36860_,
    new_n36861_, new_n36862_, new_n36863_, new_n36864_, new_n36865_,
    new_n36866_, new_n36867_, new_n36868_, new_n36869_, new_n36870_,
    new_n36871_, new_n36872_, new_n36873_, new_n36874_, new_n36875_,
    new_n36876_, new_n36877_, new_n36878_, new_n36879_, new_n36880_,
    new_n36881_, new_n36882_, new_n36883_, new_n36885_, new_n36886_,
    new_n36887_, new_n36888_, new_n36889_, new_n36890_, new_n36891_,
    new_n36892_, new_n36893_, new_n36894_, new_n36895_, new_n36896_,
    new_n36897_, new_n36898_, new_n36899_, new_n36900_, new_n36901_,
    new_n36902_, new_n36903_, new_n36904_, new_n36905_, new_n36906_,
    new_n36907_, new_n36908_, new_n36909_, new_n36910_, new_n36911_,
    new_n36912_, new_n36913_, new_n36914_, new_n36915_, new_n36917_,
    new_n36918_, new_n36919_, new_n36920_, new_n36921_, new_n36922_,
    new_n36923_, new_n36924_, new_n36925_, new_n36926_, new_n36927_,
    new_n36928_, new_n36929_, new_n36930_, new_n36931_, new_n36932_,
    new_n36933_, new_n36934_, new_n36935_, new_n36936_, new_n36937_,
    new_n36938_, new_n36939_, new_n36940_, new_n36941_, new_n36942_,
    new_n36943_, new_n36944_, new_n36945_, new_n36946_, new_n36947_,
    new_n36949_, new_n36950_, new_n36951_, new_n36952_, new_n36953_,
    new_n36954_, new_n36955_, new_n36956_, new_n36957_, new_n36958_,
    new_n36959_, new_n36960_, new_n36961_, new_n36962_, new_n36963_,
    new_n36964_, new_n36965_, new_n36966_, new_n36967_, new_n36968_,
    new_n36969_, new_n36970_, new_n36971_, new_n36972_, new_n36973_,
    new_n36974_, new_n36975_, new_n36976_, new_n36977_, new_n36978_,
    new_n36979_, new_n36981_, new_n36982_, new_n36983_, new_n36984_,
    new_n36985_, new_n36986_, new_n36987_, new_n36988_, new_n36989_,
    new_n36990_, new_n36991_, new_n36992_, new_n36993_, new_n36994_,
    new_n36995_, new_n36996_, new_n36997_, new_n36998_, new_n36999_,
    new_n37000_, new_n37001_, new_n37002_, new_n37003_, new_n37004_,
    new_n37005_, new_n37006_, new_n37007_, new_n37008_, new_n37009_,
    new_n37010_, new_n37011_, new_n37013_, new_n37014_, new_n37015_,
    new_n37016_, new_n37017_, new_n37018_, new_n37019_, new_n37020_,
    new_n37021_, new_n37022_, new_n37023_, new_n37024_, new_n37025_,
    new_n37026_, new_n37027_, new_n37028_, new_n37029_, new_n37030_,
    new_n37031_, new_n37032_, new_n37033_, new_n37034_, new_n37035_,
    new_n37037_, new_n37038_, new_n37039_, new_n37040_, new_n37041_,
    new_n37042_, new_n37043_, new_n37044_, new_n37045_, new_n37046_,
    new_n37047_, new_n37048_, new_n37049_, new_n37050_, new_n37051_,
    new_n37052_, new_n37053_, new_n37054_, new_n37055_, new_n37056_,
    new_n37057_, new_n37058_, new_n37059_, new_n37061_, new_n37062_,
    new_n37063_, new_n37064_, new_n37065_, new_n37066_, new_n37067_,
    new_n37068_, new_n37069_, new_n37070_, new_n37071_, new_n37072_,
    new_n37073_, new_n37074_, new_n37075_, new_n37076_, new_n37077_,
    new_n37078_, new_n37079_, new_n37080_, new_n37081_, new_n37082_,
    new_n37083_, new_n37085_, new_n37086_, new_n37087_, new_n37088_,
    new_n37089_, new_n37090_, new_n37091_, new_n37092_, new_n37093_,
    new_n37094_, new_n37095_, new_n37096_, new_n37097_, new_n37098_,
    new_n37099_, new_n37100_, new_n37101_, new_n37102_, new_n37103_,
    new_n37104_, new_n37105_, new_n37106_, new_n37107_, new_n37109_,
    new_n37110_, new_n37111_, new_n37112_, new_n37113_, new_n37114_,
    new_n37115_, new_n37116_, new_n37117_, new_n37118_, new_n37119_,
    new_n37120_, new_n37121_, new_n37122_, new_n37123_, new_n37124_,
    new_n37125_, new_n37126_, new_n37127_, new_n37128_, new_n37129_,
    new_n37130_, new_n37131_, new_n37133_, new_n37134_, new_n37135_,
    new_n37136_, new_n37137_, new_n37138_, new_n37139_, new_n37140_,
    new_n37141_, new_n37142_, new_n37143_, new_n37144_, new_n37145_,
    new_n37146_, new_n37147_, new_n37148_, new_n37149_, new_n37150_,
    new_n37151_, new_n37152_, new_n37153_, new_n37154_, new_n37155_,
    new_n37157_, new_n37158_, new_n37159_, new_n37160_, new_n37161_,
    new_n37162_, new_n37163_, new_n37164_, new_n37165_, new_n37166_,
    new_n37167_, new_n37168_, new_n37169_, new_n37170_, new_n37171_,
    new_n37172_, new_n37173_, new_n37174_, new_n37175_, new_n37176_,
    new_n37177_, new_n37178_, new_n37179_, new_n37181_, new_n37182_,
    new_n37183_, new_n37184_, new_n37185_, new_n37186_, new_n37187_,
    new_n37188_, new_n37189_, new_n37190_, new_n37191_, new_n37192_,
    new_n37193_, new_n37194_, new_n37195_, new_n37196_, new_n37197_,
    new_n37198_, new_n37199_, new_n37200_, new_n37201_, new_n37202_,
    new_n37203_, new_n37205_, new_n37206_, new_n37207_, new_n37208_,
    new_n37209_, new_n37210_, new_n37211_, new_n37212_, new_n37213_,
    new_n37214_, new_n37215_, new_n37216_, new_n37217_, new_n37218_,
    new_n37219_, new_n37220_, new_n37221_, new_n37222_, new_n37223_,
    new_n37224_, new_n37225_, new_n37226_, new_n37227_, new_n37229_,
    new_n37230_, new_n37231_, new_n37232_, new_n37233_, new_n37234_,
    new_n37235_, new_n37236_, new_n37237_, new_n37238_, new_n37239_,
    new_n37240_, new_n37241_, new_n37242_, new_n37243_, new_n37244_,
    new_n37245_, new_n37246_, new_n37247_, new_n37248_, new_n37249_,
    new_n37250_, new_n37251_, new_n37253_, new_n37254_, new_n37255_,
    new_n37256_, new_n37257_, new_n37258_, new_n37259_, new_n37260_,
    new_n37261_, new_n37262_, new_n37263_, new_n37264_, new_n37265_,
    new_n37266_, new_n37267_, new_n37268_, new_n37269_, new_n37270_,
    new_n37271_, new_n37272_, new_n37273_, new_n37274_, new_n37275_,
    new_n37277_, new_n37278_, new_n37279_, new_n37280_, new_n37281_,
    new_n37282_, new_n37283_, new_n37284_, new_n37285_, new_n37286_,
    new_n37287_, new_n37288_, new_n37289_, new_n37290_, new_n37291_,
    new_n37292_, new_n37293_, new_n37294_, new_n37295_, new_n37296_,
    new_n37297_, new_n37298_, new_n37299_, new_n37301_, new_n37302_,
    new_n37303_, new_n37304_, new_n37305_, new_n37306_, new_n37307_,
    new_n37308_, new_n37309_, new_n37310_, new_n37311_, new_n37312_,
    new_n37313_, new_n37314_, new_n37315_, new_n37316_, new_n37317_,
    new_n37318_, new_n37319_, new_n37320_, new_n37321_, new_n37322_,
    new_n37323_, new_n37325_, new_n37326_, new_n37327_, new_n37328_,
    new_n37329_, new_n37330_, new_n37331_, new_n37332_, new_n37333_,
    new_n37334_, new_n37335_, new_n37336_, new_n37337_, new_n37338_,
    new_n37339_, new_n37340_, new_n37341_, new_n37342_, new_n37343_,
    new_n37344_, new_n37345_, new_n37346_, new_n37347_, new_n37349_,
    new_n37350_, new_n37351_, new_n37352_, new_n37353_, new_n37354_,
    new_n37355_, new_n37356_, new_n37357_, new_n37358_, new_n37359_,
    new_n37360_, new_n37361_, new_n37362_, new_n37363_, new_n37364_,
    new_n37365_, new_n37366_, new_n37367_, new_n37368_, new_n37369_,
    new_n37370_, new_n37371_, new_n37373_, new_n37374_, new_n37375_,
    new_n37376_, new_n37377_, new_n37378_, new_n37379_, new_n37380_,
    new_n37381_, new_n37382_, new_n37383_, new_n37384_, new_n37385_,
    new_n37386_, new_n37387_, new_n37388_, new_n37389_, new_n37390_,
    new_n37391_, new_n37392_, new_n37393_, new_n37394_, new_n37395_,
    new_n37397_, new_n37398_, new_n37399_, new_n37400_, new_n37401_,
    new_n37402_, new_n37403_, new_n37404_, new_n37405_, new_n37406_,
    new_n37407_, new_n37408_, new_n37409_, new_n37410_, new_n37411_,
    new_n37412_, new_n37413_, new_n37414_, new_n37415_, new_n37416_,
    new_n37417_, new_n37418_, new_n37419_, new_n37421_, new_n37422_,
    new_n37423_, new_n37424_, new_n37425_, new_n37426_, new_n37427_,
    new_n37428_, new_n37429_, new_n37430_, new_n37431_, new_n37432_,
    new_n37433_, new_n37434_, new_n37435_, new_n37436_, new_n37437_,
    new_n37438_, new_n37439_, new_n37440_, new_n37441_, new_n37442_,
    new_n37443_, new_n37445_, new_n37446_, new_n37447_, new_n37448_,
    new_n37449_, new_n37450_, new_n37451_, new_n37452_, new_n37453_,
    new_n37454_, new_n37455_, new_n37456_, new_n37457_, new_n37458_,
    new_n37459_, new_n37460_, new_n37461_, new_n37462_, new_n37463_,
    new_n37464_, new_n37465_, new_n37466_, new_n37467_, new_n37469_,
    new_n37470_, new_n37471_, new_n37472_, new_n37473_, new_n37474_,
    new_n37475_, new_n37476_, new_n37477_, new_n37478_, new_n37479_,
    new_n37480_, new_n37481_, new_n37482_, new_n37483_, new_n37484_,
    new_n37485_, new_n37486_, new_n37487_, new_n37488_, new_n37489_,
    new_n37490_, new_n37491_, new_n37493_, new_n37494_, new_n37495_,
    new_n37496_, new_n37497_, new_n37498_, new_n37499_, new_n37500_,
    new_n37501_, new_n37502_, new_n37503_, new_n37504_, new_n37505_,
    new_n37506_, new_n37507_, new_n37508_, new_n37509_, new_n37510_,
    new_n37511_, new_n37512_, new_n37513_, new_n37514_, new_n37515_,
    new_n37517_, new_n37518_, new_n37519_, new_n37520_, new_n37521_,
    new_n37522_, new_n37523_, new_n37524_, new_n37525_, new_n37526_,
    new_n37527_, new_n37528_, new_n37529_, new_n37530_, new_n37531_,
    new_n37532_, new_n37533_, new_n37534_, new_n37535_, new_n37536_,
    new_n37537_, new_n37538_, new_n37539_, new_n37541_, new_n37542_,
    new_n37543_, new_n37544_, new_n37545_, new_n37546_, new_n37547_,
    new_n37548_, new_n37549_, new_n37550_, new_n37551_, new_n37552_,
    new_n37553_, new_n37554_, new_n37555_, new_n37556_, new_n37557_,
    new_n37558_, new_n37559_, new_n37560_, new_n37561_, new_n37562_,
    new_n37563_, new_n37565_, new_n37566_, new_n37567_, new_n37568_,
    new_n37569_, new_n37570_, new_n37571_, new_n37572_, new_n37573_,
    new_n37574_, new_n37575_, new_n37576_, new_n37577_, new_n37578_,
    new_n37579_, new_n37580_, new_n37581_, new_n37582_, new_n37583_,
    new_n37585_, new_n37586_, new_n37587_, new_n37588_, new_n37589_,
    new_n37590_, new_n37591_, new_n37592_, new_n37593_, new_n37594_,
    new_n37595_, new_n37596_, new_n37597_, new_n37599_, new_n37600_,
    new_n37601_, new_n37602_, new_n37603_, new_n37604_, new_n37605_,
    new_n37606_, new_n37607_, new_n37608_, new_n37609_, new_n37610_,
    new_n37611_, new_n37613_, new_n37614_, new_n37615_, new_n37616_,
    new_n37617_, new_n37618_, new_n37619_, new_n37620_, new_n37621_,
    new_n37622_, new_n37623_, new_n37624_, new_n37625_, new_n37627_,
    new_n37628_, new_n37629_, new_n37630_, new_n37631_, new_n37632_,
    new_n37633_, new_n37634_, new_n37635_, new_n37636_, new_n37637_,
    new_n37638_, new_n37639_, new_n37641_, new_n37642_, new_n37643_,
    new_n37644_, new_n37645_, new_n37646_, new_n37647_, new_n37648_,
    new_n37649_, new_n37650_, new_n37651_, new_n37652_, new_n37654_,
    new_n37655_, new_n37656_, new_n37657_, new_n37658_, new_n37659_,
    new_n37660_, new_n37661_, new_n37662_, new_n37663_, new_n37664_,
    new_n37665_, new_n37667_, new_n37668_, new_n37669_, new_n37670_,
    new_n37671_, new_n37672_, new_n37673_, new_n37674_, new_n37675_,
    new_n37676_, new_n37678_, new_n37679_, new_n37680_, new_n37681_,
    new_n37682_, new_n37683_, new_n37684_, new_n37685_, new_n37686_,
    new_n37687_, new_n37689_, new_n37690_, new_n37691_, new_n37692_,
    new_n37693_, new_n37694_, new_n37695_, new_n37696_, new_n37697_,
    new_n37698_, new_n37699_, new_n37700_, new_n37701_, new_n37702_,
    new_n37703_, new_n37704_, new_n37705_, new_n37706_, new_n37707_,
    new_n37708_, new_n37709_, new_n37711_, new_n37712_, new_n37713_,
    new_n37714_, new_n37715_, new_n37716_, new_n37717_, new_n37718_,
    new_n37719_, new_n37720_, new_n37721_, new_n37722_, new_n37723_,
    new_n37724_, new_n37725_, new_n37726_, new_n37727_, new_n37728_,
    new_n37729_, new_n37730_, new_n37731_, new_n37733_, new_n37734_,
    new_n37735_, new_n37736_, new_n37737_, new_n37738_, new_n37739_,
    new_n37740_, new_n37741_, new_n37742_, new_n37743_, new_n37744_,
    new_n37745_, new_n37746_, new_n37747_, new_n37748_, new_n37749_,
    new_n37750_, new_n37751_, new_n37752_, new_n37753_, new_n37755_,
    new_n37756_, new_n37757_, new_n37758_, new_n37759_, new_n37760_,
    new_n37761_, new_n37762_, new_n37763_, new_n37764_, new_n37765_,
    new_n37766_, new_n37767_, new_n37768_, new_n37769_, new_n37770_,
    new_n37771_, new_n37772_, new_n37773_, new_n37774_, new_n37775_,
    new_n37777_, new_n37778_, new_n37779_, new_n37780_, new_n37781_,
    new_n37782_, new_n37783_, new_n37784_, new_n37785_, new_n37786_,
    new_n37787_, new_n37788_, new_n37789_, new_n37790_, new_n37791_,
    new_n37792_, new_n37793_, new_n37794_, new_n37795_, new_n37796_,
    new_n37797_, new_n37799_, new_n37800_, new_n37801_, new_n37802_,
    new_n37803_, new_n37804_, new_n37805_, new_n37806_, new_n37807_,
    new_n37808_, new_n37809_, new_n37810_, new_n37811_, new_n37812_,
    new_n37813_, new_n37814_, new_n37815_, new_n37816_, new_n37817_,
    new_n37818_, new_n37819_, new_n37821_, new_n37822_, new_n37823_,
    new_n37824_, new_n37825_, new_n37826_, new_n37827_, new_n37828_,
    new_n37829_, new_n37830_, new_n37831_, new_n37832_, new_n37833_,
    new_n37834_, new_n37835_, new_n37836_, new_n37837_, new_n37838_,
    new_n37839_, new_n37840_, new_n37841_, new_n37843_, new_n37844_,
    new_n37845_, new_n37846_, new_n37847_, new_n37848_, new_n37849_,
    new_n37850_, new_n37851_, new_n37852_, new_n37853_, new_n37854_,
    new_n37855_, new_n37856_, new_n37857_, new_n37858_, new_n37859_,
    new_n37860_, new_n37861_, new_n37862_, new_n37863_, new_n37864_,
    new_n37865_, new_n37866_, new_n37867_, new_n37868_, new_n37869_,
    new_n37870_, new_n37871_, new_n37872_, new_n37873_, new_n37874_,
    new_n37875_, new_n37876_, new_n37877_, new_n37878_, new_n37879_,
    new_n37880_, new_n37881_, new_n37882_, new_n37883_, new_n37884_,
    new_n37885_, new_n37886_, new_n37887_, new_n37888_, new_n37889_,
    new_n37890_, new_n37891_, new_n37892_, new_n37894_, new_n37895_,
    new_n37896_, new_n37897_, new_n37898_, new_n37899_, new_n37900_,
    new_n37901_, new_n37902_, new_n37903_, new_n37904_, new_n37905_,
    new_n37906_, new_n37907_, new_n37909_, new_n37910_, new_n37911_,
    new_n37912_, new_n37913_, new_n37914_, new_n37915_, new_n37916_,
    new_n37917_, new_n37918_, new_n37919_, new_n37920_, new_n37921_,
    new_n37922_, new_n37924_, new_n37925_, new_n37926_, new_n37927_,
    new_n37928_, new_n37929_, new_n37930_, new_n37931_, new_n37932_,
    new_n37933_, new_n37934_, new_n37935_, new_n37936_, new_n37937_,
    new_n37939_, new_n37940_, new_n37941_, new_n37942_, new_n37943_,
    new_n37944_, new_n37945_, new_n37946_, new_n37947_, new_n37948_,
    new_n37949_, new_n37950_, new_n37951_, new_n37952_, new_n37954_,
    new_n37955_, new_n37956_, new_n37957_, new_n37958_, new_n37959_,
    new_n37960_, new_n37961_, new_n37962_, new_n37963_, new_n37964_,
    new_n37965_, new_n37966_, new_n37967_, new_n37969_, new_n37970_,
    new_n37971_, new_n37972_, new_n37973_, new_n37974_, new_n37975_,
    new_n37976_, new_n37977_, new_n37978_, new_n37979_, new_n37980_,
    new_n37981_, new_n37982_, new_n37984_, new_n37985_, new_n37986_,
    new_n37987_, new_n37988_, new_n37989_, new_n37990_, new_n37991_,
    new_n37992_, new_n37993_, new_n37994_, new_n37995_, new_n37996_,
    new_n37997_, new_n37999_, new_n38000_, new_n38001_, new_n38002_,
    new_n38003_, new_n38004_, new_n38005_, new_n38006_, new_n38007_,
    new_n38008_, new_n38009_, new_n38010_, new_n38011_, new_n38012_,
    new_n38013_, new_n38014_, new_n38015_, new_n38016_, new_n38018_,
    new_n38019_, new_n38020_, new_n38021_, new_n38022_, new_n38023_,
    new_n38024_, new_n38025_, new_n38026_, new_n38027_, new_n38028_,
    new_n38029_, new_n38030_, new_n38031_, new_n38033_, new_n38034_,
    new_n38035_, new_n38036_, new_n38037_, new_n38038_, new_n38039_,
    new_n38040_, new_n38041_, new_n38042_, new_n38043_, new_n38044_,
    new_n38045_, new_n38046_, new_n38048_, new_n38049_, new_n38050_,
    new_n38051_, new_n38052_, new_n38053_, new_n38054_, new_n38055_,
    new_n38056_, new_n38057_, new_n38058_, new_n38059_, new_n38060_,
    new_n38061_, new_n38063_, new_n38064_, new_n38065_, new_n38066_,
    new_n38067_, new_n38068_, new_n38069_, new_n38070_, new_n38071_,
    new_n38072_, new_n38073_, new_n38074_, new_n38075_, new_n38076_,
    new_n38078_, new_n38079_, new_n38080_, new_n38081_, new_n38082_,
    new_n38083_, new_n38084_, new_n38085_, new_n38086_, new_n38087_,
    new_n38088_, new_n38089_, new_n38090_, new_n38091_, new_n38093_,
    new_n38094_, new_n38095_, new_n38096_, new_n38097_, new_n38098_,
    new_n38099_, new_n38100_, new_n38101_, new_n38102_, new_n38103_,
    new_n38104_, new_n38105_, new_n38106_, new_n38108_, new_n38109_,
    new_n38110_, new_n38111_, new_n38112_, new_n38113_, new_n38114_,
    new_n38115_, new_n38116_, new_n38117_, new_n38118_, new_n38119_,
    new_n38120_, new_n38121_, new_n38123_, new_n38124_, new_n38125_,
    new_n38126_, new_n38127_, new_n38128_, new_n38129_, new_n38130_,
    new_n38131_, new_n38132_, new_n38133_, new_n38134_, new_n38135_,
    new_n38136_, new_n38138_, new_n38139_, new_n38140_, new_n38141_,
    new_n38142_, new_n38143_, new_n38144_, new_n38145_, new_n38146_,
    new_n38147_, new_n38148_, new_n38149_, new_n38150_, new_n38151_,
    new_n38153_, new_n38154_, new_n38155_, new_n38156_, new_n38157_,
    new_n38158_, new_n38159_, new_n38160_, new_n38161_, new_n38162_,
    new_n38163_, new_n38164_, new_n38165_, new_n38166_, new_n38168_,
    new_n38169_, new_n38170_, new_n38171_, new_n38172_, new_n38173_,
    new_n38174_, new_n38175_, new_n38176_, new_n38177_, new_n38178_,
    new_n38179_, new_n38180_, new_n38181_, new_n38183_, new_n38184_,
    new_n38185_, new_n38186_, new_n38187_, new_n38188_, new_n38189_,
    new_n38190_, new_n38191_, new_n38192_, new_n38193_, new_n38194_,
    new_n38195_, new_n38196_, new_n38198_, new_n38199_, new_n38200_,
    new_n38201_, new_n38202_, new_n38203_, new_n38204_, new_n38205_,
    new_n38206_, new_n38207_, new_n38208_, new_n38209_, new_n38210_,
    new_n38211_, new_n38213_, new_n38214_, new_n38215_, new_n38216_,
    new_n38217_, new_n38218_, new_n38219_, new_n38220_, new_n38221_,
    new_n38222_, new_n38223_, new_n38224_, new_n38225_, new_n38226_,
    new_n38228_, new_n38229_, new_n38230_, new_n38231_, new_n38232_,
    new_n38233_, new_n38234_, new_n38235_, new_n38236_, new_n38237_,
    new_n38238_, new_n38239_, new_n38240_, new_n38241_, new_n38243_,
    new_n38244_, new_n38245_, new_n38246_, new_n38247_, new_n38248_,
    new_n38249_, new_n38250_, new_n38251_, new_n38253_, new_n38254_,
    new_n38256_, new_n38257_, new_n38259_, new_n38260_, new_n38262_,
    new_n38263_, new_n38265_, new_n38266_, new_n38268_, new_n38269_,
    new_n38271_, new_n38272_, new_n38274_, new_n38275_, new_n38277_,
    new_n38278_, new_n38280_, new_n38281_, new_n38283_, new_n38284_,
    new_n38286_, new_n38287_, new_n38289_, new_n38290_, new_n38292_,
    new_n38293_, new_n38295_, new_n38296_, new_n38298_, new_n38299_,
    new_n38301_, new_n38302_, new_n38304_, new_n38305_, new_n38307_,
    new_n38308_, new_n38310_, new_n38311_, new_n38313_, new_n38314_,
    new_n38316_, new_n38317_, new_n38319_, new_n38320_, new_n38322_,
    new_n38323_, new_n38325_, new_n38326_, new_n38328_, new_n38329_,
    new_n38331_, new_n38332_, new_n38334_, new_n38335_, new_n38337_,
    new_n38338_, new_n38340_, new_n38341_, new_n38343_, new_n38344_,
    new_n38346_, new_n38347_, new_n38349_, new_n38350_, new_n38354_,
    new_n38355_, new_n38356_, new_n38357_, new_n38358_, new_n38367_,
    new_n38369_, new_n38370_, new_n38372_, new_n38373_, new_n38374_,
    new_n38375_, new_n38377_, new_n38378_, new_n38380_, new_n38381_,
    new_n38382_, new_n38383_, new_n38384_, new_n38385_, new_n38386_,
    new_n38387_, new_n38388_, new_n38389_, new_n38391_, new_n38392_,
    new_n38393_, new_n38394_, new_n38395_, new_n38396_, new_n38397_,
    new_n38399_, new_n38400_, new_n38401_, new_n38402_, new_n38403_,
    new_n38404_, new_n38405_, new_n38407_, new_n38408_, new_n38409_,
    new_n38410_, new_n38411_, new_n38412_, new_n38413_, new_n38415_,
    new_n38416_, new_n38417_, new_n38418_, new_n38419_, new_n38420_,
    new_n38421_, new_n38423_, new_n38424_, new_n38425_, new_n38426_,
    new_n38427_, new_n38428_, new_n38429_, new_n38431_, new_n38432_,
    new_n38433_, new_n38434_, new_n38435_, new_n38436_, new_n38437_,
    new_n38439_, new_n38440_, new_n38441_, new_n38442_, new_n38443_,
    new_n38444_, new_n38445_, new_n38447_, new_n38448_, new_n38449_,
    new_n38450_, new_n38451_, new_n38452_, new_n38453_, new_n38455_,
    new_n38456_, new_n38457_, new_n38458_, new_n38459_, new_n38460_,
    new_n38461_, new_n38463_, new_n38464_, new_n38465_, new_n38466_,
    new_n38467_, new_n38468_, new_n38469_, new_n38471_, new_n38472_,
    new_n38473_, new_n38474_, new_n38475_, new_n38476_, new_n38477_,
    new_n38479_, new_n38480_, new_n38481_, new_n38482_, new_n38483_,
    new_n38484_, new_n38485_, new_n38487_, new_n38488_, new_n38489_,
    new_n38490_, new_n38491_, new_n38492_, new_n38493_, new_n38495_,
    new_n38496_, new_n38497_, new_n38498_, new_n38499_, new_n38500_,
    new_n38501_, new_n38503_, new_n38504_, new_n38505_, new_n38506_,
    new_n38507_, new_n38508_, new_n38509_, new_n38511_, new_n38512_,
    new_n38513_, new_n38514_, new_n38515_, new_n38516_, new_n38517_,
    new_n38519_, new_n38520_, new_n38521_, new_n38522_, new_n38523_,
    new_n38524_, new_n38525_, new_n38527_, new_n38528_, new_n38529_,
    new_n38530_, new_n38531_, new_n38532_, new_n38533_, new_n38535_,
    new_n38536_, new_n38537_, new_n38538_, new_n38539_, new_n38540_,
    new_n38541_, new_n38543_, new_n38544_, new_n38545_, new_n38546_,
    new_n38547_, new_n38548_, new_n38549_, new_n38551_, new_n38552_,
    new_n38553_, new_n38554_, new_n38555_, new_n38556_, new_n38557_,
    new_n38559_, new_n38560_, new_n38561_, new_n38562_, new_n38563_,
    new_n38564_, new_n38565_, new_n38567_, new_n38568_, new_n38569_,
    new_n38570_, new_n38571_, new_n38572_, new_n38573_, new_n38575_,
    new_n38576_, new_n38577_, new_n38578_, new_n38579_, new_n38580_,
    new_n38581_, new_n38583_, new_n38584_, new_n38585_, new_n38586_,
    new_n38587_, new_n38588_, new_n38589_, new_n38591_, new_n38592_,
    new_n38593_, new_n38594_, new_n38595_, new_n38596_, new_n38597_,
    new_n38599_, new_n38600_, new_n38601_, new_n38602_, new_n38603_,
    new_n38604_, new_n38605_, new_n38607_, new_n38608_, new_n38609_,
    new_n38610_, new_n38611_, new_n38612_, new_n38613_, new_n38615_,
    new_n38616_, new_n38617_, new_n38618_, new_n38619_, new_n38620_,
    new_n38621_, new_n38623_, new_n38624_, new_n38625_, new_n38626_,
    new_n38627_, new_n38628_, new_n38629_, new_n38631_, new_n38632_,
    new_n38633_, new_n38634_, new_n38635_, new_n38636_, new_n38637_,
    new_n38639_, new_n38640_, new_n38641_, new_n38642_, new_n38643_,
    new_n38644_, new_n38645_, new_n38646_, new_n38648_, new_n38649_,
    new_n38651_, new_n38652_, new_n38654_, new_n38655_, new_n38657_,
    new_n38658_, new_n38660_, new_n38661_, new_n38663_, new_n38664_,
    new_n38666_, new_n38667_, new_n38669_, new_n38670_, new_n38672_,
    new_n38673_, new_n38675_, new_n38676_, new_n38678_, new_n38679_,
    new_n38681_, new_n38682_, new_n38684_, new_n38685_, new_n38687_,
    new_n38688_, new_n38690_, new_n38691_, new_n38693_, new_n38694_,
    new_n38696_, new_n38697_, new_n38699_, new_n38700_, new_n38702_,
    new_n38703_, new_n38705_, new_n38706_, new_n38708_, new_n38709_,
    new_n38711_, new_n38712_, new_n38714_, new_n38715_, new_n38717_,
    new_n38718_, new_n38720_, new_n38721_, new_n38723_, new_n38724_,
    new_n38726_, new_n38727_, new_n38729_, new_n38730_, new_n38732_,
    new_n38733_, new_n38735_, new_n38736_, new_n38738_, new_n38739_,
    new_n38741_, new_n38742_, new_n38744_, new_n38745_, new_n38749_,
    new_n38750_, new_n38751_, new_n38752_, new_n38761_, new_n38763_,
    new_n38764_, new_n38766_, new_n38767_, new_n38768_, new_n38769_,
    new_n38771_, new_n38772_, new_n38774_, new_n38775_, new_n38776_,
    new_n38777_, new_n38778_, new_n38779_, new_n38780_, new_n38781_,
    new_n38782_, new_n38783_, new_n38785_, new_n38786_, new_n38787_,
    new_n38788_, new_n38789_, new_n38790_, new_n38791_, new_n38793_,
    new_n38794_, new_n38795_, new_n38796_, new_n38797_, new_n38798_,
    new_n38799_, new_n38801_, new_n38802_, new_n38803_, new_n38804_,
    new_n38805_, new_n38806_, new_n38807_, new_n38809_, new_n38810_,
    new_n38811_, new_n38812_, new_n38813_, new_n38814_, new_n38815_,
    new_n38817_, new_n38818_, new_n38819_, new_n38820_, new_n38821_,
    new_n38822_, new_n38823_, new_n38825_, new_n38826_, new_n38827_,
    new_n38828_, new_n38829_, new_n38830_, new_n38831_, new_n38833_,
    new_n38834_, new_n38835_, new_n38836_, new_n38837_, new_n38838_,
    new_n38839_, new_n38841_, new_n38842_, new_n38843_, new_n38844_,
    new_n38845_, new_n38846_, new_n38847_, new_n38849_, new_n38850_,
    new_n38851_, new_n38852_, new_n38853_, new_n38854_, new_n38855_,
    new_n38857_, new_n38858_, new_n38859_, new_n38860_, new_n38861_,
    new_n38862_, new_n38863_, new_n38865_, new_n38866_, new_n38867_,
    new_n38868_, new_n38869_, new_n38870_, new_n38871_, new_n38873_,
    new_n38874_, new_n38875_, new_n38876_, new_n38877_, new_n38878_,
    new_n38879_, new_n38881_, new_n38882_, new_n38883_, new_n38884_,
    new_n38885_, new_n38886_, new_n38887_, new_n38889_, new_n38890_,
    new_n38891_, new_n38892_, new_n38893_, new_n38894_, new_n38895_,
    new_n38897_, new_n38898_, new_n38899_, new_n38900_, new_n38901_,
    new_n38902_, new_n38903_, new_n38905_, new_n38906_, new_n38907_,
    new_n38908_, new_n38909_, new_n38910_, new_n38911_, new_n38913_,
    new_n38914_, new_n38915_, new_n38916_, new_n38917_, new_n38918_,
    new_n38919_, new_n38921_, new_n38922_, new_n38923_, new_n38924_,
    new_n38925_, new_n38926_, new_n38927_, new_n38929_, new_n38930_,
    new_n38931_, new_n38932_, new_n38933_, new_n38934_, new_n38935_,
    new_n38937_, new_n38938_, new_n38939_, new_n38940_, new_n38941_,
    new_n38942_, new_n38943_, new_n38945_, new_n38946_, new_n38947_,
    new_n38948_, new_n38949_, new_n38950_, new_n38951_, new_n38953_,
    new_n38954_, new_n38955_, new_n38956_, new_n38957_, new_n38958_,
    new_n38959_, new_n38961_, new_n38962_, new_n38963_, new_n38964_,
    new_n38965_, new_n38966_, new_n38967_, new_n38969_, new_n38970_,
    new_n38971_, new_n38972_, new_n38973_, new_n38974_, new_n38975_,
    new_n38977_, new_n38978_, new_n38979_, new_n38980_, new_n38981_,
    new_n38982_, new_n38983_, new_n38985_, new_n38986_, new_n38987_,
    new_n38988_, new_n38989_, new_n38990_, new_n38991_, new_n38993_,
    new_n38994_, new_n38995_, new_n38996_, new_n38997_, new_n38998_,
    new_n38999_, new_n39001_, new_n39002_, new_n39003_, new_n39004_,
    new_n39005_, new_n39006_, new_n39007_, new_n39009_, new_n39010_,
    new_n39011_, new_n39012_, new_n39013_, new_n39014_, new_n39015_,
    new_n39017_, new_n39018_, new_n39019_, new_n39020_, new_n39021_,
    new_n39022_, new_n39023_, new_n39025_, new_n39026_, new_n39027_,
    new_n39028_, new_n39029_, new_n39030_, new_n39031_, new_n39033_,
    new_n39034_, new_n39035_, new_n39036_, new_n39037_, new_n39038_,
    new_n39039_, new_n39040_, new_n39042_, new_n39043_, new_n39045_,
    new_n39046_, new_n39048_, new_n39049_, new_n39051_, new_n39052_,
    new_n39054_, new_n39055_, new_n39057_, new_n39058_, new_n39060_,
    new_n39061_, new_n39063_, new_n39064_, new_n39066_, new_n39067_,
    new_n39069_, new_n39070_, new_n39072_, new_n39073_, new_n39075_,
    new_n39076_, new_n39078_, new_n39079_, new_n39081_, new_n39082_,
    new_n39084_, new_n39085_, new_n39087_, new_n39088_, new_n39090_,
    new_n39091_, new_n39093_, new_n39094_, new_n39096_, new_n39097_,
    new_n39099_, new_n39100_, new_n39102_, new_n39103_, new_n39105_,
    new_n39106_, new_n39108_, new_n39109_, new_n39111_, new_n39112_,
    new_n39114_, new_n39115_, new_n39117_, new_n39118_, new_n39120_,
    new_n39121_, new_n39123_, new_n39124_, new_n39126_, new_n39127_,
    new_n39129_, new_n39130_, new_n39132_, new_n39133_, new_n39135_,
    new_n39136_, new_n39138_, new_n39139_, new_n39143_, new_n39144_,
    new_n39145_, new_n39146_, new_n39155_, new_n39157_, new_n39158_,
    new_n39160_, new_n39161_, new_n39162_, new_n39163_, new_n39165_,
    new_n39166_, new_n39168_, new_n39169_, new_n39171_, new_n39172_,
    new_n39174_, new_n39176_, new_n39177_, new_n39179_, new_n39180_,
    new_n39182_, new_n39183_, new_n39185_, new_n39186_, new_n39188_,
    new_n39189_, new_n39191_, new_n39192_, new_n39194_, new_n39195_,
    new_n39197_, new_n39198_, new_n39200_, new_n39201_, new_n39203_,
    new_n39204_, new_n39206_, new_n39207_, new_n39209_, new_n39210_,
    new_n39212_, new_n39213_, new_n39215_, new_n39216_, new_n39218_,
    new_n39219_, new_n39221_, new_n39222_, new_n39224_, new_n39225_,
    new_n39227_, new_n39228_, new_n39230_, new_n39231_, new_n39233_,
    new_n39234_, new_n39236_, new_n39237_, new_n39239_, new_n39240_,
    new_n39242_, new_n39243_, new_n39245_, new_n39246_, new_n39248_,
    new_n39249_, new_n39251_, new_n39252_, new_n39254_, new_n39255_,
    new_n39257_, new_n39258_, new_n39260_, new_n39261_, new_n39263_,
    new_n39264_, new_n39266_, new_n39267_, new_n39269_, new_n39270_,
    new_n39271_, new_n39272_, new_n39273_, new_n39274_, new_n39276_,
    new_n39277_, new_n39278_, new_n39279_, new_n39280_, new_n39282_,
    new_n39283_, new_n39284_, new_n39285_, new_n39286_, new_n39288_,
    new_n39289_, new_n39290_, new_n39291_, new_n39292_, new_n39294_,
    new_n39295_, new_n39296_, new_n39297_, new_n39298_, new_n39300_,
    new_n39301_, new_n39302_, new_n39303_, new_n39304_, new_n39306_,
    new_n39307_, new_n39308_, new_n39309_, new_n39310_, new_n39312_,
    new_n39313_, new_n39314_, new_n39315_, new_n39316_, new_n39318_,
    new_n39319_, new_n39320_, new_n39321_, new_n39322_, new_n39324_,
    new_n39325_, new_n39326_, new_n39327_, new_n39328_, new_n39330_,
    new_n39331_, new_n39332_, new_n39333_, new_n39334_, new_n39336_,
    new_n39337_, new_n39338_, new_n39339_, new_n39340_, new_n39342_,
    new_n39343_, new_n39344_, new_n39345_, new_n39346_, new_n39348_,
    new_n39349_, new_n39350_, new_n39351_, new_n39352_, new_n39354_,
    new_n39355_, new_n39356_, new_n39357_, new_n39358_, new_n39360_,
    new_n39361_, new_n39362_, new_n39363_, new_n39364_, new_n39366_,
    new_n39367_, new_n39368_, new_n39369_, new_n39370_, new_n39372_,
    new_n39373_, new_n39374_, new_n39375_, new_n39376_, new_n39378_,
    new_n39379_, new_n39380_, new_n39381_, new_n39382_, new_n39384_,
    new_n39385_, new_n39386_, new_n39387_, new_n39388_, new_n39390_,
    new_n39391_, new_n39392_, new_n39393_, new_n39394_, new_n39396_,
    new_n39397_, new_n39398_, new_n39399_, new_n39400_, new_n39402_,
    new_n39403_, new_n39404_, new_n39405_, new_n39406_, new_n39408_,
    new_n39409_, new_n39410_, new_n39411_, new_n39412_, new_n39414_,
    new_n39415_, new_n39416_, new_n39417_, new_n39418_, new_n39420_,
    new_n39421_, new_n39422_, new_n39423_, new_n39424_, new_n39426_,
    new_n39427_, new_n39428_, new_n39429_, new_n39430_, new_n39432_,
    new_n39433_, new_n39434_, new_n39435_, new_n39436_, new_n39438_,
    new_n39439_, new_n39440_, new_n39441_, new_n39442_, new_n39444_,
    new_n39445_, new_n39446_, new_n39447_, new_n39448_, new_n39450_,
    new_n39451_, new_n39452_, new_n39453_, new_n39454_, new_n39456_,
    new_n39457_, new_n39458_, new_n39459_, new_n39460_, new_n39462_,
    new_n39463_, new_n39464_, new_n39467_, new_n39469_, new_n39470_,
    new_n39471_, new_n39472_, new_n39473_, new_n39474_, new_n39475_,
    new_n39476_, new_n39477_, new_n39478_, new_n39479_, new_n39480_,
    new_n39481_, new_n39482_, new_n39483_, new_n39484_, new_n39485_,
    new_n39486_, new_n39487_, new_n39488_, new_n39489_, new_n39490_,
    new_n39491_, new_n39492_, new_n39493_, new_n39494_, new_n39495_,
    new_n39496_, new_n39497_, new_n39498_, new_n39499_, new_n39500_,
    new_n39501_, new_n39502_, new_n39503_, new_n39504_, new_n39505_,
    new_n39506_, new_n39507_, new_n39508_, new_n39509_, new_n39510_,
    new_n39511_, new_n39512_, new_n39513_, new_n39514_, new_n39515_,
    new_n39516_, new_n39517_, new_n39518_, new_n39519_, new_n39520_,
    new_n39521_, new_n39522_, new_n39523_, new_n39524_, new_n39525_,
    new_n39526_, new_n39527_, new_n39528_, new_n39529_, new_n39530_,
    new_n39531_, new_n39532_, new_n39533_, new_n39534_, new_n39535_,
    new_n39536_, new_n39537_, new_n39538_, new_n39539_, new_n39540_,
    new_n39541_, new_n39542_, new_n39543_, new_n39544_, new_n39545_,
    new_n39546_, new_n39547_, new_n39548_, new_n39549_, new_n39550_,
    new_n39551_, new_n39552_, new_n39553_, new_n39554_, new_n39555_,
    new_n39556_, new_n39557_, new_n39558_, new_n39559_, new_n39560_,
    new_n39561_, new_n39562_, new_n39563_, new_n39564_, new_n39565_,
    new_n39566_, new_n39567_, new_n39568_, new_n39569_, new_n39570_,
    new_n39571_, new_n39572_, new_n39573_, new_n39574_, new_n39575_,
    new_n39576_, new_n39577_, new_n39578_, new_n39579_, new_n39580_,
    new_n39581_, new_n39582_, new_n39583_, new_n39584_, new_n39585_,
    new_n39586_, new_n39587_, new_n39588_, new_n39589_, new_n39590_,
    new_n39591_, new_n39592_, new_n39593_, new_n39594_, new_n39595_,
    new_n39596_, new_n39597_, new_n39598_, new_n39599_, new_n39600_,
    new_n39601_, new_n39602_, new_n39603_, new_n39604_, new_n39605_,
    new_n39606_, new_n39607_, new_n39608_, new_n39609_, new_n39610_,
    new_n39611_, new_n39612_, new_n39613_, new_n39614_, new_n39615_,
    new_n39616_, new_n39617_, new_n39618_, new_n39619_, new_n39620_,
    new_n39621_, new_n39622_, new_n39623_, new_n39624_, new_n39625_,
    new_n39626_, new_n39627_, new_n39628_, new_n39629_, new_n39630_,
    new_n39631_, new_n39632_, new_n39633_, new_n39634_, new_n39635_,
    new_n39636_, new_n39637_, new_n39638_, new_n39639_, new_n39640_,
    new_n39641_, new_n39642_, new_n39643_, new_n39644_, new_n39645_,
    new_n39646_, new_n39647_, new_n39648_, new_n39649_, new_n39650_,
    new_n39651_, new_n39652_, new_n39653_, new_n39654_, new_n39655_,
    new_n39656_, new_n39657_, new_n39658_, new_n39659_, new_n39660_,
    new_n39661_, new_n39662_, new_n39663_, new_n39664_, new_n39665_,
    new_n39666_, new_n39667_, new_n39668_, new_n39669_, new_n39670_,
    new_n39671_, new_n39672_, new_n39673_, new_n39674_, new_n39675_,
    new_n39676_, new_n39677_, new_n39678_, new_n39679_, new_n39680_,
    new_n39681_, new_n39682_, new_n39683_, new_n39684_, new_n39685_,
    new_n39686_, new_n39687_, new_n39688_, new_n39689_, new_n39690_,
    new_n39691_, new_n39692_, new_n39693_, new_n39694_, new_n39695_,
    new_n39696_, new_n39697_, new_n39698_, new_n39699_, new_n39700_,
    new_n39701_, new_n39702_, new_n39703_, new_n39704_, new_n39705_,
    new_n39706_, new_n39707_, new_n39708_, new_n39709_, new_n39710_,
    new_n39711_, new_n39712_, new_n39713_, new_n39714_, new_n39715_,
    new_n39716_, new_n39717_, new_n39718_, new_n39719_, new_n39720_,
    new_n39721_, new_n39722_, new_n39723_, new_n39724_, new_n39725_,
    new_n39726_, new_n39727_, new_n39728_, new_n39729_, new_n39730_,
    new_n39731_, new_n39732_, new_n39733_, new_n39734_, new_n39735_,
    new_n39736_, new_n39737_, new_n39738_, new_n39739_, new_n39740_,
    new_n39741_, new_n39742_, new_n39743_, new_n39744_, new_n39745_,
    new_n39746_, new_n39747_, new_n39748_, new_n39749_, new_n39750_,
    new_n39751_, new_n39752_, new_n39753_, new_n39754_, new_n39755_,
    new_n39756_, new_n39757_, new_n39758_, new_n39759_, new_n39760_,
    new_n39761_, new_n39762_, new_n39763_, new_n39764_, new_n39765_,
    new_n39766_, new_n39767_, new_n39768_, new_n39769_, new_n39770_,
    new_n39771_, new_n39772_, new_n39773_, new_n39774_, new_n39775_,
    new_n39776_, new_n39777_, new_n39778_, new_n39779_, new_n39780_,
    new_n39781_, new_n39782_, new_n39783_, new_n39784_, new_n39785_,
    new_n39786_, new_n39787_, new_n39788_, new_n39789_, new_n39790_,
    new_n39791_, new_n39792_, new_n39793_, new_n39794_, new_n39795_,
    new_n39796_, new_n39797_, new_n39798_, new_n39799_, new_n39800_,
    new_n39801_, new_n39802_, new_n39803_, new_n39804_, new_n39805_,
    new_n39806_, new_n39807_, new_n39808_, new_n39809_, new_n39810_,
    new_n39811_, new_n39812_, new_n39813_, new_n39814_, new_n39815_,
    new_n39816_, new_n39817_, new_n39818_, new_n39819_, new_n39820_,
    new_n39821_, new_n39822_, new_n39823_, new_n39824_, new_n39825_,
    new_n39826_, new_n39827_, new_n39828_, new_n39829_, new_n39830_,
    new_n39831_, new_n39832_, new_n39833_, new_n39834_, new_n39835_,
    new_n39836_, new_n39837_, new_n39838_, new_n39839_, new_n39840_,
    new_n39841_, new_n39842_, new_n39843_, new_n39844_, new_n39845_,
    new_n39846_, new_n39847_, new_n39848_, new_n39849_, new_n39850_,
    new_n39851_, new_n39852_, new_n39853_, new_n39854_, new_n39855_,
    new_n39856_, new_n39857_, new_n39858_, new_n39859_, new_n39860_,
    new_n39861_, new_n39862_, new_n39863_, new_n39864_, new_n39865_,
    new_n39866_, new_n39867_, new_n39868_, new_n39869_, new_n39870_,
    new_n39871_, new_n39872_, new_n39873_, new_n39874_, new_n39875_,
    new_n39876_, new_n39877_, new_n39878_, new_n39879_, new_n39880_,
    new_n39881_, new_n39882_, new_n39883_, new_n39884_, new_n39885_,
    new_n39886_, new_n39887_, new_n39888_, new_n39889_, new_n39890_,
    new_n39891_, new_n39892_, new_n39893_, new_n39894_, new_n39895_,
    new_n39896_, new_n39897_, new_n39898_, new_n39899_, new_n39900_,
    new_n39901_, new_n39902_, new_n39903_, new_n39904_, new_n39905_,
    new_n39906_, new_n39907_, new_n39908_, new_n39909_, new_n39910_,
    new_n39911_, new_n39912_, new_n39913_, new_n39914_, new_n39915_,
    new_n39916_, new_n39917_, new_n39918_, new_n39919_, new_n39920_,
    new_n39921_, new_n39922_, new_n39923_, new_n39924_, new_n39925_,
    new_n39926_, new_n39927_, new_n39928_, new_n39929_, new_n39930_,
    new_n39931_, new_n39932_, new_n39933_, new_n39934_, new_n39935_,
    new_n39936_, new_n39937_, new_n39938_, new_n39939_, new_n39940_,
    new_n39941_, new_n39942_, new_n39943_, new_n39944_, new_n39945_,
    new_n39946_, new_n39947_, new_n39948_, new_n39949_, new_n39950_,
    new_n39951_, new_n39952_, new_n39953_, new_n39954_, new_n39955_,
    new_n39956_, new_n39957_, new_n39958_, new_n39959_, new_n39960_,
    new_n39961_, new_n39962_, new_n39963_, new_n39964_, new_n39965_,
    new_n39966_, new_n39967_, new_n39968_, new_n39969_, new_n39970_,
    new_n39971_, new_n39972_, new_n39973_, new_n39974_, new_n39975_,
    new_n39976_, new_n39977_, new_n39978_, new_n39979_, new_n39980_,
    new_n39981_, new_n39982_, new_n39983_, new_n39984_, new_n39985_,
    new_n39986_, new_n39987_, new_n39988_, new_n39989_, new_n39990_,
    new_n39991_, new_n39992_, new_n39993_, new_n39994_, new_n39995_,
    new_n39996_, new_n39997_, new_n39998_, new_n39999_, new_n40000_,
    new_n40001_, new_n40002_, new_n40003_, new_n40004_, new_n40005_,
    new_n40006_, new_n40007_, new_n40008_, new_n40009_, new_n40010_,
    new_n40011_, new_n40012_, new_n40013_, new_n40014_, new_n40015_,
    new_n40016_, new_n40017_, new_n40018_, new_n40019_, new_n40020_,
    new_n40021_, new_n40022_, new_n40023_, new_n40024_, new_n40025_,
    new_n40026_, new_n40027_, new_n40028_, new_n40029_, new_n40030_,
    new_n40031_, new_n40032_, new_n40033_, new_n40034_, new_n40035_,
    new_n40036_, new_n40037_, new_n40038_, new_n40039_, new_n40040_,
    new_n40041_, new_n40042_, new_n40043_, new_n40044_, new_n40045_,
    new_n40046_, new_n40047_, new_n40048_, new_n40049_, new_n40050_,
    new_n40051_, new_n40052_, new_n40053_, new_n40054_, new_n40055_,
    new_n40056_, new_n40057_, new_n40058_, new_n40059_, new_n40060_,
    new_n40061_, new_n40062_, new_n40063_, new_n40064_, new_n40065_,
    new_n40066_, new_n40067_, new_n40068_, new_n40069_, new_n40070_,
    new_n40071_, new_n40072_, new_n40073_, new_n40074_, new_n40075_,
    new_n40076_, new_n40077_, new_n40078_, new_n40079_, new_n40080_,
    new_n40081_, new_n40082_, new_n40083_, new_n40084_, new_n40085_,
    new_n40086_, new_n40087_, new_n40088_, new_n40089_, new_n40090_,
    new_n40091_, new_n40092_, new_n40093_, new_n40094_, new_n40095_,
    new_n40096_, new_n40097_, new_n40098_, new_n40099_, new_n40100_,
    new_n40101_, new_n40102_, new_n40103_, new_n40104_, new_n40105_,
    new_n40106_, new_n40107_, new_n40108_, new_n40109_, new_n40110_,
    new_n40111_, new_n40112_, new_n40113_, new_n40114_, new_n40115_,
    new_n40116_, new_n40117_, new_n40118_, new_n40119_, new_n40120_,
    new_n40121_, new_n40122_, new_n40123_, new_n40124_, new_n40125_,
    new_n40126_, new_n40127_, new_n40128_, new_n40129_, new_n40130_,
    new_n40131_, new_n40132_, new_n40133_, new_n40134_, new_n40135_,
    new_n40136_, new_n40137_, new_n40138_, new_n40139_, new_n40140_,
    new_n40141_, new_n40142_, new_n40143_, new_n40144_, new_n40145_,
    new_n40146_, new_n40147_, new_n40148_, new_n40149_, new_n40150_,
    new_n40151_, new_n40152_, new_n40153_, new_n40154_, new_n40155_,
    new_n40156_, new_n40157_, new_n40158_, new_n40159_, new_n40160_,
    new_n40161_, new_n40162_, new_n40163_, new_n40164_, new_n40165_,
    new_n40166_, new_n40167_, new_n40168_, new_n40169_, new_n40170_,
    new_n40171_, new_n40172_, new_n40173_, new_n40174_, new_n40175_,
    new_n40176_, new_n40177_, new_n40178_, new_n40179_, new_n40180_,
    new_n40181_, new_n40182_, new_n40183_, new_n40184_, new_n40185_,
    new_n40186_, new_n40187_, new_n40188_, new_n40189_, new_n40190_,
    new_n40191_, new_n40192_, new_n40193_, new_n40194_, new_n40195_,
    new_n40196_, new_n40197_, new_n40198_, new_n40199_, new_n40200_,
    new_n40201_, new_n40202_, new_n40203_, new_n40204_, new_n40205_,
    new_n40206_, new_n40207_, new_n40208_, new_n40209_, new_n40210_,
    new_n40211_, new_n40212_, new_n40213_, new_n40214_, new_n40215_,
    new_n40216_, new_n40217_, new_n40218_, new_n40219_, new_n40220_,
    new_n40221_, new_n40222_, new_n40223_, new_n40224_, new_n40225_,
    new_n40226_, new_n40227_, new_n40228_, new_n40229_, new_n40230_,
    new_n40231_, new_n40232_, new_n40233_, new_n40234_, new_n40235_,
    new_n40236_, new_n40237_, new_n40238_, new_n40239_, new_n40240_,
    new_n40241_, new_n40242_, new_n40243_, new_n40244_, new_n40245_,
    new_n40246_, new_n40247_, new_n40248_, new_n40249_, new_n40250_,
    new_n40251_, new_n40252_, new_n40253_, new_n40254_, new_n40255_,
    new_n40256_, new_n40257_, new_n40258_, new_n40259_, new_n40260_,
    new_n40261_, new_n40262_, new_n40263_, new_n40264_, new_n40265_,
    new_n40266_, new_n40267_, new_n40268_, new_n40269_, new_n40270_,
    new_n40271_, new_n40272_, new_n40273_, new_n40274_, new_n40275_,
    new_n40276_, new_n40277_, new_n40278_, new_n40279_, new_n40280_,
    new_n40281_, new_n40282_, new_n40283_, new_n40284_, new_n40285_,
    new_n40286_, new_n40287_, new_n40288_, new_n40289_, new_n40290_,
    new_n40291_, new_n40292_, new_n40293_, new_n40294_, new_n40295_,
    new_n40296_, new_n40297_, new_n40298_, new_n40299_, new_n40300_,
    new_n40301_, new_n40302_, new_n40303_, new_n40304_, new_n40305_,
    new_n40306_, new_n40307_, new_n40308_, new_n40309_, new_n40310_,
    new_n40311_, new_n40312_, new_n40313_, new_n40314_, new_n40315_,
    new_n40316_, new_n40317_, new_n40318_, new_n40319_, new_n40320_,
    new_n40321_, new_n40322_, new_n40323_, new_n40324_, new_n40325_,
    new_n40326_, new_n40327_, new_n40328_, new_n40329_, new_n40330_,
    new_n40331_, new_n40332_, new_n40333_, new_n40334_, new_n40335_,
    new_n40336_, new_n40337_, new_n40338_, new_n40339_, new_n40340_,
    new_n40341_, new_n40342_, new_n40343_, new_n40344_, new_n40345_,
    new_n40346_, new_n40347_, new_n40348_, new_n40349_, new_n40350_,
    new_n40351_, new_n40352_, new_n40353_, new_n40354_, new_n40355_,
    new_n40356_, new_n40357_, new_n40358_, new_n40359_, new_n40360_,
    new_n40361_, new_n40362_, new_n40363_, new_n40364_, new_n40365_,
    new_n40366_, new_n40367_, new_n40368_, new_n40369_, new_n40370_,
    new_n40371_, new_n40372_, new_n40373_, new_n40374_, new_n40375_,
    new_n40376_, new_n40377_, new_n40378_, new_n40379_, new_n40380_,
    new_n40381_, new_n40382_, new_n40383_, new_n40384_, new_n40385_,
    new_n40386_, new_n40387_, new_n40388_, new_n40389_, new_n40390_,
    new_n40391_, new_n40392_, new_n40393_, new_n40394_, new_n40395_,
    new_n40396_, new_n40397_, new_n40398_, new_n40399_, new_n40400_,
    new_n40401_, new_n40402_, new_n40403_, new_n40404_, new_n40405_,
    new_n40406_, new_n40407_, new_n40408_, new_n40409_, new_n40410_,
    new_n40411_, new_n40412_, new_n40413_, new_n40414_, new_n40415_,
    new_n40416_, new_n40417_, new_n40418_, new_n40419_, new_n40420_,
    new_n40421_, new_n40422_, new_n40423_, new_n40424_, new_n40425_,
    new_n40426_, new_n40427_, new_n40428_, new_n40429_, new_n40430_,
    new_n40431_, new_n40432_, new_n40433_, new_n40434_, new_n40435_,
    new_n40436_, new_n40437_, new_n40438_, new_n40439_, new_n40440_,
    new_n40441_, new_n40442_, new_n40443_, new_n40444_, new_n40445_,
    new_n40446_, new_n40447_, new_n40448_, new_n40449_, new_n40450_,
    new_n40451_, new_n40452_, new_n40453_, new_n40454_, new_n40455_,
    new_n40456_, new_n40457_, new_n40458_, new_n40459_, new_n40460_,
    new_n40461_, new_n40462_, new_n40463_, new_n40464_, new_n40465_,
    new_n40466_, new_n40467_, new_n40468_, new_n40469_, new_n40470_,
    new_n40471_, new_n40472_, new_n40473_, new_n40474_, new_n40475_,
    new_n40476_, new_n40477_, new_n40478_, new_n40479_, new_n40480_,
    new_n40481_, new_n40482_, new_n40483_, new_n40484_, new_n40485_,
    new_n40486_, new_n40487_, new_n40488_, new_n40489_, new_n40490_,
    new_n40491_, new_n40492_, new_n40493_, new_n40494_, new_n40495_,
    new_n40496_, new_n40497_, new_n40498_, new_n40499_, new_n40500_,
    new_n40501_, new_n40502_, new_n40503_, new_n40504_, new_n40505_,
    new_n40506_, new_n40507_, new_n40508_, new_n40509_, new_n40510_,
    new_n40511_, new_n40512_, new_n40513_, new_n40514_, new_n40515_,
    new_n40516_, new_n40517_, new_n40518_, new_n40519_, new_n40520_,
    new_n40521_, new_n40522_, new_n40523_, new_n40524_, new_n40525_,
    new_n40526_, new_n40527_, new_n40528_, new_n40529_, new_n40530_,
    new_n40531_, new_n40532_, new_n40533_, new_n40534_, new_n40535_,
    new_n40536_, new_n40537_, new_n40538_, new_n40539_, new_n40540_,
    new_n40541_, new_n40542_, new_n40543_, new_n40544_, new_n40545_,
    new_n40546_, new_n40547_, new_n40548_, new_n40549_, new_n40550_,
    new_n40551_, new_n40552_, new_n40553_, new_n40554_, new_n40555_,
    new_n40556_, new_n40557_, new_n40558_, new_n40559_, new_n40560_,
    new_n40561_, new_n40562_, new_n40563_, new_n40564_, new_n40565_,
    new_n40566_, new_n40567_, new_n40568_, new_n40569_, new_n40570_,
    new_n40571_, new_n40572_, new_n40573_, new_n40574_, new_n40575_,
    new_n40576_, new_n40577_, new_n40578_, new_n40579_, new_n40580_,
    new_n40581_, new_n40582_, new_n40583_, new_n40584_, new_n40585_,
    new_n40586_, new_n40587_, new_n40588_, new_n40589_, new_n40590_,
    new_n40591_, new_n40592_, new_n40593_, new_n40594_, new_n40595_,
    new_n40596_, new_n40597_, new_n40598_, new_n40599_, new_n40600_,
    new_n40601_, new_n40602_, new_n40603_, new_n40604_, new_n40605_,
    new_n40606_, new_n40607_, new_n40608_, new_n40609_, new_n40610_,
    new_n40611_, new_n40612_, new_n40613_, new_n40614_, new_n40615_,
    new_n40616_, new_n40617_, new_n40618_, new_n40619_, new_n40620_,
    new_n40621_, new_n40622_, new_n40623_, new_n40624_, new_n40625_,
    new_n40626_, new_n40627_, new_n40628_, new_n40629_, new_n40630_,
    new_n40631_, new_n40632_, new_n40633_, new_n40634_, new_n40635_,
    new_n40636_, new_n40637_, new_n40638_, new_n40639_, new_n40640_,
    new_n40641_, new_n40642_, new_n40643_, new_n40644_, new_n40645_,
    new_n40646_, new_n40647_, new_n40648_, new_n40649_, new_n40650_,
    new_n40651_, new_n40652_, new_n40653_, new_n40654_, new_n40655_,
    new_n40656_, new_n40657_, new_n40658_, new_n40659_, new_n40660_,
    new_n40661_, new_n40662_, new_n40663_, new_n40664_, new_n40665_,
    new_n40666_, new_n40667_, new_n40668_, new_n40669_, new_n40670_,
    new_n40671_, new_n40672_, new_n40673_, new_n40674_, new_n40675_,
    new_n40676_, new_n40677_, new_n40678_, new_n40679_, new_n40680_,
    new_n40681_, new_n40682_, new_n40683_, new_n40684_, new_n40685_,
    new_n40686_, new_n40687_, new_n40688_, new_n40689_, new_n40690_,
    new_n40691_, new_n40692_, new_n40693_, new_n40694_, new_n40695_,
    new_n40696_, new_n40697_, new_n40698_, new_n40699_, new_n40700_,
    new_n40701_, new_n40702_, new_n40703_, new_n40704_, new_n40705_,
    new_n40706_, new_n40707_, new_n40708_, new_n40709_, new_n40710_,
    new_n40711_, new_n40712_, new_n40713_, new_n40714_, new_n40715_,
    new_n40716_, new_n40717_, new_n40718_, new_n40719_, new_n40720_,
    new_n40721_, new_n40722_, new_n40723_, new_n40724_, new_n40725_,
    new_n40726_, new_n40727_, new_n40728_, new_n40729_, new_n40730_,
    new_n40731_, new_n40732_, new_n40733_, new_n40734_, new_n40735_,
    new_n40736_, new_n40737_, new_n40738_, new_n40739_, new_n40740_,
    new_n40741_, new_n40742_, new_n40743_, new_n40744_, new_n40745_,
    new_n40746_, new_n40747_, new_n40748_, new_n40749_, new_n40750_,
    new_n40751_, new_n40752_, new_n40753_, new_n40754_, new_n40755_,
    new_n40756_, new_n40757_, new_n40758_, new_n40759_, new_n40760_,
    new_n40761_, new_n40762_, new_n40763_, new_n40764_, new_n40765_,
    new_n40766_, new_n40767_, new_n40768_, new_n40769_, new_n40770_,
    new_n40771_, new_n40772_, new_n40773_, new_n40774_, new_n40775_,
    new_n40776_, new_n40777_, new_n40778_, new_n40779_, new_n40780_,
    new_n40781_, new_n40782_, new_n40783_, new_n40784_, new_n40785_,
    new_n40786_, new_n40787_, new_n40788_, new_n40789_, new_n40790_,
    new_n40791_, new_n40792_, new_n40793_, new_n40794_, new_n40795_,
    new_n40796_, new_n40797_, new_n40798_, new_n40799_, new_n40800_,
    new_n40801_, new_n40802_, new_n40803_, new_n40804_, new_n40805_,
    new_n40806_, new_n40807_, new_n40808_, new_n40809_, new_n40810_,
    new_n40811_, new_n40812_, new_n40813_, new_n40814_, new_n40815_,
    new_n40816_, new_n40817_, new_n40818_, new_n40819_, new_n40820_,
    new_n40821_, new_n40822_, new_n40823_, new_n40824_, new_n40825_,
    new_n40826_, new_n40827_, new_n40828_, new_n40829_, new_n40830_,
    new_n40831_, new_n40832_, new_n40833_, new_n40834_, new_n40835_,
    new_n40836_, new_n40837_, new_n40838_, new_n40839_, new_n40840_,
    new_n40841_, new_n40842_, new_n40843_, new_n40844_, new_n40845_,
    new_n40846_, new_n40847_, new_n40848_, new_n40849_, new_n40850_,
    new_n40851_, new_n40852_, new_n40853_, new_n40854_, new_n40855_,
    new_n40856_, new_n40857_, new_n40858_, new_n40859_, new_n40860_,
    new_n40861_, new_n40862_, new_n40863_, new_n40864_, new_n40865_,
    new_n40866_, new_n40867_, new_n40868_, new_n40869_, new_n40870_,
    new_n40871_, new_n40872_, new_n40873_, new_n40874_, new_n40875_,
    new_n40876_, new_n40877_, new_n40878_, new_n40879_, new_n40880_,
    new_n40881_, new_n40882_, new_n40883_, new_n40884_, new_n40885_,
    new_n40886_, new_n40887_, new_n40888_, new_n40889_, new_n40890_,
    new_n40891_, new_n40892_, new_n40893_, new_n40894_, new_n40895_,
    new_n40896_, new_n40897_, new_n40898_, new_n40899_, new_n40900_,
    new_n40901_, new_n40902_, new_n40903_, new_n40904_, new_n40905_,
    new_n40906_, new_n40907_, new_n40908_, new_n40909_, new_n40910_,
    new_n40911_, new_n40912_, new_n40913_, new_n40914_, new_n40915_,
    new_n40916_, new_n40917_, new_n40918_, new_n40919_, new_n40920_,
    new_n40921_, new_n40922_, new_n40923_, new_n40924_, new_n40925_,
    new_n40926_, new_n40927_, new_n40928_, new_n40929_, new_n40930_,
    new_n40931_, new_n40932_, new_n40933_, new_n40934_, new_n40935_,
    new_n40936_, new_n40937_, new_n40938_, new_n40939_, new_n40940_,
    new_n40941_, new_n40942_, new_n40943_, new_n40944_, new_n40945_,
    new_n40946_, new_n40947_, new_n40948_, new_n40949_, new_n40950_,
    new_n40951_, new_n40952_, new_n40953_, new_n40954_, new_n40955_,
    new_n40956_, new_n40957_, new_n40958_, new_n40959_, new_n40960_,
    new_n40961_, new_n40962_, new_n40963_, new_n40964_, new_n40965_,
    new_n40966_, new_n40967_, new_n40968_, new_n40969_, new_n40970_,
    new_n40971_, new_n40972_, new_n40973_, new_n40974_, new_n40975_,
    new_n40976_, new_n40977_, new_n40978_, new_n40979_, new_n40980_,
    new_n40981_, new_n40982_, new_n40983_, new_n40984_, new_n40985_,
    new_n40986_, new_n40987_, new_n40988_, new_n40989_, new_n40990_,
    new_n40991_, new_n40992_, new_n40993_, new_n40994_, new_n40995_,
    new_n40996_, new_n40997_, new_n40998_, new_n40999_, new_n41000_,
    new_n41001_, new_n41002_, new_n41003_, new_n41004_, new_n41005_,
    new_n41006_, new_n41007_, new_n41008_, new_n41009_, new_n41010_,
    new_n41011_, new_n41012_, new_n41013_, new_n41014_, new_n41015_,
    new_n41016_, new_n41017_, new_n41018_, new_n41019_, new_n41020_,
    new_n41021_, new_n41022_, new_n41023_, new_n41024_, new_n41025_,
    new_n41026_, new_n41027_, new_n41028_, new_n41029_, new_n41030_,
    new_n41031_, new_n41032_, new_n41033_, new_n41034_, new_n41035_,
    new_n41036_, new_n41037_, new_n41038_, new_n41039_, new_n41040_,
    new_n41041_, new_n41042_, new_n41043_, new_n41044_, new_n41045_,
    new_n41046_, new_n41047_, new_n41048_, new_n41049_, new_n41050_,
    new_n41051_, new_n41052_, new_n41054_, new_n41055_, new_n41056_,
    new_n41057_, new_n41058_, new_n41059_, new_n41060_, new_n41061_,
    new_n41062_, new_n41063_, new_n41064_, new_n41065_, new_n41066_,
    new_n41067_, new_n41068_, new_n41069_, new_n41070_, new_n41071_,
    new_n41072_, new_n41073_, new_n41074_, new_n41075_, new_n41076_,
    new_n41077_, new_n41078_, new_n41079_, new_n41081_, new_n41082_,
    new_n41083_, new_n41084_, new_n41085_, new_n41086_, new_n41087_,
    new_n41088_, new_n41089_, new_n41090_, new_n41091_, new_n41092_,
    new_n41093_, new_n41094_, new_n41095_, new_n41096_, new_n41097_,
    new_n41098_, new_n41099_, new_n41100_, new_n41101_, new_n41102_,
    new_n41103_, new_n41104_, new_n41105_, new_n41107_, new_n41108_,
    new_n41109_, new_n41110_, new_n41111_, new_n41112_, new_n41113_,
    new_n41114_, new_n41115_, new_n41116_, new_n41117_, new_n41118_,
    new_n41119_, new_n41120_, new_n41121_, new_n41122_, new_n41123_,
    new_n41124_, new_n41125_, new_n41126_, new_n41127_, new_n41128_,
    new_n41129_, new_n41130_, new_n41131_, new_n41133_, new_n41134_,
    new_n41135_, new_n41136_, new_n41137_, new_n41138_, new_n41139_,
    new_n41140_, new_n41141_, new_n41142_, new_n41143_, new_n41144_,
    new_n41145_, new_n41146_, new_n41147_, new_n41148_, new_n41149_,
    new_n41150_, new_n41151_, new_n41152_, new_n41153_, new_n41154_,
    new_n41155_, new_n41156_, new_n41158_, new_n41159_, new_n41160_,
    new_n41161_, new_n41162_, new_n41163_, new_n41164_, new_n41165_,
    new_n41166_, new_n41167_, new_n41168_, new_n41169_, new_n41170_,
    new_n41171_, new_n41172_, new_n41173_, new_n41174_, new_n41175_,
    new_n41176_, new_n41177_, new_n41178_, new_n41179_, new_n41180_,
    new_n41181_, new_n41182_, new_n41183_, new_n41184_, new_n41186_,
    new_n41187_, new_n41188_, new_n41189_, new_n41190_, new_n41191_,
    new_n41192_, new_n41193_, new_n41194_, new_n41195_, new_n41196_,
    new_n41197_, new_n41198_, new_n41199_, new_n41200_, new_n41201_,
    new_n41202_, new_n41203_, new_n41204_, new_n41205_, new_n41206_,
    new_n41207_, new_n41208_, new_n41209_, new_n41210_, new_n41211_,
    new_n41212_, new_n41213_, new_n41215_, new_n41216_, new_n41217_,
    new_n41218_, new_n41219_, new_n41220_, new_n41221_, new_n41222_,
    new_n41223_, new_n41224_, new_n41225_, new_n41226_, new_n41227_,
    new_n41228_, new_n41229_, new_n41230_, new_n41231_, new_n41232_,
    new_n41233_, new_n41234_, new_n41235_, new_n41236_, new_n41237_,
    new_n41238_, new_n41239_, new_n41240_, new_n41241_, new_n41242_,
    new_n41244_, new_n41245_, new_n41246_, new_n41247_, new_n41248_,
    new_n41249_, new_n41250_, new_n41251_, new_n41252_, new_n41253_,
    new_n41254_, new_n41255_, new_n41256_, new_n41257_, new_n41258_,
    new_n41259_, new_n41260_, new_n41261_, new_n41262_, new_n41263_,
    new_n41264_, new_n41265_, new_n41266_, new_n41267_, new_n41268_,
    new_n41270_, new_n41271_, new_n41272_, new_n41273_, new_n41274_,
    new_n41275_, new_n41276_, new_n41277_, new_n41278_, new_n41279_,
    new_n41280_, new_n41281_, new_n41282_, new_n41283_, new_n41284_,
    new_n41285_, new_n41286_, new_n41287_, new_n41288_, new_n41289_,
    new_n41290_, new_n41291_, new_n41292_, new_n41293_, new_n41294_,
    new_n41295_, new_n41296_, new_n41298_, new_n41299_, new_n41300_,
    new_n41301_, new_n41302_, new_n41303_, new_n41304_, new_n41305_,
    new_n41306_, new_n41307_, new_n41308_, new_n41309_, new_n41310_,
    new_n41311_, new_n41312_, new_n41313_, new_n41314_, new_n41315_,
    new_n41316_, new_n41317_, new_n41318_, new_n41319_, new_n41320_,
    new_n41321_, new_n41322_, new_n41323_, new_n41324_, new_n41325_,
    new_n41327_, new_n41328_, new_n41329_, new_n41330_, new_n41331_,
    new_n41332_, new_n41333_, new_n41334_, new_n41335_, new_n41336_,
    new_n41337_, new_n41338_, new_n41339_, new_n41340_, new_n41341_,
    new_n41342_, new_n41343_, new_n41344_, new_n41345_, new_n41346_,
    new_n41347_, new_n41348_, new_n41349_, new_n41350_, new_n41351_,
    new_n41352_, new_n41353_, new_n41354_, new_n41356_, new_n41357_,
    new_n41358_, new_n41359_, new_n41360_, new_n41361_, new_n41362_,
    new_n41363_, new_n41364_, new_n41365_, new_n41366_, new_n41367_,
    new_n41368_, new_n41369_, new_n41370_, new_n41371_, new_n41372_,
    new_n41373_, new_n41374_, new_n41375_, new_n41376_, new_n41377_,
    new_n41378_, new_n41379_, new_n41380_, new_n41381_, new_n41382_,
    new_n41383_, new_n41385_, new_n41386_, new_n41387_, new_n41388_,
    new_n41389_, new_n41390_, new_n41391_, new_n41392_, new_n41393_,
    new_n41394_, new_n41395_, new_n41396_, new_n41397_, new_n41398_,
    new_n41399_, new_n41400_, new_n41401_, new_n41402_, new_n41403_,
    new_n41404_, new_n41405_, new_n41406_, new_n41407_, new_n41408_,
    new_n41409_, new_n41410_, new_n41411_, new_n41412_, new_n41414_,
    new_n41415_, new_n41416_, new_n41417_, new_n41418_, new_n41419_,
    new_n41420_, new_n41421_, new_n41422_, new_n41423_, new_n41424_,
    new_n41425_, new_n41426_, new_n41427_, new_n41428_, new_n41429_,
    new_n41430_, new_n41431_, new_n41432_, new_n41433_, new_n41434_,
    new_n41435_, new_n41436_, new_n41437_, new_n41438_, new_n41439_,
    new_n41440_, new_n41441_, new_n41443_, new_n41444_, new_n41445_,
    new_n41446_, new_n41447_, new_n41448_, new_n41449_, new_n41450_,
    new_n41451_, new_n41452_, new_n41453_, new_n41454_, new_n41455_,
    new_n41456_, new_n41457_, new_n41458_, new_n41459_, new_n41460_,
    new_n41461_, new_n41462_, new_n41463_, new_n41464_, new_n41465_,
    new_n41466_, new_n41467_, new_n41468_, new_n41469_, new_n41470_,
    new_n41472_, new_n41473_, new_n41474_, new_n41475_, new_n41476_,
    new_n41477_, new_n41478_, new_n41479_, new_n41480_, new_n41481_,
    new_n41482_, new_n41483_, new_n41484_, new_n41485_, new_n41486_,
    new_n41487_, new_n41488_, new_n41489_, new_n41490_, new_n41491_,
    new_n41492_, new_n41493_, new_n41494_, new_n41495_, new_n41496_,
    new_n41498_, new_n41499_, new_n41500_, new_n41501_, new_n41502_,
    new_n41503_, new_n41504_, new_n41505_, new_n41506_, new_n41507_,
    new_n41508_, new_n41509_, new_n41510_, new_n41511_, new_n41512_,
    new_n41513_, new_n41514_, new_n41515_, new_n41516_, new_n41517_,
    new_n41518_, new_n41519_, new_n41520_, new_n41521_, new_n41522_,
    new_n41523_, new_n41524_, new_n41525_, new_n41526_, new_n41527_,
    new_n41528_, new_n41530_, new_n41531_, new_n41532_, new_n41533_,
    new_n41534_, new_n41535_, new_n41536_, new_n41537_, new_n41538_,
    new_n41539_, new_n41540_, new_n41541_, new_n41542_, new_n41543_,
    new_n41544_, new_n41545_, new_n41546_, new_n41547_, new_n41548_,
    new_n41549_, new_n41550_, new_n41551_, new_n41552_, new_n41553_,
    new_n41554_, new_n41555_, new_n41556_, new_n41557_, new_n41558_,
    new_n41559_, new_n41560_, new_n41561_, new_n41562_, new_n41563_,
    new_n41565_, new_n41566_, new_n41567_, new_n41568_, new_n41569_,
    new_n41570_, new_n41571_, new_n41572_, new_n41573_, new_n41574_,
    new_n41575_, new_n41576_, new_n41577_, new_n41578_, new_n41579_,
    new_n41580_, new_n41581_, new_n41582_, new_n41583_, new_n41584_,
    new_n41585_, new_n41586_, new_n41587_, new_n41588_, new_n41589_,
    new_n41590_, new_n41591_, new_n41592_, new_n41593_, new_n41594_,
    new_n41595_, new_n41596_, new_n41597_, new_n41598_, new_n41600_,
    new_n41601_, new_n41602_, new_n41603_, new_n41604_, new_n41605_,
    new_n41606_, new_n41607_, new_n41608_, new_n41609_, new_n41610_,
    new_n41611_, new_n41612_, new_n41613_, new_n41614_, new_n41615_,
    new_n41616_, new_n41617_, new_n41618_, new_n41619_, new_n41620_,
    new_n41621_, new_n41622_, new_n41623_, new_n41624_, new_n41625_,
    new_n41626_, new_n41627_, new_n41628_, new_n41629_, new_n41630_,
    new_n41631_, new_n41632_, new_n41633_, new_n41635_, new_n41636_,
    new_n41637_, new_n41638_, new_n41639_, new_n41640_, new_n41641_,
    new_n41642_, new_n41643_, new_n41644_, new_n41645_, new_n41646_,
    new_n41647_, new_n41648_, new_n41649_, new_n41650_, new_n41651_,
    new_n41652_, new_n41653_, new_n41654_, new_n41655_, new_n41656_,
    new_n41657_, new_n41658_, new_n41659_, new_n41660_, new_n41661_,
    new_n41662_, new_n41663_, new_n41664_, new_n41665_, new_n41666_,
    new_n41667_, new_n41668_, new_n41669_, new_n41670_, new_n41672_,
    new_n41673_, new_n41674_, new_n41675_, new_n41676_, new_n41677_,
    new_n41678_, new_n41679_, new_n41680_, new_n41681_, new_n41682_,
    new_n41683_, new_n41684_, new_n41685_, new_n41686_, new_n41687_,
    new_n41688_, new_n41689_, new_n41690_, new_n41691_, new_n41692_,
    new_n41693_, new_n41694_, new_n41695_, new_n41696_, new_n41697_,
    new_n41698_, new_n41699_, new_n41700_, new_n41701_, new_n41702_,
    new_n41703_, new_n41704_, new_n41705_, new_n41706_, new_n41707_,
    new_n41708_, new_n41710_, new_n41711_, new_n41712_, new_n41713_,
    new_n41714_, new_n41715_, new_n41716_, new_n41717_, new_n41718_,
    new_n41719_, new_n41720_, new_n41721_, new_n41722_, new_n41723_,
    new_n41724_, new_n41725_, new_n41726_, new_n41727_, new_n41728_,
    new_n41729_, new_n41730_, new_n41731_, new_n41732_, new_n41733_,
    new_n41734_, new_n41735_, new_n41736_, new_n41737_, new_n41738_,
    new_n41739_, new_n41740_, new_n41741_, new_n41742_, new_n41743_,
    new_n41744_, new_n41745_, new_n41746_, new_n41748_, new_n41749_,
    new_n41750_, new_n41751_, new_n41752_, new_n41753_, new_n41754_,
    new_n41755_, new_n41756_, new_n41757_, new_n41758_, new_n41759_,
    new_n41760_, new_n41761_, new_n41762_, new_n41763_, new_n41764_,
    new_n41765_, new_n41766_, new_n41767_, new_n41768_, new_n41769_,
    new_n41770_, new_n41771_, new_n41772_, new_n41773_, new_n41774_,
    new_n41775_, new_n41776_, new_n41777_, new_n41778_, new_n41779_,
    new_n41780_, new_n41781_, new_n41782_, new_n41784_, new_n41785_,
    new_n41786_, new_n41787_, new_n41788_, new_n41789_, new_n41790_,
    new_n41791_, new_n41792_, new_n41793_, new_n41794_, new_n41795_,
    new_n41796_, new_n41797_, new_n41798_, new_n41799_, new_n41800_,
    new_n41801_, new_n41802_, new_n41803_, new_n41804_, new_n41805_,
    new_n41806_, new_n41807_, new_n41808_, new_n41809_, new_n41810_,
    new_n41811_, new_n41812_, new_n41813_, new_n41814_, new_n41815_,
    new_n41816_, new_n41817_, new_n41818_, new_n41819_, new_n41821_,
    new_n41822_, new_n41823_, new_n41824_, new_n41825_, new_n41826_,
    new_n41827_, new_n41828_, new_n41829_, new_n41830_, new_n41831_,
    new_n41832_, new_n41833_, new_n41834_, new_n41835_, new_n41836_,
    new_n41837_, new_n41838_, new_n41839_, new_n41840_, new_n41841_,
    new_n41842_, new_n41843_, new_n41844_, new_n41845_, new_n41846_,
    new_n41847_, new_n41848_, new_n41849_, new_n41850_, new_n41851_,
    new_n41852_, new_n41853_, new_n41854_, new_n41855_, new_n41856_,
    new_n41857_, new_n41859_, new_n41860_, new_n41861_, new_n41862_,
    new_n41863_, new_n41864_, new_n41865_, new_n41866_, new_n41867_,
    new_n41868_, new_n41869_, new_n41870_, new_n41871_, new_n41872_,
    new_n41873_, new_n41874_, new_n41875_, new_n41876_, new_n41877_,
    new_n41878_, new_n41879_, new_n41880_, new_n41881_, new_n41882_,
    new_n41883_, new_n41884_, new_n41885_, new_n41886_, new_n41887_,
    new_n41888_, new_n41889_, new_n41890_, new_n41891_, new_n41892_,
    new_n41893_, new_n41894_, new_n41895_, new_n41897_, new_n41898_,
    new_n41899_, new_n41900_, new_n41901_, new_n41902_, new_n41903_,
    new_n41904_, new_n41905_, new_n41906_, new_n41907_, new_n41908_,
    new_n41909_, new_n41910_, new_n41911_, new_n41912_, new_n41913_,
    new_n41914_, new_n41915_, new_n41916_, new_n41917_, new_n41918_,
    new_n41919_, new_n41920_, new_n41921_, new_n41922_, new_n41923_,
    new_n41924_, new_n41925_, new_n41926_, new_n41927_, new_n41928_,
    new_n41929_, new_n41930_, new_n41931_, new_n41932_, new_n41933_,
    new_n41935_, new_n41936_, new_n41937_, new_n41938_, new_n41939_,
    new_n41940_, new_n41941_, new_n41942_, new_n41943_, new_n41944_,
    new_n41945_, new_n41946_, new_n41947_, new_n41948_, new_n41949_,
    new_n41950_, new_n41951_, new_n41952_, new_n41953_, new_n41954_,
    new_n41955_, new_n41956_, new_n41957_, new_n41958_, new_n41959_,
    new_n41960_, new_n41961_, new_n41962_, new_n41963_, new_n41964_,
    new_n41965_, new_n41966_, new_n41967_, new_n41968_, new_n41969_,
    new_n41970_, new_n41972_, new_n41973_, new_n41974_, new_n41975_,
    new_n41976_, new_n41977_, new_n41978_, new_n41979_, new_n41980_,
    new_n41981_, new_n41982_, new_n41983_, new_n41984_, new_n41985_,
    new_n41986_, new_n41987_, new_n41988_, new_n41989_, new_n41990_,
    new_n41991_, new_n41992_, new_n41993_, new_n41994_, new_n41995_,
    new_n41996_, new_n41997_, new_n41998_, new_n41999_, new_n42000_,
    new_n42001_, new_n42002_, new_n42003_, new_n42004_, new_n42005_,
    new_n42006_, new_n42007_, new_n42008_, new_n42010_, new_n42011_,
    new_n42012_, new_n42013_, new_n42014_, new_n42015_, new_n42016_,
    new_n42017_, new_n42018_, new_n42019_, new_n42020_, new_n42021_,
    new_n42022_, new_n42023_, new_n42024_, new_n42025_, new_n42026_,
    new_n42027_, new_n42028_, new_n42029_, new_n42030_, new_n42031_,
    new_n42032_, new_n42033_, new_n42034_, new_n42035_, new_n42036_,
    new_n42037_, new_n42038_, new_n42039_, new_n42040_, new_n42041_,
    new_n42042_, new_n42043_, new_n42044_, new_n42045_, new_n42048_,
    new_n42049_, new_n42050_, new_n42051_, new_n42052_, new_n42053_,
    new_n42054_, new_n42055_, new_n42056_, new_n42057_, new_n42058_,
    new_n42059_, new_n42060_, new_n42061_, new_n42062_, new_n42063_,
    new_n42064_, new_n42065_, new_n42066_, new_n42068_, new_n42069_,
    new_n42070_, new_n42071_, new_n42072_, new_n42073_, new_n42074_,
    new_n42075_, new_n42076_, new_n42078_, new_n42079_, new_n42080_,
    new_n42081_, new_n42082_, new_n42083_, new_n42084_, new_n42085_,
    new_n42087_, new_n42088_, new_n42089_, new_n42090_, new_n42091_,
    new_n42093_, new_n42094_, new_n42095_, new_n42096_, new_n42097_,
    new_n42098_, new_n42099_, new_n42100_, new_n42102_, new_n42103_,
    new_n42104_, new_n42105_, new_n42106_, new_n42107_, new_n42108_,
    new_n42109_, new_n42111_, new_n42112_, new_n42113_, new_n42114_,
    new_n42115_, new_n42116_, new_n42117_, new_n42118_, new_n42119_,
    new_n42120_, new_n42121_, new_n42122_, new_n42123_, new_n42125_,
    new_n42126_, new_n42127_, new_n42128_, new_n42129_, new_n42131_,
    new_n42132_, new_n42133_, new_n42134_, new_n42135_, new_n42136_,
    new_n42137_, new_n42138_, new_n42140_, new_n42141_, new_n42142_,
    new_n42143_, new_n42144_, new_n42145_, new_n42146_, new_n42147_,
    new_n42148_, new_n42150_, new_n42151_, new_n42152_, new_n42153_,
    new_n42154_, new_n42155_, new_n42156_, new_n42157_, new_n42158_,
    new_n42159_, new_n42160_, new_n42161_, new_n42162_, new_n42163_,
    new_n42164_, new_n42165_, new_n42166_, new_n42167_, new_n42168_,
    new_n42169_, new_n42170_, new_n42171_, new_n42172_, new_n42173_,
    new_n42174_, new_n42176_, new_n42177_, new_n42178_, new_n42179_,
    new_n42180_, new_n42181_, new_n42182_, new_n42183_, new_n42185_,
    new_n42186_, new_n42187_, new_n42188_, new_n42189_, new_n42190_,
    new_n42191_, new_n42192_, new_n42193_, new_n42195_, new_n42196_,
    new_n42197_, new_n42198_, new_n42199_, new_n42200_, new_n42201_,
    new_n42202_, new_n42204_, new_n42205_, new_n42206_, new_n42207_,
    new_n42208_, new_n42209_, new_n42210_, new_n42211_, new_n42212_,
    new_n42213_, new_n42215_, new_n42216_, new_n42217_, new_n42218_,
    new_n42219_, new_n42220_, new_n42221_, new_n42222_, new_n42224_,
    new_n42225_, new_n42226_, new_n42227_, new_n42228_, new_n42229_,
    new_n42230_, new_n42231_, new_n42232_, new_n42234_, new_n42235_,
    new_n42236_, new_n42237_, new_n42238_, new_n42239_, new_n42240_,
    new_n42241_, new_n42242_, new_n42243_, new_n42244_, new_n42245_,
    new_n42246_, new_n42247_, new_n42248_, new_n42249_, new_n42250_,
    new_n42251_, new_n42252_, new_n42253_, new_n42254_, new_n42255_,
    new_n42256_, new_n42257_, new_n42258_, new_n42259_, new_n42260_,
    new_n42261_, new_n42262_, new_n42263_, new_n42264_, new_n42265_,
    new_n42266_, new_n42267_, new_n42268_, new_n42270_, new_n42271_,
    new_n42272_, new_n42273_, new_n42274_, new_n42275_, new_n42276_,
    new_n42277_, new_n42278_, new_n42280_, new_n42281_, new_n42282_,
    new_n42283_, new_n42284_, new_n42285_, new_n42286_, new_n42287_,
    new_n42288_, new_n42289_, new_n42290_, new_n42291_, new_n42293_,
    new_n42294_, new_n42295_, new_n42296_, new_n42297_, new_n42298_,
    new_n42299_, new_n42300_, new_n42301_, new_n42303_, new_n42304_,
    new_n42305_, new_n42306_, new_n42307_, new_n42308_, new_n42309_,
    new_n42310_, new_n42311_, new_n42312_, new_n42313_, new_n42314_,
    new_n42315_, new_n42316_, new_n42317_, new_n42319_, new_n42320_,
    new_n42321_, new_n42322_, new_n42323_, new_n42324_, new_n42325_,
    new_n42326_, new_n42327_, new_n42329_, new_n42330_, new_n42331_,
    new_n42332_, new_n42333_, new_n42334_, new_n42335_, new_n42336_,
    new_n42337_, new_n42338_, new_n42339_, new_n42340_, new_n42341_,
    new_n42342_, new_n42343_, new_n42345_, new_n42346_, new_n42347_,
    new_n42348_, new_n42349_, new_n42350_, new_n42351_, new_n42352_,
    new_n42353_, new_n42355_, new_n42356_, new_n42357_, new_n42358_,
    new_n42359_, new_n42360_, new_n42361_, new_n42362_, new_n42363_,
    new_n42364_, new_n42365_, new_n42366_, new_n42367_, new_n42368_,
    new_n42369_, new_n42370_, new_n42371_, new_n42372_, new_n42374_,
    new_n42375_, new_n42376_, new_n42377_, new_n42378_, new_n42379_,
    new_n42380_, new_n42381_, new_n42382_, new_n42384_, new_n42385_,
    new_n42386_, new_n42387_, new_n42388_, new_n42389_, new_n42390_,
    new_n42391_, new_n42392_, new_n42393_, new_n42394_, new_n42395_,
    new_n42396_, new_n42397_, new_n42398_, new_n42400_, new_n42401_,
    new_n42402_, new_n42403_, new_n42404_, new_n42405_, new_n42406_,
    new_n42407_, new_n42408_, new_n42410_, new_n42411_, new_n42412_,
    new_n42413_, new_n42414_, new_n42415_, new_n42416_, new_n42417_,
    new_n42418_, new_n42419_, new_n42420_, new_n42421_, new_n42422_,
    new_n42423_, new_n42424_, new_n42425_, new_n42426_, new_n42427_,
    new_n42428_, new_n42430_, new_n42431_, new_n42432_, new_n42433_,
    new_n42434_, new_n42435_, new_n42436_, new_n42437_, new_n42438_,
    new_n42440_, new_n42441_, new_n42442_, new_n42443_, new_n42444_,
    new_n42445_, new_n42446_, new_n42447_, new_n42448_, new_n42449_,
    new_n42450_, new_n42451_, new_n42452_, new_n42453_, new_n42454_,
    new_n42456_, new_n42457_, new_n42458_, new_n42459_, new_n42460_,
    new_n42461_, new_n42462_, new_n42463_, new_n42464_, new_n42466_,
    new_n42467_, new_n42468_, new_n42469_, new_n42470_, new_n42471_,
    new_n42472_, new_n42473_, new_n42474_, new_n42475_, new_n42476_,
    new_n42477_, new_n42478_, new_n42479_, new_n42480_, new_n42481_,
    new_n42482_, new_n42483_, new_n42484_, new_n42485_, new_n42486_,
    new_n42487_, new_n42488_, new_n42490_, new_n42491_, new_n42492_,
    new_n42493_, new_n42494_, new_n42495_, new_n42496_, new_n42497_,
    new_n42498_, new_n42500_, new_n42501_, new_n42502_, new_n42503_,
    new_n42504_, new_n42505_, new_n42506_, new_n42507_, new_n42508_,
    new_n42509_, new_n42510_, new_n42511_, new_n42512_, new_n42513_,
    new_n42514_, new_n42516_, new_n42517_, new_n42518_, new_n42519_,
    new_n42520_, new_n42521_, new_n42522_, new_n42523_, new_n42524_,
    new_n42526_, new_n42527_, new_n42528_, new_n42529_, new_n42530_,
    new_n42531_, new_n42532_, new_n42533_, new_n42534_, new_n42535_,
    new_n42536_, new_n42537_, new_n42538_, new_n42539_, new_n42540_,
    new_n42541_, new_n42542_, new_n42543_, new_n42544_, new_n42546_,
    new_n42547_, new_n42548_, new_n42549_, new_n42550_, new_n42551_,
    new_n42552_, new_n42553_, new_n42554_, new_n42556_, new_n42557_,
    new_n42558_, new_n42559_, new_n42560_, new_n42561_, new_n42562_,
    new_n42563_, new_n42564_, new_n42565_, new_n42566_, new_n42567_,
    new_n42568_, new_n42569_, new_n42570_, new_n42572_, new_n42573_,
    new_n42574_, new_n42575_, new_n42576_, new_n42577_, new_n42578_,
    new_n42579_, new_n42580_, new_n42582_, new_n42583_, new_n42584_,
    new_n42585_, new_n42586_, new_n42587_, new_n42588_, new_n42589_,
    new_n42590_, new_n42591_, new_n42592_, new_n42593_, new_n42594_,
    new_n42595_, new_n42596_, new_n42597_, new_n42598_, new_n42599_,
    new_n42600_, new_n42601_, new_n42602_, new_n42603_, new_n42604_,
    new_n42606_, new_n42607_, new_n42608_, new_n42609_, new_n42610_,
    new_n42611_, new_n42612_, new_n42613_, new_n42614_, new_n42616_,
    new_n42617_, new_n42618_, new_n42619_, new_n42620_, new_n42621_,
    new_n42622_, new_n42623_, new_n42624_, new_n42625_, new_n42626_,
    new_n42627_, new_n42628_, new_n42629_, new_n42630_, new_n42632_,
    new_n42633_, new_n42634_, new_n42635_, new_n42636_, new_n42637_,
    new_n42638_, new_n42639_, new_n42640_, new_n42642_, new_n42643_,
    new_n42644_, new_n42645_, new_n42646_, new_n42647_, new_n42648_,
    new_n42649_, new_n42650_, new_n42651_, new_n42652_, new_n42653_,
    new_n42654_, new_n42655_, new_n42656_, new_n42657_, new_n42658_,
    new_n42659_, new_n42660_, new_n42662_, new_n42663_, new_n42664_,
    new_n42665_, new_n42666_, new_n42667_, new_n42668_, new_n42669_,
    new_n42670_, new_n42672_, new_n42673_, new_n42674_, new_n42675_,
    new_n42676_, new_n42677_, new_n42678_, new_n42679_, new_n42680_,
    new_n42681_, new_n42682_, new_n42683_, new_n42684_, new_n42685_,
    new_n42686_, new_n42688_, new_n42689_, new_n42691_, new_n42692_,
    new_n42693_, new_n42694_, new_n42695_, new_n42696_, new_n42697_,
    new_n42698_, new_n42699_, new_n42700_, new_n42701_, new_n42702_,
    new_n42703_, new_n42704_, new_n42705_, new_n42706_, new_n42707_,
    new_n42708_, new_n42709_, new_n42710_, new_n42711_, new_n42712_,
    new_n42713_, new_n42714_, new_n42715_, new_n42716_, new_n42717_,
    new_n42719_, new_n42720_, new_n42721_, new_n42722_, new_n42723_,
    new_n42724_, new_n42725_, new_n42726_, new_n42727_, new_n42729_,
    new_n42730_, new_n42731_, new_n42732_, new_n42733_, new_n42734_,
    new_n42735_, new_n42737_, new_n42738_, new_n42740_, new_n42741_,
    new_n42743_, new_n42744_, new_n42746_, new_n42747_, new_n42749_,
    new_n42750_, new_n42752_, new_n42753_, new_n42755_, new_n42756_,
    new_n42758_, new_n42759_, new_n42761_, new_n42762_, new_n42764_,
    new_n42765_, new_n42767_, new_n42768_, new_n42770_, new_n42771_,
    new_n42773_, new_n42774_, new_n42776_, new_n42777_, new_n42779_,
    new_n42780_, new_n42782_, new_n42783_, new_n42785_, new_n42786_,
    new_n42788_, new_n42789_, new_n42790_, new_n42791_, new_n42792_,
    new_n42793_, new_n42794_, new_n42795_, new_n42796_, new_n42797_,
    new_n42798_, new_n42799_, new_n42800_, new_n42801_, new_n42802_,
    new_n42803_, new_n42804_, new_n42805_, new_n42806_, new_n42807_,
    new_n42808_, new_n42809_, new_n42810_, new_n42811_, new_n42812_,
    new_n42813_, new_n42814_, new_n42815_, new_n42816_, new_n42817_,
    new_n42818_, new_n42819_, new_n42820_, new_n42821_, new_n42822_,
    new_n42823_, new_n42824_, new_n42825_, new_n42826_, new_n42827_,
    new_n42828_, new_n42830_, new_n42831_, new_n42832_, new_n42833_,
    new_n42834_, new_n42835_, new_n42837_, new_n42838_, new_n42840_,
    new_n42841_, new_n42842_, new_n42844_, new_n42845_, new_n42846_,
    new_n42848_, new_n42849_, new_n42850_, new_n42852_, new_n42853_,
    new_n42854_, new_n42859_, new_n42865_, new_n42867_, new_n42874_,
    new_n42875_, new_n42876_, new_n42877_, new_n42878_, new_n42879_,
    new_n42880_, new_n42881_, new_n42882_, new_n42883_, new_n42884_,
    new_n42885_, new_n42886_, new_n42887_, new_n42888_, new_n42889_,
    new_n42890_, new_n42891_, new_n42892_, new_n42893_, new_n42894_,
    new_n42895_, new_n42896_, new_n42897_, new_n42898_, new_n42899_,
    new_n42900_, new_n42901_, new_n42902_, new_n42903_, new_n42905_,
    new_n42906_, new_n42907_, new_n42908_, new_n42909_, new_n42911_,
    new_n42912_, new_n42913_, new_n42914_, new_n42915_, new_n42916_,
    new_n42917_, new_n42918_, new_n42919_, new_n42920_, new_n42921_,
    new_n42922_, new_n42923_, new_n42924_, new_n42925_, new_n42926_,
    new_n42927_, new_n42928_, new_n42929_, new_n42930_, new_n42931_,
    new_n42932_, new_n42933_, new_n42934_, new_n42935_, new_n42936_,
    new_n42937_, new_n42938_, new_n42939_, new_n42940_, new_n42941_,
    new_n42942_, new_n42943_, new_n42944_, new_n42945_, new_n42947_,
    new_n42948_, new_n42949_, new_n42950_, new_n42951_, new_n42952_,
    new_n42953_, new_n42954_, new_n42955_, new_n42956_, new_n42957_,
    new_n42958_, new_n42959_, new_n42960_, new_n42961_, new_n42962_,
    new_n42963_, new_n42964_, new_n42965_, new_n42966_, new_n42967_,
    new_n42968_, new_n42969_, new_n42970_, new_n42972_, new_n42973_,
    new_n42974_, new_n42975_, new_n42976_, new_n42977_, new_n42978_,
    new_n42979_, new_n42980_, new_n42981_, new_n42982_, new_n42983_,
    new_n42984_, new_n42985_, new_n42986_, new_n42987_, new_n42988_,
    new_n42989_, new_n42990_, new_n42991_, new_n42992_, new_n42994_,
    new_n42995_, new_n42996_, new_n42997_, new_n42998_, new_n42999_,
    new_n43000_, new_n43001_, new_n43002_, new_n43003_, new_n43004_,
    new_n43005_, new_n43006_, new_n43007_, new_n43008_, new_n43009_,
    new_n43010_, new_n43011_, new_n43012_, new_n43013_, new_n43014_,
    new_n43016_, new_n43017_, new_n43018_, new_n43019_, new_n43020_,
    new_n43021_, new_n43022_, new_n43023_, new_n43024_, new_n43025_,
    new_n43026_, new_n43027_, new_n43028_, new_n43029_, new_n43030_,
    new_n43031_, new_n43032_, new_n43033_, new_n43034_, new_n43035_,
    new_n43036_, new_n43037_, new_n43039_, new_n43040_, new_n43041_,
    new_n43042_, new_n43043_, new_n43044_, new_n43045_, new_n43046_,
    new_n43047_, new_n43048_, new_n43049_, new_n43050_, new_n43051_,
    new_n43052_, new_n43053_, new_n43054_, new_n43055_, new_n43056_,
    new_n43057_, new_n43058_, new_n43059_, new_n43061_, new_n43062_,
    new_n43063_, new_n43064_, new_n43065_, new_n43066_, new_n43067_,
    new_n43068_, new_n43069_, new_n43070_, new_n43071_, new_n43072_,
    new_n43073_, new_n43074_, new_n43075_, new_n43076_, new_n43077_,
    new_n43078_, new_n43079_, new_n43080_, new_n43081_, new_n43082_,
    new_n43084_, new_n43085_, new_n43086_, new_n43087_, new_n43088_,
    new_n43089_, new_n43090_, new_n43091_, new_n43092_, new_n43093_,
    new_n43094_, new_n43095_, new_n43096_, new_n43097_, new_n43098_,
    new_n43099_, new_n43100_, new_n43101_, new_n43102_, new_n43103_,
    new_n43104_, new_n43106_, new_n43107_, new_n43108_, new_n43109_,
    new_n43110_, new_n43111_, new_n43112_, new_n43113_, new_n43114_,
    new_n43115_, new_n43116_, new_n43117_, new_n43118_, new_n43119_,
    new_n43120_, new_n43121_, new_n43122_, new_n43123_, new_n43124_,
    new_n43125_, new_n43126_, new_n43127_, new_n43128_, new_n43130_,
    new_n43131_, new_n43132_, new_n43133_, new_n43134_, new_n43135_,
    new_n43136_, new_n43137_, new_n43138_, new_n43139_, new_n43140_,
    new_n43141_, new_n43142_, new_n43143_, new_n43144_, new_n43145_,
    new_n43146_, new_n43147_, new_n43148_, new_n43149_, new_n43150_,
    new_n43152_, new_n43153_, new_n43154_, new_n43155_, new_n43156_,
    new_n43157_, new_n43158_, new_n43159_, new_n43160_, new_n43161_,
    new_n43162_, new_n43163_, new_n43164_, new_n43165_, new_n43166_,
    new_n43167_, new_n43168_, new_n43169_, new_n43170_, new_n43171_,
    new_n43172_, new_n43173_, new_n43175_, new_n43176_, new_n43177_,
    new_n43178_, new_n43179_, new_n43180_, new_n43181_, new_n43182_,
    new_n43183_, new_n43184_, new_n43185_, new_n43186_, new_n43187_,
    new_n43188_, new_n43189_, new_n43190_, new_n43191_, new_n43192_,
    new_n43193_, new_n43194_, new_n43195_, new_n43197_, new_n43198_,
    new_n43199_, new_n43200_, new_n43201_, new_n43202_, new_n43203_,
    new_n43204_, new_n43205_, new_n43206_, new_n43207_, new_n43208_,
    new_n43209_, new_n43210_, new_n43211_, new_n43212_, new_n43213_,
    new_n43214_, new_n43215_, new_n43216_, new_n43217_, new_n43218_,
    new_n43219_, new_n43221_, new_n43222_, new_n43223_, new_n43224_,
    new_n43225_, new_n43226_, new_n43227_, new_n43228_, new_n43229_,
    new_n43230_, new_n43231_, new_n43232_, new_n43233_, new_n43234_,
    new_n43235_, new_n43236_, new_n43237_, new_n43238_, new_n43239_,
    new_n43240_, new_n43241_, new_n43243_, new_n43244_, new_n43245_,
    new_n43246_, new_n43247_, new_n43248_, new_n43249_, new_n43250_,
    new_n43251_, new_n43252_, new_n43253_, new_n43254_, new_n43255_,
    new_n43256_, new_n43257_, new_n43258_, new_n43259_, new_n43260_,
    new_n43261_, new_n43262_, new_n43263_, new_n43264_, new_n43266_,
    new_n43267_, new_n43268_, new_n43269_, new_n43270_, new_n43271_,
    new_n43272_, new_n43273_, new_n43274_, new_n43275_, new_n43276_,
    new_n43277_, new_n43278_, new_n43279_, new_n43280_, new_n43281_,
    new_n43282_, new_n43283_, new_n43284_, new_n43285_, new_n43286_,
    new_n43288_, new_n43289_, new_n43290_, new_n43291_, new_n43292_,
    new_n43293_, new_n43294_, new_n43295_, new_n43296_, new_n43297_,
    new_n43298_, new_n43299_, new_n43300_, new_n43301_, new_n43302_,
    new_n43303_, new_n43304_, new_n43305_, new_n43306_, new_n43307_,
    new_n43308_, new_n43309_, new_n43310_, new_n43311_, new_n43313_,
    new_n43314_, new_n43315_, new_n43316_, new_n43317_, new_n43318_,
    new_n43319_, new_n43320_, new_n43321_, new_n43322_, new_n43323_,
    new_n43324_, new_n43325_, new_n43326_, new_n43327_, new_n43328_,
    new_n43329_, new_n43330_, new_n43331_, new_n43332_, new_n43333_,
    new_n43335_, new_n43336_, new_n43337_, new_n43338_, new_n43339_,
    new_n43340_, new_n43341_, new_n43342_, new_n43343_, new_n43344_,
    new_n43345_, new_n43346_, new_n43347_, new_n43348_, new_n43349_,
    new_n43350_, new_n43351_, new_n43352_, new_n43353_, new_n43354_,
    new_n43355_, new_n43356_, new_n43358_, new_n43359_, new_n43360_,
    new_n43361_, new_n43362_, new_n43363_, new_n43364_, new_n43365_,
    new_n43366_, new_n43367_, new_n43368_, new_n43369_, new_n43370_,
    new_n43371_, new_n43372_, new_n43373_, new_n43374_, new_n43375_,
    new_n43376_, new_n43377_, new_n43378_, new_n43380_, new_n43381_,
    new_n43382_, new_n43383_, new_n43384_, new_n43385_, new_n43386_,
    new_n43387_, new_n43388_, new_n43389_, new_n43390_, new_n43391_,
    new_n43392_, new_n43393_, new_n43394_, new_n43395_, new_n43396_,
    new_n43397_, new_n43398_, new_n43399_, new_n43400_, new_n43401_,
    new_n43402_, new_n43404_, new_n43405_, new_n43406_, new_n43407_,
    new_n43408_, new_n43409_, new_n43410_, new_n43411_, new_n43412_,
    new_n43413_, new_n43414_, new_n43415_, new_n43416_, new_n43417_,
    new_n43418_, new_n43419_, new_n43420_, new_n43421_, new_n43422_,
    new_n43423_, new_n43424_, new_n43426_, new_n43427_, new_n43428_,
    new_n43429_, new_n43430_, new_n43431_, new_n43432_, new_n43433_,
    new_n43434_, new_n43435_, new_n43436_, new_n43437_, new_n43438_,
    new_n43439_, new_n43440_, new_n43441_, new_n43442_, new_n43443_,
    new_n43444_, new_n43445_, new_n43446_, new_n43447_, new_n43449_,
    new_n43450_, new_n43451_, new_n43452_, new_n43453_, new_n43454_,
    new_n43455_, new_n43456_, new_n43457_, new_n43458_, new_n43459_,
    new_n43460_, new_n43461_, new_n43462_, new_n43463_, new_n43464_,
    new_n43465_, new_n43466_, new_n43467_, new_n43468_, new_n43469_,
    new_n43471_, new_n43472_, new_n43473_, new_n43474_, new_n43475_,
    new_n43476_, new_n43477_, new_n43478_, new_n43479_, new_n43480_,
    new_n43481_, new_n43482_, new_n43483_, new_n43484_, new_n43485_,
    new_n43486_, new_n43487_, new_n43488_, new_n43489_, new_n43490_,
    new_n43491_, new_n43492_, new_n43493_, new_n43494_, new_n43496_,
    new_n43497_, new_n43498_, new_n43499_, new_n43500_, new_n43501_,
    new_n43502_, new_n43503_, new_n43504_, new_n43505_, new_n43506_,
    new_n43507_, new_n43508_, new_n43509_, new_n43510_, new_n43511_,
    new_n43512_, new_n43513_, new_n43514_, new_n43515_, new_n43516_,
    new_n43518_, new_n43519_, new_n43520_, new_n43521_, new_n43522_,
    new_n43523_, new_n43524_, new_n43525_, new_n43526_, new_n43527_,
    new_n43528_, new_n43529_, new_n43530_, new_n43531_, new_n43532_,
    new_n43533_, new_n43534_, new_n43535_, new_n43536_, new_n43537_,
    new_n43538_, new_n43539_, new_n43541_, new_n43542_, new_n43543_,
    new_n43544_, new_n43545_, new_n43546_, new_n43547_, new_n43548_,
    new_n43549_, new_n43550_, new_n43551_, new_n43552_, new_n43553_,
    new_n43554_, new_n43555_, new_n43556_, new_n43557_, new_n43558_,
    new_n43559_, new_n43560_, new_n43561_, new_n43563_, new_n43564_,
    new_n43565_, new_n43566_, new_n43567_, new_n43568_, new_n43569_,
    new_n43570_, new_n43571_, new_n43572_, new_n43573_, new_n43574_,
    new_n43575_, new_n43576_, new_n43577_, new_n43578_, new_n43579_,
    new_n43580_, new_n43581_, new_n43582_, new_n43583_, new_n43584_,
    new_n43585_, new_n43587_, new_n43588_, new_n43589_, new_n43590_,
    new_n43591_, new_n43592_, new_n43593_, new_n43594_, new_n43595_,
    new_n43596_, new_n43597_, new_n43598_, new_n43599_, new_n43600_,
    new_n43601_, new_n43602_, new_n43603_, new_n43604_, new_n43605_,
    new_n43606_, new_n43607_, new_n43609_, new_n43610_, new_n43611_,
    new_n43612_, new_n43613_, new_n43614_, new_n43615_, new_n43616_,
    new_n43617_, new_n43618_, new_n43619_, new_n43620_, new_n43622_,
    new_n43623_, new_n43624_, new_n43625_, new_n43626_, new_n43627_,
    new_n43628_, new_n43629_, new_n43630_, new_n43632_, new_n43633_,
    new_n43634_, new_n43635_, new_n43636_, new_n43637_, new_n43638_,
    new_n43639_, new_n43640_, new_n43641_, new_n43642_, new_n43644_,
    new_n43645_, new_n43646_, new_n43647_, new_n43648_, new_n43649_,
    new_n43650_, new_n43651_, new_n43652_, new_n43654_, new_n43655_,
    new_n43656_, new_n43657_, new_n43658_, new_n43659_, new_n43660_,
    new_n43661_, new_n43663_, new_n43664_, new_n43665_, new_n43667_,
    new_n43668_, new_n43669_, new_n43671_, new_n43672_, new_n43673_,
    new_n43675_, new_n43676_, new_n43677_, new_n43679_, new_n43680_,
    new_n43681_, new_n43683_, new_n43684_, new_n43685_, new_n43687_,
    new_n43688_, new_n43689_, new_n43691_, new_n43692_, new_n43693_,
    new_n43695_, new_n43696_, new_n43697_, new_n43699_, new_n43700_,
    new_n43701_, new_n43703_, new_n43704_, new_n43705_, new_n43707_,
    new_n43708_, new_n43709_, new_n43711_, new_n43712_, new_n43713_,
    new_n43715_, new_n43716_, new_n43717_, new_n43719_, new_n43720_,
    new_n43721_, new_n43723_, new_n43724_, new_n43725_, new_n43727_,
    new_n43728_, new_n43729_, new_n43731_, new_n43732_, new_n43733_,
    new_n43735_, new_n43736_, new_n43737_, new_n43739_, new_n43740_,
    new_n43741_, new_n43743_, new_n43744_, new_n43745_, new_n43747_,
    new_n43748_, new_n43749_, new_n43751_, new_n43752_, new_n43753_,
    new_n43755_, new_n43756_, new_n43757_, new_n43759_, new_n43760_,
    new_n43761_, new_n43763_, new_n43764_, new_n43765_, new_n43767_,
    new_n43768_, new_n43769_, new_n43771_, new_n43772_, new_n43773_,
    new_n43775_, new_n43776_, new_n43777_, new_n43779_, new_n43780_,
    new_n43781_, new_n43783_, new_n43784_, new_n43785_, new_n43787_,
    new_n43788_, new_n43789_, new_n43791_, new_n43792_, new_n43793_,
    new_n43795_, new_n43796_, new_n43797_, new_n43799_, new_n43800_,
    new_n43801_, new_n43802_, new_n43803_, new_n43804_, new_n43805_,
    new_n43806_, new_n43808_, new_n43809_, new_n43810_, new_n43812_,
    new_n43813_, new_n43814_, new_n43816_, new_n43817_, new_n43818_,
    new_n43820_, new_n43821_, new_n43822_, new_n43824_, new_n43825_,
    new_n43826_, new_n43828_, new_n43829_, new_n43830_, new_n43832_,
    new_n43833_, new_n43834_, new_n43836_, new_n43837_, new_n43838_,
    new_n43840_, new_n43841_, new_n43842_, new_n43844_, new_n43845_,
    new_n43846_, new_n43848_, new_n43849_, new_n43850_, new_n43852_,
    new_n43853_, new_n43854_, new_n43856_, new_n43857_, new_n43858_,
    new_n43860_, new_n43861_, new_n43862_, new_n43864_, new_n43865_,
    new_n43866_, new_n43868_, new_n43869_, new_n43870_, new_n43872_,
    new_n43873_, new_n43874_, new_n43876_, new_n43877_, new_n43878_,
    new_n43880_, new_n43881_, new_n43882_, new_n43884_, new_n43885_,
    new_n43886_, new_n43888_, new_n43889_, new_n43890_, new_n43892_,
    new_n43893_, new_n43894_, new_n43896_, new_n43897_, new_n43898_,
    new_n43900_, new_n43901_, new_n43902_, new_n43904_, new_n43905_,
    new_n43906_, new_n43908_, new_n43909_, new_n43910_, new_n43912_,
    new_n43913_, new_n43914_, new_n43916_, new_n43917_, new_n43918_,
    new_n43920_, new_n43921_, new_n43922_, new_n43924_, new_n43925_,
    new_n43926_, new_n43928_, new_n43929_, new_n43930_, new_n43932_,
    new_n43933_, new_n43934_, new_n43936_, new_n43937_, new_n43938_,
    new_n43940_, new_n43941_, new_n43942_, new_n43944_, new_n43945_,
    new_n43946_, new_n43947_, new_n43948_, new_n43949_, new_n43950_,
    new_n43951_, new_n43953_, new_n43954_, new_n43955_, new_n43957_,
    new_n43958_, new_n43959_, new_n43961_, new_n43962_, new_n43963_,
    new_n43965_, new_n43966_, new_n43967_, new_n43969_, new_n43970_,
    new_n43971_, new_n43973_, new_n43974_, new_n43975_, new_n43977_,
    new_n43978_, new_n43979_, new_n43981_, new_n43982_, new_n43983_,
    new_n43985_, new_n43986_, new_n43987_, new_n43989_, new_n43990_,
    new_n43991_, new_n43993_, new_n43994_, new_n43995_, new_n43997_,
    new_n43998_, new_n43999_, new_n44001_, new_n44002_, new_n44003_,
    new_n44005_, new_n44006_, new_n44007_, new_n44009_, new_n44010_,
    new_n44011_, new_n44013_, new_n44014_, new_n44015_, new_n44017_,
    new_n44018_, new_n44019_, new_n44021_, new_n44022_, new_n44023_,
    new_n44025_, new_n44026_, new_n44027_, new_n44029_, new_n44030_,
    new_n44031_, new_n44033_, new_n44034_, new_n44035_, new_n44037_,
    new_n44038_, new_n44039_, new_n44041_, new_n44042_, new_n44043_,
    new_n44045_, new_n44046_, new_n44047_, new_n44049_, new_n44050_,
    new_n44051_, new_n44053_, new_n44054_, new_n44055_, new_n44057_,
    new_n44058_, new_n44059_, new_n44061_, new_n44062_, new_n44063_,
    new_n44065_, new_n44066_, new_n44067_, new_n44069_, new_n44070_,
    new_n44071_, new_n44073_, new_n44074_, new_n44075_, new_n44077_,
    new_n44078_, new_n44079_, new_n44081_, new_n44082_, new_n44083_,
    new_n44085_, new_n44086_, new_n44087_, new_n44089_, new_n44090_,
    new_n44091_, new_n44092_, new_n44093_, new_n44094_, new_n44095_,
    new_n44096_, new_n44097_, new_n44098_, new_n44099_, new_n44100_,
    new_n44102_, new_n44103_, new_n44104_, new_n44105_, new_n44106_,
    new_n44107_, new_n44108_, new_n44109_, new_n44110_, new_n44111_,
    new_n44112_, new_n44113_, new_n44114_, new_n44115_, new_n44116_,
    new_n44117_, new_n44118_, new_n44119_, new_n44120_, new_n44121_,
    new_n44122_, new_n44124_, new_n44125_, new_n44126_, new_n44127_,
    new_n44128_, new_n44129_, new_n44130_, new_n44132_, new_n44133_,
    new_n44134_, new_n44135_, new_n44136_, new_n44137_, new_n44138_,
    new_n44140_, new_n44141_, new_n44142_, new_n44144_, new_n44145_,
    new_n44146_, new_n44147_, new_n44148_, new_n44149_, new_n44150_,
    new_n44152_, new_n44153_, new_n44154_, new_n44156_, new_n44157_,
    new_n44158_, new_n44160_, new_n44161_, new_n44162_, new_n44164_,
    new_n44165_, new_n44166_, new_n44168_, new_n44169_, new_n44170_,
    new_n44172_, new_n44173_, new_n44174_, new_n44175_, new_n44176_,
    new_n44177_, new_n44178_, new_n44179_, new_n44181_, new_n44182_,
    new_n44183_, new_n44185_, new_n44186_, new_n44187_, new_n44189_,
    new_n44190_, new_n44191_, new_n44193_, new_n44194_, new_n44195_,
    new_n44197_, new_n44198_, new_n44199_, new_n44201_, new_n44202_,
    new_n44203_, new_n44205_, new_n44206_, new_n44207_, new_n44209_,
    new_n44210_, new_n44211_, new_n44213_, new_n44214_, new_n44215_,
    new_n44217_, new_n44218_, new_n44219_, new_n44221_, new_n44222_,
    new_n44223_, new_n44225_, new_n44226_, new_n44227_, new_n44229_,
    new_n44230_, new_n44231_, new_n44233_, new_n44234_, new_n44235_,
    new_n44237_, new_n44238_, new_n44239_, new_n44241_, new_n44242_,
    new_n44243_, new_n44245_, new_n44246_, new_n44247_, new_n44249_,
    new_n44250_, new_n44251_, new_n44253_, new_n44254_, new_n44255_,
    new_n44257_, new_n44258_, new_n44259_, new_n44261_, new_n44262_,
    new_n44263_, new_n44265_, new_n44266_, new_n44267_, new_n44269_,
    new_n44270_, new_n44271_, new_n44273_, new_n44274_, new_n44275_,
    new_n44277_, new_n44278_, new_n44279_, new_n44281_, new_n44282_,
    new_n44283_, new_n44285_, new_n44286_, new_n44287_, new_n44289_,
    new_n44290_, new_n44291_, new_n44293_, new_n44294_, new_n44295_,
    new_n44297_, new_n44298_, new_n44299_, new_n44301_, new_n44302_,
    new_n44303_, new_n44305_, new_n44306_, new_n44307_, new_n44309_,
    new_n44310_, new_n44311_, new_n44313_, new_n44314_, new_n44315_,
    new_n44317_, new_n44318_, new_n44319_, new_n44320_, new_n44321_,
    new_n44322_, new_n44323_, new_n44324_, new_n44326_, new_n44327_,
    new_n44328_, new_n44330_, new_n44331_, new_n44332_, new_n44334_,
    new_n44335_, new_n44336_, new_n44338_, new_n44339_, new_n44340_,
    new_n44342_, new_n44343_, new_n44344_, new_n44346_, new_n44347_,
    new_n44348_, new_n44350_, new_n44351_, new_n44352_, new_n44354_,
    new_n44355_, new_n44356_, new_n44358_, new_n44359_, new_n44360_,
    new_n44362_, new_n44363_, new_n44364_, new_n44366_, new_n44367_,
    new_n44368_, new_n44370_, new_n44371_, new_n44372_, new_n44374_,
    new_n44375_, new_n44376_, new_n44378_, new_n44379_, new_n44380_,
    new_n44382_, new_n44383_, new_n44384_, new_n44386_, new_n44387_,
    new_n44388_, new_n44390_, new_n44391_, new_n44392_, new_n44394_,
    new_n44395_, new_n44396_, new_n44398_, new_n44399_, new_n44400_,
    new_n44402_, new_n44403_, new_n44404_, new_n44406_, new_n44407_,
    new_n44408_, new_n44410_, new_n44411_, new_n44412_, new_n44414_,
    new_n44415_, new_n44416_, new_n44418_, new_n44419_, new_n44420_,
    new_n44422_, new_n44423_, new_n44424_, new_n44426_, new_n44427_,
    new_n44428_, new_n44430_, new_n44431_, new_n44432_, new_n44434_,
    new_n44435_, new_n44436_, new_n44438_, new_n44439_, new_n44440_,
    new_n44442_, new_n44443_, new_n44444_, new_n44446_, new_n44447_,
    new_n44448_, new_n44450_, new_n44451_, new_n44452_, new_n44454_,
    new_n44455_, new_n44456_, new_n44458_, new_n44459_, new_n44460_,
    new_n44462_, new_n44463_, new_n44464_, new_n44465_, new_n44466_,
    new_n44467_, new_n44468_, new_n44469_, new_n44471_, new_n44472_,
    new_n44473_, new_n44475_, new_n44476_, new_n44477_, new_n44479_,
    new_n44480_, new_n44481_, new_n44483_, new_n44484_, new_n44485_,
    new_n44487_, new_n44488_, new_n44489_, new_n44491_, new_n44492_,
    new_n44493_, new_n44495_, new_n44496_, new_n44497_, new_n44499_,
    new_n44500_, new_n44501_, new_n44503_, new_n44504_, new_n44505_,
    new_n44507_, new_n44508_, new_n44509_, new_n44511_, new_n44512_,
    new_n44513_, new_n44515_, new_n44516_, new_n44517_, new_n44519_,
    new_n44520_, new_n44521_, new_n44523_, new_n44524_, new_n44525_,
    new_n44527_, new_n44528_, new_n44529_, new_n44531_, new_n44532_,
    new_n44533_, new_n44535_, new_n44536_, new_n44537_, new_n44539_,
    new_n44540_, new_n44541_, new_n44543_, new_n44544_, new_n44545_,
    new_n44547_, new_n44548_, new_n44549_, new_n44551_, new_n44552_,
    new_n44553_, new_n44555_, new_n44556_, new_n44557_, new_n44559_,
    new_n44560_, new_n44561_, new_n44563_, new_n44564_, new_n44565_,
    new_n44567_, new_n44568_, new_n44569_, new_n44571_, new_n44572_,
    new_n44573_, new_n44575_, new_n44576_, new_n44577_, new_n44579_,
    new_n44580_, new_n44581_, new_n44583_, new_n44584_, new_n44585_,
    new_n44587_, new_n44588_, new_n44589_, new_n44591_, new_n44592_,
    new_n44593_, new_n44595_, new_n44596_, new_n44597_, new_n44599_,
    new_n44600_, new_n44601_, new_n44603_, new_n44604_, new_n44605_,
    new_n44607_, new_n44608_, new_n44609_, new_n44610_, new_n44611_,
    new_n44612_, new_n44613_, new_n44614_, new_n44615_, new_n44616_,
    new_n44617_, new_n44618_, new_n44620_, new_n44621_, new_n44622_,
    new_n44624_, new_n44625_, new_n44626_, new_n44627_, new_n44628_,
    new_n44629_, new_n44630_, new_n44632_, new_n44634_, new_n44636_,
    new_n44637_, new_n44638_, new_n44639_, new_n44641_, new_n44642_,
    new_n44643_, new_n44644_, new_n44645_, new_n44646_, new_n44647_,
    new_n44648_, new_n44650_, new_n44651_, new_n44652_, new_n44654_,
    new_n44655_, new_n44656_, new_n44658_, new_n44659_, new_n44660_,
    new_n44662_, new_n44663_, new_n44664_, new_n44666_, new_n44667_,
    new_n44668_, new_n44670_, new_n44671_, new_n44672_, new_n44674_,
    new_n44675_, new_n44676_, new_n44678_, new_n44679_, new_n44680_,
    new_n44682_, new_n44683_, new_n44684_, new_n44686_, new_n44687_,
    new_n44688_, new_n44690_, new_n44691_, new_n44692_, new_n44694_,
    new_n44695_, new_n44696_, new_n44698_, new_n44699_, new_n44700_,
    new_n44702_, new_n44703_, new_n44704_, new_n44706_, new_n44707_,
    new_n44708_, new_n44710_, new_n44711_, new_n44712_, new_n44714_,
    new_n44715_, new_n44716_, new_n44718_, new_n44719_, new_n44720_,
    new_n44722_, new_n44723_, new_n44724_, new_n44726_, new_n44727_,
    new_n44728_, new_n44730_, new_n44731_, new_n44732_, new_n44734_,
    new_n44735_, new_n44736_, new_n44738_, new_n44739_, new_n44740_,
    new_n44742_, new_n44743_, new_n44744_, new_n44746_, new_n44747_,
    new_n44748_, new_n44750_, new_n44751_, new_n44752_, new_n44754_,
    new_n44755_, new_n44756_, new_n44758_, new_n44759_, new_n44760_,
    new_n44762_, new_n44763_, new_n44764_, new_n44766_, new_n44767_,
    new_n44768_, new_n44770_, new_n44771_, new_n44772_, new_n44774_,
    new_n44775_, new_n44776_, new_n44778_, new_n44779_, new_n44780_,
    new_n44782_, new_n44783_, new_n44784_, new_n44786_, new_n44787_,
    new_n44788_, new_n44789_, new_n44790_, new_n44791_, new_n44792_,
    new_n44793_, new_n44795_, new_n44796_, new_n44797_, new_n44799_,
    new_n44800_, new_n44801_, new_n44803_, new_n44804_, new_n44805_,
    new_n44807_, new_n44808_, new_n44809_, new_n44811_, new_n44812_,
    new_n44813_, new_n44815_, new_n44816_, new_n44817_, new_n44819_,
    new_n44820_, new_n44821_, new_n44823_, new_n44824_, new_n44825_,
    new_n44827_, new_n44828_, new_n44829_, new_n44831_, new_n44832_,
    new_n44833_, new_n44835_, new_n44836_, new_n44837_, new_n44839_,
    new_n44840_, new_n44841_, new_n44843_, new_n44844_, new_n44845_,
    new_n44847_, new_n44848_, new_n44849_, new_n44851_, new_n44852_,
    new_n44853_, new_n44855_, new_n44856_, new_n44857_, new_n44859_,
    new_n44860_, new_n44861_, new_n44863_, new_n44864_, new_n44865_,
    new_n44867_, new_n44868_, new_n44869_, new_n44871_, new_n44872_,
    new_n44873_, new_n44875_, new_n44876_, new_n44877_, new_n44879_,
    new_n44880_, new_n44881_, new_n44883_, new_n44884_, new_n44885_,
    new_n44887_, new_n44888_, new_n44889_, new_n44891_, new_n44892_,
    new_n44893_, new_n44895_, new_n44896_, new_n44897_, new_n44899_,
    new_n44900_, new_n44901_, new_n44903_, new_n44904_, new_n44905_,
    new_n44907_, new_n44908_, new_n44909_, new_n44911_, new_n44912_,
    new_n44913_, new_n44915_, new_n44916_, new_n44917_, new_n44919_,
    new_n44920_, new_n44921_, new_n44923_, new_n44924_, new_n44925_,
    new_n44927_, new_n44928_, new_n44929_, new_n44931_, new_n44932_,
    new_n44933_, new_n44934_, new_n44935_, new_n44936_, new_n44937_,
    new_n44938_, new_n44940_, new_n44941_, new_n44942_, new_n44944_,
    new_n44945_, new_n44946_, new_n44948_, new_n44949_, new_n44950_,
    new_n44952_, new_n44953_, new_n44954_, new_n44956_, new_n44957_,
    new_n44958_, new_n44960_, new_n44961_, new_n44962_, new_n44964_,
    new_n44965_, new_n44966_, new_n44968_, new_n44969_, new_n44970_,
    new_n44972_, new_n44973_, new_n44974_, new_n44976_, new_n44977_,
    new_n44978_, new_n44980_, new_n44981_, new_n44982_, new_n44984_,
    new_n44985_, new_n44986_, new_n44988_, new_n44989_, new_n44990_,
    new_n44992_, new_n44993_, new_n44994_, new_n44996_, new_n44997_,
    new_n44998_, new_n45000_, new_n45001_, new_n45002_, new_n45004_,
    new_n45005_, new_n45006_, new_n45008_, new_n45009_, new_n45010_,
    new_n45012_, new_n45013_, new_n45014_, new_n45016_, new_n45017_,
    new_n45018_, new_n45020_, new_n45021_, new_n45022_, new_n45024_,
    new_n45025_, new_n45026_, new_n45028_, new_n45029_, new_n45030_,
    new_n45032_, new_n45033_, new_n45034_, new_n45036_, new_n45037_,
    new_n45038_, new_n45040_, new_n45041_, new_n45042_, new_n45044_,
    new_n45045_, new_n45046_, new_n45048_, new_n45049_, new_n45050_,
    new_n45052_, new_n45053_, new_n45054_, new_n45056_, new_n45057_,
    new_n45058_, new_n45060_, new_n45061_, new_n45062_, new_n45064_,
    new_n45065_, new_n45066_, new_n45068_, new_n45069_, new_n45070_,
    new_n45072_, new_n45073_, new_n45074_, new_n45076_, new_n45077_,
    new_n45078_, new_n45079_, new_n45080_, new_n45081_, new_n45082_,
    new_n45083_, new_n45085_, new_n45086_, new_n45087_, new_n45089_,
    new_n45090_, new_n45091_, new_n45093_, new_n45094_, new_n45095_,
    new_n45097_, new_n45098_, new_n45099_, new_n45101_, new_n45102_,
    new_n45103_, new_n45105_, new_n45106_, new_n45107_, new_n45109_,
    new_n45110_, new_n45111_, new_n45113_, new_n45114_, new_n45115_,
    new_n45117_, new_n45118_, new_n45119_, new_n45121_, new_n45122_,
    new_n45123_, new_n45125_, new_n45126_, new_n45127_, new_n45129_,
    new_n45130_, new_n45131_, new_n45133_, new_n45134_, new_n45135_,
    new_n45137_, new_n45138_, new_n45139_, new_n45141_, new_n45142_,
    new_n45143_, new_n45145_, new_n45146_, new_n45147_, new_n45149_,
    new_n45150_, new_n45151_, new_n45153_, new_n45154_, new_n45155_,
    new_n45157_, new_n45158_, new_n45159_, new_n45161_, new_n45162_,
    new_n45163_, new_n45165_, new_n45166_, new_n45167_, new_n45169_,
    new_n45170_, new_n45171_, new_n45173_, new_n45174_, new_n45175_,
    new_n45177_, new_n45178_, new_n45179_, new_n45181_, new_n45182_,
    new_n45183_, new_n45185_, new_n45186_, new_n45187_, new_n45189_,
    new_n45190_, new_n45191_, new_n45193_, new_n45194_, new_n45195_,
    new_n45197_, new_n45198_, new_n45199_, new_n45201_, new_n45202_,
    new_n45203_, new_n45205_, new_n45206_, new_n45207_, new_n45209_,
    new_n45210_, new_n45211_, new_n45213_, new_n45214_, new_n45215_,
    new_n45217_, new_n45218_, new_n45219_, new_n45221_, new_n45222_,
    new_n45223_, new_n45224_, new_n45225_, new_n45226_, new_n45227_,
    new_n45228_, new_n45230_, new_n45231_, new_n45232_, new_n45234_,
    new_n45235_, new_n45236_, new_n45238_, new_n45239_, new_n45240_,
    new_n45242_, new_n45243_, new_n45244_, new_n45246_, new_n45247_,
    new_n45248_, new_n45250_, new_n45251_, new_n45252_, new_n45254_,
    new_n45255_, new_n45256_, new_n45258_, new_n45259_, new_n45260_,
    new_n45262_, new_n45263_, new_n45264_, new_n45266_, new_n45267_,
    new_n45268_, new_n45270_, new_n45271_, new_n45272_, new_n45274_,
    new_n45275_, new_n45276_, new_n45278_, new_n45279_, new_n45280_,
    new_n45282_, new_n45283_, new_n45284_, new_n45286_, new_n45287_,
    new_n45288_, new_n45290_, new_n45291_, new_n45292_, new_n45294_,
    new_n45295_, new_n45296_, new_n45298_, new_n45299_, new_n45300_,
    new_n45302_, new_n45303_, new_n45304_, new_n45306_, new_n45307_,
    new_n45308_, new_n45310_, new_n45311_, new_n45312_, new_n45314_,
    new_n45315_, new_n45316_, new_n45318_, new_n45319_, new_n45320_,
    new_n45322_, new_n45323_, new_n45324_, new_n45326_, new_n45327_,
    new_n45328_, new_n45330_, new_n45331_, new_n45332_, new_n45334_,
    new_n45335_, new_n45336_, new_n45338_, new_n45339_, new_n45340_,
    new_n45342_, new_n45343_, new_n45344_, new_n45346_, new_n45347_,
    new_n45348_, new_n45350_, new_n45351_, new_n45352_, new_n45354_,
    new_n45355_, new_n45356_, new_n45358_, new_n45359_, new_n45360_,
    new_n45362_, new_n45363_, new_n45364_, new_n45366_, new_n45367_,
    new_n45368_, new_n45369_, new_n45370_, new_n45371_, new_n45372_,
    new_n45373_, new_n45375_, new_n45376_, new_n45377_, new_n45379_,
    new_n45380_, new_n45381_, new_n45383_, new_n45384_, new_n45385_,
    new_n45387_, new_n45388_, new_n45389_, new_n45391_, new_n45392_,
    new_n45393_, new_n45395_, new_n45396_, new_n45397_, new_n45399_,
    new_n45400_, new_n45401_, new_n45403_, new_n45404_, new_n45405_,
    new_n45407_, new_n45408_, new_n45409_, new_n45411_, new_n45412_,
    new_n45413_, new_n45415_, new_n45416_, new_n45417_, new_n45419_,
    new_n45420_, new_n45421_, new_n45423_, new_n45424_, new_n45425_,
    new_n45427_, new_n45428_, new_n45429_, new_n45431_, new_n45432_,
    new_n45433_, new_n45435_, new_n45436_, new_n45437_, new_n45439_,
    new_n45440_, new_n45441_, new_n45443_, new_n45444_, new_n45445_,
    new_n45447_, new_n45448_, new_n45449_, new_n45451_, new_n45452_,
    new_n45453_, new_n45455_, new_n45456_, new_n45457_, new_n45459_,
    new_n45460_, new_n45461_, new_n45463_, new_n45464_, new_n45465_,
    new_n45467_, new_n45468_, new_n45469_, new_n45471_, new_n45472_,
    new_n45473_, new_n45475_, new_n45476_, new_n45477_, new_n45479_,
    new_n45480_, new_n45481_, new_n45483_, new_n45484_, new_n45485_,
    new_n45487_, new_n45488_, new_n45489_, new_n45491_, new_n45492_,
    new_n45493_, new_n45495_, new_n45496_, new_n45497_, new_n45499_,
    new_n45500_, new_n45501_, new_n45503_, new_n45504_, new_n45505_,
    new_n45507_, new_n45508_, new_n45509_, new_n45511_, new_n45512_,
    new_n45513_, new_n45514_, new_n45515_, new_n45516_, new_n45517_,
    new_n45518_, new_n45519_, new_n45520_, new_n45521_, new_n45522_,
    new_n45523_, new_n45524_, new_n45525_, new_n45526_, new_n45527_,
    new_n45528_, new_n45529_, new_n45530_, new_n45531_, new_n45532_,
    new_n45533_, new_n45534_, new_n45535_, new_n45536_, new_n45537_,
    new_n45538_, new_n45539_, new_n45540_, new_n45541_, new_n45542_,
    new_n45543_, new_n45544_, new_n45545_, new_n45546_, new_n45547_,
    new_n45548_, new_n45549_, new_n45550_, new_n45551_, new_n45552_,
    new_n45553_, new_n45554_, new_n45555_, new_n45556_, new_n45557_,
    new_n45558_, new_n45559_, new_n45560_, new_n45561_, new_n45562_,
    new_n45563_, new_n45564_, new_n45565_, new_n45566_, new_n45567_,
    new_n45568_, new_n45569_, new_n45570_, new_n45571_, new_n45572_,
    new_n45573_, new_n45574_, new_n45575_, new_n45576_, new_n45577_,
    new_n45578_, new_n45579_, new_n45580_, new_n45581_, new_n45582_,
    new_n45583_, new_n45584_, new_n45585_, new_n45586_, new_n45587_,
    new_n45588_, new_n45589_, new_n45590_, new_n45591_, new_n45592_,
    new_n45593_, new_n45594_, new_n45595_, new_n45596_, new_n45597_,
    new_n45598_, new_n45599_, new_n45601_, new_n45602_, new_n45603_,
    new_n45604_, new_n45605_, new_n45606_, new_n45607_, new_n45608_,
    new_n45609_, new_n45610_, new_n45611_, new_n45612_, new_n45613_,
    new_n45614_, new_n45615_, new_n45616_, new_n45617_, new_n45618_,
    new_n45619_, new_n45620_, new_n45621_, new_n45622_, new_n45623_,
    new_n45624_, new_n45625_, new_n45626_, new_n45627_, new_n45628_,
    new_n45629_, new_n45630_, new_n45631_, new_n45632_, new_n45633_,
    new_n45634_, new_n45635_, new_n45637_, new_n45638_, new_n45639_,
    new_n45640_, new_n45641_, new_n45642_, new_n45643_, new_n45644_,
    new_n45645_, new_n45646_, new_n45648_, new_n45649_, new_n45650_,
    new_n45651_, new_n45652_, new_n45653_, new_n45654_, new_n45655_,
    new_n45656_, new_n45658_, new_n45659_, new_n45660_, new_n45661_,
    new_n45662_, new_n45663_, new_n45664_, new_n45665_, new_n45666_,
    new_n45667_, new_n45668_, new_n45670_, new_n45671_, new_n45672_,
    new_n45673_, new_n45674_, new_n45675_, new_n45676_, new_n45677_,
    new_n45678_, new_n45679_, new_n45681_, new_n45682_, new_n45683_,
    new_n45684_, new_n45685_, new_n45686_, new_n45687_, new_n45688_,
    new_n45689_, new_n45690_, new_n45692_, new_n45693_, new_n45694_,
    new_n45695_, new_n45696_, new_n45697_, new_n45698_, new_n45699_,
    new_n45700_, new_n45701_, new_n45703_, new_n45704_, new_n45705_,
    new_n45706_, new_n45707_, new_n45708_, new_n45709_, new_n45710_,
    new_n45711_, new_n45712_, new_n45713_, new_n45714_, new_n45716_,
    new_n45717_, new_n45718_, new_n45719_, new_n45720_, new_n45721_,
    new_n45722_, new_n45723_, new_n45724_, new_n45725_, new_n45727_,
    new_n45728_, new_n45729_, new_n45730_, new_n45731_, new_n45732_,
    new_n45733_, new_n45734_, new_n45735_, new_n45736_, new_n45737_,
    new_n45738_, new_n45740_, new_n45741_, new_n45752_, new_n45753_,
    new_n45755_, new_n45756_, new_n45758_, new_n45759_, new_n45760_,
    new_n45761_, new_n45763_, new_n45764_, new_n45765_, new_n45766_,
    new_n45769_, new_n45770_, new_n45772_, new_n45774_, new_n45776_,
    new_n45778_, new_n45779_, new_n45780_, new_n45781_, new_n45782_,
    new_n45783_, new_n45784_, new_n45785_, new_n45786_, new_n45787_,
    new_n45788_, new_n45789_, new_n45790_, new_n45791_, new_n45792_,
    new_n45793_, new_n45794_, new_n45795_, new_n45796_, new_n45797_,
    new_n45798_, new_n45799_, new_n45800_, new_n45801_, new_n45802_,
    new_n45803_, new_n45807_, new_n45808_, new_n45809_, new_n45811_,
    new_n45812_, new_n45813_, new_n45815_, new_n45816_, new_n45817_,
    new_n45819_, new_n45820_, new_n45821_, new_n45823_, new_n45824_,
    new_n45825_, new_n45827_, new_n45828_, new_n45829_, new_n45831_,
    new_n45832_, new_n45833_, new_n45835_, new_n45836_, new_n45837_,
    new_n45839_, new_n45840_, new_n45841_, new_n45843_, new_n45844_,
    new_n45845_, new_n45847_, new_n45848_, new_n45849_, new_n45851_,
    new_n45852_, new_n45853_, new_n45855_, new_n45856_, new_n45857_,
    new_n45859_, new_n45860_, new_n45861_, new_n45863_, new_n45864_,
    new_n45865_, new_n45867_, new_n45868_, new_n45869_, new_n45871_,
    new_n45872_, new_n45873_, new_n45875_, new_n45876_, new_n45877_,
    new_n45879_, new_n45880_, new_n45881_, new_n45883_, new_n45884_,
    new_n45885_, new_n45887_, new_n45888_, new_n45889_, new_n45891_,
    new_n45892_, new_n45893_, new_n45895_, new_n45896_, new_n45897_,
    new_n45899_, new_n45900_, new_n45901_, new_n45903_, new_n45904_,
    new_n45905_, new_n45907_, new_n45908_, new_n45909_, new_n45911_,
    new_n45912_, new_n45913_, new_n45915_, new_n45916_, new_n45917_,
    new_n45919_, new_n45920_, new_n45921_, new_n45923_, new_n45924_,
    new_n45925_, new_n45927_, new_n45928_, new_n45929_, new_n45931_,
    new_n45932_, new_n45933_, new_n45935_, new_n45936_, new_n45937_,
    new_n45938_, new_n45939_, new_n45940_, new_n45941_, new_n45942_,
    new_n45943_, new_n45944_, new_n45945_, new_n45946_, new_n45947_,
    new_n45948_, new_n45949_, new_n45951_, new_n45952_, new_n45953_,
    new_n45954_, new_n45955_, new_n45956_, new_n45957_, new_n45959_,
    new_n45960_, new_n45961_, new_n45962_, new_n45963_, new_n45964_,
    new_n45965_, new_n45967_, new_n45968_, new_n45969_, new_n45970_,
    new_n45971_, new_n45972_, new_n45973_, new_n45975_, new_n45976_,
    new_n45977_, new_n45978_, new_n45979_, new_n45980_, new_n45981_,
    new_n45983_, new_n45984_, new_n45985_, new_n45986_, new_n45987_,
    new_n45988_, new_n45989_, new_n45991_, new_n45992_, new_n45993_,
    new_n45994_, new_n45995_, new_n45996_, new_n45997_, new_n45999_,
    new_n46000_, new_n46001_, new_n46002_, new_n46003_, new_n46004_,
    new_n46005_, new_n46007_, new_n46008_, new_n46009_, new_n46010_,
    new_n46011_, new_n46012_, new_n46013_, new_n46015_, new_n46016_,
    new_n46017_, new_n46018_, new_n46019_, new_n46020_, new_n46021_,
    new_n46023_, new_n46024_, new_n46025_, new_n46026_, new_n46027_,
    new_n46028_, new_n46029_, new_n46031_, new_n46032_, new_n46033_,
    new_n46034_, new_n46035_, new_n46036_, new_n46037_, new_n46039_,
    new_n46040_, new_n46041_, new_n46042_, new_n46043_, new_n46044_,
    new_n46045_, new_n46047_, new_n46048_, new_n46049_, new_n46050_,
    new_n46051_, new_n46052_, new_n46053_, new_n46055_, new_n46056_,
    new_n46057_, new_n46058_, new_n46059_, new_n46060_, new_n46061_,
    new_n46063_, new_n46064_, new_n46065_, new_n46066_, new_n46067_,
    new_n46068_, new_n46069_, new_n46071_, new_n46072_, new_n46073_,
    new_n46074_, new_n46075_, new_n46076_, new_n46077_, new_n46079_,
    new_n46080_, new_n46081_, new_n46082_, new_n46083_, new_n46084_,
    new_n46085_, new_n46087_, new_n46088_, new_n46089_, new_n46090_,
    new_n46091_, new_n46092_, new_n46093_, new_n46095_, new_n46096_,
    new_n46097_, new_n46098_, new_n46099_, new_n46100_, new_n46101_,
    new_n46103_, new_n46104_, new_n46105_, new_n46106_, new_n46107_,
    new_n46108_, new_n46109_, new_n46111_, new_n46112_, new_n46113_,
    new_n46114_, new_n46115_, new_n46116_, new_n46117_, new_n46119_,
    new_n46120_, new_n46121_, new_n46122_, new_n46123_, new_n46124_,
    new_n46125_, new_n46127_, new_n46128_, new_n46129_, new_n46130_,
    new_n46131_, new_n46132_, new_n46133_, new_n46135_, new_n46136_,
    new_n46137_, new_n46138_, new_n46139_, new_n46140_, new_n46141_,
    new_n46143_, new_n46144_, new_n46145_, new_n46146_, new_n46147_,
    new_n46148_, new_n46149_, new_n46151_, new_n46152_, new_n46153_,
    new_n46154_, new_n46155_, new_n46156_, new_n46157_, new_n46159_,
    new_n46160_, new_n46161_, new_n46162_, new_n46163_, new_n46164_,
    new_n46165_, new_n46167_, new_n46168_, new_n46169_, new_n46170_,
    new_n46171_, new_n46172_, new_n46173_, new_n46175_, new_n46176_,
    new_n46177_, new_n46178_, new_n46179_, new_n46180_, new_n46181_,
    new_n46183_, new_n46184_, new_n46185_, new_n46186_, new_n46187_,
    new_n46188_, new_n46189_, new_n46191_, new_n46192_, new_n46193_,
    new_n46194_, new_n46195_, new_n46196_, new_n46197_, new_n46199_,
    new_n46200_, new_n46201_, new_n46202_, new_n46203_, new_n46204_,
    new_n46205_, new_n46206_, new_n46207_, new_n46208_, new_n46209_,
    new_n46210_, new_n46211_, new_n46212_, new_n46213_, new_n46214_,
    new_n46215_, new_n46216_, new_n46217_, new_n46218_, new_n46219_,
    new_n46220_, new_n46221_, new_n46222_, new_n46223_, new_n46224_,
    new_n46225_, new_n46226_, new_n46227_, new_n46228_, new_n46229_,
    new_n46230_, new_n46231_, new_n46232_, new_n46233_, new_n46234_,
    new_n46235_, new_n46236_, new_n46237_, new_n46238_, new_n46239_,
    new_n46240_, new_n46241_, new_n46242_, new_n46243_, new_n46244_,
    new_n46245_, new_n46246_, new_n46247_, new_n46248_, new_n46249_,
    new_n46250_, new_n46251_, new_n46252_, new_n46253_, new_n46254_,
    new_n46255_, new_n46256_, new_n46257_, new_n46258_, new_n46259_,
    new_n46260_, new_n46261_, new_n46262_, new_n46263_, new_n46264_,
    new_n46265_, new_n46266_, new_n46267_, new_n46269_, new_n46270_,
    new_n46271_, new_n46272_, new_n46273_, new_n46274_, new_n46275_,
    new_n46276_, new_n46277_, new_n46278_, new_n46279_, new_n46280_,
    new_n46281_, new_n46282_, new_n46283_, new_n46284_, new_n46285_,
    new_n46286_, new_n46287_, new_n46288_, new_n46289_, new_n46290_,
    new_n46291_, new_n46292_, new_n46293_, new_n46294_, new_n46295_,
    new_n46296_, new_n46297_, new_n46298_, new_n46299_, new_n46300_,
    new_n46301_, new_n46302_, new_n46303_, new_n46304_, new_n46306_,
    new_n46307_, new_n46308_, new_n46309_, new_n46310_, new_n46311_,
    new_n46312_, new_n46313_, new_n46314_, new_n46315_, new_n46316_,
    new_n46317_, new_n46318_, new_n46319_, new_n46320_, new_n46321_,
    new_n46322_, new_n46323_, new_n46324_, new_n46325_, new_n46326_,
    new_n46327_, new_n46328_, new_n46329_, new_n46330_, new_n46331_,
    new_n46332_, new_n46333_, new_n46334_, new_n46335_, new_n46336_,
    new_n46337_, new_n46338_, new_n46339_, new_n46340_, new_n46341_,
    new_n46342_, new_n46343_, new_n46345_, new_n46346_, new_n46347_,
    new_n46348_, new_n46349_, new_n46350_, new_n46351_, new_n46352_,
    new_n46353_, new_n46354_, new_n46355_, new_n46356_, new_n46357_,
    new_n46358_, new_n46359_, new_n46360_, new_n46361_, new_n46362_,
    new_n46363_, new_n46364_, new_n46365_, new_n46366_, new_n46367_,
    new_n46368_, new_n46369_, new_n46370_, new_n46371_, new_n46372_,
    new_n46373_, new_n46374_, new_n46375_, new_n46376_, new_n46377_,
    new_n46378_, new_n46379_, new_n46380_, new_n46381_, new_n46382_,
    new_n46384_, new_n46385_, new_n46386_, new_n46387_, new_n46388_,
    new_n46389_, new_n46390_, new_n46391_, new_n46392_, new_n46393_,
    new_n46394_, new_n46395_, new_n46396_, new_n46397_, new_n46398_,
    new_n46399_, new_n46400_, new_n46401_, new_n46402_, new_n46403_,
    new_n46404_, new_n46405_, new_n46406_, new_n46407_, new_n46408_,
    new_n46409_, new_n46410_, new_n46411_, new_n46412_, new_n46413_,
    new_n46414_, new_n46415_, new_n46416_, new_n46417_, new_n46418_,
    new_n46419_, new_n46421_, new_n46422_, new_n46423_, new_n46424_,
    new_n46425_, new_n46426_, new_n46427_, new_n46428_, new_n46429_,
    new_n46430_, new_n46431_, new_n46432_, new_n46433_, new_n46434_,
    new_n46435_, new_n46436_, new_n46437_, new_n46438_, new_n46439_,
    new_n46440_, new_n46441_, new_n46442_, new_n46443_, new_n46444_,
    new_n46445_, new_n46446_, new_n46447_, new_n46448_, new_n46449_,
    new_n46450_, new_n46452_, new_n46453_, new_n46454_, new_n46455_,
    new_n46456_, new_n46457_, new_n46458_, new_n46459_, new_n46460_,
    new_n46461_, new_n46462_, new_n46463_, new_n46464_, new_n46465_,
    new_n46466_, new_n46467_, new_n46468_, new_n46469_, new_n46470_,
    new_n46471_, new_n46472_, new_n46473_, new_n46474_, new_n46475_,
    new_n46476_, new_n46477_, new_n46478_, new_n46479_, new_n46480_,
    new_n46481_, new_n46483_, new_n46484_, new_n46485_, new_n46486_,
    new_n46487_, new_n46488_, new_n46489_, new_n46490_, new_n46491_,
    new_n46492_, new_n46493_, new_n46494_, new_n46495_, new_n46496_,
    new_n46497_, new_n46498_, new_n46499_, new_n46500_, new_n46501_,
    new_n46502_, new_n46503_, new_n46504_, new_n46505_, new_n46506_,
    new_n46507_, new_n46508_, new_n46509_, new_n46510_, new_n46511_,
    new_n46512_, new_n46514_, new_n46515_, new_n46516_, new_n46517_,
    new_n46518_, new_n46519_, new_n46520_, new_n46521_, new_n46522_,
    new_n46523_, new_n46524_, new_n46525_, new_n46526_, new_n46527_,
    new_n46528_, new_n46529_, new_n46530_, new_n46531_, new_n46532_,
    new_n46533_, new_n46534_, new_n46535_, new_n46536_, new_n46537_,
    new_n46538_, new_n46539_, new_n46540_, new_n46541_, new_n46542_,
    new_n46543_, new_n46545_, new_n46546_, new_n46547_, new_n46548_,
    new_n46549_, new_n46550_, new_n46551_, new_n46552_, new_n46553_,
    new_n46554_, new_n46555_, new_n46556_, new_n46557_, new_n46558_,
    new_n46559_, new_n46560_, new_n46561_, new_n46562_, new_n46563_,
    new_n46564_, new_n46565_, new_n46566_, new_n46567_, new_n46568_,
    new_n46569_, new_n46570_, new_n46571_, new_n46572_, new_n46573_,
    new_n46574_, new_n46576_, new_n46577_, new_n46578_, new_n46579_,
    new_n46580_, new_n46581_, new_n46582_, new_n46583_, new_n46584_,
    new_n46585_, new_n46586_, new_n46587_, new_n46588_, new_n46589_,
    new_n46590_, new_n46591_, new_n46592_, new_n46593_, new_n46594_,
    new_n46595_, new_n46596_, new_n46597_, new_n46598_, new_n46599_,
    new_n46600_, new_n46601_, new_n46602_, new_n46603_, new_n46604_,
    new_n46605_, new_n46607_, new_n46608_, new_n46609_, new_n46610_,
    new_n46611_, new_n46612_, new_n46613_, new_n46614_, new_n46615_,
    new_n46616_, new_n46617_, new_n46618_, new_n46619_, new_n46620_,
    new_n46621_, new_n46622_, new_n46623_, new_n46624_, new_n46625_,
    new_n46626_, new_n46627_, new_n46628_, new_n46629_, new_n46630_,
    new_n46631_, new_n46632_, new_n46633_, new_n46634_, new_n46635_,
    new_n46636_, new_n46638_, new_n46639_, new_n46640_, new_n46641_,
    new_n46642_, new_n46643_, new_n46644_, new_n46645_, new_n46646_,
    new_n46647_, new_n46648_, new_n46649_, new_n46650_, new_n46651_,
    new_n46652_, new_n46653_, new_n46654_, new_n46655_, new_n46656_,
    new_n46657_, new_n46658_, new_n46659_, new_n46660_, new_n46661_,
    new_n46662_, new_n46663_, new_n46664_, new_n46665_, new_n46666_,
    new_n46667_, new_n46669_, new_n46670_, new_n46671_, new_n46672_,
    new_n46673_, new_n46674_, new_n46675_, new_n46676_, new_n46677_,
    new_n46678_, new_n46679_, new_n46680_, new_n46681_, new_n46682_,
    new_n46683_, new_n46684_, new_n46685_, new_n46686_, new_n46687_,
    new_n46688_, new_n46689_, new_n46690_, new_n46691_, new_n46692_,
    new_n46693_, new_n46694_, new_n46695_, new_n46696_, new_n46697_,
    new_n46698_, new_n46700_, new_n46701_, new_n46702_, new_n46703_,
    new_n46704_, new_n46705_, new_n46706_, new_n46707_, new_n46708_,
    new_n46709_, new_n46710_, new_n46711_, new_n46712_, new_n46713_,
    new_n46714_, new_n46715_, new_n46716_, new_n46717_, new_n46718_,
    new_n46719_, new_n46720_, new_n46721_, new_n46722_, new_n46723_,
    new_n46724_, new_n46725_, new_n46726_, new_n46727_, new_n46728_,
    new_n46729_, new_n46731_, new_n46732_, new_n46733_, new_n46734_,
    new_n46735_, new_n46736_, new_n46737_, new_n46738_, new_n46739_,
    new_n46740_, new_n46741_, new_n46742_, new_n46743_, new_n46744_,
    new_n46745_, new_n46746_, new_n46747_, new_n46748_, new_n46749_,
    new_n46750_, new_n46751_, new_n46752_, new_n46753_, new_n46754_,
    new_n46755_, new_n46756_, new_n46757_, new_n46758_, new_n46759_,
    new_n46760_, new_n46762_, new_n46763_, new_n46764_, new_n46765_,
    new_n46766_, new_n46767_, new_n46768_, new_n46769_, new_n46770_,
    new_n46771_, new_n46772_, new_n46773_, new_n46774_, new_n46775_,
    new_n46776_, new_n46777_, new_n46778_, new_n46779_, new_n46780_,
    new_n46781_, new_n46782_, new_n46783_, new_n46784_, new_n46785_,
    new_n46786_, new_n46787_, new_n46788_, new_n46789_, new_n46790_,
    new_n46791_, new_n46793_, new_n46794_, new_n46795_, new_n46796_,
    new_n46797_, new_n46798_, new_n46799_, new_n46800_, new_n46801_,
    new_n46802_, new_n46803_, new_n46804_, new_n46805_, new_n46806_,
    new_n46807_, new_n46808_, new_n46809_, new_n46810_, new_n46811_,
    new_n46812_, new_n46813_, new_n46814_, new_n46815_, new_n46816_,
    new_n46817_, new_n46818_, new_n46819_, new_n46820_, new_n46821_,
    new_n46822_, new_n46824_, new_n46825_, new_n46826_, new_n46827_,
    new_n46828_, new_n46829_, new_n46830_, new_n46831_, new_n46832_,
    new_n46833_, new_n46834_, new_n46835_, new_n46836_, new_n46837_,
    new_n46838_, new_n46839_, new_n46840_, new_n46841_, new_n46842_,
    new_n46843_, new_n46844_, new_n46845_, new_n46846_, new_n46847_,
    new_n46848_, new_n46849_, new_n46850_, new_n46851_, new_n46852_,
    new_n46853_, new_n46855_, new_n46856_, new_n46857_, new_n46858_,
    new_n46859_, new_n46860_, new_n46861_, new_n46862_, new_n46863_,
    new_n46864_, new_n46865_, new_n46866_, new_n46867_, new_n46868_,
    new_n46869_, new_n46870_, new_n46871_, new_n46872_, new_n46873_,
    new_n46874_, new_n46875_, new_n46876_, new_n46877_, new_n46878_,
    new_n46879_, new_n46880_, new_n46881_, new_n46882_, new_n46883_,
    new_n46884_, new_n46886_, new_n46887_, new_n46888_, new_n46889_,
    new_n46890_, new_n46891_, new_n46892_, new_n46893_, new_n46894_,
    new_n46895_, new_n46896_, new_n46897_, new_n46898_, new_n46899_,
    new_n46900_, new_n46901_, new_n46902_, new_n46903_, new_n46904_,
    new_n46905_, new_n46906_, new_n46907_, new_n46908_, new_n46909_,
    new_n46910_, new_n46911_, new_n46912_, new_n46913_, new_n46914_,
    new_n46915_, new_n46917_, new_n46918_, new_n46919_, new_n46920_,
    new_n46921_, new_n46922_, new_n46923_, new_n46924_, new_n46925_,
    new_n46926_, new_n46927_, new_n46928_, new_n46929_, new_n46930_,
    new_n46931_, new_n46932_, new_n46933_, new_n46934_, new_n46935_,
    new_n46936_, new_n46937_, new_n46938_, new_n46939_, new_n46940_,
    new_n46941_, new_n46942_, new_n46943_, new_n46944_, new_n46945_,
    new_n46946_, new_n46948_, new_n46949_, new_n46950_, new_n46951_,
    new_n46952_, new_n46953_, new_n46954_, new_n46955_, new_n46956_,
    new_n46957_, new_n46958_, new_n46959_, new_n46960_, new_n46961_,
    new_n46962_, new_n46963_, new_n46964_, new_n46965_, new_n46966_,
    new_n46967_, new_n46968_, new_n46969_, new_n46970_, new_n46971_,
    new_n46972_, new_n46973_, new_n46974_, new_n46975_, new_n46976_,
    new_n46977_, new_n46979_, new_n46980_, new_n46981_, new_n46982_,
    new_n46983_, new_n46984_, new_n46985_, new_n46986_, new_n46987_,
    new_n46988_, new_n46989_, new_n46990_, new_n46991_, new_n46992_,
    new_n46993_, new_n46994_, new_n46995_, new_n46996_, new_n46997_,
    new_n46998_, new_n46999_, new_n47000_, new_n47001_, new_n47002_,
    new_n47003_, new_n47004_, new_n47005_, new_n47006_, new_n47007_,
    new_n47008_, new_n47010_, new_n47011_, new_n47012_, new_n47013_,
    new_n47014_, new_n47015_, new_n47016_, new_n47017_, new_n47018_,
    new_n47019_, new_n47020_, new_n47021_, new_n47022_, new_n47023_,
    new_n47024_, new_n47025_, new_n47026_, new_n47027_, new_n47028_,
    new_n47029_, new_n47030_, new_n47031_, new_n47032_, new_n47033_,
    new_n47034_, new_n47035_, new_n47036_, new_n47037_, new_n47038_,
    new_n47039_, new_n47041_, new_n47042_, new_n47043_, new_n47044_,
    new_n47045_, new_n47046_, new_n47047_, new_n47048_, new_n47049_,
    new_n47050_, new_n47051_, new_n47052_, new_n47053_, new_n47054_,
    new_n47055_, new_n47056_, new_n47057_, new_n47058_, new_n47059_,
    new_n47060_, new_n47061_, new_n47062_, new_n47063_, new_n47064_,
    new_n47065_, new_n47066_, new_n47067_, new_n47068_, new_n47069_,
    new_n47070_, new_n47072_, new_n47073_, new_n47074_, new_n47075_,
    new_n47076_, new_n47077_, new_n47078_, new_n47079_, new_n47080_,
    new_n47081_, new_n47082_, new_n47083_, new_n47084_, new_n47085_,
    new_n47086_, new_n47087_, new_n47088_, new_n47089_, new_n47090_,
    new_n47091_, new_n47092_, new_n47093_, new_n47094_, new_n47095_,
    new_n47096_, new_n47097_, new_n47098_, new_n47099_, new_n47100_,
    new_n47101_, new_n47103_, new_n47104_, new_n47105_, new_n47106_,
    new_n47107_, new_n47108_, new_n47109_, new_n47110_, new_n47111_,
    new_n47112_, new_n47113_, new_n47114_, new_n47115_, new_n47116_,
    new_n47117_, new_n47118_, new_n47119_, new_n47120_, new_n47121_,
    new_n47122_, new_n47123_, new_n47124_, new_n47125_, new_n47126_,
    new_n47127_, new_n47128_, new_n47129_, new_n47130_, new_n47131_,
    new_n47132_, new_n47134_, new_n47135_, new_n47136_, new_n47137_,
    new_n47138_, new_n47139_, new_n47140_, new_n47141_, new_n47142_,
    new_n47143_, new_n47144_, new_n47145_, new_n47146_, new_n47147_,
    new_n47148_, new_n47149_, new_n47150_, new_n47151_, new_n47152_,
    new_n47153_, new_n47154_, new_n47155_, new_n47156_, new_n47157_,
    new_n47158_, new_n47159_, new_n47160_, new_n47161_, new_n47162_,
    new_n47163_, new_n47165_, new_n47166_, new_n47167_, new_n47168_,
    new_n47169_, new_n47170_, new_n47171_, new_n47172_, new_n47173_,
    new_n47174_, new_n47175_, new_n47176_, new_n47177_, new_n47178_,
    new_n47179_, new_n47180_, new_n47181_, new_n47182_, new_n47183_,
    new_n47184_, new_n47185_, new_n47186_, new_n47187_, new_n47188_,
    new_n47189_, new_n47190_, new_n47191_, new_n47192_, new_n47193_,
    new_n47194_, new_n47196_, new_n47197_, new_n47198_, new_n47199_,
    new_n47200_, new_n47201_, new_n47202_, new_n47203_, new_n47204_,
    new_n47205_, new_n47206_, new_n47207_, new_n47208_, new_n47209_,
    new_n47210_, new_n47211_, new_n47212_, new_n47213_, new_n47214_,
    new_n47215_, new_n47216_, new_n47217_, new_n47218_, new_n47219_,
    new_n47220_, new_n47221_, new_n47222_, new_n47223_, new_n47224_,
    new_n47225_, new_n47227_, new_n47228_, new_n47229_, new_n47230_,
    new_n47231_, new_n47232_, new_n47233_, new_n47234_, new_n47235_,
    new_n47236_, new_n47237_, new_n47238_, new_n47239_, new_n47240_,
    new_n47241_, new_n47242_, new_n47243_, new_n47244_, new_n47245_,
    new_n47246_, new_n47247_, new_n47248_, new_n47249_, new_n47250_,
    new_n47251_, new_n47252_, new_n47253_, new_n47254_, new_n47255_,
    new_n47256_, new_n47258_, new_n47259_, new_n47261_, new_n47262_,
    new_n47263_, new_n47264_, new_n47265_, new_n47267_, new_n47268_,
    new_n47269_, new_n47270_, new_n47271_, new_n47272_, new_n47273_,
    new_n47274_, new_n47276_, new_n47277_, new_n47278_, new_n47280_,
    new_n47281_, new_n47282_, new_n47284_, new_n47285_, new_n47286_,
    new_n47288_, new_n47289_, new_n47290_, new_n47292_, new_n47293_,
    new_n47294_, new_n47296_, new_n47297_, new_n47298_, new_n47300_,
    new_n47301_, new_n47302_, new_n47304_, new_n47305_, new_n47306_,
    new_n47308_, new_n47309_, new_n47310_, new_n47312_, new_n47313_,
    new_n47314_, new_n47316_, new_n47317_, new_n47318_, new_n47320_,
    new_n47321_, new_n47322_, new_n47324_, new_n47325_, new_n47326_,
    new_n47328_, new_n47329_, new_n47330_, new_n47332_, new_n47333_,
    new_n47334_, new_n47336_, new_n47337_, new_n47338_, new_n47340_,
    new_n47341_, new_n47342_, new_n47344_, new_n47345_, new_n47346_,
    new_n47348_, new_n47349_, new_n47350_, new_n47352_, new_n47353_,
    new_n47354_, new_n47356_, new_n47357_, new_n47358_, new_n47360_,
    new_n47361_, new_n47362_, new_n47364_, new_n47365_, new_n47366_,
    new_n47368_, new_n47369_, new_n47370_, new_n47372_, new_n47373_,
    new_n47374_, new_n47376_, new_n47377_, new_n47378_, new_n47380_,
    new_n47381_, new_n47382_, new_n47384_, new_n47385_, new_n47386_,
    new_n47388_, new_n47389_, new_n47390_, new_n47392_, new_n47393_,
    new_n47394_, new_n47396_, new_n47397_, new_n47398_, new_n47400_,
    new_n47401_, new_n47402_, new_n47404_, new_n47405_, new_n47406_,
    new_n47408_, new_n47409_, new_n47410_, new_n47411_, new_n47412_,
    new_n47413_, new_n47414_, new_n47415_, new_n47417_, new_n47418_,
    new_n47419_, new_n47421_, new_n47422_, new_n47423_, new_n47425_,
    new_n47426_, new_n47427_, new_n47429_, new_n47430_, new_n47431_,
    new_n47433_, new_n47434_, new_n47435_, new_n47437_, new_n47438_,
    new_n47439_, new_n47441_, new_n47442_, new_n47443_, new_n47445_,
    new_n47446_, new_n47447_, new_n47449_, new_n47450_, new_n47451_,
    new_n47453_, new_n47454_, new_n47455_, new_n47457_, new_n47458_,
    new_n47459_, new_n47461_, new_n47462_, new_n47463_, new_n47465_,
    new_n47466_, new_n47467_, new_n47469_, new_n47470_, new_n47471_,
    new_n47473_, new_n47474_, new_n47475_, new_n47477_, new_n47478_,
    new_n47479_, new_n47481_, new_n47482_, new_n47483_, new_n47485_,
    new_n47486_, new_n47487_, new_n47489_, new_n47490_, new_n47491_,
    new_n47493_, new_n47494_, new_n47495_, new_n47497_, new_n47498_,
    new_n47499_, new_n47501_, new_n47502_, new_n47503_, new_n47505_,
    new_n47506_, new_n47507_, new_n47509_, new_n47510_, new_n47511_,
    new_n47513_, new_n47514_, new_n47515_, new_n47517_, new_n47518_,
    new_n47519_, new_n47521_, new_n47522_, new_n47523_, new_n47525_,
    new_n47526_, new_n47527_, new_n47529_, new_n47530_, new_n47531_,
    new_n47533_, new_n47534_, new_n47535_, new_n47537_, new_n47538_,
    new_n47539_, new_n47541_, new_n47542_, new_n47543_, new_n47545_,
    new_n47546_, new_n47547_, new_n47549_, new_n47550_, new_n47551_,
    new_n47552_, new_n47553_, new_n47554_, new_n47555_, new_n47556_,
    new_n47558_, new_n47559_, new_n47560_, new_n47562_, new_n47563_,
    new_n47564_, new_n47566_, new_n47567_, new_n47568_, new_n47570_,
    new_n47571_, new_n47572_, new_n47574_, new_n47575_, new_n47576_,
    new_n47578_, new_n47579_, new_n47580_, new_n47582_, new_n47583_,
    new_n47584_, new_n47586_, new_n47587_, new_n47588_, new_n47590_,
    new_n47591_, new_n47592_, new_n47594_, new_n47595_, new_n47596_,
    new_n47598_, new_n47599_, new_n47600_, new_n47602_, new_n47603_,
    new_n47604_, new_n47606_, new_n47607_, new_n47608_, new_n47610_,
    new_n47611_, new_n47612_, new_n47614_, new_n47615_, new_n47616_,
    new_n47618_, new_n47619_, new_n47620_, new_n47622_, new_n47623_,
    new_n47624_, new_n47626_, new_n47627_, new_n47628_, new_n47630_,
    new_n47631_, new_n47632_, new_n47634_, new_n47635_, new_n47636_,
    new_n47638_, new_n47639_, new_n47640_, new_n47642_, new_n47643_,
    new_n47644_, new_n47646_, new_n47647_, new_n47648_, new_n47650_,
    new_n47651_, new_n47652_, new_n47654_, new_n47655_, new_n47656_,
    new_n47658_, new_n47659_, new_n47660_, new_n47662_, new_n47663_,
    new_n47664_, new_n47666_, new_n47667_, new_n47668_, new_n47670_,
    new_n47671_, new_n47672_, new_n47674_, new_n47675_, new_n47676_,
    new_n47678_, new_n47679_, new_n47680_, new_n47682_, new_n47683_,
    new_n47684_, new_n47686_, new_n47687_, new_n47688_, new_n47690_,
    new_n47691_, new_n47692_, new_n47693_, new_n47694_, new_n47695_,
    new_n47696_, new_n47697_, new_n47699_, new_n47700_, new_n47701_,
    new_n47703_, new_n47704_, new_n47705_, new_n47707_, new_n47708_,
    new_n47709_, new_n47711_, new_n47712_, new_n47713_, new_n47715_,
    new_n47716_, new_n47717_, new_n47719_, new_n47720_, new_n47721_,
    new_n47723_, new_n47724_, new_n47725_, new_n47727_, new_n47728_,
    new_n47729_, new_n47731_, new_n47732_, new_n47733_, new_n47735_,
    new_n47736_, new_n47737_, new_n47739_, new_n47740_, new_n47741_,
    new_n47743_, new_n47744_, new_n47745_, new_n47747_, new_n47748_,
    new_n47749_, new_n47751_, new_n47752_, new_n47753_, new_n47755_,
    new_n47756_, new_n47757_, new_n47759_, new_n47760_, new_n47761_,
    new_n47763_, new_n47764_, new_n47765_, new_n47767_, new_n47768_,
    new_n47769_, new_n47771_, new_n47772_, new_n47773_, new_n47775_,
    new_n47776_, new_n47777_, new_n47779_, new_n47780_, new_n47781_,
    new_n47783_, new_n47784_, new_n47785_, new_n47787_, new_n47788_,
    new_n47789_, new_n47791_, new_n47792_, new_n47793_, new_n47795_,
    new_n47796_, new_n47797_, new_n47799_, new_n47800_, new_n47801_,
    new_n47803_, new_n47804_, new_n47805_, new_n47807_, new_n47808_,
    new_n47809_, new_n47811_, new_n47812_, new_n47813_, new_n47815_,
    new_n47816_, new_n47817_, new_n47819_, new_n47820_, new_n47821_,
    new_n47823_, new_n47824_, new_n47825_, new_n47827_, new_n47828_,
    new_n47829_, new_n47831_, new_n47832_, new_n47833_, new_n47834_,
    new_n47835_, new_n47836_, new_n47837_, new_n47838_, new_n47840_,
    new_n47841_, new_n47842_, new_n47844_, new_n47845_, new_n47846_,
    new_n47848_, new_n47849_, new_n47850_, new_n47852_, new_n47853_,
    new_n47854_, new_n47856_, new_n47857_, new_n47858_, new_n47860_,
    new_n47861_, new_n47862_, new_n47864_, new_n47865_, new_n47866_,
    new_n47868_, new_n47869_, new_n47870_, new_n47872_, new_n47873_,
    new_n47874_, new_n47876_, new_n47877_, new_n47878_, new_n47880_,
    new_n47881_, new_n47882_, new_n47884_, new_n47885_, new_n47886_,
    new_n47888_, new_n47889_, new_n47890_, new_n47892_, new_n47893_,
    new_n47894_, new_n47896_, new_n47897_, new_n47898_, new_n47900_,
    new_n47901_, new_n47902_, new_n47904_, new_n47905_, new_n47906_,
    new_n47908_, new_n47909_, new_n47910_, new_n47912_, new_n47913_,
    new_n47914_, new_n47916_, new_n47917_, new_n47918_, new_n47920_,
    new_n47921_, new_n47922_, new_n47924_, new_n47925_, new_n47926_,
    new_n47928_, new_n47929_, new_n47930_, new_n47932_, new_n47933_,
    new_n47934_, new_n47936_, new_n47937_, new_n47938_, new_n47940_,
    new_n47941_, new_n47942_, new_n47944_, new_n47945_, new_n47946_,
    new_n47948_, new_n47949_, new_n47950_, new_n47952_, new_n47953_,
    new_n47954_, new_n47956_, new_n47957_, new_n47958_, new_n47960_,
    new_n47961_, new_n47962_, new_n47964_, new_n47965_, new_n47966_,
    new_n47968_, new_n47969_, new_n47970_, new_n47972_, new_n47973_,
    new_n47974_, new_n47975_, new_n47976_, new_n47977_, new_n47978_,
    new_n47979_, new_n47981_, new_n47982_, new_n47983_, new_n47985_,
    new_n47986_, new_n47987_, new_n47989_, new_n47990_, new_n47991_,
    new_n47993_, new_n47994_, new_n47995_, new_n47997_, new_n47998_,
    new_n47999_, new_n48001_, new_n48002_, new_n48003_, new_n48005_,
    new_n48006_, new_n48007_, new_n48009_, new_n48010_, new_n48011_,
    new_n48013_, new_n48014_, new_n48015_, new_n48017_, new_n48018_,
    new_n48019_, new_n48021_, new_n48022_, new_n48023_, new_n48025_,
    new_n48026_, new_n48027_, new_n48029_, new_n48030_, new_n48031_,
    new_n48033_, new_n48034_, new_n48035_, new_n48037_, new_n48038_,
    new_n48039_, new_n48041_, new_n48042_, new_n48043_, new_n48045_,
    new_n48046_, new_n48047_, new_n48049_, new_n48050_, new_n48051_,
    new_n48053_, new_n48054_, new_n48055_, new_n48057_, new_n48058_,
    new_n48059_, new_n48061_, new_n48062_, new_n48063_, new_n48065_,
    new_n48066_, new_n48067_, new_n48069_, new_n48070_, new_n48071_,
    new_n48073_, new_n48074_, new_n48075_, new_n48077_, new_n48078_,
    new_n48079_, new_n48081_, new_n48082_, new_n48083_, new_n48085_,
    new_n48086_, new_n48087_, new_n48089_, new_n48090_, new_n48091_,
    new_n48093_, new_n48094_, new_n48095_, new_n48097_, new_n48098_,
    new_n48099_, new_n48101_, new_n48102_, new_n48103_, new_n48105_,
    new_n48106_, new_n48107_, new_n48109_, new_n48110_, new_n48111_,
    new_n48113_, new_n48114_, new_n48115_, new_n48116_, new_n48117_,
    new_n48118_, new_n48119_, new_n48120_, new_n48122_, new_n48123_,
    new_n48124_, new_n48126_, new_n48127_, new_n48128_, new_n48130_,
    new_n48131_, new_n48132_, new_n48134_, new_n48135_, new_n48136_,
    new_n48138_, new_n48139_, new_n48140_, new_n48142_, new_n48143_,
    new_n48144_, new_n48146_, new_n48147_, new_n48148_, new_n48150_,
    new_n48151_, new_n48152_, new_n48154_, new_n48155_, new_n48156_,
    new_n48158_, new_n48159_, new_n48160_, new_n48162_, new_n48163_,
    new_n48164_, new_n48166_, new_n48167_, new_n48168_, new_n48170_,
    new_n48171_, new_n48172_, new_n48174_, new_n48175_, new_n48176_,
    new_n48178_, new_n48179_, new_n48180_, new_n48182_, new_n48183_,
    new_n48184_, new_n48186_, new_n48187_, new_n48188_, new_n48190_,
    new_n48191_, new_n48192_, new_n48194_, new_n48195_, new_n48196_,
    new_n48198_, new_n48199_, new_n48200_, new_n48202_, new_n48203_,
    new_n48204_, new_n48206_, new_n48207_, new_n48208_, new_n48210_,
    new_n48211_, new_n48212_, new_n48214_, new_n48215_, new_n48216_,
    new_n48218_, new_n48219_, new_n48220_, new_n48222_, new_n48223_,
    new_n48224_, new_n48226_, new_n48227_, new_n48228_, new_n48230_,
    new_n48231_, new_n48232_, new_n48234_, new_n48235_, new_n48236_,
    new_n48238_, new_n48239_, new_n48240_, new_n48242_, new_n48243_,
    new_n48244_, new_n48246_, new_n48247_, new_n48248_, new_n48250_,
    new_n48251_, new_n48252_, new_n48254_, new_n48255_, new_n48256_,
    new_n48257_, new_n48258_, new_n48259_, new_n48260_, new_n48261_,
    new_n48263_, new_n48264_, new_n48265_, new_n48267_, new_n48268_,
    new_n48269_, new_n48271_, new_n48272_, new_n48273_, new_n48275_,
    new_n48276_, new_n48277_, new_n48279_, new_n48280_, new_n48281_,
    new_n48283_, new_n48284_, new_n48285_, new_n48287_, new_n48288_,
    new_n48289_, new_n48291_, new_n48292_, new_n48293_, new_n48295_,
    new_n48296_, new_n48297_, new_n48299_, new_n48300_, new_n48301_,
    new_n48303_, new_n48304_, new_n48305_, new_n48307_, new_n48308_,
    new_n48309_, new_n48311_, new_n48312_, new_n48313_, new_n48315_,
    new_n48316_, new_n48317_, new_n48319_, new_n48320_, new_n48321_,
    new_n48323_, new_n48324_, new_n48325_, new_n48327_, new_n48328_,
    new_n48329_, new_n48331_, new_n48332_, new_n48333_, new_n48335_,
    new_n48336_, new_n48337_, new_n48339_, new_n48340_, new_n48341_,
    new_n48343_, new_n48344_, new_n48345_, new_n48347_, new_n48348_,
    new_n48349_, new_n48351_, new_n48352_, new_n48353_, new_n48355_,
    new_n48356_, new_n48357_, new_n48359_, new_n48360_, new_n48361_,
    new_n48363_, new_n48364_, new_n48365_, new_n48367_, new_n48368_,
    new_n48369_, new_n48371_, new_n48372_, new_n48373_, new_n48375_,
    new_n48376_, new_n48377_, new_n48379_, new_n48380_, new_n48381_,
    new_n48383_, new_n48384_, new_n48385_, new_n48387_, new_n48388_,
    new_n48389_, new_n48390_, new_n48391_, new_n48392_, new_n48393_,
    new_n48394_, new_n48396_, new_n48397_, new_n48398_, new_n48400_,
    new_n48401_, new_n48402_, new_n48404_, new_n48405_, new_n48406_,
    new_n48408_, new_n48409_, new_n48410_, new_n48412_, new_n48413_,
    new_n48414_, new_n48416_, new_n48417_, new_n48418_, new_n48420_,
    new_n48421_, new_n48422_, new_n48424_, new_n48425_, new_n48426_,
    new_n48428_, new_n48429_, new_n48430_, new_n48432_, new_n48433_,
    new_n48434_, new_n48436_, new_n48437_, new_n48438_, new_n48440_,
    new_n48441_, new_n48442_, new_n48444_, new_n48445_, new_n48446_,
    new_n48448_, new_n48449_, new_n48450_, new_n48452_, new_n48453_,
    new_n48454_, new_n48456_, new_n48457_, new_n48458_, new_n48460_,
    new_n48461_, new_n48462_, new_n48464_, new_n48465_, new_n48466_,
    new_n48468_, new_n48469_, new_n48470_, new_n48472_, new_n48473_,
    new_n48474_, new_n48476_, new_n48477_, new_n48478_, new_n48480_,
    new_n48481_, new_n48482_, new_n48484_, new_n48485_, new_n48486_,
    new_n48488_, new_n48489_, new_n48490_, new_n48492_, new_n48493_,
    new_n48494_, new_n48496_, new_n48497_, new_n48498_, new_n48500_,
    new_n48501_, new_n48502_, new_n48504_, new_n48505_, new_n48506_,
    new_n48508_, new_n48509_, new_n48510_, new_n48512_, new_n48513_,
    new_n48514_, new_n48516_, new_n48517_, new_n48518_, new_n48520_,
    new_n48521_, new_n48522_, new_n48523_, new_n48524_, new_n48525_,
    new_n48526_, new_n48527_, new_n48529_, new_n48530_, new_n48531_,
    new_n48533_, new_n48534_, new_n48535_, new_n48537_, new_n48538_,
    new_n48539_, new_n48541_, new_n48542_, new_n48543_, new_n48545_,
    new_n48546_, new_n48547_, new_n48549_, new_n48550_, new_n48551_,
    new_n48553_, new_n48554_, new_n48555_, new_n48557_, new_n48558_,
    new_n48559_, new_n48561_, new_n48562_, new_n48563_, new_n48565_,
    new_n48566_, new_n48567_, new_n48569_, new_n48570_, new_n48571_,
    new_n48573_, new_n48574_, new_n48575_, new_n48577_, new_n48578_,
    new_n48579_, new_n48581_, new_n48582_, new_n48583_, new_n48585_,
    new_n48586_, new_n48587_, new_n48589_, new_n48590_, new_n48591_,
    new_n48593_, new_n48594_, new_n48595_, new_n48597_, new_n48598_,
    new_n48599_, new_n48601_, new_n48602_, new_n48603_, new_n48605_,
    new_n48606_, new_n48607_, new_n48609_, new_n48610_, new_n48611_,
    new_n48613_, new_n48614_, new_n48615_, new_n48617_, new_n48618_,
    new_n48619_, new_n48621_, new_n48622_, new_n48623_, new_n48625_,
    new_n48626_, new_n48627_, new_n48629_, new_n48630_, new_n48631_,
    new_n48633_, new_n48634_, new_n48635_, new_n48637_, new_n48638_,
    new_n48639_, new_n48641_, new_n48642_, new_n48643_, new_n48645_,
    new_n48646_, new_n48647_, new_n48649_, new_n48650_, new_n48651_,
    new_n48653_, new_n48654_, new_n48655_, new_n48657_, new_n48658_,
    new_n48659_, new_n48661_, new_n48662_, new_n48663_, new_n48665_,
    new_n48666_, new_n48667_, new_n48669_, new_n48670_, new_n48671_,
    new_n48673_, new_n48674_, new_n48675_, new_n48677_, new_n48678_,
    new_n48679_, new_n48681_, new_n48682_, new_n48683_, new_n48685_,
    new_n48686_, new_n48687_, new_n48689_, new_n48690_, new_n48691_,
    new_n48693_, new_n48694_, new_n48695_, new_n48697_, new_n48698_,
    new_n48699_, new_n48701_, new_n48702_, new_n48703_, new_n48705_,
    new_n48706_, new_n48707_, new_n48709_, new_n48710_, new_n48711_,
    new_n48713_, new_n48714_, new_n48715_, new_n48717_, new_n48718_,
    new_n48719_, new_n48721_, new_n48722_, new_n48723_, new_n48725_,
    new_n48726_, new_n48727_, new_n48729_, new_n48730_, new_n48731_,
    new_n48733_, new_n48734_, new_n48735_, new_n48737_, new_n48738_,
    new_n48739_, new_n48741_, new_n48742_, new_n48743_, new_n48745_,
    new_n48746_, new_n48747_, new_n48749_, new_n48750_, new_n48751_,
    new_n48753_, new_n48754_, new_n48755_, new_n48757_, new_n48758_,
    new_n48759_, new_n48761_, new_n48762_, new_n48763_, new_n48765_,
    new_n48766_, new_n48767_, new_n48769_, new_n48770_, new_n48771_,
    new_n48773_, new_n48774_, new_n48775_, new_n48777_, new_n48778_,
    new_n48779_, new_n48781_, new_n48782_, new_n48783_, new_n48785_,
    new_n48786_, new_n48787_, new_n48789_, new_n48790_, new_n48791_,
    new_n48793_, new_n48794_, new_n48795_, new_n48797_, new_n48798_,
    new_n48799_, new_n48801_, new_n48802_, new_n48803_, new_n48805_,
    new_n48806_, new_n48807_, new_n48809_, new_n48810_, new_n48811_,
    new_n48813_, new_n48814_, new_n48815_, new_n48817_, new_n48818_,
    new_n48819_, new_n48821_, new_n48822_, new_n48823_, new_n48825_,
    new_n48826_, new_n48827_, new_n48829_, new_n48830_, new_n48831_,
    new_n48833_, new_n48834_, new_n48835_, new_n48837_, new_n48838_,
    new_n48839_, new_n48841_, new_n48842_, new_n48843_, new_n48845_,
    new_n48846_, new_n48847_, new_n48849_, new_n48850_, new_n48851_,
    new_n48853_, new_n48854_, new_n48855_, new_n48857_, new_n48858_,
    new_n48859_, new_n48861_, new_n48862_, new_n48863_, new_n48865_,
    new_n48866_, new_n48867_, new_n48869_, new_n48870_, new_n48871_,
    new_n48873_, new_n48874_, new_n48875_, new_n48877_, new_n48878_,
    new_n48879_, new_n48881_, new_n48882_, new_n48883_, new_n48885_,
    new_n48886_, new_n48887_, new_n48889_, new_n48890_, new_n48891_,
    new_n48893_, new_n48894_, new_n48895_, new_n48897_, new_n48898_,
    new_n48899_, new_n48901_, new_n48902_, new_n48903_, new_n48905_,
    new_n48906_, new_n48907_, new_n48909_, new_n48910_, new_n48911_,
    new_n48913_, new_n48914_, new_n48915_, new_n48917_, new_n48918_,
    new_n48919_, new_n48921_, new_n48922_, new_n48923_, new_n48925_,
    new_n48926_, new_n48927_, new_n48929_, new_n48930_, new_n48931_,
    new_n48933_, new_n48934_, new_n48935_, new_n48937_, new_n48938_,
    new_n48939_, new_n48941_, new_n48942_, new_n48943_, new_n48945_,
    new_n48946_, new_n48947_, new_n48949_, new_n48950_, new_n48951_,
    new_n48953_, new_n48954_, new_n48955_, new_n48957_, new_n48958_,
    new_n48959_, new_n48961_, new_n48962_, new_n48963_, new_n48965_,
    new_n48966_, new_n48967_, new_n48969_, new_n48970_, new_n48971_,
    new_n48973_, new_n48974_, new_n48975_, new_n48977_, new_n48978_,
    new_n48979_, new_n48981_, new_n48982_, new_n48983_, new_n48985_,
    new_n48986_, new_n48987_, new_n48989_, new_n48990_, new_n48991_,
    new_n48993_, new_n48994_, new_n48995_, new_n48997_, new_n48998_,
    new_n48999_, new_n49001_, new_n49002_, new_n49003_, new_n49005_,
    new_n49006_, new_n49007_, new_n49009_, new_n49010_, new_n49011_,
    new_n49013_, new_n49014_, new_n49015_, new_n49017_, new_n49018_,
    new_n49019_, new_n49021_, new_n49022_, new_n49023_, new_n49025_,
    new_n49026_, new_n49027_, new_n49029_, new_n49030_, new_n49031_,
    new_n49033_, new_n49034_, new_n49035_, new_n49037_, new_n49038_,
    new_n49039_, new_n49041_, new_n49042_, new_n49043_, new_n49045_,
    new_n49046_, new_n49047_, new_n49049_, new_n49050_, new_n49051_,
    new_n49053_, new_n49054_, new_n49055_, new_n49057_, new_n49058_,
    new_n49059_, new_n49061_, new_n49062_, new_n49063_, new_n49065_,
    new_n49066_, new_n49067_, new_n49069_, new_n49070_, new_n49071_,
    new_n49073_, new_n49074_, new_n49075_, new_n49077_, new_n49078_,
    new_n49079_, new_n49081_, new_n49082_, new_n49083_, new_n49085_,
    new_n49086_, new_n49087_, new_n49089_, new_n49090_, new_n49091_,
    new_n49093_, new_n49094_, new_n49095_, new_n49097_, new_n49098_,
    new_n49099_, new_n49101_, new_n49102_, new_n49103_, new_n49105_,
    new_n49106_, new_n49107_, new_n49109_, new_n49110_, new_n49111_,
    new_n49113_, new_n49114_, new_n49115_, new_n49117_, new_n49118_,
    new_n49119_, new_n49121_, new_n49122_, new_n49123_, new_n49125_,
    new_n49126_, new_n49127_, new_n49129_, new_n49130_, new_n49131_,
    new_n49133_, new_n49134_, new_n49135_, new_n49137_, new_n49138_,
    new_n49139_, new_n49141_, new_n49142_, new_n49143_, new_n49145_,
    new_n49146_, new_n49147_, new_n49149_, new_n49150_, new_n49151_,
    new_n49153_, new_n49154_, new_n49155_, new_n49157_, new_n49158_,
    new_n49159_, new_n49161_, new_n49162_, new_n49163_, new_n49165_,
    new_n49166_, new_n49167_, new_n49169_, new_n49170_, new_n49171_,
    new_n49173_, new_n49174_, new_n49175_, new_n49177_, new_n49178_,
    new_n49179_, new_n49181_, new_n49182_, new_n49183_, new_n49185_,
    new_n49186_, new_n49187_, new_n49189_, new_n49190_, new_n49191_,
    new_n49193_, new_n49194_, new_n49195_, new_n49197_, new_n49198_,
    new_n49199_, new_n49201_, new_n49202_, new_n49203_, new_n49205_,
    new_n49206_, new_n49207_, new_n49209_, new_n49210_, new_n49211_,
    new_n49213_, new_n49214_, new_n49215_, new_n49217_, new_n49218_,
    new_n49219_, new_n49221_, new_n49222_, new_n49223_, new_n49225_,
    new_n49226_, new_n49227_, new_n49229_, new_n49230_, new_n49231_,
    new_n49233_, new_n49234_, new_n49235_, new_n49237_, new_n49238_,
    new_n49239_, new_n49241_, new_n49242_, new_n49243_, new_n49245_,
    new_n49246_, new_n49247_, new_n49249_, new_n49250_, new_n49251_,
    new_n49253_, new_n49254_, new_n49255_, new_n49257_, new_n49258_,
    new_n49259_, new_n49261_, new_n49262_, new_n49263_, new_n49265_,
    new_n49266_, new_n49267_, new_n49269_, new_n49270_, new_n49271_,
    new_n49273_, new_n49274_, new_n49275_, new_n49277_, new_n49278_,
    new_n49279_, new_n49281_, new_n49282_, new_n49283_, new_n49285_,
    new_n49286_, new_n49287_, new_n49289_, new_n49290_, new_n49291_,
    new_n49293_, new_n49294_, new_n49295_, new_n49297_, new_n49298_,
    new_n49299_, new_n49301_, new_n49302_, new_n49303_, new_n49305_,
    new_n49306_, new_n49307_, new_n49309_, new_n49310_, new_n49311_,
    new_n49313_, new_n49314_, new_n49315_, new_n49317_, new_n49318_,
    new_n49319_, new_n49321_, new_n49322_, new_n49323_, new_n49325_,
    new_n49326_, new_n49327_, new_n49329_, new_n49330_, new_n49331_,
    new_n49333_, new_n49334_, new_n49335_, new_n49337_, new_n49338_,
    new_n49339_, new_n49341_, new_n49342_, new_n49343_, new_n49345_,
    new_n49346_, new_n49347_, new_n49349_, new_n49350_, new_n49351_,
    new_n49353_, new_n49354_, new_n49355_, new_n49357_, new_n49358_,
    new_n49359_, new_n49361_, new_n49362_, new_n49363_, new_n49365_,
    new_n49366_, new_n49367_, new_n49369_, new_n49370_, new_n49371_,
    new_n49373_, new_n49374_, new_n49375_, new_n49377_, new_n49378_,
    new_n49379_, new_n49381_, new_n49382_, new_n49383_, new_n49385_,
    new_n49386_, new_n49387_, new_n49389_, new_n49390_, new_n49391_,
    new_n49393_, new_n49394_, new_n49395_, new_n49397_, new_n49398_,
    new_n49399_, new_n49401_, new_n49402_, new_n49403_, new_n49405_,
    new_n49406_, new_n49407_, new_n49409_, new_n49410_, new_n49411_,
    new_n49413_, new_n49414_, new_n49415_, new_n49417_, new_n49418_,
    new_n49419_, new_n49421_, new_n49422_, new_n49423_, new_n49425_,
    new_n49426_, new_n49427_, new_n49429_, new_n49430_, new_n49431_,
    new_n49433_, new_n49434_, new_n49435_, new_n49437_, new_n49438_,
    new_n49439_, new_n49441_, new_n49442_, new_n49443_, new_n49445_,
    new_n49446_, new_n49447_, new_n49449_, new_n49450_, new_n49451_,
    new_n49453_, new_n49454_, new_n49455_, new_n49457_, new_n49458_,
    new_n49459_, new_n49461_, new_n49462_, new_n49463_, new_n49465_,
    new_n49466_, new_n49467_, new_n49469_, new_n49470_, new_n49471_,
    new_n49473_, new_n49474_, new_n49475_, new_n49477_, new_n49478_,
    new_n49479_, new_n49481_, new_n49482_, new_n49483_, new_n49485_,
    new_n49486_, new_n49487_, new_n49489_, new_n49490_, new_n49491_,
    new_n49493_, new_n49494_, new_n49495_, new_n49497_, new_n49498_,
    new_n49499_, new_n49501_, new_n49502_, new_n49503_, new_n49505_,
    new_n49506_, new_n49507_, new_n49509_, new_n49510_, new_n49511_,
    new_n49513_, new_n49514_, new_n49515_, new_n49517_, new_n49518_,
    new_n49519_, new_n49521_, new_n49522_, new_n49523_, new_n49525_,
    new_n49526_, new_n49527_, new_n49529_, new_n49530_, new_n49531_,
    new_n49533_, new_n49534_, new_n49535_, new_n49537_, new_n49538_,
    new_n49539_, new_n49541_, new_n49542_, new_n49543_, new_n49545_,
    new_n49546_, new_n49547_, new_n49549_, new_n49550_, new_n49551_,
    new_n49553_, new_n49554_, new_n49555_, new_n49557_, new_n49558_,
    new_n49559_, new_n49561_, new_n49562_, new_n49563_, new_n49565_,
    new_n49566_, new_n49567_, new_n49569_, new_n49570_, new_n49571_,
    new_n49573_, new_n49574_, new_n49575_, new_n49577_, new_n49578_,
    new_n49579_, new_n49581_, new_n49582_, new_n49583_, new_n49585_,
    new_n49586_, new_n49587_, new_n49589_, new_n49590_, new_n49591_,
    new_n49593_, new_n49594_, new_n49595_, new_n49597_, new_n49598_,
    new_n49599_, new_n49601_, new_n49602_, new_n49603_, new_n49605_,
    new_n49606_, new_n49607_, new_n49609_, new_n49610_, new_n49611_,
    new_n49613_, new_n49614_, new_n49615_, new_n49617_, new_n49618_,
    new_n49619_, new_n49621_, new_n49622_, new_n49623_, new_n49625_,
    new_n49626_, new_n49627_, new_n49629_, new_n49630_, new_n49631_,
    new_n49633_, new_n49634_, new_n49635_, new_n49637_, new_n49638_,
    new_n49639_, new_n49641_, new_n49642_, new_n49643_, new_n49645_,
    new_n49646_, new_n49647_, new_n49649_, new_n49650_, new_n49651_,
    new_n49653_, new_n49654_, new_n49655_, new_n49657_, new_n49658_,
    new_n49659_, new_n49661_, new_n49662_, new_n49663_, new_n49665_,
    new_n49666_, new_n49667_, new_n49669_, new_n49670_, new_n49671_,
    new_n49673_, new_n49674_, new_n49675_, new_n49677_, new_n49678_,
    new_n49679_, new_n49681_, new_n49682_, new_n49683_, new_n49685_,
    new_n49686_, new_n49687_, new_n49689_, new_n49690_, new_n49691_,
    new_n49693_, new_n49694_, new_n49695_, new_n49697_, new_n49698_,
    new_n49699_, new_n49701_, new_n49702_, new_n49703_, new_n49705_,
    new_n49706_, new_n49707_, new_n49709_, new_n49710_, new_n49711_,
    new_n49713_, new_n49714_, new_n49715_, new_n49717_, new_n49718_,
    new_n49719_, new_n49721_, new_n49722_, new_n49723_, new_n49725_,
    new_n49726_, new_n49727_, new_n49729_, new_n49730_, new_n49731_,
    new_n49733_, new_n49734_, new_n49735_, new_n49737_, new_n49738_,
    new_n49739_, new_n49741_, new_n49742_, new_n49743_, new_n49745_,
    new_n49746_, new_n49747_, new_n49749_, new_n49750_, new_n49751_,
    new_n49753_, new_n49754_, new_n49755_, new_n49757_, new_n49758_,
    new_n49759_, new_n49761_, new_n49762_, new_n49763_, new_n49765_,
    new_n49766_, new_n49767_, new_n49769_, new_n49770_, new_n49771_,
    new_n49773_, new_n49774_, new_n49775_, new_n49777_, new_n49778_,
    new_n49779_, new_n49781_, new_n49782_, new_n49783_, new_n49785_,
    new_n49786_, new_n49787_, new_n49789_, new_n49790_, new_n49791_,
    new_n49793_, new_n49794_, new_n49795_, new_n49797_, new_n49798_,
    new_n49799_, new_n49801_, new_n49802_, new_n49803_, new_n49805_,
    new_n49806_, new_n49807_, new_n49809_, new_n49810_, new_n49811_,
    new_n49813_, new_n49814_, new_n49815_, new_n49817_, new_n49818_,
    new_n49819_, new_n49821_, new_n49822_, new_n49823_, new_n49825_,
    new_n49826_, new_n49827_, new_n49829_, new_n49830_, new_n49831_,
    new_n49833_, new_n49834_, new_n49835_, new_n49837_, new_n49838_,
    new_n49839_, new_n49841_, new_n49842_, new_n49843_, new_n49845_,
    new_n49846_, new_n49847_, new_n49849_, new_n49850_, new_n49851_,
    new_n49853_, new_n49854_, new_n49855_, new_n49857_, new_n49858_,
    new_n49859_, new_n49861_, new_n49862_, new_n49863_, new_n49865_,
    new_n49866_, new_n49867_, new_n49869_, new_n49870_, new_n49871_,
    new_n49873_, new_n49874_, new_n49875_, new_n49877_, new_n49878_,
    new_n49879_, new_n49881_, new_n49882_, new_n49883_, new_n49885_,
    new_n49886_, new_n49887_, new_n49889_, new_n49890_, new_n49891_,
    new_n49893_, new_n49894_, new_n49895_, new_n49897_, new_n49898_,
    new_n49899_, new_n49901_, new_n49902_, new_n49903_, new_n49905_,
    new_n49906_, new_n49907_, new_n49909_, new_n49910_, new_n49911_,
    new_n49913_, new_n49914_, new_n49915_, new_n49917_, new_n49918_,
    new_n49919_, new_n49921_, new_n49922_, new_n49923_, new_n49925_,
    new_n49926_, new_n49927_, new_n49929_, new_n49930_, new_n49931_,
    new_n49933_, new_n49934_, new_n49935_, new_n49937_, new_n49938_,
    new_n49939_, new_n49941_, new_n49942_, new_n49943_, new_n49945_,
    new_n49946_, new_n49947_, new_n49949_, new_n49950_, new_n49951_,
    new_n49953_, new_n49954_, new_n49955_, new_n49957_, new_n49958_,
    new_n49959_, new_n49961_, new_n49962_, new_n49963_, new_n49965_,
    new_n49966_, new_n49967_, new_n49969_, new_n49970_, new_n49971_,
    new_n49973_, new_n49974_, new_n49975_, new_n49977_, new_n49978_,
    new_n49979_, new_n49981_, new_n49982_, new_n49983_, new_n49985_,
    new_n49986_, new_n49987_, new_n49989_, new_n49990_, new_n49991_,
    new_n49993_, new_n49994_, new_n49995_, new_n49997_, new_n49998_,
    new_n49999_, new_n50001_, new_n50002_, new_n50003_, new_n50005_,
    new_n50006_, new_n50007_, new_n50009_, new_n50010_, new_n50011_,
    new_n50013_, new_n50014_, new_n50015_, new_n50017_, new_n50018_,
    new_n50019_, new_n50021_, new_n50022_, new_n50023_, new_n50025_,
    new_n50026_, new_n50027_, new_n50029_, new_n50030_, new_n50031_,
    new_n50033_, new_n50034_, new_n50035_, new_n50037_, new_n50038_,
    new_n50039_, new_n50041_, new_n50042_, new_n50043_, new_n50045_,
    new_n50046_, new_n50047_, new_n50049_, new_n50050_, new_n50051_,
    new_n50053_, new_n50054_, new_n50055_, new_n50057_, new_n50058_,
    new_n50059_, new_n50061_, new_n50062_, new_n50063_, new_n50065_,
    new_n50066_, new_n50067_, new_n50069_, new_n50070_, new_n50071_,
    new_n50073_, new_n50074_, new_n50075_, new_n50077_, new_n50078_,
    new_n50079_, new_n50081_, new_n50082_, new_n50083_, new_n50085_,
    new_n50086_, new_n50087_, new_n50089_, new_n50090_, new_n50091_,
    new_n50093_, new_n50094_, new_n50095_, new_n50097_, new_n50098_,
    new_n50099_, new_n50101_, new_n50102_, new_n50103_, new_n50105_,
    new_n50106_, new_n50107_, new_n50109_, new_n50110_, new_n50111_,
    new_n50113_, new_n50114_, new_n50115_, new_n50117_, new_n50118_,
    new_n50119_, new_n50121_, new_n50122_, new_n50123_, new_n50125_,
    new_n50126_, new_n50127_, new_n50129_, new_n50130_, new_n50131_,
    new_n50133_, new_n50134_, new_n50135_, new_n50137_, new_n50138_,
    new_n50139_, new_n50141_, new_n50142_, new_n50143_, new_n50145_,
    new_n50146_, new_n50147_, new_n50149_, new_n50150_, new_n50151_,
    new_n50153_, new_n50154_, new_n50155_, new_n50157_, new_n50158_,
    new_n50159_, new_n50161_, new_n50162_, new_n50163_, new_n50165_,
    new_n50166_, new_n50167_, new_n50169_, new_n50170_, new_n50171_,
    new_n50173_, new_n50174_, new_n50175_, new_n50177_, new_n50178_,
    new_n50179_, new_n50181_, new_n50182_, new_n50183_, new_n50185_,
    new_n50186_, new_n50187_, new_n50189_, new_n50190_, new_n50191_,
    new_n50193_, new_n50194_, new_n50195_, new_n50197_, new_n50198_,
    new_n50199_, new_n50201_, new_n50202_, new_n50203_, new_n50205_,
    new_n50206_, new_n50207_, new_n50209_, new_n50210_, new_n50211_,
    new_n50213_, new_n50214_, new_n50215_, new_n50217_, new_n50218_,
    new_n50219_, new_n50221_, new_n50222_, new_n50223_, new_n50225_,
    new_n50226_, new_n50227_, new_n50229_, new_n50230_, new_n50231_,
    new_n50233_, new_n50234_, new_n50235_, new_n50237_, new_n50238_,
    new_n50239_, new_n50241_, new_n50242_, new_n50243_, new_n50245_,
    new_n50246_, new_n50247_, new_n50249_, new_n50250_, new_n50251_,
    new_n50253_, new_n50254_, new_n50255_, new_n50257_, new_n50258_,
    new_n50259_, new_n50261_, new_n50262_, new_n50263_, new_n50265_,
    new_n50266_, new_n50267_, new_n50269_, new_n50270_, new_n50271_,
    new_n50273_, new_n50274_, new_n50275_, new_n50277_, new_n50278_,
    new_n50279_, new_n50281_, new_n50282_, new_n50283_, new_n50285_,
    new_n50286_, new_n50287_, new_n50289_, new_n50290_, new_n50291_,
    new_n50293_, new_n50294_, new_n50295_, new_n50297_, new_n50298_,
    new_n50299_, new_n50301_, new_n50302_, new_n50303_, new_n50305_,
    new_n50306_, new_n50307_, new_n50309_, new_n50310_, new_n50311_,
    new_n50313_, new_n50314_, new_n50315_, new_n50317_, new_n50318_,
    new_n50319_, new_n50321_, new_n50322_, new_n50323_, new_n50325_,
    new_n50326_, new_n50327_, new_n50329_, new_n50330_, new_n50331_,
    new_n50333_, new_n50334_, new_n50335_, new_n50337_, new_n50338_,
    new_n50339_, new_n50341_, new_n50342_, new_n50343_, new_n50345_,
    new_n50346_, new_n50347_, new_n50349_, new_n50350_, new_n50351_,
    new_n50353_, new_n50354_, new_n50355_, new_n50357_, new_n50358_,
    new_n50359_, new_n50361_, new_n50362_, new_n50363_, new_n50365_,
    new_n50366_, new_n50367_, new_n50369_, new_n50370_, new_n50371_,
    new_n50373_, new_n50374_, new_n50375_, new_n50377_, new_n50378_,
    new_n50379_, new_n50381_, new_n50382_, new_n50383_, new_n50385_,
    new_n50386_, new_n50387_, new_n50389_, new_n50390_, new_n50391_,
    new_n50393_, new_n50394_, new_n50395_, new_n50397_, new_n50398_,
    new_n50399_, new_n50401_, new_n50402_, new_n50403_, new_n50405_,
    new_n50406_, new_n50407_, new_n50409_, new_n50410_, new_n50411_,
    new_n50413_, new_n50414_, new_n50415_, new_n50417_, new_n50418_,
    new_n50419_, new_n50421_, new_n50422_, new_n50423_, new_n50425_,
    new_n50426_, new_n50427_, new_n50429_, new_n50430_, new_n50431_,
    new_n50433_, new_n50434_, new_n50435_, new_n50437_, new_n50438_,
    new_n50439_, new_n50441_, new_n50442_, new_n50443_, new_n50445_,
    new_n50446_, new_n50447_, new_n50449_, new_n50450_, new_n50451_,
    new_n50453_, new_n50454_, new_n50455_, new_n50457_, new_n50458_,
    new_n50459_, new_n50461_, new_n50462_, new_n50463_, new_n50465_,
    new_n50466_, new_n50467_, new_n50469_, new_n50470_, new_n50471_,
    new_n50473_, new_n50474_, new_n50475_, new_n50477_, new_n50478_,
    new_n50479_, new_n50481_, new_n50482_, new_n50483_, new_n50485_,
    new_n50486_, new_n50487_, new_n50489_, new_n50490_, new_n50491_,
    new_n50493_, new_n50494_, new_n50495_, new_n50497_, new_n50498_,
    new_n50499_, new_n50501_, new_n50502_, new_n50503_, new_n50505_,
    new_n50506_, new_n50507_, new_n50509_, new_n50510_, new_n50511_,
    new_n50513_, new_n50514_, new_n50515_, new_n50517_, new_n50518_,
    new_n50519_, new_n50521_, new_n50522_, new_n50523_, new_n50525_,
    new_n50526_, new_n50527_, new_n50529_, new_n50530_, new_n50531_,
    new_n50533_, new_n50534_, new_n50535_, new_n50537_, new_n50538_,
    new_n50539_, new_n50541_, new_n50542_, new_n50543_, new_n50545_,
    new_n50546_, new_n50547_, new_n50549_, new_n50550_, new_n50551_,
    new_n50553_, new_n50554_, new_n50555_, new_n50557_, new_n50558_,
    new_n50559_, new_n50561_, new_n50562_, new_n50563_, new_n50565_,
    new_n50566_, new_n50567_, new_n50569_, new_n50570_, new_n50571_,
    new_n50573_, new_n50574_, new_n50575_, new_n50577_, new_n50578_,
    new_n50579_, new_n50581_, new_n50582_, new_n50583_, new_n50585_,
    new_n50586_, new_n50587_, new_n50589_, new_n50590_, new_n50591_,
    new_n50593_, new_n50594_, new_n50595_, new_n50597_, new_n50598_,
    new_n50599_, new_n50601_, new_n50602_, new_n50603_, new_n50605_,
    new_n50606_, new_n50607_, new_n50609_, new_n50610_, new_n50611_,
    new_n50613_, new_n50614_, new_n50615_, new_n50617_, new_n50618_,
    new_n50619_, new_n50621_, new_n50622_, new_n50623_, new_n50625_,
    new_n50626_, new_n50627_, new_n50629_, new_n50630_, new_n50631_,
    new_n50633_, new_n50634_, new_n50635_, new_n50637_, new_n50638_,
    new_n50639_, new_n50641_, new_n50642_, new_n50643_, new_n50645_,
    new_n50646_, new_n50647_, new_n50649_, new_n50650_, new_n50651_,
    new_n50653_, new_n50654_, new_n50655_, new_n50657_, new_n50658_,
    new_n50659_, new_n50661_, new_n50662_, new_n50663_, new_n50665_,
    new_n50666_, new_n50667_, new_n50670_, new_n50671_, new_n50672_,
    new_n50673_, new_n50674_, new_n50675_, new_n50676_, new_n50677_,
    new_n50678_, new_n50679_, new_n50680_, new_n50681_, new_n50682_,
    new_n50683_, new_n50684_, new_n50685_, new_n50686_, new_n50688_,
    new_n50689_, new_n50690_, new_n50691_, new_n50692_, new_n50693_,
    new_n50694_, new_n50695_, new_n50696_, new_n50697_, new_n50698_,
    new_n50699_, new_n50701_, new_n50702_, new_n50703_, new_n50704_,
    new_n50705_, new_n50706_, new_n50707_, new_n50708_, new_n50709_,
    new_n50710_, new_n50711_, new_n50712_, new_n50714_, new_n50715_,
    new_n50716_, new_n50717_, new_n50718_, new_n50719_, new_n50720_,
    new_n50721_, new_n50722_, new_n50723_, new_n50724_, new_n50725_,
    new_n50727_, new_n50728_, new_n50729_, new_n50730_, new_n50731_,
    new_n50732_, new_n50733_, new_n50734_, new_n50735_, new_n50736_,
    new_n50737_, new_n50738_, new_n50740_, new_n50741_, new_n50742_,
    new_n50743_, new_n50744_, new_n50745_, new_n50746_, new_n50747_,
    new_n50748_, new_n50749_, new_n50750_, new_n50751_, new_n50753_,
    new_n50754_, new_n50755_, new_n50756_, new_n50757_, new_n50758_,
    new_n50759_, new_n50760_, new_n50761_, new_n50762_, new_n50763_,
    new_n50764_, new_n50766_, new_n50767_, new_n50768_, new_n50769_,
    new_n50770_, new_n50771_, new_n50772_, new_n50773_, new_n50774_,
    new_n50775_, new_n50776_, new_n50777_, new_n50779_, new_n50780_,
    new_n50781_, new_n50782_, new_n50783_, new_n50784_, new_n50785_,
    new_n50786_, new_n50787_, new_n50788_, new_n50789_, new_n50790_,
    new_n50792_, new_n50793_, new_n50794_, new_n50795_, new_n50796_,
    new_n50797_, new_n50798_, new_n50799_, new_n50800_, new_n50801_,
    new_n50802_, new_n50803_, new_n50805_, new_n50806_, new_n50807_,
    new_n50808_, new_n50809_, new_n50810_, new_n50811_, new_n50812_,
    new_n50813_, new_n50814_, new_n50815_, new_n50816_, new_n50818_,
    new_n50819_, new_n50820_, new_n50821_, new_n50822_, new_n50823_,
    new_n50824_, new_n50825_, new_n50826_, new_n50827_, new_n50828_,
    new_n50829_, new_n50831_, new_n50832_, new_n50833_, new_n50834_,
    new_n50835_, new_n50836_, new_n50837_, new_n50838_, new_n50839_,
    new_n50840_, new_n50841_, new_n50842_, new_n50844_, new_n50845_,
    new_n50846_, new_n50847_, new_n50848_, new_n50849_, new_n50850_,
    new_n50851_, new_n50852_, new_n50853_, new_n50854_, new_n50855_,
    new_n50857_, new_n50858_, new_n50859_, new_n50860_, new_n50861_,
    new_n50862_, new_n50863_, new_n50864_, new_n50865_, new_n50866_,
    new_n50867_, new_n50868_, new_n50870_, new_n50871_, new_n50872_,
    new_n50873_, new_n50874_, new_n50875_, new_n50876_, new_n50877_,
    new_n50878_, new_n50879_, new_n50880_, new_n50881_, new_n50883_,
    new_n50884_, new_n50885_, new_n50886_, new_n50887_, new_n50888_,
    new_n50889_, new_n50890_, new_n50891_, new_n50892_, new_n50893_,
    new_n50894_, new_n50896_, new_n50897_, new_n50898_, new_n50899_,
    new_n50900_, new_n50901_, new_n50902_, new_n50903_, new_n50904_,
    new_n50905_, new_n50906_, new_n50907_, new_n50909_, new_n50910_,
    new_n50911_, new_n50912_, new_n50913_, new_n50914_, new_n50915_,
    new_n50916_, new_n50917_, new_n50918_, new_n50919_, new_n50920_,
    new_n50922_, new_n50923_, new_n50924_, new_n50925_, new_n50926_,
    new_n50927_, new_n50928_, new_n50929_, new_n50930_, new_n50931_,
    new_n50932_, new_n50933_, new_n50935_, new_n50936_, new_n50937_,
    new_n50938_, new_n50939_, new_n50940_, new_n50941_, new_n50942_,
    new_n50943_, new_n50944_, new_n50945_, new_n50946_, new_n50948_,
    new_n50949_, new_n50950_, new_n50951_, new_n50953_, new_n50954_,
    new_n50955_, new_n50956_, new_n50957_, new_n50958_, new_n50959_,
    new_n50960_, new_n50961_, new_n50962_, new_n50963_, new_n50964_,
    new_n50965_, new_n50967_, new_n50968_, new_n50969_, new_n50970_,
    new_n50971_, new_n50972_, new_n50973_, new_n50974_, new_n50975_,
    new_n50977_, new_n50978_, new_n50979_, new_n50980_, new_n50981_,
    new_n50982_, new_n50983_, new_n50984_, new_n50985_, new_n50987_,
    new_n50988_, new_n50989_, new_n50990_, new_n50991_, new_n50992_,
    new_n50993_, new_n50994_, new_n50995_, new_n50997_, new_n50998_,
    new_n50999_, new_n51000_, new_n51001_, new_n51002_, new_n51003_,
    new_n51004_, new_n51005_, new_n51007_, new_n51008_, new_n51009_,
    new_n51010_, new_n51011_, new_n51012_, new_n51013_, new_n51014_,
    new_n51015_, new_n51017_, new_n51018_, new_n51019_, new_n51020_,
    new_n51021_, new_n51022_, new_n51023_, new_n51024_, new_n51025_,
    new_n51027_, new_n51028_, new_n51029_, new_n51030_, new_n51031_,
    new_n51032_, new_n51033_, new_n51034_, new_n51035_, new_n51037_,
    new_n51038_, new_n51039_, new_n51040_, new_n51041_, new_n51042_,
    new_n51043_, new_n51044_, new_n51045_, new_n51047_, new_n51048_,
    new_n51049_, new_n51050_, new_n51051_, new_n51052_, new_n51053_,
    new_n51054_, new_n51055_, new_n51057_, new_n51058_, new_n51059_,
    new_n51060_, new_n51061_, new_n51062_, new_n51063_, new_n51064_,
    new_n51065_, new_n51067_, new_n51068_, new_n51069_, new_n51070_,
    new_n51071_, new_n51072_, new_n51073_, new_n51074_, new_n51075_,
    new_n51077_, new_n51078_, new_n51079_, new_n51080_, new_n51081_,
    new_n51082_, new_n51083_, new_n51084_, new_n51085_, new_n51087_,
    new_n51088_, new_n51089_, new_n51090_, new_n51091_, new_n51092_,
    new_n51093_, new_n51094_, new_n51095_, new_n51097_, new_n51098_,
    new_n51099_, new_n51100_, new_n51101_, new_n51102_, new_n51103_,
    new_n51104_, new_n51105_, new_n51107_, new_n51108_, new_n51109_,
    new_n51110_, new_n51111_, new_n51112_, new_n51113_, new_n51114_,
    new_n51115_, new_n51117_, new_n51118_, new_n51119_, new_n51120_,
    new_n51121_, new_n51122_, new_n51123_, new_n51124_, new_n51125_,
    new_n51127_, new_n51128_, new_n51129_, new_n51130_, new_n51131_,
    new_n51132_, new_n51133_, new_n51134_, new_n51135_, new_n51137_,
    new_n51138_, new_n51139_, new_n51140_, new_n51141_, new_n51142_,
    new_n51143_, new_n51144_, new_n51145_, new_n51147_, new_n51148_,
    new_n51149_, new_n51150_, new_n51151_, new_n51152_, new_n51153_,
    new_n51154_, new_n51155_, new_n51157_, new_n51158_, new_n51159_,
    new_n51160_, new_n51161_, new_n51162_, new_n51163_, new_n51164_,
    new_n51165_, new_n51167_, new_n51168_, new_n51169_, new_n51170_,
    new_n51172_, new_n51173_, new_n51174_, new_n51175_, new_n51176_,
    new_n51177_, new_n51178_, new_n51179_, new_n51180_, new_n51181_,
    new_n51182_, new_n51183_, new_n51184_, new_n51186_, new_n51187_,
    new_n51188_, new_n51189_, new_n51190_, new_n51191_, new_n51192_,
    new_n51193_, new_n51194_, new_n51196_, new_n51197_, new_n51198_,
    new_n51199_, new_n51200_, new_n51201_, new_n51202_, new_n51203_,
    new_n51204_, new_n51206_, new_n51207_, new_n51208_, new_n51209_,
    new_n51210_, new_n51211_, new_n51212_, new_n51213_, new_n51214_,
    new_n51216_, new_n51217_, new_n51218_, new_n51219_, new_n51220_,
    new_n51221_, new_n51222_, new_n51223_, new_n51224_, new_n51226_,
    new_n51227_, new_n51228_, new_n51229_, new_n51230_, new_n51231_,
    new_n51232_, new_n51233_, new_n51234_, new_n51236_, new_n51237_,
    new_n51238_, new_n51239_, new_n51240_, new_n51241_, new_n51242_,
    new_n51243_, new_n51244_, new_n51246_, new_n51247_, new_n51248_,
    new_n51249_, new_n51250_, new_n51251_, new_n51252_, new_n51253_,
    new_n51254_, new_n51256_, new_n51257_, new_n51258_, new_n51259_,
    new_n51260_, new_n51261_, new_n51262_, new_n51263_, new_n51264_,
    new_n51266_, new_n51267_, new_n51268_, new_n51269_, new_n51270_,
    new_n51271_, new_n51272_, new_n51273_, new_n51274_, new_n51276_,
    new_n51277_, new_n51278_, new_n51279_, new_n51280_, new_n51281_,
    new_n51282_, new_n51283_, new_n51284_, new_n51286_, new_n51287_,
    new_n51288_, new_n51289_, new_n51290_, new_n51291_, new_n51292_,
    new_n51293_, new_n51294_, new_n51296_, new_n51297_, new_n51298_,
    new_n51299_, new_n51300_, new_n51301_, new_n51302_, new_n51303_,
    new_n51304_, new_n51306_, new_n51307_, new_n51308_, new_n51309_,
    new_n51310_, new_n51311_, new_n51312_, new_n51313_, new_n51314_,
    new_n51316_, new_n51317_, new_n51318_, new_n51319_, new_n51320_,
    new_n51321_, new_n51322_, new_n51323_, new_n51324_, new_n51326_,
    new_n51327_, new_n51328_, new_n51329_, new_n51330_, new_n51331_,
    new_n51332_, new_n51333_, new_n51334_, new_n51336_, new_n51337_,
    new_n51338_, new_n51339_, new_n51340_, new_n51341_, new_n51342_,
    new_n51343_, new_n51344_, new_n51346_, new_n51347_, new_n51348_,
    new_n51349_, new_n51350_, new_n51351_, new_n51352_, new_n51353_,
    new_n51354_, new_n51356_, new_n51357_, new_n51358_, new_n51359_,
    new_n51360_, new_n51361_, new_n51362_, new_n51363_, new_n51364_,
    new_n51366_, new_n51367_, new_n51368_, new_n51369_, new_n51370_,
    new_n51371_, new_n51372_, new_n51373_, new_n51374_, new_n51376_,
    new_n51377_, new_n51378_, new_n51379_, new_n51380_, new_n51381_,
    new_n51382_, new_n51383_, new_n51384_, new_n51386_, new_n51387_,
    new_n51388_, new_n51390_, new_n51391_, new_n51392_, new_n51393_,
    new_n51394_, new_n51395_, new_n51397_, new_n51398_, new_n51399_,
    new_n51400_, new_n51401_, new_n51402_, new_n51404_, new_n51405_,
    new_n51406_, new_n51407_, new_n51408_, new_n51409_, new_n51411_,
    new_n51412_, new_n51413_, new_n51414_, new_n51415_, new_n51416_,
    new_n51418_, new_n51419_, new_n51420_, new_n51421_, new_n51422_,
    new_n51423_, new_n51425_, new_n51426_, new_n51427_, new_n51428_,
    new_n51429_, new_n51430_, new_n51432_, new_n51433_, new_n51434_,
    new_n51435_, new_n51436_, new_n51437_, new_n51439_, new_n51440_,
    new_n51441_, new_n51442_, new_n51443_, new_n51444_, new_n51446_,
    new_n51447_, new_n51448_, new_n51449_, new_n51450_, new_n51451_,
    new_n51453_, new_n51454_, new_n51455_, new_n51456_, new_n51457_,
    new_n51458_, new_n51460_, new_n51461_, new_n51462_, new_n51463_,
    new_n51464_, new_n51465_, new_n51467_, new_n51468_, new_n51469_,
    new_n51470_, new_n51471_, new_n51472_, new_n51474_, new_n51475_,
    new_n51476_, new_n51477_, new_n51478_, new_n51479_, new_n51481_,
    new_n51482_, new_n51483_, new_n51484_, new_n51485_, new_n51486_,
    new_n51488_, new_n51489_, new_n51490_, new_n51491_, new_n51492_,
    new_n51493_, new_n51495_, new_n51496_, new_n51497_, new_n51498_,
    new_n51499_, new_n51500_, new_n51502_, new_n51503_, new_n51504_,
    new_n51505_, new_n51506_, new_n51507_, new_n51509_, new_n51510_,
    new_n51511_, new_n51512_, new_n51513_, new_n51514_, new_n51516_,
    new_n51517_, new_n51518_, new_n51519_, new_n51520_, new_n51521_,
    new_n51523_, new_n51524_, new_n51525_, new_n51526_, new_n51527_,
    new_n51528_, new_n51530_, new_n51531_, new_n51532_, new_n51533_,
    new_n51534_, new_n51535_, new_n51537_, new_n51538_, new_n51539_,
    new_n51540_, new_n51541_, new_n51542_, new_n51544_, new_n51545_,
    new_n51546_, new_n51547_, new_n51548_, new_n51549_, new_n51551_,
    new_n51552_, new_n51553_, new_n51554_, new_n51555_, new_n51556_,
    new_n51558_, new_n51559_, new_n51560_, new_n51561_, new_n51562_,
    new_n51563_, new_n51565_, new_n51566_, new_n51567_, new_n51568_,
    new_n51569_, new_n51570_, new_n51572_, new_n51573_, new_n51574_,
    new_n51575_, new_n51576_, new_n51577_, new_n51579_, new_n51580_,
    new_n51581_, new_n51582_, new_n51583_, new_n51584_, new_n51586_,
    new_n51587_, new_n51588_, new_n51589_, new_n51590_, new_n51591_,
    new_n51593_, new_n51594_, new_n51595_, new_n51596_, new_n51597_,
    new_n51598_, new_n51600_, new_n51601_, new_n51602_, new_n51603_,
    new_n51604_, new_n51605_, new_n51607_, new_n51608_, new_n51609_,
    new_n51610_, new_n51612_, new_n51615_, new_n51616_, new_n51617_,
    new_n51618_, new_n51619_, new_n51620_, new_n51621_, new_n51622_,
    new_n51623_, new_n51624_, new_n51625_, new_n51627_, new_n51628_,
    new_n51629_, new_n51630_, new_n51631_, new_n51635_, new_n51637_,
    new_n51638_, new_n51639_, new_n51640_, new_n51642_, new_n51643_,
    new_n51645_, new_n51646_, new_n51647_, new_n51649_, new_n51650_,
    new_n51651_, new_n51653_, new_n51654_, new_n51655_, new_n51656_,
    new_n51658_, new_n51659_, new_n51660_, new_n51662_, new_n51663_,
    new_n51664_, new_n51665_, new_n51667_, new_n51668_, new_n51669_,
    new_n51671_, new_n51672_, new_n51673_, new_n51674_, new_n51675_,
    new_n51677_, new_n51678_, new_n51679_, new_n51681_, new_n51682_,
    new_n51683_, new_n51684_, new_n51686_, new_n51687_, new_n51688_,
    new_n51690_, new_n51691_, new_n51692_, new_n51693_, new_n51694_,
    new_n51696_, new_n51697_, new_n51698_, new_n51700_, new_n51701_,
    new_n51702_, new_n51703_, new_n51705_, new_n51706_, new_n51707_,
    new_n51709_, new_n51710_, new_n51711_, new_n51712_, new_n51713_,
    new_n51714_, new_n51716_, new_n51717_, new_n51718_, new_n51720_,
    new_n51721_, new_n51722_, new_n51723_, new_n51725_, new_n51726_,
    new_n51727_, new_n51729_, new_n51730_, new_n51731_, new_n51732_,
    new_n51733_, new_n51735_, new_n51736_, new_n51737_, new_n51739_,
    new_n51740_, new_n51741_, new_n51742_, new_n51744_, new_n51745_,
    new_n51746_, new_n51748_, new_n51749_, new_n51750_, new_n51751_,
    new_n51752_, new_n51753_, new_n51755_, new_n51756_, new_n51757_,
    new_n51759_, new_n51760_, new_n51761_, new_n51762_, new_n51764_,
    new_n51765_, new_n51766_, new_n51768_, new_n51769_, new_n51770_,
    new_n51771_, new_n51772_, new_n51774_, new_n51775_, new_n51776_,
    new_n51778_, new_n51779_, new_n51780_, new_n51781_, new_n51783_,
    new_n51784_, new_n51785_, new_n51787_, new_n51788_, new_n51789_,
    new_n51790_, new_n51791_, new_n51792_, new_n51793_, new_n51795_,
    new_n51796_, new_n51798_, new_n51799_, new_n51801_, new_n51802_,
    new_n51803_, new_n51805_, new_n51806_, new_n51808_, new_n51809_,
    new_n51810_, new_n51812_, new_n51813_, new_n51814_, new_n51816_,
    new_n51817_, new_n51819_, new_n51820_, new_n51822_, new_n51823_,
    new_n51824_, new_n51826_, new_n51827_, new_n51829_, new_n51830_,
    new_n51831_, new_n51833_, new_n51834_, new_n51835_, new_n51837_,
    new_n51838_, new_n51842_, new_n51843_, new_n51845_, new_n51846_,
    new_n51847_, new_n51849_, new_n51850_, new_n51851_, new_n51852_,
    new_n51854_, new_n51855_, new_n51860_, new_n51861_, new_n51862_,
    new_n51863_, new_n51864_, new_n51865_, new_n51867_, new_n51868_,
    new_n51870_, new_n51871_, new_n51872_, new_n51874_, new_n51875_,
    new_n51876_, new_n51877_, new_n51878_, new_n51879_, new_n51880_,
    new_n51881_, new_n51882_, new_n51883_, new_n51884_, new_n51885_,
    new_n51886_, new_n51887_, new_n51888_, new_n51889_, new_n51890_,
    new_n51891_, new_n51892_, new_n51895_, new_n51896_, new_n51897_,
    new_n51898_, new_n51899_, new_n51903_, new_n51904_, new_n51905_,
    new_n51906_, new_n51907_, new_n51908_, new_n51909_, new_n51910_,
    new_n51911_, new_n51912_, new_n51913_, new_n51914_, new_n51916_,
    new_n51917_, new_n51918_, new_n51919_, new_n51920_, new_n51921_,
    new_n51922_, new_n51923_, new_n51924_, new_n51925_, new_n51926_,
    new_n51927_, new_n51928_, new_n51929_, new_n51930_, new_n51931_,
    new_n51932_, new_n51933_, new_n51934_, new_n51935_, new_n51936_,
    new_n51937_, new_n51938_, new_n51939_, new_n51940_, new_n51941_,
    new_n51942_, new_n51943_, new_n51944_, new_n51945_, new_n51946_,
    new_n51947_, new_n51948_, new_n51949_, new_n51950_, new_n51951_,
    new_n51952_, new_n51953_, new_n51954_, new_n51955_, new_n51956_,
    new_n51957_, new_n51958_, new_n51959_, new_n51960_, new_n51961_,
    new_n51962_, new_n51963_, new_n51964_, new_n51965_, new_n51966_,
    new_n51967_, new_n51968_, new_n51969_, new_n51970_, new_n51971_,
    new_n51972_, new_n51973_, new_n51974_, new_n51975_, new_n51976_,
    new_n51977_, new_n51978_, new_n51979_, new_n51980_, new_n51981_,
    new_n51982_, new_n51983_, new_n51984_, new_n51985_, new_n51986_,
    new_n51987_, new_n51988_, new_n51989_, new_n51990_, new_n51991_,
    new_n51992_, new_n51993_, new_n51994_, new_n51995_, new_n51996_,
    new_n51997_, new_n51998_, new_n51999_, new_n52000_, new_n52001_,
    new_n52002_, new_n52003_, new_n52004_, new_n52005_, new_n52006_,
    new_n52007_, new_n52008_, new_n52009_, new_n52010_, new_n52011_,
    new_n52012_, new_n52013_, new_n52014_, new_n52015_, new_n52016_,
    new_n52017_, new_n52018_, new_n52019_, new_n52020_, new_n52021_,
    new_n52022_, new_n52023_, new_n52024_, new_n52025_, new_n52026_,
    new_n52027_, new_n52028_, new_n52029_, new_n52030_, new_n52031_,
    new_n52032_, new_n52033_, new_n52034_, new_n52035_, new_n52036_,
    new_n52037_, new_n52038_, new_n52039_, new_n52040_, new_n52041_,
    new_n52042_, new_n52043_, new_n52044_, new_n52045_, new_n52046_,
    new_n52047_, new_n52048_, new_n52049_, new_n52050_, new_n52051_,
    new_n52052_, new_n52053_, new_n52054_, new_n52055_, new_n52056_,
    new_n52057_, new_n52058_, new_n52059_, new_n52060_, new_n52061_,
    new_n52062_, new_n52063_, new_n52064_, new_n52065_, new_n52066_,
    new_n52067_, new_n52068_, new_n52069_, new_n52070_, new_n52071_,
    new_n52072_, new_n52073_, new_n52074_, new_n52075_, new_n52076_,
    new_n52077_, new_n52078_, new_n52079_, new_n52080_, new_n52081_,
    new_n52082_, new_n52083_, new_n52084_, new_n52085_, new_n52086_,
    new_n52087_, new_n52088_, new_n52089_, new_n52090_, new_n52091_,
    new_n52092_, new_n52093_, new_n52094_, new_n52095_, new_n52096_,
    new_n52097_, new_n52098_, new_n52099_, new_n52100_, new_n52101_,
    new_n52102_, new_n52103_, new_n52104_, new_n52105_, new_n52106_,
    new_n52107_, new_n52108_, new_n52109_, new_n52110_, new_n52111_,
    new_n52112_, new_n52113_, new_n52114_, new_n52115_, new_n52116_,
    new_n52117_, new_n52118_, new_n52119_, new_n52120_, new_n52121_,
    new_n52122_, new_n52123_, new_n52124_, new_n52125_, new_n52126_,
    new_n52127_, new_n52128_, new_n52129_, new_n52130_, new_n52131_,
    new_n52132_, new_n52133_, new_n52134_, new_n52135_, new_n52136_,
    new_n52137_, new_n52138_, new_n52139_, new_n52140_, new_n52141_,
    new_n52142_, new_n52143_, new_n52144_, new_n52145_, new_n52146_,
    new_n52147_, new_n52148_, new_n52149_, new_n52150_, new_n52151_,
    new_n52152_, new_n52153_, new_n52154_, new_n52155_, new_n52156_,
    new_n52157_, new_n52158_, new_n52159_, new_n52160_, new_n52161_,
    new_n52162_, new_n52163_, new_n52164_, new_n52165_, new_n52166_,
    new_n52167_, new_n52168_, new_n52169_, new_n52170_, new_n52171_,
    new_n52172_, new_n52173_, new_n52174_, new_n52175_, new_n52176_,
    new_n52177_, new_n52178_, new_n52179_, new_n52180_, new_n52181_,
    new_n52182_, new_n52183_, new_n52184_, new_n52185_, new_n52186_,
    new_n52187_, new_n52188_, new_n52189_, new_n52190_, new_n52191_,
    new_n52192_, new_n52193_, new_n52194_, new_n52195_, new_n52196_,
    new_n52197_, new_n52198_, new_n52199_, new_n52200_, new_n52201_,
    new_n52202_, new_n52203_, new_n52204_, new_n52205_, new_n52206_,
    new_n52207_, new_n52208_, new_n52209_, new_n52210_, new_n52211_,
    new_n52212_, new_n52213_, new_n52214_, new_n52215_, new_n52216_,
    new_n52217_, new_n52218_, new_n52219_, new_n52220_, new_n52221_,
    new_n52222_, new_n52223_, new_n52224_, new_n52225_, new_n52226_,
    new_n52227_, new_n52228_, new_n52229_, new_n52230_, new_n52231_,
    new_n52232_, new_n52233_, new_n52234_, new_n52235_, new_n52236_,
    new_n52237_, new_n52238_, new_n52239_, new_n52240_, new_n52241_,
    new_n52242_, new_n52243_, new_n52244_, new_n52245_, new_n52246_,
    new_n52247_, new_n52248_, new_n52249_, new_n52250_, new_n52251_,
    new_n52252_, new_n52253_, new_n52254_, new_n52255_, new_n52256_,
    new_n52257_, new_n52258_, new_n52259_, new_n52260_, new_n52261_,
    new_n52262_, new_n52263_, new_n52264_, new_n52265_, new_n52266_,
    new_n52267_, new_n52268_, new_n52269_, new_n52270_, new_n52271_,
    new_n52272_, new_n52273_, new_n52274_, new_n52275_, new_n52276_,
    new_n52277_, new_n52278_, new_n52279_, new_n52280_, new_n52281_,
    new_n52282_, new_n52283_, new_n52284_, new_n52285_, new_n52286_,
    new_n52287_, new_n52288_, new_n52289_, new_n52290_, new_n52291_,
    new_n52292_, new_n52293_, new_n52294_, new_n52295_, new_n52296_,
    new_n52297_, new_n52298_, new_n52299_, new_n52300_, new_n52301_,
    new_n52302_, new_n52303_, new_n52304_, new_n52305_, new_n52306_,
    new_n52307_, new_n52308_, new_n52309_, new_n52310_, new_n52311_,
    new_n52312_, new_n52313_, new_n52314_, new_n52315_, new_n52316_,
    new_n52317_, new_n52318_, new_n52319_, new_n52320_, new_n52321_,
    new_n52322_, new_n52323_, new_n52324_, new_n52325_, new_n52326_,
    new_n52327_, new_n52328_, new_n52329_, new_n52330_, new_n52331_,
    new_n52332_, new_n52333_, new_n52334_, new_n52335_, new_n52336_,
    new_n52337_, new_n52338_, new_n52339_, new_n52340_, new_n52341_,
    new_n52342_, new_n52343_, new_n52344_, new_n52345_, new_n52346_,
    new_n52347_, new_n52348_, new_n52349_, new_n52350_, new_n52351_,
    new_n52352_, new_n52353_, new_n52354_, new_n52355_, new_n52356_,
    new_n52357_, new_n52358_, new_n52359_, new_n52360_, new_n52361_,
    new_n52362_, new_n52363_, new_n52364_, new_n52365_, new_n52366_,
    new_n52367_, new_n52368_, new_n52369_, new_n52370_, new_n52371_,
    new_n52372_, new_n52373_, new_n52374_, new_n52375_, new_n52376_,
    new_n52377_, new_n52378_, new_n52379_, new_n52380_, new_n52381_,
    new_n52382_, new_n52383_, new_n52384_, new_n52385_, new_n52386_,
    new_n52387_, new_n52388_, new_n52389_, new_n52390_, new_n52391_,
    new_n52392_, new_n52393_, new_n52394_, new_n52395_, new_n52396_,
    new_n52397_, new_n52398_, new_n52399_, new_n52400_, new_n52401_,
    new_n52402_, new_n52403_, new_n52404_, new_n52405_, new_n52406_,
    new_n52407_, new_n52408_, new_n52409_, new_n52410_, new_n52411_,
    new_n52412_, new_n52413_, new_n52414_, new_n52415_, new_n52416_,
    new_n52417_, new_n52418_, new_n52419_, new_n52420_, new_n52421_,
    new_n52422_, new_n52423_, new_n52424_, new_n52425_, new_n52426_,
    new_n52427_, new_n52428_, new_n52429_, new_n52430_, new_n52431_,
    new_n52432_, new_n52433_, new_n52434_, new_n52435_, new_n52436_,
    new_n52437_, new_n52438_, new_n52439_, new_n52440_, new_n52441_,
    new_n52442_, new_n52443_, new_n52444_, new_n52445_, new_n52446_,
    new_n52447_, new_n52448_, new_n52449_, new_n52450_, new_n52451_,
    new_n52452_, new_n52453_, new_n52454_, new_n52455_, new_n52456_,
    new_n52457_, new_n52458_, new_n52459_, new_n52460_, new_n52461_,
    new_n52462_, new_n52463_, new_n52464_, new_n52465_, new_n52466_,
    new_n52467_, new_n52468_, new_n52469_, new_n52470_, new_n52471_,
    new_n52472_, new_n52473_, new_n52474_, new_n52475_, new_n52476_,
    new_n52477_, new_n52478_, new_n52479_, new_n52480_, new_n52481_,
    new_n52482_, new_n52483_, new_n52484_, new_n52485_, new_n52486_,
    new_n52487_, new_n52488_, new_n52489_, new_n52490_, new_n52491_,
    new_n52492_, new_n52493_, new_n52494_, new_n52495_, new_n52496_,
    new_n52497_, new_n52498_, new_n52499_, new_n52500_, new_n52501_,
    new_n52502_, new_n52503_, new_n52504_, new_n52505_, new_n52506_,
    new_n52507_, new_n52508_, new_n52509_, new_n52510_, new_n52511_,
    new_n52512_, new_n52513_, new_n52514_, new_n52515_, new_n52516_,
    new_n52517_, new_n52518_, new_n52519_, new_n52520_, new_n52521_,
    new_n52522_, new_n52523_, new_n52524_, new_n52525_, new_n52526_,
    new_n52527_, new_n52528_, new_n52529_, new_n52530_, new_n52531_,
    new_n52532_, new_n52533_, new_n52534_, new_n52535_, new_n52536_,
    new_n52537_, new_n52538_, new_n52539_, new_n52540_, new_n52541_,
    new_n52542_, new_n52543_, new_n52545_, new_n52546_, new_n52547_,
    new_n52548_, new_n52549_, new_n52550_, new_n52551_, new_n52552_,
    new_n52553_, new_n52556_, new_n52557_, new_n52558_, new_n52559_,
    new_n52560_, new_n52561_, new_n52562_, new_n52563_, new_n52564_,
    new_n52565_, new_n52566_, new_n52567_, new_n52568_, new_n52573_,
    new_n52578_, new_n52580_, new_n52582_, new_n52583_, new_n52584_,
    new_n52586_, new_n52587_, new_n52588_, new_n52591_, new_n52596_,
    new_n52597_, new_n52598_, new_n52599_, new_n52600_, new_n52601_,
    new_n52603_, new_n52605_, new_n52606_, new_n52607_, new_n52608_,
    new_n52609_, new_n52611_, new_n52612_, new_n52613_, new_n52614_,
    new_n52615_, new_n52616_, new_n52617_, new_n52618_, new_n52619_,
    new_n52620_, new_n52621_, new_n52623_, new_n52624_, new_n52625_,
    new_n52626_, new_n52627_, new_n52628_, new_n52629_, new_n52630_,
    new_n52631_, new_n52632_, new_n52633_, new_n52634_, new_n52635_,
    new_n52636_, new_n52637_, new_n52638_, new_n52639_, new_n52640_,
    new_n52641_, new_n52642_, new_n52643_, new_n52644_, new_n52645_,
    new_n52646_, new_n52650_, new_n52651_, new_n52652_, new_n52656_,
    new_n52658_, new_n52659_, new_n52661_, new_n52662_, new_n52663_,
    new_n52665_, new_n52667_, new_n52668_, new_n52669_, new_n52671_,
    new_n52672_, new_n52674_, new_n52676_, new_n52677_, new_n52678_,
    new_n52679_, new_n52680_, new_n52681_, new_n52682_, new_n52683_,
    new_n52684_, new_n52686_, new_n52687_, new_n52688_, new_n52689_,
    new_n52690_, new_n52691_, new_n52692_, new_n52693_, new_n52694_,
    new_n52696_, new_n52697_, new_n52698_, new_n52699_, new_n52702_,
    new_n52703_, new_n52704_, new_n52705_, new_n52706_, new_n52707_,
    new_n52708_, new_n52709_, new_n52710_, new_n52711_, new_n52712_,
    new_n52713_, new_n52714_, new_n52715_, new_n52716_, new_n52717_,
    new_n52718_, new_n52719_, new_n52720_, new_n52722_, new_n52723_,
    new_n52724_, new_n52726_, new_n52728_, new_n52729_, new_n52730_,
    new_n52731_, new_n52732_, new_n52733_, new_n52734_, new_n52736_,
    new_n52737_, new_n52738_, new_n52739_, new_n52740_, new_n52742_,
    new_n52743_, new_n52744_, new_n52745_, new_n52746_, new_n52748_,
    new_n52749_, new_n52750_, new_n52751_, new_n52752_, new_n52753_,
    new_n52754_, new_n52755_, new_n52756_, new_n52757_, new_n52758_,
    new_n52759_, new_n52760_, new_n52762_, new_n52763_, new_n52764_,
    new_n52765_, new_n52766_, new_n52767_, new_n52768_, new_n52769_,
    new_n52770_, new_n52771_, new_n52773_, new_n52774_, new_n52775_,
    new_n52777_, new_n52778_, new_n52779_, new_n52780_, new_n52781_,
    new_n52782_, new_n52783_, new_n52784_, new_n52785_, new_n52786_,
    new_n52787_, new_n52788_, new_n52789_, new_n52790_, new_n52791_,
    new_n52792_, new_n52793_, new_n52794_, new_n52795_, new_n52796_,
    new_n52797_, new_n52798_, new_n52799_, new_n52800_, new_n52801_,
    new_n52802_, new_n52803_, new_n52804_, new_n52805_, new_n52806_,
    new_n52807_, new_n52808_, new_n52809_, new_n52810_, new_n52811_,
    new_n52812_, new_n52813_, new_n52814_, new_n52815_, new_n52816_,
    new_n52817_, new_n52818_, new_n52819_, new_n52820_, new_n52821_,
    new_n52822_, new_n52823_, new_n52824_, new_n52825_, new_n52826_,
    new_n52827_, new_n52828_, new_n52829_, new_n52830_, new_n52831_,
    new_n52832_, new_n52833_, new_n52834_, new_n52835_, new_n52836_,
    new_n52837_, new_n52838_, new_n52839_, new_n52840_, new_n52841_,
    new_n52842_, new_n52843_, new_n52844_, new_n52845_, new_n52846_,
    new_n52847_, new_n52848_, new_n52849_, new_n52850_, new_n52851_,
    new_n52852_, new_n52853_, new_n52854_, new_n52855_, new_n52856_,
    new_n52857_, new_n52858_, new_n52859_, new_n52860_, new_n52861_,
    new_n52862_, new_n52863_, new_n52864_, new_n52865_, new_n52866_,
    new_n52867_, new_n52868_, new_n52869_, new_n52870_, new_n52871_,
    new_n52872_, new_n52875_, new_n52876_, new_n52877_, new_n52879_,
    new_n52880_, new_n52881_, new_n52882_, new_n52883_, new_n52884_,
    new_n52886_, new_n52887_, new_n52888_, new_n52890_, new_n52891_,
    new_n52892_, new_n52894_, new_n52895_, new_n52896_, new_n52898_,
    new_n52899_, new_n52900_, new_n52902_, new_n52903_, new_n52904_,
    new_n52906_, new_n52907_, new_n52908_, new_n52910_, new_n52911_,
    new_n52912_, new_n52914_, new_n52915_, new_n52916_, new_n52918_,
    new_n52919_, new_n52920_, new_n52922_, new_n52923_, new_n52924_,
    new_n52932_, new_n52933_, new_n52934_, new_n52935_, new_n52936_,
    new_n52937_, new_n52938_, new_n52939_, new_n52940_, new_n52942_,
    new_n52943_, new_n52944_, new_n52945_, new_n52946_, new_n52948_,
    new_n52949_, new_n52950_, new_n52951_, new_n52952_, new_n52954_,
    new_n52955_, new_n52956_, new_n52957_, new_n52958_, new_n52960_,
    new_n52961_, new_n52962_, new_n52963_, new_n52965_, new_n52966_,
    new_n52967_, new_n52968_, new_n52969_, new_n52971_, new_n52972_,
    new_n52973_, new_n52974_, new_n52975_, new_n52976_, new_n52977_,
    new_n52979_, new_n52980_, new_n52981_, new_n52982_, new_n52983_,
    new_n52984_, new_n52985_, new_n52986_, new_n52987_, new_n52988_,
    new_n52989_, new_n52990_, new_n52991_, new_n52992_, new_n52993_,
    new_n52994_, new_n52996_, new_n52997_, new_n52998_, new_n52999_,
    new_n53000_, new_n53001_, new_n53003_, new_n53004_, new_n53005_,
    new_n53006_, new_n53008_, new_n53009_, new_n53010_, new_n53011_,
    new_n53012_, new_n53013_, new_n53014_, new_n53015_, new_n53016_,
    new_n53017_, new_n53018_, new_n53019_, new_n53020_, new_n53021_,
    new_n53022_, new_n53023_, new_n53024_, new_n53025_, new_n53026_,
    new_n53027_, new_n53028_, new_n53029_, new_n53030_, new_n53031_,
    new_n53032_, new_n53033_, new_n53034_, new_n53035_, new_n53036_,
    new_n53037_, new_n53038_, new_n53039_, new_n53040_, new_n53042_,
    new_n53043_, new_n53044_, new_n53045_, new_n53046_, new_n53047_,
    new_n53048_, new_n53049_, new_n53050_, new_n53051_, new_n53053_,
    new_n53054_, new_n53055_, new_n53056_, new_n53057_, new_n53058_,
    new_n53059_, new_n53060_, new_n53061_, new_n53062_, new_n53063_,
    new_n53064_, new_n53065_, new_n53066_, new_n53070_, new_n53071_,
    new_n53073_, new_n53075_, new_n53078_, new_n53080_, new_n53082_,
    new_n53084_, new_n53085_, new_n53086_, new_n53088_, new_n53089_,
    new_n53092_, new_n53093_, new_n53095_, new_n53096_, new_n53097_,
    new_n53098_, new_n53099_, new_n53100_, new_n53101_, new_n53104_,
    new_n53106_, new_n53108_, new_n53110_, new_n53111_, new_n53112_,
    new_n53113_, new_n53114_, new_n53115_, new_n53116_, new_n53117_,
    new_n53118_, new_n53120_, new_n53121_, new_n53122_, new_n53123_,
    new_n53124_, new_n53125_, new_n53128_, new_n53129_, new_n53133_,
    new_n53134_, new_n53135_, new_n53136_, new_n53137_, new_n53138_,
    new_n53139_, new_n53140_, new_n53141_, new_n53144_, new_n53147_,
    new_n53148_, new_n53149_, new_n53151_, new_n53152_, new_n53153_,
    new_n53155_, new_n53157_, new_n53158_, new_n53159_, new_n53160_,
    new_n53161_, new_n53162_, new_n53163_, new_n53164_, new_n53165_,
    new_n53166_, new_n53167_, new_n53169_, new_n53170_, new_n53173_,
    new_n53174_, new_n53175_, new_n53176_, new_n53177_, new_n53178_,
    new_n53179_, new_n53180_, new_n53181_, new_n53182_, new_n53183_,
    new_n53184_, new_n53185_, new_n53186_, new_n53187_, new_n53189_,
    new_n53190_, new_n53191_, new_n53192_, new_n53193_, new_n53195_,
    new_n53196_, new_n53197_, new_n53198_, new_n53199_, new_n53200_,
    new_n53201_, new_n53202_, new_n53203_, new_n53204_, new_n53205_,
    new_n53207_, new_n53208_, new_n53209_, new_n53210_, new_n53211_,
    new_n53213_, new_n53214_, new_n53215_, new_n53216_, new_n53217_,
    new_n53218_, new_n53219_, new_n53220_, new_n53222_, new_n53223_,
    new_n53224_, new_n53225_, new_n53226_, new_n53228_, new_n53229_,
    new_n53230_, new_n53231_, new_n53232_, new_n53233_, new_n53234_,
    new_n53235_, new_n53236_, new_n53237_, new_n53238_, new_n53239_,
    new_n53240_, new_n53241_, new_n53242_, new_n53243_, new_n53244_,
    new_n53245_, new_n53246_, new_n53247_, new_n53248_, new_n53249_,
    new_n53250_, new_n53251_, new_n53252_, new_n53253_, new_n53254_,
    new_n53255_, new_n53257_, new_n53258_, new_n53259_, new_n53260_,
    new_n53261_, new_n53262_, new_n53263_, new_n53265_, new_n53266_,
    new_n53267_, new_n53268_, new_n53269_, new_n53270_, new_n53271_,
    new_n53272_, new_n53273_, new_n53274_, new_n53275_, new_n53276_,
    new_n53278_, new_n53279_, new_n53280_, new_n53281_, new_n53282_,
    new_n53283_, new_n53284_, new_n53285_, new_n53286_, new_n53287_,
    new_n53288_, new_n53289_, new_n53290_, new_n53292_, new_n53293_,
    new_n53294_, new_n53295_, new_n53296_, new_n53297_, new_n53298_,
    new_n53299_, new_n53301_, new_n53302_, new_n53304_, new_n53305_,
    new_n53306_, new_n53307_, new_n53308_, new_n53310_, new_n53311_,
    new_n53312_, new_n53313_, new_n53314_, new_n53315_, new_n53316_,
    new_n53317_, new_n53318_, new_n53320_, new_n53321_, new_n53322_,
    new_n53323_, new_n53324_, new_n53326_, new_n53327_, new_n53328_,
    new_n53329_, new_n53330_, new_n53331_, new_n53332_, new_n53333_,
    new_n53335_, new_n53336_, new_n53337_, new_n53338_, new_n53339_,
    new_n53341_, new_n53342_, new_n53343_, new_n53344_, new_n53345_,
    new_n53346_, new_n53347_, new_n53348_, new_n53349_, new_n53350_,
    new_n53351_, new_n53352_, new_n53353_, new_n53355_, new_n53356_,
    new_n53357_, new_n53358_, new_n53359_, new_n53360_, new_n53361_,
    new_n53362_, new_n53363_, new_n53364_, new_n53365_, new_n53366_,
    new_n53368_, new_n53369_, new_n53370_, new_n53371_, new_n53372_,
    new_n53373_, new_n53374_, new_n53375_, new_n53376_, new_n53377_,
    new_n53378_, new_n53379_, new_n53380_, new_n53382_, new_n53383_,
    new_n53384_, new_n53385_, new_n53386_, new_n53387_, new_n53388_,
    new_n53389_, new_n53391_, new_n53392_, new_n53394_, new_n53395_,
    new_n53396_, new_n53397_, new_n53398_, new_n53400_, new_n53401_,
    new_n53402_, new_n53403_, new_n53404_, new_n53405_, new_n53406_,
    new_n53407_, new_n53408_, new_n53410_, new_n53411_, new_n53412_,
    new_n53413_, new_n53414_, new_n53416_, new_n53417_, new_n53418_,
    new_n53419_, new_n53420_, new_n53421_, new_n53422_, new_n53423_,
    new_n53425_, new_n53426_, new_n53427_, new_n53428_, new_n53429_,
    new_n53431_, new_n53432_, new_n53433_, new_n53434_, new_n53435_,
    new_n53436_, new_n53437_, new_n53438_, new_n53439_, new_n53440_,
    new_n53441_, new_n53442_, new_n53443_, new_n53445_, new_n53446_,
    new_n53447_, new_n53448_, new_n53449_, new_n53450_, new_n53451_,
    new_n53452_, new_n53453_, new_n53454_, new_n53455_, new_n53456_,
    new_n53458_, new_n53459_, new_n53460_, new_n53461_, new_n53462_,
    new_n53463_, new_n53464_, new_n53465_, new_n53466_, new_n53467_,
    new_n53468_, new_n53469_, new_n53470_, new_n53472_, new_n53473_,
    new_n53474_, new_n53475_, new_n53476_, new_n53477_, new_n53478_,
    new_n53479_, new_n53481_, new_n53482_, new_n53484_, new_n53485_,
    new_n53486_, new_n53487_, new_n53488_, new_n53490_, new_n53491_,
    new_n53492_, new_n53493_, new_n53494_, new_n53495_, new_n53496_,
    new_n53497_, new_n53498_, new_n53500_, new_n53501_, new_n53502_,
    new_n53503_, new_n53504_, new_n53506_, new_n53507_, new_n53508_,
    new_n53509_, new_n53510_, new_n53511_, new_n53512_, new_n53513_,
    new_n53515_, new_n53516_, new_n53517_, new_n53518_, new_n53519_,
    new_n53521_, new_n53522_, new_n53523_, new_n53524_, new_n53525_,
    new_n53526_, new_n53527_, new_n53528_, new_n53529_, new_n53530_,
    new_n53531_, new_n53532_, new_n53533_, new_n53535_, new_n53536_,
    new_n53537_, new_n53538_, new_n53539_, new_n53540_, new_n53541_,
    new_n53542_, new_n53543_, new_n53544_, new_n53545_, new_n53546_,
    new_n53548_, new_n53549_, new_n53550_, new_n53551_, new_n53552_,
    new_n53553_, new_n53554_, new_n53555_, new_n53556_, new_n53557_,
    new_n53558_, new_n53559_, new_n53560_, new_n53562_, new_n53563_,
    new_n53564_, new_n53565_, new_n53566_, new_n53567_, new_n53568_,
    new_n53569_, new_n53571_, new_n53572_, new_n53574_, new_n53575_,
    new_n53576_, new_n53577_, new_n53578_, new_n53580_, new_n53581_,
    new_n53582_, new_n53583_, new_n53584_, new_n53585_, new_n53586_,
    new_n53587_, new_n53588_, new_n53590_, new_n53591_, new_n53592_,
    new_n53593_, new_n53594_, new_n53596_, new_n53597_, new_n53598_,
    new_n53599_, new_n53600_, new_n53601_, new_n53602_, new_n53603_,
    new_n53605_, new_n53606_, new_n53607_, new_n53608_, new_n53609_,
    new_n53611_, new_n53612_, new_n53613_, new_n53614_, new_n53615_,
    new_n53616_, new_n53617_, new_n53618_, new_n53619_, new_n53620_,
    new_n53621_, new_n53622_, new_n53623_, new_n53625_, new_n53626_,
    new_n53627_, new_n53628_, new_n53629_, new_n53630_, new_n53631_,
    new_n53632_, new_n53633_, new_n53634_, new_n53635_, new_n53636_,
    new_n53638_, new_n53639_, new_n53640_, new_n53641_, new_n53642_,
    new_n53643_, new_n53644_, new_n53645_, new_n53646_, new_n53647_,
    new_n53648_, new_n53649_, new_n53650_, new_n53652_, new_n53653_,
    new_n53654_, new_n53655_, new_n53656_, new_n53657_, new_n53658_,
    new_n53659_, new_n53662_, new_n53663_, new_n53664_, new_n53665_,
    new_n53666_, new_n53667_, new_n53668_, new_n53670_, new_n53671_,
    new_n53672_, new_n53673_, new_n53674_, new_n53675_, new_n53676_,
    new_n53677_, new_n53678_, new_n53679_, new_n53680_, new_n53681_,
    new_n53682_, new_n53683_, new_n53684_, new_n53685_, new_n53686_,
    new_n53687_, new_n53689_, new_n53690_, new_n53691_, new_n53692_,
    new_n53693_, new_n53694_, new_n53695_, new_n53696_, new_n53697_,
    new_n53698_, new_n53699_, new_n53700_, new_n53702_, new_n53703_,
    new_n53704_, new_n53705_, new_n53706_, new_n53707_, new_n53708_,
    new_n53709_, new_n53710_, new_n53711_, new_n53712_, new_n53713_,
    new_n53714_, new_n53716_, new_n53717_, new_n53718_, new_n53719_,
    new_n53720_, new_n53722_, new_n53723_, new_n53724_, new_n53725_,
    new_n53726_, new_n53727_, new_n53728_, new_n53729_, new_n53730_,
    new_n53731_, new_n53732_, new_n53733_, new_n53734_, new_n53735_,
    new_n53736_, new_n53737_, new_n53738_, new_n53739_, new_n53740_,
    new_n53741_, new_n53742_, new_n53743_, new_n53744_, new_n53745_,
    new_n53746_, new_n53747_, new_n53748_, new_n53749_, new_n53752_,
    new_n53753_, new_n53754_, new_n53755_, new_n53756_, new_n53757_,
    new_n53758_, new_n53759_, new_n53760_, new_n53761_, new_n53762_,
    new_n53763_, new_n53764_, new_n53765_, new_n53766_, new_n53767_,
    new_n53768_, new_n53769_, new_n53770_, new_n53771_, new_n53772_,
    new_n53773_, new_n53774_, new_n53775_, new_n53776_, new_n53777_,
    new_n53778_, new_n53779_, new_n53780_, new_n53781_, new_n53782_,
    new_n53783_, new_n53784_, new_n53785_, new_n53786_, new_n53787_,
    new_n53788_, new_n53789_, new_n53790_, new_n53791_, new_n53792_,
    new_n53793_, new_n53794_, new_n53795_, new_n53796_, new_n53797_,
    new_n53798_, new_n53799_, new_n53800_, new_n53801_, new_n53802_,
    new_n53803_, new_n53804_, new_n53805_, new_n53806_, new_n53807_,
    new_n53808_, new_n53809_, new_n53810_, new_n53811_, new_n53812_,
    new_n53813_, new_n53814_, new_n53815_, new_n53816_, new_n53817_,
    new_n53818_, new_n53819_, new_n53820_, new_n53821_, new_n53822_,
    new_n53823_, new_n53824_, new_n53825_, new_n53826_, new_n53827_,
    new_n53828_, new_n53829_, new_n53830_, new_n53831_, new_n53832_,
    new_n53833_, new_n53834_, new_n53835_, new_n53836_, new_n53837_,
    new_n53838_, new_n53839_, new_n53840_, new_n53841_, new_n53842_,
    new_n53843_, new_n53844_, new_n53845_, new_n53846_, new_n53847_,
    new_n53848_, new_n53849_, new_n53850_, new_n53851_, new_n53852_,
    new_n53853_, new_n53854_, new_n53855_, new_n53856_, new_n53857_,
    new_n53858_, new_n53859_, new_n53860_, new_n53861_, new_n53862_,
    new_n53863_, new_n53864_, new_n53865_, new_n53866_, new_n53867_,
    new_n53868_, new_n53869_, new_n53870_, new_n53871_, new_n53872_,
    new_n53873_, new_n53874_, new_n53875_, new_n53876_, new_n53877_,
    new_n53878_, new_n53879_, new_n53880_, new_n53881_, new_n53882_,
    new_n53883_, new_n53884_, new_n53885_, new_n53886_, new_n53887_,
    new_n53888_, new_n53889_, new_n53890_, new_n53891_, new_n53892_,
    new_n53893_, new_n53894_, new_n53895_, new_n53896_, new_n53897_,
    new_n53898_, new_n53899_, new_n53900_, new_n53901_, new_n53902_,
    new_n53903_, new_n53904_, new_n53905_, new_n53906_, new_n53907_,
    new_n53908_, new_n53909_, new_n53910_, new_n53911_, new_n53912_,
    new_n53913_, new_n53914_, new_n53915_, new_n53916_, new_n53917_,
    new_n53918_, new_n53919_, new_n53920_, new_n53921_, new_n53922_,
    new_n53923_, new_n53924_, new_n53925_, new_n53926_, new_n53927_,
    new_n53928_, new_n53929_, new_n53930_, new_n53931_, new_n53932_,
    new_n53933_, new_n53934_, new_n53935_, new_n53936_, new_n53937_,
    new_n53938_, new_n53939_, new_n53940_, new_n53941_, new_n53942_,
    new_n53943_, new_n53944_, new_n53945_, new_n53946_, new_n53947_,
    new_n53948_, new_n53949_, new_n53950_, new_n53951_, new_n53952_,
    new_n53953_, new_n53954_, new_n53955_, new_n53956_, new_n53957_,
    new_n53958_, new_n53959_, new_n53960_, new_n53961_, new_n53962_,
    new_n53964_, new_n53965_, new_n53966_, new_n53967_, new_n53968_,
    new_n53969_, new_n53970_, new_n53971_, new_n53972_, new_n53973_,
    new_n53974_, new_n53975_, new_n53976_, new_n53977_, new_n53978_,
    new_n53979_, new_n53980_, new_n53981_, new_n53982_, new_n53983_,
    new_n53984_, new_n53985_, new_n53986_, new_n53987_, new_n53988_,
    new_n53989_, new_n53990_, new_n53991_, new_n53992_, new_n53993_,
    new_n53994_, new_n53995_, new_n53996_, new_n53997_, new_n53998_,
    new_n53999_, new_n54000_, new_n54001_, new_n54002_, new_n54003_,
    new_n54004_, new_n54005_, new_n54006_, new_n54007_, new_n54008_,
    new_n54009_, new_n54010_, new_n54011_, new_n54012_, new_n54013_,
    new_n54014_, new_n54015_, new_n54016_, new_n54018_, new_n54019_,
    new_n54020_, new_n54021_, new_n54022_, new_n54023_, new_n54024_,
    new_n54025_, new_n54026_, new_n54028_, new_n54029_, new_n54030_,
    new_n54031_, new_n54032_, new_n54033_, new_n54034_, new_n54035_,
    new_n54036_, new_n54037_, new_n54038_, new_n54039_, new_n54040_,
    new_n54041_, new_n54042_, new_n54043_, new_n54044_, new_n54045_,
    new_n54046_, new_n54047_, new_n54048_, new_n54049_, new_n54050_,
    new_n54051_, new_n54052_, new_n54053_, new_n54054_, new_n54055_,
    new_n54056_, new_n54057_, new_n54058_, new_n54059_, new_n54060_,
    new_n54061_, new_n54062_, new_n54063_, new_n54064_, new_n54065_,
    new_n54066_, new_n54067_, new_n54068_, new_n54069_, new_n54070_,
    new_n54071_, new_n54072_, new_n54073_, new_n54074_, new_n54075_,
    new_n54076_, new_n54077_, new_n54078_, new_n54080_, new_n54081_,
    new_n54082_, new_n54083_, new_n54084_, new_n54085_, new_n54086_,
    new_n54087_, new_n54088_, new_n54090_, new_n54091_, new_n54092_,
    new_n54093_, new_n54094_, new_n54095_, new_n54096_, new_n54097_,
    new_n54098_, new_n54099_, new_n54100_, new_n54101_, new_n54102_,
    new_n54103_, new_n54104_, new_n54105_, new_n54106_, new_n54107_,
    new_n54108_, new_n54109_, new_n54110_, new_n54111_, new_n54112_,
    new_n54113_, new_n54114_, new_n54115_, new_n54116_, new_n54117_,
    new_n54118_, new_n54119_, new_n54120_, new_n54121_, new_n54122_,
    new_n54123_, new_n54124_, new_n54125_, new_n54126_, new_n54127_,
    new_n54128_, new_n54129_, new_n54130_, new_n54131_, new_n54132_,
    new_n54133_, new_n54134_, new_n54135_, new_n54136_, new_n54137_,
    new_n54138_, new_n54139_, new_n54140_, new_n54141_, new_n54142_,
    new_n54143_, new_n54145_, new_n54146_, new_n54147_, new_n54148_,
    new_n54149_, new_n54150_, new_n54151_, new_n54152_, new_n54153_,
    new_n54155_, new_n54156_, new_n54157_, new_n54158_, new_n54159_,
    new_n54160_, new_n54161_, new_n54162_, new_n54163_, new_n54164_,
    new_n54165_, new_n54166_, new_n54167_, new_n54168_, new_n54169_,
    new_n54170_, new_n54171_, new_n54172_, new_n54173_, new_n54174_,
    new_n54175_, new_n54176_, new_n54177_, new_n54178_, new_n54179_,
    new_n54180_, new_n54181_, new_n54182_, new_n54183_, new_n54184_,
    new_n54185_, new_n54186_, new_n54187_, new_n54188_, new_n54189_,
    new_n54190_, new_n54191_, new_n54192_, new_n54193_, new_n54194_,
    new_n54195_, new_n54196_, new_n54197_, new_n54198_, new_n54199_,
    new_n54200_, new_n54201_, new_n54202_, new_n54203_, new_n54204_,
    new_n54205_, new_n54206_, new_n54207_, new_n54208_, new_n54209_,
    new_n54210_, new_n54211_, new_n54212_, new_n54213_, new_n54214_,
    new_n54215_, new_n54216_, new_n54217_, new_n54218_, new_n54219_,
    new_n54220_, new_n54221_, new_n54222_, new_n54224_, new_n54225_,
    new_n54226_, new_n54227_, new_n54228_, new_n54229_, new_n54230_,
    new_n54231_, new_n54232_, new_n54234_, new_n54235_, new_n54236_,
    new_n54237_, new_n54238_, new_n54239_, new_n54240_, new_n54241_,
    new_n54242_, new_n54243_, new_n54244_, new_n54245_, new_n54246_,
    new_n54247_, new_n54248_, new_n54249_, new_n54250_, new_n54251_,
    new_n54252_, new_n54253_, new_n54254_, new_n54255_, new_n54256_,
    new_n54257_, new_n54258_, new_n54259_, new_n54260_, new_n54261_,
    new_n54262_, new_n54263_, new_n54264_, new_n54265_, new_n54266_,
    new_n54267_, new_n54268_, new_n54269_, new_n54270_, new_n54271_,
    new_n54272_, new_n54273_, new_n54274_, new_n54275_, new_n54276_,
    new_n54277_, new_n54278_, new_n54279_, new_n54280_, new_n54281_,
    new_n54282_, new_n54283_, new_n54284_, new_n54285_, new_n54286_,
    new_n54287_, new_n54288_, new_n54289_, new_n54290_, new_n54291_,
    new_n54292_, new_n54293_, new_n54294_, new_n54295_, new_n54296_,
    new_n54297_, new_n54298_, new_n54299_, new_n54301_, new_n54302_,
    new_n54303_, new_n54304_, new_n54305_, new_n54306_, new_n54307_,
    new_n54308_, new_n54309_, new_n54311_, new_n54312_, new_n54313_,
    new_n54314_, new_n54315_, new_n54316_, new_n54317_, new_n54318_,
    new_n54319_, new_n54320_, new_n54321_, new_n54322_, new_n54323_,
    new_n54324_, new_n54325_, new_n54326_, new_n54327_, new_n54328_,
    new_n54329_, new_n54330_, new_n54331_, new_n54332_, new_n54333_,
    new_n54334_, new_n54335_, new_n54336_, new_n54337_, new_n54338_,
    new_n54339_, new_n54340_, new_n54341_, new_n54342_, new_n54343_,
    new_n54344_, new_n54345_, new_n54346_, new_n54347_, new_n54348_,
    new_n54349_, new_n54350_, new_n54351_, new_n54352_, new_n54353_,
    new_n54354_, new_n54355_, new_n54356_, new_n54357_, new_n54358_,
    new_n54359_, new_n54360_, new_n54361_, new_n54362_, new_n54363_,
    new_n54364_, new_n54365_, new_n54366_, new_n54367_, new_n54368_,
    new_n54369_, new_n54370_, new_n54371_, new_n54372_, new_n54373_,
    new_n54374_, new_n54375_, new_n54376_, new_n54377_, new_n54378_,
    new_n54379_, new_n54381_, new_n54382_, new_n54383_, new_n54384_,
    new_n54385_, new_n54386_, new_n54387_, new_n54388_, new_n54389_,
    new_n54391_, new_n54392_, new_n54393_, new_n54394_, new_n54395_,
    new_n54396_, new_n54397_, new_n54398_, new_n54399_, new_n54400_,
    new_n54401_, new_n54402_, new_n54403_, new_n54404_, new_n54405_,
    new_n54406_, new_n54407_, new_n54408_, new_n54409_, new_n54410_,
    new_n54411_, new_n54412_, new_n54413_, new_n54414_, new_n54415_,
    new_n54416_, new_n54417_, new_n54418_, new_n54419_, new_n54420_,
    new_n54421_, new_n54422_, new_n54423_, new_n54424_, new_n54425_,
    new_n54426_, new_n54427_, new_n54428_, new_n54429_, new_n54430_,
    new_n54431_, new_n54432_, new_n54433_, new_n54434_, new_n54435_,
    new_n54436_, new_n54437_, new_n54438_, new_n54439_, new_n54440_,
    new_n54441_, new_n54442_, new_n54443_, new_n54444_, new_n54445_,
    new_n54446_, new_n54447_, new_n54448_, new_n54449_, new_n54450_,
    new_n54451_, new_n54452_, new_n54453_, new_n54454_, new_n54455_,
    new_n54456_, new_n54457_, new_n54458_, new_n54459_, new_n54460_,
    new_n54461_, new_n54462_, new_n54463_, new_n54464_, new_n54465_,
    new_n54466_, new_n54467_, new_n54468_, new_n54469_, new_n54470_,
    new_n54471_, new_n54472_, new_n54473_, new_n54474_, new_n54475_,
    new_n54476_, new_n54477_, new_n54479_, new_n54480_, new_n54481_,
    new_n54482_, new_n54483_, new_n54484_, new_n54485_, new_n54486_,
    new_n54487_, new_n54489_, new_n54490_, new_n54491_, new_n54492_,
    new_n54493_, new_n54494_, new_n54495_, new_n54496_, new_n54497_,
    new_n54498_, new_n54499_, new_n54500_, new_n54501_, new_n54502_,
    new_n54503_, new_n54504_, new_n54505_, new_n54506_, new_n54507_,
    new_n54508_, new_n54509_, new_n54510_, new_n54511_, new_n54512_,
    new_n54513_, new_n54514_, new_n54515_, new_n54516_, new_n54517_,
    new_n54518_, new_n54519_, new_n54520_, new_n54521_, new_n54522_,
    new_n54523_, new_n54524_, new_n54525_, new_n54526_, new_n54527_,
    new_n54528_, new_n54529_, new_n54530_, new_n54531_, new_n54532_,
    new_n54533_, new_n54534_, new_n54535_, new_n54536_, new_n54537_,
    new_n54538_, new_n54539_, new_n54540_, new_n54541_, new_n54542_,
    new_n54543_, new_n54544_, new_n54545_, new_n54546_, new_n54547_,
    new_n54548_, new_n54549_, new_n54550_, new_n54551_, new_n54552_,
    new_n54553_, new_n54554_, new_n54555_, new_n54556_, new_n54557_,
    new_n54558_, new_n54559_, new_n54560_, new_n54561_, new_n54562_,
    new_n54563_, new_n54564_, new_n54565_, new_n54566_, new_n54567_,
    new_n54568_, new_n54569_, new_n54570_, new_n54571_, new_n54572_,
    new_n54573_, new_n54575_, new_n54576_, new_n54577_, new_n54578_,
    new_n54579_, new_n54580_, new_n54581_, new_n54582_, new_n54583_,
    new_n54585_, new_n54586_, new_n54587_, new_n54588_, new_n54589_,
    new_n54590_, new_n54591_, new_n54592_, new_n54593_, new_n54594_,
    new_n54595_, new_n54596_, new_n54597_, new_n54598_, new_n54599_,
    new_n54600_, new_n54601_, new_n54602_, new_n54603_, new_n54604_,
    new_n54605_, new_n54606_, new_n54607_, new_n54608_, new_n54609_,
    new_n54610_, new_n54611_, new_n54612_, new_n54613_, new_n54614_,
    new_n54615_, new_n54616_, new_n54617_, new_n54618_, new_n54619_,
    new_n54620_, new_n54621_, new_n54622_, new_n54623_, new_n54624_,
    new_n54625_, new_n54626_, new_n54627_, new_n54628_, new_n54629_,
    new_n54630_, new_n54631_, new_n54632_, new_n54633_, new_n54634_,
    new_n54635_, new_n54636_, new_n54637_, new_n54638_, new_n54639_,
    new_n54640_, new_n54641_, new_n54642_, new_n54643_, new_n54644_,
    new_n54645_, new_n54646_, new_n54647_, new_n54648_, new_n54649_,
    new_n54650_, new_n54651_, new_n54652_, new_n54653_, new_n54654_,
    new_n54655_, new_n54656_, new_n54657_, new_n54658_, new_n54659_,
    new_n54660_, new_n54661_, new_n54662_, new_n54663_, new_n54664_,
    new_n54665_, new_n54666_, new_n54667_, new_n54668_, new_n54669_,
    new_n54670_, new_n54671_, new_n54672_, new_n54673_, new_n54674_,
    new_n54675_, new_n54676_, new_n54677_, new_n54678_, new_n54679_,
    new_n54680_, new_n54681_, new_n54682_, new_n54684_, new_n54685_,
    new_n54686_, new_n54687_, new_n54688_, new_n54689_, new_n54690_,
    new_n54691_, new_n54692_, new_n54694_, new_n54695_, new_n54696_,
    new_n54697_, new_n54698_, new_n54699_, new_n54700_, new_n54701_,
    new_n54702_, new_n54703_, new_n54704_, new_n54705_, new_n54706_,
    new_n54707_, new_n54708_, new_n54709_, new_n54710_, new_n54711_,
    new_n54712_, new_n54713_, new_n54714_, new_n54715_, new_n54716_,
    new_n54717_, new_n54718_, new_n54719_, new_n54720_, new_n54721_,
    new_n54722_, new_n54723_, new_n54724_, new_n54725_, new_n54726_,
    new_n54727_, new_n54728_, new_n54729_, new_n54730_, new_n54731_,
    new_n54732_, new_n54733_, new_n54734_, new_n54735_, new_n54736_,
    new_n54737_, new_n54738_, new_n54739_, new_n54740_, new_n54741_,
    new_n54742_, new_n54743_, new_n54744_, new_n54745_, new_n54746_,
    new_n54747_, new_n54748_, new_n54749_, new_n54750_, new_n54751_,
    new_n54752_, new_n54753_, new_n54754_, new_n54755_, new_n54756_,
    new_n54757_, new_n54758_, new_n54759_, new_n54760_, new_n54761_,
    new_n54762_, new_n54763_, new_n54764_, new_n54765_, new_n54766_,
    new_n54767_, new_n54768_, new_n54769_, new_n54770_, new_n54771_,
    new_n54772_, new_n54773_, new_n54774_, new_n54775_, new_n54776_,
    new_n54777_, new_n54778_, new_n54779_, new_n54780_, new_n54781_,
    new_n54782_, new_n54783_, new_n54784_, new_n54785_, new_n54786_,
    new_n54787_, new_n54788_, new_n54789_, new_n54790_, new_n54791_,
    new_n54792_, new_n54793_, new_n54794_, new_n54795_, new_n54796_,
    new_n54797_, new_n54798_, new_n54799_, new_n54800_, new_n54801_,
    new_n54802_, new_n54803_, new_n54804_, new_n54805_, new_n54806_,
    new_n54808_, new_n54809_, new_n54810_, new_n54811_, new_n54812_,
    new_n54813_, new_n54814_, new_n54815_, new_n54816_, new_n54818_,
    new_n54819_, new_n54820_, new_n54821_, new_n54822_, new_n54823_,
    new_n54824_, new_n54825_, new_n54826_, new_n54827_, new_n54828_,
    new_n54829_, new_n54830_, new_n54831_, new_n54832_, new_n54833_,
    new_n54834_, new_n54835_, new_n54836_, new_n54837_, new_n54838_,
    new_n54839_, new_n54840_, new_n54841_, new_n54842_, new_n54843_,
    new_n54844_, new_n54845_, new_n54846_, new_n54847_, new_n54848_,
    new_n54849_, new_n54850_, new_n54851_, new_n54852_, new_n54853_,
    new_n54854_, new_n54855_, new_n54856_, new_n54857_, new_n54858_,
    new_n54859_, new_n54860_, new_n54861_, new_n54862_, new_n54863_,
    new_n54864_, new_n54865_, new_n54866_, new_n54867_, new_n54868_,
    new_n54869_, new_n54870_, new_n54871_, new_n54872_, new_n54873_,
    new_n54874_, new_n54875_, new_n54876_, new_n54877_, new_n54878_,
    new_n54879_, new_n54880_, new_n54881_, new_n54882_, new_n54883_,
    new_n54884_, new_n54885_, new_n54886_, new_n54887_, new_n54888_,
    new_n54889_, new_n54890_, new_n54891_, new_n54892_, new_n54893_,
    new_n54894_, new_n54895_, new_n54896_, new_n54897_, new_n54898_,
    new_n54899_, new_n54900_, new_n54901_, new_n54902_, new_n54903_,
    new_n54904_, new_n54905_, new_n54906_, new_n54907_, new_n54908_,
    new_n54909_, new_n54910_, new_n54911_, new_n54912_, new_n54913_,
    new_n54914_, new_n54915_, new_n54916_, new_n54917_, new_n54918_,
    new_n54919_, new_n54920_, new_n54921_, new_n54922_, new_n54923_,
    new_n54924_, new_n54925_, new_n54926_, new_n54927_, new_n54928_,
    new_n54930_, new_n54931_, new_n54932_, new_n54933_, new_n54934_,
    new_n54935_, new_n54936_, new_n54937_, new_n54938_, new_n54940_,
    new_n54941_, new_n54942_, new_n54943_, new_n54944_, new_n54945_,
    new_n54946_, new_n54947_, new_n54948_, new_n54949_, new_n54950_,
    new_n54951_, new_n54952_, new_n54953_, new_n54954_, new_n54955_,
    new_n54956_, new_n54957_, new_n54958_, new_n54959_, new_n54960_,
    new_n54961_, new_n54962_, new_n54963_, new_n54964_, new_n54965_,
    new_n54966_, new_n54967_, new_n54968_, new_n54969_, new_n54970_,
    new_n54971_, new_n54972_, new_n54973_, new_n54974_, new_n54975_,
    new_n54976_, new_n54977_, new_n54978_, new_n54979_, new_n54980_,
    new_n54981_, new_n54982_, new_n54983_, new_n54984_, new_n54985_,
    new_n54986_, new_n54987_, new_n54988_, new_n54989_, new_n54990_,
    new_n54991_, new_n54992_, new_n54993_, new_n54994_, new_n54995_,
    new_n54996_, new_n54997_, new_n54998_, new_n54999_, new_n55000_,
    new_n55001_, new_n55002_, new_n55003_, new_n55004_, new_n55005_,
    new_n55006_, new_n55007_, new_n55008_, new_n55009_, new_n55010_,
    new_n55011_, new_n55012_, new_n55013_, new_n55014_, new_n55015_,
    new_n55016_, new_n55017_, new_n55018_, new_n55019_, new_n55020_,
    new_n55021_, new_n55022_, new_n55023_, new_n55024_, new_n55025_,
    new_n55026_, new_n55027_, new_n55028_, new_n55029_, new_n55030_,
    new_n55031_, new_n55032_, new_n55033_, new_n55034_, new_n55035_,
    new_n55036_, new_n55037_, new_n55038_, new_n55039_, new_n55040_,
    new_n55041_, new_n55042_, new_n55043_, new_n55044_, new_n55045_,
    new_n55046_, new_n55047_, new_n55048_, new_n55049_, new_n55050_,
    new_n55051_, new_n55052_, new_n55053_, new_n55055_, new_n55056_,
    new_n55057_, new_n55058_, new_n55059_, new_n55060_, new_n55061_,
    new_n55062_, new_n55063_, new_n55065_, new_n55066_, new_n55067_,
    new_n55068_, new_n55069_, new_n55070_, new_n55071_, new_n55072_,
    new_n55073_, new_n55074_, new_n55075_, new_n55076_, new_n55077_,
    new_n55078_, new_n55079_, new_n55080_, new_n55081_, new_n55082_,
    new_n55083_, new_n55084_, new_n55085_, new_n55086_, new_n55087_,
    new_n55088_, new_n55089_, new_n55090_, new_n55091_, new_n55092_,
    new_n55093_, new_n55094_, new_n55095_, new_n55096_, new_n55097_,
    new_n55098_, new_n55099_, new_n55100_, new_n55101_, new_n55102_,
    new_n55103_, new_n55104_, new_n55105_, new_n55106_, new_n55107_,
    new_n55108_, new_n55109_, new_n55110_, new_n55111_, new_n55112_,
    new_n55113_, new_n55114_, new_n55115_, new_n55116_, new_n55117_,
    new_n55118_, new_n55119_, new_n55120_, new_n55121_, new_n55122_,
    new_n55123_, new_n55124_, new_n55125_, new_n55126_, new_n55127_,
    new_n55128_, new_n55129_, new_n55130_, new_n55131_, new_n55132_,
    new_n55133_, new_n55134_, new_n55135_, new_n55136_, new_n55137_,
    new_n55138_, new_n55139_, new_n55140_, new_n55141_, new_n55142_,
    new_n55143_, new_n55144_, new_n55145_, new_n55146_, new_n55147_,
    new_n55148_, new_n55149_, new_n55150_, new_n55151_, new_n55152_,
    new_n55153_, new_n55154_, new_n55155_, new_n55156_, new_n55157_,
    new_n55158_, new_n55159_, new_n55160_, new_n55161_, new_n55162_,
    new_n55163_, new_n55164_, new_n55165_, new_n55166_, new_n55167_,
    new_n55168_, new_n55169_, new_n55170_, new_n55171_, new_n55172_,
    new_n55173_, new_n55174_, new_n55175_, new_n55176_, new_n55177_,
    new_n55178_, new_n55179_, new_n55180_, new_n55181_, new_n55182_,
    new_n55183_, new_n55184_, new_n55185_, new_n55186_, new_n55187_,
    new_n55188_, new_n55189_, new_n55190_, new_n55191_, new_n55192_,
    new_n55194_, new_n55195_, new_n55196_, new_n55197_, new_n55198_,
    new_n55199_, new_n55200_, new_n55201_, new_n55202_, new_n55204_,
    new_n55205_, new_n55206_, new_n55207_, new_n55208_, new_n55209_,
    new_n55210_, new_n55211_, new_n55212_, new_n55213_, new_n55214_,
    new_n55215_, new_n55216_, new_n55217_, new_n55218_, new_n55219_,
    new_n55220_, new_n55221_, new_n55222_, new_n55223_, new_n55224_,
    new_n55225_, new_n55226_, new_n55227_, new_n55228_, new_n55229_,
    new_n55230_, new_n55231_, new_n55232_, new_n55233_, new_n55234_,
    new_n55235_, new_n55236_, new_n55237_, new_n55238_, new_n55239_,
    new_n55240_, new_n55241_, new_n55242_, new_n55243_, new_n55244_,
    new_n55245_, new_n55246_, new_n55247_, new_n55248_, new_n55249_,
    new_n55250_, new_n55251_, new_n55252_, new_n55253_, new_n55254_,
    new_n55255_, new_n55256_, new_n55257_, new_n55258_, new_n55259_,
    new_n55260_, new_n55261_, new_n55262_, new_n55263_, new_n55264_,
    new_n55265_, new_n55266_, new_n55267_, new_n55268_, new_n55269_,
    new_n55270_, new_n55271_, new_n55272_, new_n55273_, new_n55274_,
    new_n55275_, new_n55276_, new_n55277_, new_n55278_, new_n55279_,
    new_n55280_, new_n55281_, new_n55282_, new_n55283_, new_n55284_,
    new_n55285_, new_n55286_, new_n55287_, new_n55288_, new_n55289_,
    new_n55290_, new_n55291_, new_n55292_, new_n55293_, new_n55294_,
    new_n55295_, new_n55296_, new_n55297_, new_n55298_, new_n55299_,
    new_n55300_, new_n55301_, new_n55302_, new_n55303_, new_n55304_,
    new_n55305_, new_n55306_, new_n55307_, new_n55308_, new_n55309_,
    new_n55310_, new_n55311_, new_n55312_, new_n55313_, new_n55314_,
    new_n55315_, new_n55316_, new_n55317_, new_n55318_, new_n55319_,
    new_n55320_, new_n55321_, new_n55322_, new_n55323_, new_n55324_,
    new_n55325_, new_n55326_, new_n55327_, new_n55328_, new_n55329_,
    new_n55331_, new_n55332_, new_n55333_, new_n55334_, new_n55335_,
    new_n55336_, new_n55337_, new_n55338_, new_n55339_, new_n55341_,
    new_n55342_, new_n55343_, new_n55344_, new_n55345_, new_n55346_,
    new_n55347_, new_n55348_, new_n55349_, new_n55350_, new_n55351_,
    new_n55352_, new_n55353_, new_n55354_, new_n55355_, new_n55356_,
    new_n55357_, new_n55358_, new_n55359_, new_n55360_, new_n55361_,
    new_n55362_, new_n55363_, new_n55364_, new_n55365_, new_n55366_,
    new_n55367_, new_n55368_, new_n55369_, new_n55370_, new_n55371_,
    new_n55372_, new_n55373_, new_n55374_, new_n55375_, new_n55376_,
    new_n55377_, new_n55378_, new_n55379_, new_n55380_, new_n55381_,
    new_n55382_, new_n55383_, new_n55384_, new_n55385_, new_n55386_,
    new_n55387_, new_n55388_, new_n55389_, new_n55390_, new_n55391_,
    new_n55392_, new_n55393_, new_n55394_, new_n55395_, new_n55396_,
    new_n55397_, new_n55398_, new_n55399_, new_n55400_, new_n55401_,
    new_n55402_, new_n55403_, new_n55404_, new_n55405_, new_n55406_,
    new_n55407_, new_n55408_, new_n55409_, new_n55410_, new_n55411_,
    new_n55412_, new_n55413_, new_n55414_, new_n55415_, new_n55416_,
    new_n55417_, new_n55418_, new_n55419_, new_n55420_, new_n55421_,
    new_n55422_, new_n55423_, new_n55424_, new_n55425_, new_n55426_,
    new_n55427_, new_n55428_, new_n55429_, new_n55430_, new_n55431_,
    new_n55432_, new_n55433_, new_n55434_, new_n55435_, new_n55436_,
    new_n55437_, new_n55438_, new_n55439_, new_n55440_, new_n55441_,
    new_n55442_, new_n55443_, new_n55444_, new_n55445_, new_n55446_,
    new_n55447_, new_n55448_, new_n55449_, new_n55450_, new_n55451_,
    new_n55452_, new_n55453_, new_n55454_, new_n55455_, new_n55456_,
    new_n55457_, new_n55458_, new_n55459_, new_n55460_, new_n55461_,
    new_n55462_, new_n55463_, new_n55464_, new_n55465_, new_n55466_,
    new_n55467_, new_n55468_, new_n55469_, new_n55471_, new_n55472_,
    new_n55473_, new_n55474_, new_n55475_, new_n55476_, new_n55477_,
    new_n55478_, new_n55479_, new_n55481_, new_n55482_, new_n55483_,
    new_n55484_, new_n55485_, new_n55486_, new_n55487_, new_n55488_,
    new_n55489_, new_n55490_, new_n55491_, new_n55492_, new_n55493_,
    new_n55494_, new_n55495_, new_n55496_, new_n55497_, new_n55498_,
    new_n55499_, new_n55500_, new_n55501_, new_n55502_, new_n55503_,
    new_n55504_, new_n55505_, new_n55506_, new_n55507_, new_n55508_,
    new_n55509_, new_n55510_, new_n55511_, new_n55512_, new_n55513_,
    new_n55514_, new_n55515_, new_n55516_, new_n55517_, new_n55518_,
    new_n55519_, new_n55520_, new_n55521_, new_n55522_, new_n55523_,
    new_n55524_, new_n55525_, new_n55526_, new_n55527_, new_n55528_,
    new_n55529_, new_n55530_, new_n55531_, new_n55532_, new_n55533_,
    new_n55534_, new_n55535_, new_n55536_, new_n55537_, new_n55538_,
    new_n55539_, new_n55540_, new_n55541_, new_n55542_, new_n55543_,
    new_n55544_, new_n55545_, new_n55546_, new_n55547_, new_n55548_,
    new_n55549_, new_n55550_, new_n55551_, new_n55552_, new_n55553_,
    new_n55554_, new_n55555_, new_n55556_, new_n55557_, new_n55558_,
    new_n55559_, new_n55560_, new_n55561_, new_n55562_, new_n55563_,
    new_n55564_, new_n55565_, new_n55566_, new_n55567_, new_n55568_,
    new_n55569_, new_n55570_, new_n55571_, new_n55572_, new_n55573_,
    new_n55574_, new_n55575_, new_n55576_, new_n55577_, new_n55578_,
    new_n55579_, new_n55580_, new_n55581_, new_n55582_, new_n55583_,
    new_n55584_, new_n55585_, new_n55586_, new_n55587_, new_n55588_,
    new_n55589_, new_n55590_, new_n55591_, new_n55592_, new_n55593_,
    new_n55594_, new_n55595_, new_n55596_, new_n55597_, new_n55598_,
    new_n55599_, new_n55600_, new_n55601_, new_n55602_, new_n55603_,
    new_n55604_, new_n55605_, new_n55606_, new_n55607_, new_n55608_,
    new_n55609_, new_n55610_, new_n55611_, new_n55613_, new_n55614_,
    new_n55615_, new_n55616_, new_n55617_, new_n55618_, new_n55619_,
    new_n55620_, new_n55621_, new_n55623_, new_n55624_, new_n55625_,
    new_n55626_, new_n55627_, new_n55628_, new_n55629_, new_n55630_,
    new_n55631_, new_n55632_, new_n55633_, new_n55634_, new_n55635_,
    new_n55636_, new_n55637_, new_n55638_, new_n55639_, new_n55640_,
    new_n55641_, new_n55642_, new_n55643_, new_n55644_, new_n55645_,
    new_n55646_, new_n55647_, new_n55648_, new_n55649_, new_n55650_,
    new_n55651_, new_n55652_, new_n55653_, new_n55654_, new_n55655_,
    new_n55656_, new_n55657_, new_n55658_, new_n55659_, new_n55660_,
    new_n55661_, new_n55662_, new_n55663_, new_n55664_, new_n55665_,
    new_n55666_, new_n55667_, new_n55668_, new_n55669_, new_n55670_,
    new_n55671_, new_n55672_, new_n55673_, new_n55674_, new_n55675_,
    new_n55676_, new_n55677_, new_n55678_, new_n55679_, new_n55680_,
    new_n55681_, new_n55682_, new_n55683_, new_n55684_, new_n55685_,
    new_n55686_, new_n55687_, new_n55688_, new_n55689_, new_n55690_,
    new_n55691_, new_n55692_, new_n55693_, new_n55694_, new_n55695_,
    new_n55696_, new_n55697_, new_n55698_, new_n55699_, new_n55700_,
    new_n55701_, new_n55702_, new_n55703_, new_n55704_, new_n55705_,
    new_n55706_, new_n55707_, new_n55708_, new_n55709_, new_n55710_,
    new_n55711_, new_n55712_, new_n55713_, new_n55714_, new_n55715_,
    new_n55716_, new_n55717_, new_n55718_, new_n55719_, new_n55720_,
    new_n55721_, new_n55722_, new_n55723_, new_n55724_, new_n55725_,
    new_n55726_, new_n55727_, new_n55728_, new_n55729_, new_n55730_,
    new_n55731_, new_n55732_, new_n55733_, new_n55734_, new_n55735_,
    new_n55736_, new_n55737_, new_n55738_, new_n55739_, new_n55740_,
    new_n55741_, new_n55742_, new_n55743_, new_n55744_, new_n55745_,
    new_n55746_, new_n55747_, new_n55748_, new_n55749_, new_n55750_,
    new_n55751_, new_n55752_, new_n55753_, new_n55755_, new_n55756_,
    new_n55757_, new_n55758_, new_n55759_, new_n55760_, new_n55761_,
    new_n55762_, new_n55763_, new_n55765_, new_n55766_, new_n55767_,
    new_n55768_, new_n55769_, new_n55770_, new_n55771_, new_n55772_,
    new_n55773_, new_n55774_, new_n55775_, new_n55776_, new_n55777_,
    new_n55778_, new_n55779_, new_n55780_, new_n55781_, new_n55782_,
    new_n55783_, new_n55784_, new_n55785_, new_n55786_, new_n55787_,
    new_n55788_, new_n55789_, new_n55790_, new_n55791_, new_n55792_,
    new_n55793_, new_n55794_, new_n55795_, new_n55796_, new_n55797_,
    new_n55798_, new_n55799_, new_n55800_, new_n55801_, new_n55802_,
    new_n55803_, new_n55804_, new_n55805_, new_n55806_, new_n55807_,
    new_n55808_, new_n55809_, new_n55810_, new_n55811_, new_n55812_,
    new_n55813_, new_n55814_, new_n55815_, new_n55816_, new_n55817_,
    new_n55818_, new_n55819_, new_n55820_, new_n55821_, new_n55822_,
    new_n55823_, new_n55824_, new_n55825_, new_n55826_, new_n55827_,
    new_n55828_, new_n55829_, new_n55830_, new_n55831_, new_n55832_,
    new_n55833_, new_n55834_, new_n55835_, new_n55836_, new_n55837_,
    new_n55838_, new_n55839_, new_n55840_, new_n55841_, new_n55842_,
    new_n55843_, new_n55844_, new_n55845_, new_n55846_, new_n55847_,
    new_n55848_, new_n55849_, new_n55850_, new_n55851_, new_n55852_,
    new_n55853_, new_n55854_, new_n55855_, new_n55856_, new_n55857_,
    new_n55858_, new_n55859_, new_n55860_, new_n55861_, new_n55862_,
    new_n55863_, new_n55864_, new_n55865_, new_n55866_, new_n55867_,
    new_n55868_, new_n55869_, new_n55870_, new_n55871_, new_n55872_,
    new_n55873_, new_n55874_, new_n55875_, new_n55876_, new_n55877_,
    new_n55878_, new_n55879_, new_n55880_, new_n55881_, new_n55882_,
    new_n55883_, new_n55884_, new_n55885_, new_n55886_, new_n55887_,
    new_n55888_, new_n55889_, new_n55890_, new_n55891_, new_n55892_,
    new_n55893_, new_n55894_, new_n55895_, new_n55897_, new_n55898_,
    new_n55899_, new_n55900_, new_n55901_, new_n55902_, new_n55903_,
    new_n55904_, new_n55905_, new_n55907_, new_n55908_, new_n55909_,
    new_n55910_, new_n55911_, new_n55912_, new_n55913_, new_n55914_,
    new_n55915_, new_n55916_, new_n55917_, new_n55918_, new_n55919_,
    new_n55920_, new_n55921_, new_n55922_, new_n55923_, new_n55924_,
    new_n55925_, new_n55926_, new_n55927_, new_n55928_, new_n55929_,
    new_n55930_, new_n55931_, new_n55932_, new_n55933_, new_n55934_,
    new_n55935_, new_n55936_, new_n55937_, new_n55938_, new_n55939_,
    new_n55940_, new_n55941_, new_n55942_, new_n55943_, new_n55944_,
    new_n55945_, new_n55946_, new_n55947_, new_n55948_, new_n55949_,
    new_n55950_, new_n55951_, new_n55952_, new_n55953_, new_n55954_,
    new_n55955_, new_n55956_, new_n55957_, new_n55958_, new_n55959_,
    new_n55960_, new_n55961_, new_n55962_, new_n55963_, new_n55964_,
    new_n55965_, new_n55966_, new_n55967_, new_n55968_, new_n55969_,
    new_n55970_, new_n55971_, new_n55972_, new_n55973_, new_n55974_,
    new_n55975_, new_n55976_, new_n55977_, new_n55978_, new_n55979_,
    new_n55980_, new_n55981_, new_n55982_, new_n55983_, new_n55984_,
    new_n55985_, new_n55986_, new_n55987_, new_n55988_, new_n55989_,
    new_n55990_, new_n55991_, new_n55992_, new_n55993_, new_n55994_,
    new_n55995_, new_n55996_, new_n55997_, new_n55998_, new_n55999_,
    new_n56000_, new_n56001_, new_n56002_, new_n56003_, new_n56004_,
    new_n56005_, new_n56006_, new_n56007_, new_n56008_, new_n56009_,
    new_n56010_, new_n56011_, new_n56012_, new_n56013_, new_n56014_,
    new_n56015_, new_n56016_, new_n56017_, new_n56018_, new_n56019_,
    new_n56020_, new_n56021_, new_n56022_, new_n56023_, new_n56024_,
    new_n56025_, new_n56026_, new_n56027_, new_n56028_, new_n56029_,
    new_n56030_, new_n56031_, new_n56032_, new_n56033_, new_n56034_,
    new_n56035_, new_n56036_, new_n56037_, new_n56039_, new_n56040_,
    new_n56041_, new_n56042_, new_n56043_, new_n56044_, new_n56045_,
    new_n56046_, new_n56047_, new_n56049_, new_n56050_, new_n56051_,
    new_n56052_, new_n56053_, new_n56054_, new_n56055_, new_n56056_,
    new_n56057_, new_n56058_, new_n56059_, new_n56060_, new_n56061_,
    new_n56062_, new_n56063_, new_n56064_, new_n56065_, new_n56066_,
    new_n56067_, new_n56068_, new_n56069_, new_n56070_, new_n56071_,
    new_n56072_, new_n56073_, new_n56074_, new_n56075_, new_n56076_,
    new_n56077_, new_n56078_, new_n56079_, new_n56080_, new_n56081_,
    new_n56082_, new_n56083_, new_n56084_, new_n56085_, new_n56086_,
    new_n56087_, new_n56088_, new_n56089_, new_n56090_, new_n56091_,
    new_n56092_, new_n56093_, new_n56094_, new_n56095_, new_n56096_,
    new_n56097_, new_n56098_, new_n56099_, new_n56100_, new_n56101_,
    new_n56102_, new_n56103_, new_n56104_, new_n56105_, new_n56106_,
    new_n56107_, new_n56108_, new_n56109_, new_n56110_, new_n56111_,
    new_n56112_, new_n56113_, new_n56114_, new_n56115_, new_n56116_,
    new_n56117_, new_n56118_, new_n56119_, new_n56120_, new_n56121_,
    new_n56122_, new_n56123_, new_n56124_, new_n56125_, new_n56126_,
    new_n56127_, new_n56128_, new_n56129_, new_n56130_, new_n56131_,
    new_n56132_, new_n56133_, new_n56134_, new_n56135_, new_n56136_,
    new_n56137_, new_n56138_, new_n56139_, new_n56140_, new_n56141_,
    new_n56142_, new_n56143_, new_n56144_, new_n56145_, new_n56146_,
    new_n56147_, new_n56148_, new_n56149_, new_n56150_, new_n56151_,
    new_n56152_, new_n56153_, new_n56154_, new_n56155_, new_n56156_,
    new_n56157_, new_n56158_, new_n56159_, new_n56160_, new_n56161_,
    new_n56162_, new_n56163_, new_n56164_, new_n56165_, new_n56166_,
    new_n56167_, new_n56168_, new_n56169_, new_n56170_, new_n56171_,
    new_n56172_, new_n56173_, new_n56174_, new_n56175_, new_n56176_,
    new_n56177_, new_n56178_, new_n56179_, new_n56181_, new_n56182_,
    new_n56183_, new_n56184_, new_n56185_, new_n56186_, new_n56187_,
    new_n56188_, new_n56189_, new_n56191_, new_n56192_, new_n56193_,
    new_n56194_, new_n56195_, new_n56196_, new_n56197_, new_n56198_,
    new_n56199_, new_n56200_, new_n56201_, new_n56202_, new_n56203_,
    new_n56204_, new_n56205_, new_n56206_, new_n56207_, new_n56208_,
    new_n56209_, new_n56210_, new_n56211_, new_n56212_, new_n56213_,
    new_n56214_, new_n56215_, new_n56216_, new_n56217_, new_n56218_,
    new_n56219_, new_n56220_, new_n56221_, new_n56222_, new_n56223_,
    new_n56224_, new_n56225_, new_n56226_, new_n56227_, new_n56228_,
    new_n56229_, new_n56230_, new_n56231_, new_n56232_, new_n56233_,
    new_n56234_, new_n56235_, new_n56236_, new_n56237_, new_n56238_,
    new_n56239_, new_n56240_, new_n56241_, new_n56242_, new_n56243_,
    new_n56244_, new_n56245_, new_n56246_, new_n56247_, new_n56248_,
    new_n56249_, new_n56250_, new_n56251_, new_n56252_, new_n56253_,
    new_n56254_, new_n56255_, new_n56256_, new_n56257_, new_n56258_,
    new_n56259_, new_n56260_, new_n56261_, new_n56262_, new_n56263_,
    new_n56264_, new_n56265_, new_n56266_, new_n56267_, new_n56268_,
    new_n56269_, new_n56270_, new_n56271_, new_n56272_, new_n56273_,
    new_n56274_, new_n56275_, new_n56276_, new_n56277_, new_n56278_,
    new_n56279_, new_n56280_, new_n56281_, new_n56282_, new_n56283_,
    new_n56284_, new_n56285_, new_n56286_, new_n56287_, new_n56288_,
    new_n56289_, new_n56290_, new_n56291_, new_n56292_, new_n56293_,
    new_n56294_, new_n56295_, new_n56296_, new_n56297_, new_n56298_,
    new_n56299_, new_n56300_, new_n56301_, new_n56302_, new_n56303_,
    new_n56304_, new_n56305_, new_n56306_, new_n56307_, new_n56308_,
    new_n56309_, new_n56310_, new_n56311_, new_n56312_, new_n56313_,
    new_n56314_, new_n56315_, new_n56316_, new_n56317_, new_n56318_,
    new_n56319_, new_n56320_, new_n56321_, new_n56323_, new_n56324_,
    new_n56325_, new_n56326_, new_n56327_, new_n56328_, new_n56329_,
    new_n56330_, new_n56331_, new_n56333_, new_n56334_, new_n56335_,
    new_n56336_, new_n56337_, new_n56338_, new_n56339_, new_n56340_,
    new_n56341_, new_n56342_, new_n56343_, new_n56344_, new_n56345_,
    new_n56346_, new_n56347_, new_n56348_, new_n56349_, new_n56350_,
    new_n56351_, new_n56352_, new_n56353_, new_n56354_, new_n56355_,
    new_n56356_, new_n56357_, new_n56358_, new_n56359_, new_n56360_,
    new_n56361_, new_n56362_, new_n56363_, new_n56364_, new_n56365_,
    new_n56366_, new_n56367_, new_n56368_, new_n56369_, new_n56370_,
    new_n56371_, new_n56372_, new_n56373_, new_n56374_, new_n56375_,
    new_n56376_, new_n56377_, new_n56378_, new_n56379_, new_n56380_,
    new_n56381_, new_n56382_, new_n56383_, new_n56384_, new_n56385_,
    new_n56386_, new_n56387_, new_n56388_, new_n56389_, new_n56390_,
    new_n56391_, new_n56392_, new_n56393_, new_n56394_, new_n56395_,
    new_n56396_, new_n56397_, new_n56398_, new_n56399_, new_n56400_,
    new_n56401_, new_n56402_, new_n56403_, new_n56404_, new_n56405_,
    new_n56406_, new_n56407_, new_n56408_, new_n56409_, new_n56410_,
    new_n56411_, new_n56412_, new_n56413_, new_n56414_, new_n56415_,
    new_n56416_, new_n56417_, new_n56418_, new_n56419_, new_n56420_,
    new_n56421_, new_n56422_, new_n56423_, new_n56424_, new_n56425_,
    new_n56426_, new_n56427_, new_n56428_, new_n56429_, new_n56430_,
    new_n56431_, new_n56432_, new_n56433_, new_n56434_, new_n56435_,
    new_n56436_, new_n56437_, new_n56438_, new_n56439_, new_n56440_,
    new_n56441_, new_n56442_, new_n56443_, new_n56444_, new_n56445_,
    new_n56446_, new_n56447_, new_n56448_, new_n56449_, new_n56450_,
    new_n56451_, new_n56452_, new_n56453_, new_n56454_, new_n56455_,
    new_n56456_, new_n56457_, new_n56458_, new_n56459_, new_n56460_,
    new_n56461_, new_n56462_, new_n56463_, new_n56465_, new_n56466_,
    new_n56467_, new_n56468_, new_n56469_, new_n56470_, new_n56471_,
    new_n56472_, new_n56473_, new_n56475_, new_n56476_, new_n56477_,
    new_n56478_, new_n56479_, new_n56480_, new_n56481_, new_n56482_,
    new_n56483_, new_n56484_, new_n56485_, new_n56486_, new_n56487_,
    new_n56488_, new_n56489_, new_n56490_, new_n56491_, new_n56492_,
    new_n56493_, new_n56494_, new_n56495_, new_n56496_, new_n56497_,
    new_n56498_, new_n56499_, new_n56500_, new_n56501_, new_n56502_,
    new_n56503_, new_n56504_, new_n56505_, new_n56506_, new_n56507_,
    new_n56508_, new_n56509_, new_n56510_, new_n56511_, new_n56512_,
    new_n56513_, new_n56514_, new_n56515_, new_n56516_, new_n56517_,
    new_n56518_, new_n56519_, new_n56520_, new_n56521_, new_n56522_,
    new_n56523_, new_n56524_, new_n56525_, new_n56526_, new_n56527_,
    new_n56528_, new_n56529_, new_n56530_, new_n56531_, new_n56532_,
    new_n56533_, new_n56534_, new_n56535_, new_n56536_, new_n56537_,
    new_n56538_, new_n56539_, new_n56540_, new_n56541_, new_n56542_,
    new_n56543_, new_n56544_, new_n56545_, new_n56546_, new_n56547_,
    new_n56548_, new_n56549_, new_n56550_, new_n56551_, new_n56552_,
    new_n56553_, new_n56554_, new_n56555_, new_n56556_, new_n56557_,
    new_n56558_, new_n56559_, new_n56560_, new_n56561_, new_n56562_,
    new_n56563_, new_n56564_, new_n56565_, new_n56566_, new_n56567_,
    new_n56568_, new_n56569_, new_n56570_, new_n56571_, new_n56572_,
    new_n56573_, new_n56574_, new_n56575_, new_n56576_, new_n56577_,
    new_n56578_, new_n56579_, new_n56580_, new_n56581_, new_n56582_,
    new_n56583_, new_n56584_, new_n56585_, new_n56586_, new_n56587_,
    new_n56588_, new_n56589_, new_n56590_, new_n56591_, new_n56592_,
    new_n56593_, new_n56594_, new_n56595_, new_n56596_, new_n56597_,
    new_n56598_, new_n56599_, new_n56600_, new_n56601_, new_n56602_,
    new_n56603_, new_n56604_, new_n56605_, new_n56607_, new_n56608_,
    new_n56609_, new_n56610_, new_n56611_, new_n56612_, new_n56613_,
    new_n56614_, new_n56615_, new_n56617_, new_n56618_, new_n56619_,
    new_n56620_, new_n56621_, new_n56622_, new_n56623_, new_n56624_,
    new_n56625_, new_n56626_, new_n56627_, new_n56628_, new_n56629_,
    new_n56630_, new_n56631_, new_n56632_, new_n56633_, new_n56634_,
    new_n56635_, new_n56636_, new_n56637_, new_n56638_, new_n56639_,
    new_n56640_, new_n56641_, new_n56642_, new_n56643_, new_n56644_,
    new_n56645_, new_n56646_, new_n56647_, new_n56648_, new_n56649_,
    new_n56650_, new_n56651_, new_n56652_, new_n56653_, new_n56654_,
    new_n56655_, new_n56656_, new_n56657_, new_n56658_, new_n56659_,
    new_n56660_, new_n56661_, new_n56662_, new_n56663_, new_n56664_,
    new_n56665_, new_n56666_, new_n56667_, new_n56668_, new_n56669_,
    new_n56670_, new_n56671_, new_n56672_, new_n56673_, new_n56674_,
    new_n56675_, new_n56676_, new_n56677_, new_n56678_, new_n56679_,
    new_n56680_, new_n56681_, new_n56682_, new_n56683_, new_n56684_,
    new_n56685_, new_n56686_, new_n56687_, new_n56688_, new_n56689_,
    new_n56690_, new_n56691_, new_n56692_, new_n56693_, new_n56694_,
    new_n56695_, new_n56696_, new_n56697_, new_n56698_, new_n56699_,
    new_n56700_, new_n56701_, new_n56702_, new_n56703_, new_n56704_,
    new_n56705_, new_n56706_, new_n56707_, new_n56708_, new_n56709_,
    new_n56710_, new_n56711_, new_n56712_, new_n56713_, new_n56714_,
    new_n56715_, new_n56716_, new_n56717_, new_n56718_, new_n56719_,
    new_n56720_, new_n56721_, new_n56722_, new_n56723_, new_n56724_,
    new_n56725_, new_n56726_, new_n56727_, new_n56728_, new_n56729_,
    new_n56730_, new_n56731_, new_n56732_, new_n56733_, new_n56734_,
    new_n56735_, new_n56736_, new_n56737_, new_n56738_, new_n56739_,
    new_n56740_, new_n56741_, new_n56742_, new_n56743_, new_n56744_,
    new_n56745_, new_n56746_, new_n56747_, new_n56749_, new_n56750_,
    new_n56751_, new_n56752_, new_n56753_, new_n56754_, new_n56755_,
    new_n56756_, new_n56757_, new_n56759_, new_n56760_, new_n56761_,
    new_n56762_, new_n56763_, new_n56764_, new_n56765_, new_n56766_,
    new_n56767_, new_n56768_, new_n56769_, new_n56770_, new_n56771_,
    new_n56772_, new_n56773_, new_n56774_, new_n56775_, new_n56776_,
    new_n56777_, new_n56778_, new_n56779_, new_n56780_, new_n56781_,
    new_n56782_, new_n56783_, new_n56784_, new_n56785_, new_n56786_,
    new_n56787_, new_n56788_, new_n56789_, new_n56790_, new_n56791_,
    new_n56792_, new_n56793_, new_n56794_, new_n56795_, new_n56796_,
    new_n56797_, new_n56798_, new_n56799_, new_n56800_, new_n56801_,
    new_n56802_, new_n56803_, new_n56804_, new_n56805_, new_n56806_,
    new_n56807_, new_n56808_, new_n56809_, new_n56810_, new_n56811_,
    new_n56812_, new_n56813_, new_n56814_, new_n56815_, new_n56816_,
    new_n56817_, new_n56818_, new_n56819_, new_n56820_, new_n56821_,
    new_n56822_, new_n56823_, new_n56824_, new_n56825_, new_n56826_,
    new_n56827_, new_n56828_, new_n56829_, new_n56830_, new_n56831_,
    new_n56832_, new_n56833_, new_n56834_, new_n56835_, new_n56836_,
    new_n56837_, new_n56838_, new_n56839_, new_n56840_, new_n56841_,
    new_n56842_, new_n56843_, new_n56844_, new_n56845_, new_n56846_,
    new_n56847_, new_n56848_, new_n56849_, new_n56850_, new_n56851_,
    new_n56852_, new_n56853_, new_n56854_, new_n56855_, new_n56856_,
    new_n56857_, new_n56858_, new_n56859_, new_n56860_, new_n56861_,
    new_n56862_, new_n56863_, new_n56864_, new_n56865_, new_n56866_,
    new_n56867_, new_n56868_, new_n56869_, new_n56870_, new_n56871_,
    new_n56872_, new_n56873_, new_n56874_, new_n56875_, new_n56876_,
    new_n56877_, new_n56878_, new_n56879_, new_n56880_, new_n56881_,
    new_n56882_, new_n56883_, new_n56884_, new_n56885_, new_n56886_,
    new_n56887_, new_n56888_, new_n56889_, new_n56891_, new_n56892_,
    new_n56893_, new_n56894_, new_n56895_, new_n56896_, new_n56897_,
    new_n56898_, new_n56899_, new_n56901_, new_n56902_, new_n56903_,
    new_n56904_, new_n56905_, new_n56906_, new_n56907_, new_n56908_,
    new_n56909_, new_n56910_, new_n56911_, new_n56912_, new_n56913_,
    new_n56914_, new_n56915_, new_n56916_, new_n56917_, new_n56918_,
    new_n56919_, new_n56920_, new_n56921_, new_n56922_, new_n56923_,
    new_n56924_, new_n56925_, new_n56926_, new_n56927_, new_n56928_,
    new_n56929_, new_n56930_, new_n56931_, new_n56932_, new_n56933_,
    new_n56934_, new_n56935_, new_n56936_, new_n56937_, new_n56938_,
    new_n56939_, new_n56940_, new_n56941_, new_n56942_, new_n56943_,
    new_n56944_, new_n56945_, new_n56946_, new_n56947_, new_n56948_,
    new_n56949_, new_n56950_, new_n56951_, new_n56952_, new_n56953_,
    new_n56954_, new_n56955_, new_n56956_, new_n56957_, new_n56958_,
    new_n56959_, new_n56960_, new_n56961_, new_n56962_, new_n56963_,
    new_n56964_, new_n56965_, new_n56966_, new_n56967_, new_n56968_,
    new_n56969_, new_n56970_, new_n56971_, new_n56972_, new_n56973_,
    new_n56974_, new_n56975_, new_n56976_, new_n56977_, new_n56978_,
    new_n56979_, new_n56980_, new_n56981_, new_n56982_, new_n56983_,
    new_n56984_, new_n56985_, new_n56986_, new_n56987_, new_n56988_,
    new_n56989_, new_n56990_, new_n56991_, new_n56992_, new_n56993_,
    new_n56994_, new_n56995_, new_n56996_, new_n56997_, new_n56998_,
    new_n56999_, new_n57000_, new_n57001_, new_n57002_, new_n57003_,
    new_n57004_, new_n57005_, new_n57006_, new_n57007_, new_n57008_,
    new_n57009_, new_n57010_, new_n57011_, new_n57012_, new_n57013_,
    new_n57014_, new_n57015_, new_n57016_, new_n57017_, new_n57018_,
    new_n57019_, new_n57020_, new_n57021_, new_n57022_, new_n57023_,
    new_n57024_, new_n57025_, new_n57026_, new_n57027_, new_n57028_,
    new_n57029_, new_n57030_, new_n57031_, new_n57033_, new_n57034_,
    new_n57035_, new_n57036_, new_n57037_, new_n57038_, new_n57039_,
    new_n57040_, new_n57041_, new_n57043_, new_n57044_, new_n57045_,
    new_n57046_, new_n57047_, new_n57048_, new_n57049_, new_n57050_,
    new_n57051_, new_n57052_, new_n57053_, new_n57054_, new_n57055_,
    new_n57056_, new_n57057_, new_n57058_, new_n57059_, new_n57060_,
    new_n57061_, new_n57062_, new_n57063_, new_n57064_, new_n57065_,
    new_n57066_, new_n57067_, new_n57068_, new_n57069_, new_n57070_,
    new_n57071_, new_n57072_, new_n57073_, new_n57074_, new_n57075_,
    new_n57076_, new_n57077_, new_n57078_, new_n57079_, new_n57080_,
    new_n57081_, new_n57082_, new_n57083_, new_n57084_, new_n57085_,
    new_n57086_, new_n57087_, new_n57088_, new_n57089_, new_n57090_,
    new_n57091_, new_n57092_, new_n57093_, new_n57094_, new_n57095_,
    new_n57096_, new_n57097_, new_n57098_, new_n57099_, new_n57100_,
    new_n57101_, new_n57102_, new_n57103_, new_n57104_, new_n57105_,
    new_n57106_, new_n57107_, new_n57108_, new_n57109_, new_n57110_,
    new_n57111_, new_n57112_, new_n57113_, new_n57114_, new_n57115_,
    new_n57116_, new_n57117_, new_n57118_, new_n57119_, new_n57120_,
    new_n57121_, new_n57122_, new_n57123_, new_n57124_, new_n57125_,
    new_n57126_, new_n57127_, new_n57128_, new_n57129_, new_n57130_,
    new_n57131_, new_n57132_, new_n57133_, new_n57134_, new_n57135_,
    new_n57136_, new_n57137_, new_n57138_, new_n57139_, new_n57140_,
    new_n57141_, new_n57142_, new_n57143_, new_n57144_, new_n57145_,
    new_n57146_, new_n57147_, new_n57148_, new_n57149_, new_n57150_,
    new_n57151_, new_n57152_, new_n57153_, new_n57154_, new_n57155_,
    new_n57156_, new_n57157_, new_n57158_, new_n57159_, new_n57160_,
    new_n57161_, new_n57162_, new_n57163_, new_n57164_, new_n57165_,
    new_n57166_, new_n57167_, new_n57168_, new_n57169_, new_n57170_,
    new_n57171_, new_n57172_, new_n57173_, new_n57175_, new_n57176_,
    new_n57177_, new_n57178_, new_n57179_, new_n57180_, new_n57181_,
    new_n57182_, new_n57183_, new_n57185_, new_n57186_, new_n57187_,
    new_n57188_, new_n57189_, new_n57190_, new_n57191_, new_n57192_,
    new_n57193_, new_n57194_, new_n57195_, new_n57196_, new_n57197_,
    new_n57198_, new_n57199_, new_n57200_, new_n57201_, new_n57202_,
    new_n57203_, new_n57204_, new_n57205_, new_n57206_, new_n57207_,
    new_n57208_, new_n57209_, new_n57210_, new_n57211_, new_n57212_,
    new_n57213_, new_n57214_, new_n57215_, new_n57216_, new_n57217_,
    new_n57218_, new_n57219_, new_n57220_, new_n57221_, new_n57222_,
    new_n57223_, new_n57224_, new_n57225_, new_n57226_, new_n57227_,
    new_n57228_, new_n57229_, new_n57230_, new_n57231_, new_n57232_,
    new_n57233_, new_n57234_, new_n57235_, new_n57236_, new_n57237_,
    new_n57238_, new_n57239_, new_n57240_, new_n57241_, new_n57242_,
    new_n57243_, new_n57244_, new_n57245_, new_n57246_, new_n57247_,
    new_n57248_, new_n57249_, new_n57250_, new_n57251_, new_n57252_,
    new_n57253_, new_n57254_, new_n57255_, new_n57256_, new_n57257_,
    new_n57258_, new_n57259_, new_n57260_, new_n57261_, new_n57262_,
    new_n57263_, new_n57264_, new_n57265_, new_n57266_, new_n57267_,
    new_n57268_, new_n57269_, new_n57270_, new_n57271_, new_n57272_,
    new_n57273_, new_n57274_, new_n57275_, new_n57276_, new_n57277_,
    new_n57278_, new_n57279_, new_n57280_, new_n57281_, new_n57282_,
    new_n57283_, new_n57284_, new_n57285_, new_n57286_, new_n57287_,
    new_n57288_, new_n57289_, new_n57290_, new_n57291_, new_n57292_,
    new_n57293_, new_n57294_, new_n57295_, new_n57296_, new_n57297_,
    new_n57298_, new_n57299_, new_n57300_, new_n57301_, new_n57302_,
    new_n57303_, new_n57304_, new_n57305_, new_n57306_, new_n57307_,
    new_n57308_, new_n57309_, new_n57310_, new_n57311_, new_n57312_,
    new_n57313_, new_n57314_, new_n57315_, new_n57317_, new_n57318_,
    new_n57319_, new_n57320_, new_n57321_, new_n57322_, new_n57323_,
    new_n57324_, new_n57325_, new_n57327_, new_n57328_, new_n57329_,
    new_n57330_, new_n57331_, new_n57332_, new_n57333_, new_n57334_,
    new_n57335_, new_n57336_, new_n57337_, new_n57338_, new_n57339_,
    new_n57340_, new_n57341_, new_n57342_, new_n57343_, new_n57344_,
    new_n57345_, new_n57346_, new_n57347_, new_n57348_, new_n57349_,
    new_n57350_, new_n57351_, new_n57352_, new_n57353_, new_n57354_,
    new_n57355_, new_n57356_, new_n57357_, new_n57358_, new_n57359_,
    new_n57360_, new_n57361_, new_n57362_, new_n57363_, new_n57364_,
    new_n57365_, new_n57366_, new_n57367_, new_n57368_, new_n57369_,
    new_n57370_, new_n57371_, new_n57372_, new_n57373_, new_n57374_,
    new_n57375_, new_n57376_, new_n57377_, new_n57378_, new_n57379_,
    new_n57380_, new_n57381_, new_n57382_, new_n57383_, new_n57384_,
    new_n57385_, new_n57386_, new_n57387_, new_n57388_, new_n57389_,
    new_n57390_, new_n57391_, new_n57392_, new_n57393_, new_n57394_,
    new_n57395_, new_n57396_, new_n57397_, new_n57398_, new_n57399_,
    new_n57400_, new_n57401_, new_n57402_, new_n57403_, new_n57404_,
    new_n57405_, new_n57406_, new_n57407_, new_n57408_, new_n57409_,
    new_n57410_, new_n57411_, new_n57412_, new_n57413_, new_n57414_,
    new_n57415_, new_n57416_, new_n57417_, new_n57418_, new_n57419_,
    new_n57420_, new_n57421_, new_n57422_, new_n57423_, new_n57424_,
    new_n57425_, new_n57426_, new_n57427_, new_n57428_, new_n57429_,
    new_n57430_, new_n57431_, new_n57432_, new_n57433_, new_n57434_,
    new_n57435_, new_n57436_, new_n57437_, new_n57438_, new_n57439_,
    new_n57440_, new_n57441_, new_n57442_, new_n57443_, new_n57444_,
    new_n57445_, new_n57446_, new_n57447_, new_n57448_, new_n57449_,
    new_n57450_, new_n57451_, new_n57452_, new_n57453_, new_n57454_,
    new_n57455_, new_n57456_, new_n57457_, new_n57459_, new_n57460_,
    new_n57461_, new_n57462_, new_n57463_, new_n57464_, new_n57465_,
    new_n57466_, new_n57467_, new_n57469_, new_n57470_, new_n57471_,
    new_n57472_, new_n57473_, new_n57474_, new_n57475_, new_n57476_,
    new_n57477_, new_n57478_, new_n57479_, new_n57480_, new_n57481_,
    new_n57482_, new_n57483_, new_n57484_, new_n57485_, new_n57486_,
    new_n57487_, new_n57488_, new_n57489_, new_n57490_, new_n57491_,
    new_n57492_, new_n57493_, new_n57494_, new_n57495_, new_n57496_,
    new_n57497_, new_n57498_, new_n57499_, new_n57500_, new_n57501_,
    new_n57502_, new_n57503_, new_n57504_, new_n57505_, new_n57506_,
    new_n57507_, new_n57508_, new_n57509_, new_n57510_, new_n57511_,
    new_n57512_, new_n57513_, new_n57514_, new_n57515_, new_n57516_,
    new_n57517_, new_n57518_, new_n57519_, new_n57520_, new_n57521_,
    new_n57522_, new_n57523_, new_n57524_, new_n57525_, new_n57526_,
    new_n57527_, new_n57528_, new_n57529_, new_n57530_, new_n57531_,
    new_n57532_, new_n57533_, new_n57534_, new_n57535_, new_n57536_,
    new_n57537_, new_n57538_, new_n57539_, new_n57540_, new_n57541_,
    new_n57542_, new_n57543_, new_n57544_, new_n57545_, new_n57546_,
    new_n57547_, new_n57548_, new_n57549_, new_n57550_, new_n57551_,
    new_n57552_, new_n57553_, new_n57554_, new_n57555_, new_n57556_,
    new_n57557_, new_n57558_, new_n57559_, new_n57560_, new_n57561_,
    new_n57562_, new_n57563_, new_n57564_, new_n57565_, new_n57566_,
    new_n57567_, new_n57568_, new_n57569_, new_n57570_, new_n57571_,
    new_n57572_, new_n57573_, new_n57574_, new_n57575_, new_n57576_,
    new_n57577_, new_n57578_, new_n57579_, new_n57580_, new_n57581_,
    new_n57582_, new_n57583_, new_n57584_, new_n57585_, new_n57586_,
    new_n57587_, new_n57588_, new_n57589_, new_n57590_, new_n57591_,
    new_n57592_, new_n57593_, new_n57594_, new_n57595_, new_n57596_,
    new_n57597_, new_n57598_, new_n57599_, new_n57601_, new_n57602_,
    new_n57603_, new_n57604_, new_n57605_, new_n57606_, new_n57607_,
    new_n57608_, new_n57609_, new_n57611_, new_n57612_, new_n57613_,
    new_n57614_, new_n57615_, new_n57616_, new_n57617_, new_n57618_,
    new_n57619_, new_n57620_, new_n57621_, new_n57622_, new_n57623_,
    new_n57624_, new_n57625_, new_n57626_, new_n57627_, new_n57628_,
    new_n57629_, new_n57630_, new_n57631_, new_n57632_, new_n57633_,
    new_n57634_, new_n57635_, new_n57636_, new_n57637_, new_n57638_,
    new_n57639_, new_n57640_, new_n57641_, new_n57642_, new_n57643_,
    new_n57644_, new_n57645_, new_n57646_, new_n57647_, new_n57648_,
    new_n57649_, new_n57650_, new_n57651_, new_n57652_, new_n57653_,
    new_n57654_, new_n57655_, new_n57656_, new_n57657_, new_n57658_,
    new_n57659_, new_n57660_, new_n57661_, new_n57662_, new_n57663_,
    new_n57664_, new_n57665_, new_n57666_, new_n57667_, new_n57668_,
    new_n57669_, new_n57670_, new_n57671_, new_n57672_, new_n57673_,
    new_n57674_, new_n57675_, new_n57676_, new_n57677_, new_n57678_,
    new_n57679_, new_n57680_, new_n57681_, new_n57682_, new_n57683_,
    new_n57684_, new_n57685_, new_n57686_, new_n57687_, new_n57688_,
    new_n57689_, new_n57690_, new_n57691_, new_n57692_, new_n57693_,
    new_n57694_, new_n57695_, new_n57696_, new_n57697_, new_n57698_,
    new_n57699_, new_n57700_, new_n57701_, new_n57702_, new_n57703_,
    new_n57704_, new_n57705_, new_n57706_, new_n57707_, new_n57708_,
    new_n57709_, new_n57710_, new_n57711_, new_n57712_, new_n57713_,
    new_n57714_, new_n57715_, new_n57716_, new_n57717_, new_n57718_,
    new_n57719_, new_n57720_, new_n57721_, new_n57722_, new_n57723_,
    new_n57724_, new_n57725_, new_n57726_, new_n57727_, new_n57728_,
    new_n57729_, new_n57730_, new_n57731_, new_n57732_, new_n57733_,
    new_n57734_, new_n57735_, new_n57736_, new_n57737_, new_n57738_,
    new_n57739_, new_n57740_, new_n57741_, new_n57743_, new_n57744_,
    new_n57745_, new_n57746_, new_n57747_, new_n57748_, new_n57749_,
    new_n57750_, new_n57751_, new_n57753_, new_n57754_, new_n57755_,
    new_n57756_, new_n57757_, new_n57758_, new_n57759_, new_n57760_,
    new_n57761_, new_n57762_, new_n57763_, new_n57764_, new_n57765_,
    new_n57766_, new_n57767_, new_n57768_, new_n57769_, new_n57770_,
    new_n57771_, new_n57772_, new_n57773_, new_n57774_, new_n57775_,
    new_n57776_, new_n57777_, new_n57778_, new_n57779_, new_n57780_,
    new_n57781_, new_n57782_, new_n57783_, new_n57784_, new_n57785_,
    new_n57786_, new_n57787_, new_n57788_, new_n57789_, new_n57790_,
    new_n57791_, new_n57792_, new_n57793_, new_n57794_, new_n57795_,
    new_n57796_, new_n57797_, new_n57798_, new_n57799_, new_n57800_,
    new_n57801_, new_n57802_, new_n57803_, new_n57804_, new_n57805_,
    new_n57806_, new_n57807_, new_n57808_, new_n57809_, new_n57810_,
    new_n57811_, new_n57812_, new_n57813_, new_n57814_, new_n57815_,
    new_n57816_, new_n57817_, new_n57818_, new_n57819_, new_n57820_,
    new_n57821_, new_n57822_, new_n57823_, new_n57824_, new_n57825_,
    new_n57826_, new_n57827_, new_n57828_, new_n57829_, new_n57830_,
    new_n57831_, new_n57832_, new_n57833_, new_n57834_, new_n57835_,
    new_n57836_, new_n57837_, new_n57838_, new_n57839_, new_n57840_,
    new_n57841_, new_n57842_, new_n57843_, new_n57844_, new_n57845_,
    new_n57846_, new_n57847_, new_n57848_, new_n57849_, new_n57850_,
    new_n57851_, new_n57852_, new_n57853_, new_n57854_, new_n57855_,
    new_n57856_, new_n57857_, new_n57858_, new_n57859_, new_n57860_,
    new_n57861_, new_n57862_, new_n57863_, new_n57864_, new_n57865_,
    new_n57866_, new_n57867_, new_n57868_, new_n57869_, new_n57870_,
    new_n57871_, new_n57872_, new_n57873_, new_n57874_, new_n57875_,
    new_n57876_, new_n57877_, new_n57878_, new_n57879_, new_n57881_,
    new_n57882_, new_n57883_, new_n57884_, new_n57885_, new_n57886_,
    new_n57887_, new_n57888_, new_n57889_, new_n57891_, new_n57892_,
    new_n57893_, new_n57894_, new_n57895_, new_n57896_, new_n57897_,
    new_n57898_, new_n57899_, new_n57900_, new_n57901_, new_n57902_,
    new_n57903_, new_n57904_, new_n57905_, new_n57906_, new_n57907_,
    new_n57908_, new_n57909_, new_n57910_, new_n57911_, new_n57912_,
    new_n57913_, new_n57914_, new_n57915_, new_n57916_, new_n57917_,
    new_n57918_, new_n57919_, new_n57920_, new_n57921_, new_n57922_,
    new_n57923_, new_n57924_, new_n57925_, new_n57926_, new_n57927_,
    new_n57928_, new_n57929_, new_n57930_, new_n57931_, new_n57932_,
    new_n57933_, new_n57934_, new_n57935_, new_n57936_, new_n57937_,
    new_n57938_, new_n57939_, new_n57940_, new_n57941_, new_n57942_,
    new_n57943_, new_n57944_, new_n57945_, new_n57946_, new_n57947_,
    new_n57948_, new_n57949_, new_n57950_, new_n57951_, new_n57952_,
    new_n57953_, new_n57954_, new_n57955_, new_n57956_, new_n57957_,
    new_n57958_, new_n57959_, new_n57960_, new_n57961_, new_n57962_,
    new_n57963_, new_n57964_, new_n57965_, new_n57966_, new_n57967_,
    new_n57968_, new_n57969_, new_n57970_, new_n57971_, new_n57972_,
    new_n57973_, new_n57974_, new_n57975_, new_n57976_, new_n57977_,
    new_n57978_, new_n57979_, new_n57980_, new_n57981_, new_n57982_,
    new_n57983_, new_n57984_, new_n57985_, new_n57986_, new_n57987_,
    new_n57988_, new_n57989_, new_n57990_, new_n57991_, new_n57992_,
    new_n57993_, new_n57994_, new_n57995_, new_n57996_, new_n57997_,
    new_n57998_, new_n57999_, new_n58000_, new_n58001_, new_n58002_,
    new_n58003_, new_n58004_, new_n58005_, new_n58006_, new_n58007_,
    new_n58008_, new_n58009_, new_n58010_, new_n58012_, new_n58013_,
    new_n58014_, new_n58015_, new_n58016_, new_n58017_, new_n58018_,
    new_n58019_, new_n58020_, new_n58022_, new_n58023_, new_n58024_,
    new_n58025_, new_n58026_, new_n58027_, new_n58028_, new_n58029_,
    new_n58030_, new_n58031_, new_n58032_, new_n58033_, new_n58034_,
    new_n58035_, new_n58036_, new_n58037_, new_n58038_, new_n58039_,
    new_n58040_, new_n58041_, new_n58042_, new_n58043_, new_n58044_,
    new_n58045_, new_n58046_, new_n58047_, new_n58048_, new_n58049_,
    new_n58050_, new_n58051_, new_n58052_, new_n58053_, new_n58054_,
    new_n58055_, new_n58056_, new_n58057_, new_n58058_, new_n58059_,
    new_n58060_, new_n58061_, new_n58062_, new_n58063_, new_n58064_,
    new_n58065_, new_n58066_, new_n58067_, new_n58068_, new_n58069_,
    new_n58070_, new_n58071_, new_n58072_, new_n58073_, new_n58074_,
    new_n58075_, new_n58076_, new_n58077_, new_n58078_, new_n58079_,
    new_n58080_, new_n58081_, new_n58082_, new_n58083_, new_n58084_,
    new_n58085_, new_n58086_, new_n58087_, new_n58088_, new_n58089_,
    new_n58090_, new_n58091_, new_n58092_, new_n58093_, new_n58094_,
    new_n58095_, new_n58096_, new_n58097_, new_n58098_, new_n58099_,
    new_n58100_, new_n58101_, new_n58102_, new_n58103_, new_n58104_,
    new_n58105_, new_n58106_, new_n58107_, new_n58108_, new_n58109_,
    new_n58110_, new_n58111_, new_n58112_, new_n58113_, new_n58114_,
    new_n58115_, new_n58116_, new_n58117_, new_n58118_, new_n58119_,
    new_n58120_, new_n58121_, new_n58122_, new_n58123_, new_n58124_,
    new_n58125_, new_n58126_, new_n58127_, new_n58128_, new_n58129_,
    new_n58130_, new_n58132_, new_n58133_, new_n58134_, new_n58135_,
    new_n58136_, new_n58137_, new_n58138_, new_n58139_, new_n58140_,
    new_n58142_, new_n58143_, new_n58144_, new_n58145_, new_n58146_,
    new_n58147_, new_n58148_, new_n58149_, new_n58150_, new_n58151_,
    new_n58152_, new_n58153_, new_n58154_, new_n58155_, new_n58156_,
    new_n58157_, new_n58158_, new_n58159_, new_n58160_, new_n58161_,
    new_n58162_, new_n58163_, new_n58164_, new_n58165_, new_n58166_,
    new_n58167_, new_n58168_, new_n58169_, new_n58170_, new_n58171_,
    new_n58172_, new_n58173_, new_n58174_, new_n58175_, new_n58176_,
    new_n58177_, new_n58178_, new_n58179_, new_n58180_, new_n58181_,
    new_n58182_, new_n58183_, new_n58184_, new_n58185_, new_n58186_,
    new_n58187_, new_n58188_, new_n58189_, new_n58190_, new_n58191_,
    new_n58192_, new_n58193_, new_n58194_, new_n58195_, new_n58196_,
    new_n58197_, new_n58198_, new_n58199_, new_n58200_, new_n58201_,
    new_n58202_, new_n58203_, new_n58204_, new_n58205_, new_n58206_,
    new_n58207_, new_n58208_, new_n58209_, new_n58210_, new_n58211_,
    new_n58212_, new_n58213_, new_n58214_, new_n58215_, new_n58216_,
    new_n58217_, new_n58218_, new_n58219_, new_n58220_, new_n58221_,
    new_n58222_, new_n58223_, new_n58224_, new_n58225_, new_n58226_,
    new_n58227_, new_n58228_, new_n58229_, new_n58230_, new_n58231_,
    new_n58232_, new_n58233_, new_n58234_, new_n58235_, new_n58236_,
    new_n58237_, new_n58238_, new_n58239_, new_n58240_, new_n58241_,
    new_n58242_, new_n58243_, new_n58244_, new_n58245_, new_n58246_,
    new_n58247_, new_n58248_, new_n58249_, new_n58250_, new_n58252_,
    new_n58253_, new_n58254_, new_n58255_, new_n58256_, new_n58257_,
    new_n58258_, new_n58259_, new_n58260_, new_n58262_, new_n58263_,
    new_n58264_, new_n58265_, new_n58266_, new_n58267_, new_n58268_,
    new_n58269_, new_n58270_, new_n58271_, new_n58272_, new_n58273_,
    new_n58274_, new_n58275_, new_n58276_, new_n58277_, new_n58278_,
    new_n58279_, new_n58280_, new_n58281_, new_n58282_, new_n58283_,
    new_n58284_, new_n58285_, new_n58286_, new_n58287_, new_n58288_,
    new_n58289_, new_n58290_, new_n58291_, new_n58292_, new_n58293_,
    new_n58294_, new_n58295_, new_n58296_, new_n58297_, new_n58298_,
    new_n58299_, new_n58300_, new_n58301_, new_n58302_, new_n58303_,
    new_n58304_, new_n58305_, new_n58306_, new_n58307_, new_n58308_,
    new_n58309_, new_n58310_, new_n58311_, new_n58312_, new_n58313_,
    new_n58314_, new_n58315_, new_n58316_, new_n58317_, new_n58318_,
    new_n58319_, new_n58320_, new_n58321_, new_n58322_, new_n58323_,
    new_n58324_, new_n58325_, new_n58326_, new_n58327_, new_n58328_,
    new_n58329_, new_n58330_, new_n58331_, new_n58332_, new_n58333_,
    new_n58334_, new_n58335_, new_n58336_, new_n58337_, new_n58338_,
    new_n58339_, new_n58340_, new_n58341_, new_n58342_, new_n58343_,
    new_n58344_, new_n58345_, new_n58346_, new_n58348_, new_n58349_,
    new_n58350_, new_n58351_, new_n58352_, new_n58353_, new_n58354_,
    new_n58355_, new_n58356_, new_n58358_, new_n58359_, new_n58360_,
    new_n58361_, new_n58362_, new_n58363_, new_n58364_, new_n58365_,
    new_n58366_, new_n58367_, new_n58368_, new_n58369_, new_n58370_,
    new_n58371_, new_n58372_, new_n58373_, new_n58374_, new_n58375_,
    new_n58376_, new_n58377_, new_n58378_, new_n58379_, new_n58380_,
    new_n58381_, new_n58382_, new_n58383_, new_n58384_, new_n58385_,
    new_n58386_, new_n58387_, new_n58388_, new_n58389_, new_n58390_,
    new_n58391_, new_n58392_, new_n58393_, new_n58394_, new_n58395_,
    new_n58396_, new_n58397_, new_n58398_, new_n58399_, new_n58400_,
    new_n58401_, new_n58402_, new_n58403_, new_n58404_, new_n58405_,
    new_n58406_, new_n58407_, new_n58408_, new_n58409_, new_n58410_,
    new_n58411_, new_n58412_, new_n58413_, new_n58414_, new_n58415_,
    new_n58416_, new_n58417_, new_n58418_, new_n58419_, new_n58420_,
    new_n58421_, new_n58422_, new_n58423_, new_n58424_, new_n58425_,
    new_n58426_, new_n58427_, new_n58428_, new_n58429_, new_n58430_,
    new_n58431_, new_n58432_, new_n58433_, new_n58434_, new_n58435_,
    new_n58436_, new_n58437_, new_n58438_, new_n58439_, new_n58440_,
    new_n58442_, new_n58443_, new_n58444_, new_n58445_, new_n58446_,
    new_n58447_, new_n58448_, new_n58449_, new_n58450_, new_n58452_,
    new_n58453_, new_n58454_, new_n58455_, new_n58456_, new_n58457_,
    new_n58458_, new_n58459_, new_n58460_, new_n58461_, new_n58462_,
    new_n58463_, new_n58464_, new_n58465_, new_n58466_, new_n58467_,
    new_n58468_, new_n58469_, new_n58470_, new_n58471_, new_n58472_,
    new_n58473_, new_n58474_, new_n58475_, new_n58476_, new_n58477_,
    new_n58478_, new_n58479_, new_n58480_, new_n58481_, new_n58482_,
    new_n58483_, new_n58484_, new_n58485_, new_n58486_, new_n58487_,
    new_n58488_, new_n58489_, new_n58490_, new_n58491_, new_n58492_,
    new_n58493_, new_n58494_, new_n58495_, new_n58496_, new_n58497_,
    new_n58498_, new_n58499_, new_n58500_, new_n58501_, new_n58502_,
    new_n58503_, new_n58504_, new_n58505_, new_n58506_, new_n58507_,
    new_n58508_, new_n58509_, new_n58510_, new_n58511_, new_n58512_,
    new_n58513_, new_n58514_, new_n58515_, new_n58516_, new_n58517_,
    new_n58518_, new_n58519_, new_n58520_, new_n58521_, new_n58522_,
    new_n58523_, new_n58524_, new_n58525_, new_n58526_, new_n58527_,
    new_n58528_, new_n58529_, new_n58530_, new_n58531_, new_n58532_,
    new_n58533_, new_n58534_, new_n58535_, new_n58536_, new_n58537_,
    new_n58538_, new_n58539_, new_n58540_, new_n58541_, new_n58542_,
    new_n58544_, new_n58545_, new_n58546_, new_n58547_, new_n58548_,
    new_n58549_, new_n58550_, new_n58551_, new_n58552_, new_n58554_,
    new_n58555_, new_n58556_, new_n58557_, new_n58558_, new_n58559_,
    new_n58560_, new_n58561_, new_n58562_, new_n58563_, new_n58564_,
    new_n58565_, new_n58566_, new_n58567_, new_n58568_, new_n58569_,
    new_n58570_, new_n58571_, new_n58572_, new_n58573_, new_n58574_,
    new_n58575_, new_n58576_, new_n58577_, new_n58578_, new_n58579_,
    new_n58580_, new_n58581_, new_n58582_, new_n58583_, new_n58584_,
    new_n58585_, new_n58586_, new_n58587_, new_n58588_, new_n58589_,
    new_n58590_, new_n58591_, new_n58592_, new_n58593_, new_n58594_,
    new_n58595_, new_n58596_, new_n58597_, new_n58598_, new_n58599_,
    new_n58600_, new_n58601_, new_n58602_, new_n58603_, new_n58604_,
    new_n58605_, new_n58606_, new_n58607_, new_n58608_, new_n58609_,
    new_n58610_, new_n58611_, new_n58612_, new_n58613_, new_n58614_,
    new_n58615_, new_n58616_, new_n58617_, new_n58618_, new_n58619_,
    new_n58620_, new_n58621_, new_n58622_, new_n58623_, new_n58624_,
    new_n58625_, new_n58626_, new_n58627_, new_n58628_, new_n58629_,
    new_n58630_, new_n58631_, new_n58633_, new_n58634_, new_n58635_,
    new_n58636_, new_n58637_, new_n58638_, new_n58639_, new_n58640_,
    new_n58641_, new_n58643_, new_n58644_, new_n58645_, new_n58646_,
    new_n58647_, new_n58648_, new_n58649_, new_n58650_, new_n58651_,
    new_n58652_, new_n58653_, new_n58654_, new_n58655_, new_n58657_,
    new_n58658_, new_n58660_, new_n58661_, new_n58662_, new_n58663_,
    new_n58664_, new_n58665_, new_n58666_, new_n58667_, new_n58668_,
    new_n58669_, new_n58670_, new_n58671_, new_n58672_, new_n58673_,
    new_n58674_, new_n58675_, new_n58676_, new_n58677_, new_n58678_,
    new_n58679_, new_n58680_, new_n58681_, new_n58682_, new_n58683_,
    new_n58684_, new_n58685_, new_n58686_, new_n58687_, new_n58688_,
    new_n58689_, new_n58690_, new_n58691_, new_n58692_, new_n58693_,
    new_n58694_, new_n58695_, new_n58696_, new_n58697_, new_n58698_,
    new_n58699_, new_n58700_, new_n58701_, new_n58702_, new_n58703_,
    new_n58704_, new_n58705_, new_n58706_, new_n58707_, new_n58708_,
    new_n58709_, new_n58710_, new_n58711_, new_n58712_, new_n58713_,
    new_n58714_, new_n58715_, new_n58717_, new_n58718_, new_n58720_,
    new_n58721_, new_n58722_, new_n58723_, new_n58724_, new_n58725_,
    new_n58726_, new_n58727_, new_n58728_, new_n58729_, new_n58730_,
    new_n58731_, new_n58732_, new_n58733_, new_n58734_, new_n58735_,
    new_n58736_, new_n58737_, new_n58738_, new_n58739_, new_n58740_,
    new_n58741_, new_n58742_, new_n58743_, new_n58744_, new_n58745_,
    new_n58746_, new_n58747_, new_n58748_, new_n58749_, new_n58750_,
    new_n58751_, new_n58752_, new_n58753_, new_n58754_, new_n58755_,
    new_n58756_, new_n58757_, new_n58758_, new_n58759_, new_n58760_,
    new_n58761_, new_n58762_, new_n58763_, new_n58764_, new_n58765_,
    new_n58766_, new_n58767_, new_n58768_, new_n58769_, new_n58770_,
    new_n58771_, new_n58772_, new_n58773_, new_n58774_, new_n58775_,
    new_n58776_, new_n58777_, new_n58778_, new_n58779_, new_n58780_,
    new_n58781_, new_n58782_, new_n58783_, new_n58784_, new_n58785_,
    new_n58786_, new_n58787_, new_n58788_, new_n58789_, new_n58790_,
    new_n58791_, new_n58792_, new_n58793_, new_n58794_, new_n58795_,
    new_n58796_, new_n58797_, new_n58798_, new_n58799_, new_n58800_,
    new_n58801_, new_n58802_, new_n58803_, new_n58804_, new_n58805_,
    new_n58806_, new_n58807_, new_n58809_, new_n58810_, new_n58811_,
    new_n58812_, new_n58813_, new_n58814_, new_n58815_, new_n58816_,
    new_n58817_, new_n58819_, new_n58820_, new_n58821_, new_n58822_,
    new_n58823_, new_n58824_, new_n58825_, new_n58826_, new_n58827_,
    new_n58828_, new_n58829_, new_n58830_, new_n58831_, new_n58833_,
    new_n58834_, new_n58836_, new_n58837_, new_n58838_, new_n58839_,
    new_n58840_, new_n58841_, new_n58842_, new_n58843_, new_n58844_,
    new_n58845_, new_n58846_, new_n58847_, new_n58848_, new_n58849_,
    new_n58850_, new_n58851_, new_n58852_, new_n58853_, new_n58854_,
    new_n58855_, new_n58856_, new_n58857_, new_n58858_, new_n58859_,
    new_n58860_, new_n58861_, new_n58862_, new_n58863_, new_n58864_,
    new_n58865_, new_n58867_, new_n58868_, new_n58870_, new_n58871_,
    new_n58872_, new_n58873_, new_n58874_, new_n58875_, new_n58876_,
    new_n58877_, new_n58878_, new_n58879_, new_n58880_, new_n58881_,
    new_n58882_, new_n58883_, new_n58884_, new_n58885_, new_n58886_,
    new_n58887_, new_n58888_, new_n58889_, new_n58890_, new_n58891_,
    new_n58892_, new_n58893_, new_n58894_, new_n58895_, new_n58896_,
    new_n58897_, new_n58898_, new_n58899_, new_n58901_, new_n58902_,
    new_n58904_, new_n58905_, new_n58906_, new_n58907_, new_n58908_,
    new_n58909_, new_n58910_, new_n58911_, new_n58912_, new_n58914_,
    new_n58915_, new_n58916_, new_n58917_, new_n58918_, new_n58919_,
    new_n58920_, new_n58921_, new_n58922_, new_n58923_, new_n58924_,
    new_n58925_, new_n58926_, new_n58927_, new_n58928_, new_n58929_,
    new_n58930_, new_n58931_, new_n58932_, new_n58934_, new_n58935_,
    new_n58937_, new_n58938_, new_n58940_, new_n58941_, new_n58945_,
    new_n58946_, new_n58947_, new_n58948_, new_n58949_, new_n58952_,
    new_n58953_, new_n58954_, new_n58955_, new_n58956_, new_n58957_,
    new_n58958_, new_n58959_, new_n58960_, new_n58964_, new_n58965_,
    new_n58966_, new_n58967_, new_n58968_, new_n58969_, new_n58970_,
    new_n58971_, new_n58972_, new_n58973_, new_n58974_, new_n58975_,
    new_n58977_, new_n58978_, new_n58981_, new_n58982_, new_n58983_,
    new_n58984_, new_n58985_, new_n58987_, new_n58989_, new_n58990_,
    new_n58991_, new_n58992_, new_n58993_, new_n58994_, new_n58995_,
    new_n58996_, new_n58997_, new_n58998_, new_n58999_, new_n59000_,
    new_n59001_, new_n59002_, new_n59003_, new_n59004_, new_n59005_,
    new_n59006_, new_n59007_, new_n59008_, new_n59009_, new_n59010_,
    new_n59011_, new_n59012_, new_n59013_, new_n59014_, new_n59015_,
    new_n59016_, new_n59017_, new_n59018_, new_n59019_, new_n59020_,
    new_n59021_, new_n59022_, new_n59023_, new_n59024_, new_n59025_,
    new_n59026_, new_n59027_, new_n59028_, new_n59029_, new_n59030_,
    new_n59031_, new_n59032_, new_n59033_, new_n59034_, new_n59035_,
    new_n59036_, new_n59037_, new_n59038_, new_n59039_, new_n59040_,
    new_n59041_, new_n59042_, new_n59043_, new_n59044_, new_n59045_,
    new_n59046_, new_n59047_, new_n59048_, new_n59049_, new_n59050_,
    new_n59051_, new_n59052_, new_n59053_, new_n59054_, new_n59055_,
    new_n59056_, new_n59057_, new_n59058_, new_n59059_, new_n59060_,
    new_n59061_, new_n59062_, new_n59063_, new_n59064_, new_n59065_,
    new_n59066_, new_n59067_, new_n59068_, new_n59069_, new_n59070_,
    new_n59071_, new_n59072_, new_n59073_, new_n59074_, new_n59075_,
    new_n59076_, new_n59077_, new_n59078_, new_n59079_, new_n59080_,
    new_n59081_, new_n59082_, new_n59083_, new_n59087_, new_n59088_,
    new_n59089_, new_n59090_, new_n59091_, new_n59092_, new_n59094_,
    new_n59096_, new_n59097_, new_n59099_, new_n59101_, new_n59103_,
    new_n59105_, new_n59107_, new_n59108_, new_n59109_, new_n59110_,
    new_n59111_, new_n59113_, new_n59114_, new_n59115_, new_n59117_,
    new_n59119_, new_n59120_, new_n59121_, new_n59122_, new_n59123_,
    new_n59125_, new_n59126_, new_n59127_, new_n59128_, new_n59129_,
    new_n59131_, new_n59133_, new_n59134_, new_n59136_, new_n59137_,
    new_n59139_, new_n59140_, new_n59141_, new_n59142_, new_n59143_,
    new_n59145_, new_n59146_, new_n59147_, new_n59148_, new_n59150_,
    new_n59151_, new_n59153_, new_n59154_, new_n59156_, new_n59157_,
    new_n59158_, new_n59159_, new_n59160_, new_n59162_, new_n59163_,
    new_n59164_, new_n59165_, new_n59166_, new_n59168_, new_n59169_,
    new_n59171_, new_n59172_, new_n59174_, new_n59175_, new_n59176_,
    new_n59177_, new_n59178_, new_n59180_, new_n59181_, new_n59182_,
    new_n59183_, new_n59184_, new_n59186_, new_n59187_, new_n59189_,
    new_n59190_, new_n59192_, new_n59193_, new_n59194_, new_n59195_,
    new_n59196_, new_n59198_, new_n59199_, new_n59200_, new_n59201_,
    new_n59202_, new_n59204_, new_n59205_, new_n59207_, new_n59208_,
    new_n59211_, new_n59213_, new_n59214_, new_n59216_, new_n59217_,
    new_n59219_, new_n59220_, new_n59221_, new_n59223_, new_n59224_,
    new_n59226_, new_n59227_, new_n59228_, new_n59230_, new_n59231_,
    new_n59232_, new_n59234_, new_n59235_, new_n59237_, new_n59238_,
    new_n59239_, new_n59240_, new_n59242_, new_n59243_, new_n59245_,
    new_n59246_, new_n59247_, new_n59248_, new_n59250_, new_n59251_,
    new_n59252_, new_n59253_, new_n59255_, new_n59256_, new_n59257_,
    new_n59258_, new_n59260_, new_n59261_, new_n59263_, new_n59264_,
    new_n59265_, new_n59266_, new_n59268_, new_n59269_, new_n59270_,
    new_n59271_, new_n59273_, new_n59274_, new_n59275_, new_n59276_,
    new_n59278_, new_n59279_, new_n59280_, new_n59281_, new_n59283_,
    new_n59284_, new_n59285_, new_n59286_, new_n59288_, new_n59289_,
    new_n59290_, new_n59291_, new_n59293_, new_n59294_, new_n59295_,
    new_n59296_;
  assign new_n11532_ = ~ys__n35124 & ~ys__n35727;
  assign new_n11533_ = ys__n35124 & ys__n35727;
  assign new_n11534_ = ~new_n11532_ & ~new_n11533_;
  assign new_n11535_ = ~ys__n35122 & ~ys__n35725;
  assign new_n11536_ = ys__n35122 & ys__n35725;
  assign new_n11537_ = ~new_n11535_ & ~new_n11536_;
  assign new_n11538_ = ~new_n11534_ & ~new_n11537_;
  assign new_n11539_ = ~ys__n35120 & ~ys__n35723;
  assign new_n11540_ = ys__n35120 & ys__n35723;
  assign new_n11541_ = ~new_n11539_ & ~new_n11540_;
  assign new_n11542_ = ~ys__n35118 & ~ys__n35721;
  assign new_n11543_ = ys__n35118 & ys__n35721;
  assign new_n11544_ = ~new_n11542_ & ~new_n11543_;
  assign new_n11545_ = ~new_n11541_ & ~new_n11544_;
  assign new_n11546_ = new_n11538_ & new_n11545_;
  assign new_n11547_ = ~ys__n35116 & ~ys__n35719;
  assign new_n11548_ = ys__n35116 & ys__n35719;
  assign new_n11549_ = ~new_n11547_ & ~new_n11548_;
  assign new_n11550_ = ~ys__n35114 & ~ys__n35717;
  assign new_n11551_ = ys__n35114 & ys__n35717;
  assign new_n11552_ = ~new_n11550_ & ~new_n11551_;
  assign new_n11553_ = ~new_n11549_ & ~new_n11552_;
  assign new_n11554_ = ~ys__n24207 & ~ys__n35112;
  assign new_n11555_ = ys__n24207 & ys__n35112;
  assign new_n11556_ = ~new_n11554_ & ~new_n11555_;
  assign new_n11557_ = ~ys__n24205 & ~ys__n35110;
  assign new_n11558_ = ys__n24205 & ys__n35110;
  assign new_n11559_ = ~new_n11557_ & ~new_n11558_;
  assign new_n11560_ = ~new_n11556_ & ~new_n11559_;
  assign new_n11561_ = new_n11553_ & new_n11560_;
  assign new_n11562_ = ~ys__n24203 & ~ys__n35108;
  assign new_n11563_ = ys__n24203 & ys__n35108;
  assign new_n11564_ = ~new_n11562_ & ~new_n11563_;
  assign new_n11565_ = ~ys__n24201 & ~ys__n35106;
  assign new_n11566_ = ys__n24201 & ys__n35106;
  assign new_n11567_ = ~new_n11565_ & ~new_n11566_;
  assign new_n11568_ = ~new_n11564_ & ~new_n11567_;
  assign new_n11569_ = ys__n24199 & ~ys__n35104;
  assign new_n11570_ = ~ys__n24199 & ~ys__n35104;
  assign new_n11571_ = ys__n24199 & ys__n35104;
  assign new_n11572_ = ~new_n11570_ & ~new_n11571_;
  assign new_n11573_ = ys__n24197 & ~ys__n35102;
  assign new_n11574_ = ~ys__n24197 & ~ys__n35102;
  assign new_n11575_ = ys__n24197 & ys__n35102;
  assign new_n11576_ = ~new_n11574_ & ~new_n11575_;
  assign new_n11577_ = ~new_n11573_ & new_n11576_;
  assign new_n11578_ = ~new_n11572_ & ~new_n11577_;
  assign new_n11579_ = ~new_n11569_ & ~new_n11578_;
  assign new_n11580_ = new_n11568_ & ~new_n11579_;
  assign new_n11581_ = ys__n24203 & ~ys__n35108;
  assign new_n11582_ = ys__n24201 & ~ys__n35106;
  assign new_n11583_ = ~new_n11564_ & new_n11582_;
  assign new_n11584_ = ~new_n11581_ & ~new_n11583_;
  assign new_n11585_ = ~new_n11580_ & new_n11584_;
  assign new_n11586_ = new_n11561_ & ~new_n11585_;
  assign new_n11587_ = ys__n24207 & ~ys__n35112;
  assign new_n11588_ = ys__n24205 & ~ys__n35110;
  assign new_n11589_ = ~new_n11556_ & new_n11588_;
  assign new_n11590_ = ~new_n11587_ & ~new_n11589_;
  assign new_n11591_ = new_n11553_ & ~new_n11590_;
  assign new_n11592_ = ~ys__n35116 & ys__n35719;
  assign new_n11593_ = ~ys__n35114 & ys__n35717;
  assign new_n11594_ = ~new_n11549_ & new_n11593_;
  assign new_n11595_ = ~new_n11592_ & ~new_n11594_;
  assign new_n11596_ = ~new_n11591_ & new_n11595_;
  assign new_n11597_ = ~new_n11586_ & new_n11596_;
  assign new_n11598_ = new_n11546_ & ~new_n11597_;
  assign new_n11599_ = ~ys__n35120 & ys__n35723;
  assign new_n11600_ = ~ys__n35118 & ys__n35721;
  assign new_n11601_ = ~new_n11541_ & new_n11600_;
  assign new_n11602_ = ~new_n11599_ & ~new_n11601_;
  assign new_n11603_ = new_n11538_ & ~new_n11602_;
  assign new_n11604_ = ~ys__n35124 & ys__n35727;
  assign new_n11605_ = ~ys__n35122 & ys__n35725;
  assign new_n11606_ = ~new_n11534_ & new_n11605_;
  assign new_n11607_ = ~new_n11604_ & ~new_n11606_;
  assign new_n11608_ = ~new_n11603_ & new_n11607_;
  assign new_n11609_ = ~new_n11598_ & new_n11608_;
  assign new_n11610_ = ~new_n11572_ & ~new_n11576_;
  assign new_n11611_ = new_n11568_ & new_n11610_;
  assign new_n11612_ = new_n11546_ & new_n11611_;
  assign new_n11613_ = new_n11561_ & new_n11612_;
  assign new_n11614_ = ~new_n11609_ & ~new_n11613_;
  assign new_n11615_ = ~ys__n33265 & ~ys__n35723;
  assign new_n11616_ = ys__n33265 & ys__n35723;
  assign new_n11617_ = ~new_n11615_ & ~new_n11616_;
  assign new_n11618_ = ~ys__n33263 & ~ys__n35721;
  assign new_n11619_ = ys__n33263 & ys__n35721;
  assign new_n11620_ = ~new_n11618_ & ~new_n11619_;
  assign new_n11621_ = ~new_n11617_ & ~new_n11620_;
  assign new_n11622_ = ~ys__n33269 & ~ys__n35727;
  assign new_n11623_ = ys__n33269 & ys__n35727;
  assign new_n11624_ = ~new_n11622_ & ~new_n11623_;
  assign new_n11625_ = ~ys__n33267 & ~ys__n35725;
  assign new_n11626_ = ys__n33267 & ys__n35725;
  assign new_n11627_ = ~new_n11625_ & ~new_n11626_;
  assign new_n11628_ = ~new_n11624_ & ~new_n11627_;
  assign new_n11629_ = ~ys__n33261 & ~ys__n35719;
  assign new_n11630_ = ys__n33261 & ys__n35719;
  assign new_n11631_ = ~new_n11629_ & ~new_n11630_;
  assign new_n11632_ = ~ys__n33259 & ~ys__n35717;
  assign new_n11633_ = ys__n33259 & ys__n35717;
  assign new_n11634_ = ~new_n11632_ & ~new_n11633_;
  assign new_n11635_ = ~new_n11631_ & ~new_n11634_;
  assign new_n11636_ = new_n11628_ & new_n11635_;
  assign new_n11637_ = new_n11621_ & new_n11636_;
  assign new_n11638_ = ~ys__n33261 & ys__n35719;
  assign new_n11639_ = ~ys__n33259 & ys__n35717;
  assign new_n11640_ = new_n11634_ & ~new_n11639_;
  assign new_n11641_ = ~new_n11631_ & ~new_n11640_;
  assign new_n11642_ = ~new_n11638_ & ~new_n11641_;
  assign new_n11643_ = new_n11621_ & ~new_n11642_;
  assign new_n11644_ = ~ys__n33265 & ys__n35723;
  assign new_n11645_ = ~ys__n33263 & ys__n35721;
  assign new_n11646_ = ~new_n11617_ & new_n11645_;
  assign new_n11647_ = ~new_n11644_ & ~new_n11646_;
  assign new_n11648_ = ~new_n11643_ & new_n11647_;
  assign new_n11649_ = new_n11628_ & ~new_n11648_;
  assign new_n11650_ = ~ys__n33269 & ys__n35727;
  assign new_n11651_ = ~ys__n33267 & ys__n35725;
  assign new_n11652_ = ~new_n11624_ & new_n11651_;
  assign new_n11653_ = ~new_n11650_ & ~new_n11652_;
  assign new_n11654_ = ~new_n11649_ & new_n11653_;
  assign new_n11655_ = ~new_n11637_ & ~new_n11654_;
  assign new_n11656_ = ~new_n11637_ & ~new_n11655_;
  assign new_n11657_ = ys__n128 & ~ys__n38605;
  assign new_n11658_ = ~ys__n38606 & ys__n38607;
  assign new_n11659_ = ~new_n11657_ & ~new_n11658_;
  assign new_n11660_ = ys__n38606 & ~ys__n38607;
  assign new_n11661_ = ~ys__n38608 & ys__n38609;
  assign new_n11662_ = ~new_n11660_ & ~new_n11661_;
  assign new_n11663_ = new_n11659_ & new_n11662_;
  assign new_n11664_ = ys__n132 & ~ys__n38603;
  assign new_n11665_ = ~ys__n130 & ys__n38604;
  assign new_n11666_ = ~new_n11664_ & ~new_n11665_;
  assign new_n11667_ = ys__n130 & ~ys__n38604;
  assign new_n11668_ = ~ys__n128 & ys__n38605;
  assign new_n11669_ = ~new_n11667_ & ~new_n11668_;
  assign new_n11670_ = new_n11666_ & new_n11669_;
  assign new_n11671_ = new_n11663_ & new_n11670_;
  assign new_n11672_ = ys__n130 & ys__n132;
  assign new_n11673_ = ys__n134 & ys__n136;
  assign new_n11674_ = new_n11672_ & new_n11673_;
  assign new_n11675_ = ys__n122 & ys__n124;
  assign new_n11676_ = ys__n126 & ys__n128;
  assign new_n11677_ = new_n11675_ & new_n11676_;
  assign new_n11678_ = new_n11674_ & new_n11677_;
  assign new_n11679_ = ys__n38610 & ~ys__n38611;
  assign new_n11680_ = ys__n38608 & ~ys__n38609;
  assign new_n11681_ = ~ys__n38610 & ys__n38611;
  assign new_n11682_ = ~new_n11680_ & ~new_n11681_;
  assign new_n11683_ = ~new_n11679_ & new_n11682_;
  assign new_n11684_ = ~new_n11678_ & new_n11683_;
  assign new_n11685_ = new_n11671_ & new_n11684_;
  assign new_n11686_ = ~ys__n38585 & ys__n38586;
  assign new_n11687_ = ~ys__n38557 & ~new_n11686_;
  assign new_n11688_ = ys__n38585 & ~ys__n38586;
  assign new_n11689_ = ~ys__n38587 & ys__n38588;
  assign new_n11690_ = ~new_n11688_ & ~new_n11689_;
  assign new_n11691_ = ys__n38587 & ~ys__n38588;
  assign new_n11692_ = ~ys__n38589 & ys__n38590;
  assign new_n11693_ = ~new_n11691_ & ~new_n11692_;
  assign new_n11694_ = new_n11690_ & new_n11693_;
  assign new_n11695_ = new_n11687_ & new_n11694_;
  assign new_n11696_ = ys__n38593 & ~ys__n38594;
  assign new_n11697_ = ~ys__n38595 & ys__n38596;
  assign new_n11698_ = ~new_n11696_ & ~new_n11697_;
  assign new_n11699_ = ys__n38595 & ~ys__n38596;
  assign new_n11700_ = ~ys__n38597 & ys__n38598;
  assign new_n11701_ = ~new_n11699_ & ~new_n11700_;
  assign new_n11702_ = new_n11698_ & new_n11701_;
  assign new_n11703_ = ys__n38589 & ~ys__n38590;
  assign new_n11704_ = ~ys__n38591 & ys__n38592;
  assign new_n11705_ = ~new_n11703_ & ~new_n11704_;
  assign new_n11706_ = ys__n38591 & ~ys__n38592;
  assign new_n11707_ = ~ys__n38593 & ys__n38594;
  assign new_n11708_ = ~new_n11706_ & ~new_n11707_;
  assign new_n11709_ = new_n11705_ & new_n11708_;
  assign new_n11710_ = new_n11702_ & new_n11709_;
  assign new_n11711_ = ys__n136 & ~ys__n38601;
  assign new_n11712_ = ~ys__n134 & ys__n38602;
  assign new_n11713_ = ~new_n11711_ & ~new_n11712_;
  assign new_n11714_ = ys__n134 & ~ys__n38602;
  assign new_n11715_ = ~ys__n132 & ys__n38603;
  assign new_n11716_ = ~new_n11714_ & ~new_n11715_;
  assign new_n11717_ = new_n11713_ & new_n11716_;
  assign new_n11718_ = ys__n38597 & ~ys__n38598;
  assign new_n11719_ = ~ys__n38599 & ys__n38600;
  assign new_n11720_ = ~new_n11718_ & ~new_n11719_;
  assign new_n11721_ = ys__n38599 & ~ys__n38600;
  assign new_n11722_ = ~ys__n136 & ys__n38601;
  assign new_n11723_ = ~new_n11721_ & ~new_n11722_;
  assign new_n11724_ = new_n11720_ & new_n11723_;
  assign new_n11725_ = new_n11717_ & new_n11724_;
  assign new_n11726_ = new_n11710_ & new_n11725_;
  assign new_n11727_ = new_n11695_ & new_n11726_;
  assign new_n11728_ = new_n11685_ & new_n11727_;
  assign new_n11729_ = ~new_n11656_ & new_n11728_;
  assign new_n11730_ = ~new_n11614_ & new_n11729_;
  assign new_n11731_ = ys__n1072 & new_n11730_;
  assign new_n11732_ = ~ys__n4613 & ~new_n11731_;
  assign new_n11733_ = ~ys__n4185 & ~new_n11732_;
  assign new_n11734_ = ys__n1029 & ~ys__n24131;
  assign new_n11735_ = ~new_n11733_ & new_n11734_;
  assign new_n11736_ = ys__n1072 & ~ys__n4185;
  assign new_n11737_ = new_n11730_ & new_n11736_;
  assign new_n11738_ = ys__n29897 & ~new_n11737_;
  assign new_n11739_ = ~new_n11735_ & new_n11738_;
  assign ys__n4192 = ys__n4185 | ys__n4613;
  assign new_n11741_ = ~ys__n4184 & ~ys__n4190;
  assign new_n11742_ = ~ys__n4192 & new_n11741_;
  assign new_n11743_ = ~ys__n4625 & ~ys__n4627;
  assign new_n11744_ = ~ys__n4176 & ~ys__n4698;
  assign new_n11745_ = new_n11743_ & new_n11744_;
  assign new_n11746_ = new_n11742_ & new_n11745_;
  assign new_n11747_ = ~ys__n846 & ~ys__n4177;
  assign ys__n738 = ~new_n11746_ | ~new_n11747_;
  assign new_n11749_ = ys__n23339 & ~ys__n738;
  assign new_n11750_ = ys__n23763 & ys__n738;
  assign ys__n23764 = new_n11749_ | new_n11750_;
  assign new_n11752_ = new_n11739_ & ~ys__n23764;
  assign new_n11753_ = ys__n29913 & ~new_n11737_;
  assign new_n11754_ = ~new_n11735_ & new_n11753_;
  assign new_n11755_ = ys__n22464 & ~ys__n738;
  assign new_n11756_ = ys__n22465 & ys__n738;
  assign ys__n22466 = new_n11755_ | new_n11756_;
  assign new_n11758_ = new_n11754_ & ~ys__n22466;
  assign new_n11759_ = new_n11739_ & ys__n22466;
  assign new_n11760_ = ~new_n11758_ & ~new_n11759_;
  assign new_n11761_ = ys__n23764 & ~new_n11760_;
  assign new_n11762_ = ~new_n11752_ & ~new_n11761_;
  assign new_n11763_ = ~ys__n532 & ~ys__n746;
  assign new_n11764_ = ys__n742 & ys__n744;
  assign new_n11765_ = new_n11763_ & new_n11764_;
  assign new_n11766_ = ~ys__n748 & ~ys__n750;
  assign new_n11767_ = new_n11765_ & new_n11766_;
  assign new_n11768_ = ys__n518 & ~ys__n548;
  assign new_n11769_ = ~ys__n550 & new_n11768_;
  assign new_n11770_ = ~ys__n518 & ~ys__n548;
  assign new_n11771_ = ~ys__n550 & new_n11770_;
  assign new_n11772_ = ~new_n11769_ & ~new_n11771_;
  assign new_n11773_ = ~ys__n23730 & ~new_n11772_;
  assign new_n11774_ = new_n11767_ & new_n11773_;
  assign new_n11775_ = ~ys__n742 & ys__n744;
  assign new_n11776_ = new_n11763_ & new_n11775_;
  assign new_n11777_ = new_n11766_ & new_n11776_;
  assign new_n11778_ = ys__n532 & ~ys__n746;
  assign new_n11779_ = new_n11775_ & new_n11778_;
  assign new_n11780_ = new_n11766_ & new_n11779_;
  assign new_n11781_ = ~new_n11777_ & ~new_n11780_;
  assign new_n11782_ = ~ys__n532 & ys__n746;
  assign new_n11783_ = ~ys__n742 & ~ys__n744;
  assign new_n11784_ = new_n11782_ & new_n11783_;
  assign new_n11785_ = new_n11766_ & new_n11784_;
  assign new_n11786_ = new_n11781_ & ~new_n11785_;
  assign new_n11787_ = ~ys__n23730 & ~new_n11786_;
  assign new_n11788_ = ~new_n11774_ & ~new_n11787_;
  assign new_n11789_ = ~new_n11767_ & new_n11786_;
  assign new_n11790_ = ~new_n11788_ & ~new_n11789_;
  assign new_n11791_ = new_n11763_ & new_n11783_;
  assign new_n11792_ = ys__n748 & ~ys__n750;
  assign new_n11793_ = new_n11791_ & new_n11792_;
  assign new_n11794_ = new_n11776_ & new_n11792_;
  assign new_n11795_ = ~new_n11793_ & ~new_n11794_;
  assign new_n11796_ = new_n11778_ & new_n11783_;
  assign new_n11797_ = new_n11792_ & new_n11796_;
  assign new_n11798_ = new_n11779_ & new_n11792_;
  assign new_n11799_ = ~new_n11797_ & ~new_n11798_;
  assign new_n11800_ = new_n11795_ & new_n11799_;
  assign new_n11801_ = ys__n532 & ys__n746;
  assign new_n11802_ = new_n11783_ & new_n11801_;
  assign new_n11803_ = new_n11792_ & new_n11802_;
  assign new_n11804_ = new_n11784_ & new_n11792_;
  assign new_n11805_ = ~new_n11803_ & ~new_n11804_;
  assign new_n11806_ = new_n11775_ & new_n11782_;
  assign new_n11807_ = new_n11792_ & new_n11806_;
  assign new_n11808_ = new_n11805_ & ~new_n11807_;
  assign new_n11809_ = new_n11800_ & new_n11808_;
  assign new_n11810_ = ~ys__n23730 & ~new_n11809_;
  assign new_n11811_ = ~new_n11790_ & ~new_n11810_;
  assign new_n11812_ = ys__n28243 & ~new_n11811_;
  assign new_n11813_ = ys__n23332 & ys__n38438;
  assign new_n11814_ = ~ys__n23332 & ys__n38449;
  assign new_n11815_ = ys__n23332 & ys__n38448;
  assign new_n11816_ = ~new_n11814_ & ~new_n11815_;
  assign new_n11817_ = ~new_n11813_ & new_n11816_;
  assign new_n11818_ = ~ys__n38437 & ~ys__n38438;
  assign new_n11819_ = new_n11817_ & new_n11818_;
  assign new_n11820_ = ys__n23627 & ~new_n11819_;
  assign new_n11821_ = ~ys__n23310 & ys__n28019;
  assign new_n11822_ = ys__n23310 & ~ys__n28019;
  assign new_n11823_ = ~new_n11821_ & ~new_n11822_;
  assign new_n11824_ = ~ys__n23312 & ys__n28020;
  assign new_n11825_ = ys__n23312 & ~ys__n28020;
  assign new_n11826_ = ~new_n11824_ & ~new_n11825_;
  assign new_n11827_ = new_n11823_ & new_n11826_;
  assign new_n11828_ = ~ys__n23314 & ys__n28021;
  assign new_n11829_ = ys__n23314 & ~ys__n28021;
  assign new_n11830_ = ~new_n11828_ & ~new_n11829_;
  assign new_n11831_ = ~ys__n23316 & ys__n28022;
  assign new_n11832_ = ys__n23316 & ~ys__n28022;
  assign new_n11833_ = ~new_n11831_ & ~new_n11832_;
  assign new_n11834_ = new_n11830_ & new_n11833_;
  assign new_n11835_ = new_n11827_ & new_n11834_;
  assign new_n11836_ = ~ys__n23302 & ys__n28015;
  assign new_n11837_ = ys__n23302 & ~ys__n28015;
  assign new_n11838_ = ~new_n11836_ & ~new_n11837_;
  assign new_n11839_ = ~ys__n23304 & ys__n28016;
  assign new_n11840_ = ys__n23304 & ~ys__n28016;
  assign new_n11841_ = ~new_n11839_ & ~new_n11840_;
  assign new_n11842_ = new_n11838_ & new_n11841_;
  assign new_n11843_ = ~ys__n23306 & ys__n28017;
  assign new_n11844_ = ys__n23306 & ~ys__n28017;
  assign new_n11845_ = ~new_n11843_ & ~new_n11844_;
  assign new_n11846_ = ~ys__n23308 & ys__n28018;
  assign new_n11847_ = ys__n23308 & ~ys__n28018;
  assign new_n11848_ = ~new_n11846_ & ~new_n11847_;
  assign new_n11849_ = new_n11845_ & new_n11848_;
  assign new_n11850_ = new_n11842_ & new_n11849_;
  assign new_n11851_ = new_n11835_ & new_n11850_;
  assign new_n11852_ = ~ys__n23326 & ys__n28027;
  assign new_n11853_ = ys__n23326 & ~ys__n28027;
  assign new_n11854_ = ~new_n11852_ & ~new_n11853_;
  assign new_n11855_ = ~ys__n23328 & ys__n28028;
  assign new_n11856_ = ys__n23328 & ~ys__n28028;
  assign new_n11857_ = ~new_n11855_ & ~new_n11856_;
  assign new_n11858_ = new_n11854_ & new_n11857_;
  assign new_n11859_ = ~ys__n23330 & ys__n28029;
  assign new_n11860_ = ys__n23330 & ~ys__n28029;
  assign new_n11861_ = ~new_n11859_ & ~new_n11860_;
  assign new_n11862_ = ~ys__n23332 & ys__n28030;
  assign new_n11863_ = ys__n23332 & ~ys__n28030;
  assign new_n11864_ = ~new_n11862_ & ~new_n11863_;
  assign new_n11865_ = new_n11861_ & new_n11864_;
  assign new_n11866_ = new_n11858_ & new_n11865_;
  assign new_n11867_ = ~ys__n23318 & ys__n28023;
  assign new_n11868_ = ys__n23318 & ~ys__n28023;
  assign new_n11869_ = ~new_n11867_ & ~new_n11868_;
  assign new_n11870_ = ~ys__n23320 & ys__n28024;
  assign new_n11871_ = ys__n23320 & ~ys__n28024;
  assign new_n11872_ = ~new_n11870_ & ~new_n11871_;
  assign new_n11873_ = new_n11869_ & new_n11872_;
  assign new_n11874_ = ~ys__n23322 & ys__n28025;
  assign new_n11875_ = ys__n23322 & ~ys__n28025;
  assign new_n11876_ = ~new_n11874_ & ~new_n11875_;
  assign new_n11877_ = ~ys__n23324 & ys__n28026;
  assign new_n11878_ = ys__n23324 & ~ys__n28026;
  assign new_n11879_ = ~new_n11877_ & ~new_n11878_;
  assign new_n11880_ = new_n11876_ & new_n11879_;
  assign new_n11881_ = new_n11873_ & new_n11880_;
  assign new_n11882_ = new_n11866_ & new_n11881_;
  assign new_n11883_ = new_n11851_ & new_n11882_;
  assign new_n11884_ = ~ys__n23278 & ys__n27863;
  assign new_n11885_ = ys__n23278 & ~ys__n27863;
  assign new_n11886_ = ~new_n11884_ & ~new_n11885_;
  assign new_n11887_ = ~ys__n23280 & ys__n27865;
  assign new_n11888_ = ys__n23280 & ~ys__n27865;
  assign new_n11889_ = ~new_n11887_ & ~new_n11888_;
  assign new_n11890_ = new_n11886_ & new_n11889_;
  assign new_n11891_ = ~ys__n23282 & ys__n27867;
  assign new_n11892_ = ys__n23282 & ~ys__n27867;
  assign new_n11893_ = ~new_n11891_ & ~new_n11892_;
  assign new_n11894_ = ~ys__n23284 & ys__n27869;
  assign new_n11895_ = ys__n23284 & ~ys__n27869;
  assign new_n11896_ = ~new_n11894_ & ~new_n11895_;
  assign new_n11897_ = new_n11893_ & new_n11896_;
  assign new_n11898_ = new_n11890_ & new_n11897_;
  assign new_n11899_ = ~ys__n23335 & ys__n27855;
  assign new_n11900_ = ys__n23335 & ~ys__n27855;
  assign new_n11901_ = ~new_n11899_ & ~new_n11900_;
  assign new_n11902_ = ~ys__n23272 & ys__n27857;
  assign new_n11903_ = ys__n23272 & ~ys__n27857;
  assign new_n11904_ = ~new_n11902_ & ~new_n11903_;
  assign new_n11905_ = new_n11901_ & new_n11904_;
  assign new_n11906_ = ~ys__n23274 & ys__n27859;
  assign new_n11907_ = ys__n23274 & ~ys__n27859;
  assign new_n11908_ = ~new_n11906_ & ~new_n11907_;
  assign new_n11909_ = ~ys__n23276 & ys__n27861;
  assign new_n11910_ = ys__n23276 & ~ys__n27861;
  assign new_n11911_ = ~new_n11909_ & ~new_n11910_;
  assign new_n11912_ = new_n11908_ & new_n11911_;
  assign new_n11913_ = new_n11905_ & new_n11912_;
  assign new_n11914_ = new_n11898_ & new_n11913_;
  assign new_n11915_ = ~ys__n23294 & ys__n27879;
  assign new_n11916_ = ys__n23294 & ~ys__n27879;
  assign new_n11917_ = ~new_n11915_ & ~new_n11916_;
  assign new_n11918_ = ~ys__n23296 & ys__n27881;
  assign new_n11919_ = ys__n23296 & ~ys__n27881;
  assign new_n11920_ = ~new_n11918_ & ~new_n11919_;
  assign new_n11921_ = new_n11917_ & new_n11920_;
  assign new_n11922_ = ~ys__n23298 & ys__n27883;
  assign new_n11923_ = ys__n23298 & ~ys__n27883;
  assign new_n11924_ = ~new_n11922_ & ~new_n11923_;
  assign new_n11925_ = ~ys__n23300 & ys__n27885;
  assign new_n11926_ = ys__n23300 & ~ys__n27885;
  assign new_n11927_ = ~new_n11925_ & ~new_n11926_;
  assign new_n11928_ = new_n11924_ & new_n11927_;
  assign new_n11929_ = new_n11921_ & new_n11928_;
  assign new_n11930_ = ~ys__n23286 & ys__n27871;
  assign new_n11931_ = ys__n23286 & ~ys__n27871;
  assign new_n11932_ = ~new_n11930_ & ~new_n11931_;
  assign new_n11933_ = ~ys__n23288 & ys__n27873;
  assign new_n11934_ = ys__n23288 & ~ys__n27873;
  assign new_n11935_ = ~new_n11933_ & ~new_n11934_;
  assign new_n11936_ = new_n11932_ & new_n11935_;
  assign new_n11937_ = ~ys__n23290 & ys__n27875;
  assign new_n11938_ = ys__n23290 & ~ys__n27875;
  assign new_n11939_ = ~new_n11937_ & ~new_n11938_;
  assign new_n11940_ = ~ys__n23292 & ys__n27877;
  assign new_n11941_ = ys__n23292 & ~ys__n27877;
  assign new_n11942_ = ~new_n11940_ & ~new_n11941_;
  assign new_n11943_ = new_n11939_ & new_n11942_;
  assign new_n11944_ = new_n11936_ & new_n11943_;
  assign new_n11945_ = new_n11929_ & new_n11944_;
  assign new_n11946_ = new_n11914_ & new_n11945_;
  assign new_n11947_ = new_n11883_ & new_n11946_;
  assign new_n11948_ = new_n11820_ & new_n11947_;
  assign new_n11949_ = ~ys__n23332 & ys__n38443;
  assign new_n11950_ = ~ys__n38441 & ~new_n11949_;
  assign new_n11951_ = new_n11817_ & new_n11950_;
  assign new_n11952_ = ys__n23627 & ~new_n11951_;
  assign new_n11953_ = ~new_n11947_ & new_n11952_;
  assign new_n11954_ = ~new_n11948_ & ~new_n11953_;
  assign new_n11955_ = ~ys__n23641 & ~ys__n23645;
  assign new_n11956_ = ~ys__n23652 & ~ys__n38413;
  assign new_n11957_ = new_n11955_ & new_n11956_;
  assign new_n11958_ = ys__n935 & ys__n33340;
  assign new_n11959_ = ~ys__n33380 & ~ys__n33384;
  assign new_n11960_ = ~ys__n33386 & new_n11959_;
  assign new_n11961_ = ~new_n11958_ & new_n11960_;
  assign ys__n478 = ~new_n11957_ & new_n11961_;
  assign ys__n4566 = ys__n935 | ys__n478;
  assign new_n11964_ = ys__n23627 & ~ys__n23717;
  assign new_n11965_ = ~ys__n4566 & new_n11964_;
  assign new_n11966_ = new_n11954_ & new_n11965_;
  assign ys__n18120 = new_n11812_ | ~new_n11966_;
  assign new_n11968_ = ys__n19245 & ~ys__n19253;
  assign new_n11969_ = ~ys__n738 & new_n11968_;
  assign new_n11970_ = ~ys__n18120 & new_n11969_;
  assign new_n11971_ = ~ys__n306 & ys__n38567;
  assign new_n11972_ = ys__n306 & ~ys__n38567;
  assign new_n11973_ = ~new_n11971_ & ~new_n11972_;
  assign new_n11974_ = ~ys__n38568 & ys__n38569;
  assign new_n11975_ = ys__n38568 & ~ys__n38569;
  assign new_n11976_ = ~new_n11974_ & ~new_n11975_;
  assign new_n11977_ = new_n11973_ & new_n11976_;
  assign ys__n1073 = ys__n18124 & ys__n24177;
  assign new_n11979_ = new_n11977_ & ys__n1073;
  assign new_n11980_ = ~ys__n418 & ys__n38528;
  assign new_n11981_ = ys__n18121 & ys__n18124;
  assign new_n11982_ = ~new_n11980_ & new_n11981_;
  assign new_n11983_ = ys__n35704 & ~ys__n38529;
  assign new_n11984_ = ys__n418 & ~ys__n38528;
  assign new_n11985_ = ~ys__n35704 & ys__n38529;
  assign new_n11986_ = ~new_n11984_ & ~new_n11985_;
  assign new_n11987_ = ~new_n11983_ & new_n11986_;
  assign new_n11988_ = new_n11982_ & new_n11987_;
  assign new_n11989_ = ys__n18122 & ys__n18124;
  assign new_n11990_ = ~new_n11988_ & ~new_n11989_;
  assign ys__n30223 = new_n11979_ | ~new_n11990_;
  assign new_n11992_ = ys__n19253 & ys__n30223;
  assign new_n11993_ = ~new_n11970_ & ~new_n11992_;
  assign new_n11994_ = ys__n140 & ~ys__n19245;
  assign new_n11995_ = ~ys__n738 & new_n11994_;
  assign new_n11996_ = ys__n19245 & ~ys__n738;
  assign new_n11997_ = ys__n18120 & new_n11996_;
  assign new_n11998_ = ~new_n11995_ & ~new_n11997_;
  assign new_n11999_ = new_n11993_ & new_n11998_;
  assign new_n12000_ = ~new_n11993_ & ~new_n11999_;
  assign ys__n25436 = ~new_n11762_ & new_n12000_;
  assign new_n12002_ = ys__n738 & new_n11994_;
  assign new_n12003_ = ys__n19245 & ys__n738;
  assign new_n12004_ = ~new_n12002_ & ~new_n12003_;
  assign new_n12005_ = ~ys__n19253 & ~new_n12004_;
  assign new_n12006_ = ys__n19253 & ~ys__n30223;
  assign ys__n19256 = new_n12005_ | new_n12006_;
  assign new_n12008_ = ys__n25436 & ~ys__n19256;
  assign new_n12009_ = ys__n642 & ys__n19256;
  assign new_n12010_ = ~new_n12008_ & ~new_n12009_;
  assign ys__n2 = ys__n874 & ~new_n12010_;
  assign new_n12012_ = ~ys__n4299 & ~ys__n4300;
  assign new_n12013_ = ~ys__n4305 & ys__n19263;
  assign new_n12014_ = new_n12012_ & new_n12013_;
  assign new_n12015_ = ys__n244 & ~ys__n4291;
  assign new_n12016_ = ~ys__n4292 & ~ys__n4294;
  assign new_n12017_ = ~ys__n4296 & ~ys__n4297;
  assign new_n12018_ = new_n12016_ & new_n12017_;
  assign new_n12019_ = new_n12015_ & new_n12018_;
  assign new_n12020_ = new_n12014_ & new_n12019_;
  assign new_n12021_ = ys__n20273 & ~ys__n28243;
  assign new_n12022_ = ~ys__n738 & new_n12021_;
  assign ys__n246 = ~new_n12020_ & new_n12022_;
  assign new_n12024_ = ys__n28243 & ~ys__n38203;
  assign new_n12025_ = ys__n28243 & ~ys__n38202;
  assign new_n12026_ = ~ys__n28243 & ys__n38203;
  assign new_n12027_ = ~new_n12025_ & ~new_n12026_;
  assign new_n12028_ = ~new_n12024_ & new_n12027_;
  assign new_n12029_ = ~ys__n28243 & ys__n38199;
  assign new_n12030_ = ys__n38183 & ~ys__n38200;
  assign new_n12031_ = ~new_n12029_ & new_n12030_;
  assign new_n12032_ = ys__n28243 & ~ys__n38199;
  assign new_n12033_ = ~ys__n28243 & ys__n38201;
  assign new_n12034_ = ~new_n12032_ & ~new_n12033_;
  assign new_n12035_ = ys__n28243 & ~ys__n38201;
  assign new_n12036_ = ~ys__n28243 & ys__n38202;
  assign new_n12037_ = ~new_n12035_ & ~new_n12036_;
  assign new_n12038_ = new_n12034_ & new_n12037_;
  assign new_n12039_ = new_n12031_ & new_n12038_;
  assign new_n12040_ = new_n12028_ & new_n12039_;
  assign new_n12041_ = ys__n20273 & ys__n28243;
  assign new_n12042_ = ~ys__n738 & new_n12041_;
  assign new_n12043_ = ~new_n12020_ & new_n12042_;
  assign ys__n250 = new_n12040_ & new_n12043_;
  assign new_n12045_ = ~ys__n19263 & ys__n20279;
  assign new_n12046_ = ~ys__n738 & new_n12045_;
  assign new_n12047_ = ~ys__n19263 & ~new_n12046_;
  assign new_n12048_ = ~ys__n19263 & ys__n20273;
  assign new_n12049_ = ys__n20280 & new_n12048_;
  assign new_n12050_ = ~ys__n738 & new_n12049_;
  assign new_n12051_ = ys__n738 & new_n12048_;
  assign new_n12052_ = ys__n20273 & ~new_n12051_;
  assign new_n12053_ = ~new_n12050_ & new_n12052_;
  assign new_n12054_ = ~new_n12047_ & new_n12053_;
  assign new_n12055_ = ~ys__n766 & ys__n28243;
  assign new_n12056_ = ~ys__n764 & ys__n28243;
  assign new_n12057_ = ys__n766 & ~ys__n28243;
  assign new_n12058_ = ~new_n12056_ & ~new_n12057_;
  assign new_n12059_ = ~new_n12055_ & new_n12058_;
  assign new_n12060_ = ys__n758 & ~ys__n28243;
  assign new_n12061_ = ~ys__n760 & ys__n38198;
  assign new_n12062_ = ~new_n12060_ & new_n12061_;
  assign new_n12063_ = ~ys__n758 & ys__n28243;
  assign new_n12064_ = ys__n762 & ~ys__n28243;
  assign new_n12065_ = ~new_n12063_ & ~new_n12064_;
  assign new_n12066_ = ~ys__n762 & ys__n28243;
  assign new_n12067_ = ys__n764 & ~ys__n28243;
  assign new_n12068_ = ~new_n12066_ & ~new_n12067_;
  assign new_n12069_ = new_n12065_ & new_n12068_;
  assign new_n12070_ = new_n12062_ & new_n12069_;
  assign new_n12071_ = new_n12059_ & new_n12070_;
  assign new_n12072_ = ~new_n12040_ & new_n12071_;
  assign new_n12073_ = new_n12043_ & new_n12072_;
  assign ys__n252 = ~new_n12054_ & new_n12073_;
  assign new_n12075_ = ys__n28243 & ~ys__n738;
  assign new_n12076_ = ~new_n12020_ & new_n12075_;
  assign new_n12077_ = new_n12072_ & new_n12076_;
  assign new_n12078_ = new_n12054_ & new_n12077_;
  assign new_n12079_ = ~new_n12020_ & ~new_n12078_;
  assign ys__n254 = ys__n20273 & ~new_n12079_;
  assign new_n12081_ = ys__n28243 & ~ys__n38197;
  assign new_n12082_ = ys__n28243 & ~ys__n38196;
  assign new_n12083_ = ~ys__n28243 & ys__n38197;
  assign new_n12084_ = ~new_n12082_ & ~new_n12083_;
  assign new_n12085_ = ~new_n12081_ & new_n12084_;
  assign new_n12086_ = ~ys__n28243 & ys__n38193;
  assign new_n12087_ = ys__n38192 & ~ys__n38194;
  assign new_n12088_ = ~new_n12086_ & new_n12087_;
  assign new_n12089_ = ys__n28243 & ~ys__n38193;
  assign new_n12090_ = ~ys__n28243 & ys__n38195;
  assign new_n12091_ = ~new_n12089_ & ~new_n12090_;
  assign new_n12092_ = ys__n28243 & ~ys__n38195;
  assign new_n12093_ = ~ys__n28243 & ys__n38196;
  assign new_n12094_ = ~new_n12092_ & ~new_n12093_;
  assign new_n12095_ = new_n12091_ & new_n12094_;
  assign new_n12096_ = new_n12088_ & new_n12095_;
  assign new_n12097_ = new_n12085_ & new_n12096_;
  assign new_n12098_ = ~new_n12040_ & ~new_n12071_;
  assign new_n12099_ = new_n12097_ & new_n12098_;
  assign ys__n270 = new_n12043_ & new_n12099_;
  assign new_n12101_ = ~new_n12097_ & new_n12098_;
  assign ys__n278 = new_n12043_ & new_n12101_;
  assign ys__n404 = ys__n17849 & ~ys__n18156;
  assign new_n12104_ = ~ys__n33384 & ys__n38315;
  assign new_n12105_ = ys__n38323 & new_n12104_;
  assign new_n12106_ = ~ys__n38320 & ~new_n12105_;
  assign new_n12107_ = ys__n38217 & ~new_n12106_;
  assign new_n12108_ = ys__n38215 & ~new_n12106_;
  assign new_n12109_ = ~new_n12107_ & new_n12108_;
  assign new_n12110_ = ~new_n12107_ & ~new_n12109_;
  assign new_n12111_ = ~ys__n23641 & ~new_n12110_;
  assign new_n12112_ = ~ys__n23641 & ~new_n12111_;
  assign new_n12113_ = ~ys__n23645 & ~ys__n23652;
  assign new_n12114_ = ~new_n12112_ & new_n12113_;
  assign ys__n480 = ys__n23652 | new_n12114_;
  assign new_n12116_ = new_n11955_ & new_n12109_;
  assign new_n12117_ = ys__n23644 & ys__n23645;
  assign new_n12118_ = ~new_n12116_ & ~new_n12117_;
  assign ys__n482 = ~ys__n23652 & ~new_n12118_;
  assign new_n12120_ = ~ys__n206 & ~ys__n208;
  assign new_n12121_ = ~ys__n190 & ~ys__n192;
  assign new_n12122_ = ~ys__n204 & ~ys__n860;
  assign new_n12123_ = new_n12121_ & new_n12122_;
  assign new_n12124_ = new_n12120_ & new_n12123_;
  assign new_n12125_ = ys__n33403 & ~new_n12124_;
  assign new_n12126_ = ys__n30863 & ~ys__n33384;
  assign new_n12127_ = ys__n176 & ~ys__n178;
  assign new_n12128_ = new_n12126_ & new_n12127_;
  assign new_n12129_ = ~new_n12125_ & new_n12128_;
  assign new_n12130_ = ~ys__n176 & ys__n178;
  assign new_n12131_ = new_n12126_ & new_n12130_;
  assign new_n12132_ = new_n12124_ & new_n12131_;
  assign new_n12133_ = ~new_n12129_ & ~new_n12132_;
  assign new_n12134_ = ~ys__n176 & ~ys__n178;
  assign new_n12135_ = ys__n176 & ys__n178;
  assign new_n12136_ = ~new_n12134_ & ~new_n12135_;
  assign new_n12137_ = ~new_n12127_ & ~new_n12130_;
  assign new_n12138_ = new_n12136_ & new_n12137_;
  assign new_n12139_ = ~new_n12133_ & ~new_n12138_;
  assign new_n12140_ = ~ys__n738 & ~ys__n4566;
  assign ys__n502 = new_n12139_ & new_n12140_;
  assign new_n12142_ = ys__n568 & ~ys__n572;
  assign new_n12143_ = ~ys__n566 & ys__n570;
  assign new_n12144_ = new_n12142_ & new_n12143_;
  assign new_n12145_ = ~ys__n568 & ~ys__n572;
  assign new_n12146_ = new_n12143_ & new_n12145_;
  assign new_n12147_ = ys__n568 & ys__n572;
  assign new_n12148_ = ys__n566 & ~ys__n570;
  assign new_n12149_ = new_n12147_ & new_n12148_;
  assign new_n12150_ = ~new_n12146_ & ~new_n12149_;
  assign new_n12151_ = ~new_n12144_ & new_n12150_;
  assign new_n12152_ = ~ys__n568 & ys__n572;
  assign new_n12153_ = new_n12148_ & new_n12152_;
  assign new_n12154_ = new_n12142_ & new_n12148_;
  assign new_n12155_ = ~new_n12153_ & ~new_n12154_;
  assign new_n12156_ = new_n12145_ & new_n12148_;
  assign new_n12157_ = ~ys__n566 & ~ys__n570;
  assign new_n12158_ = new_n12147_ & new_n12157_;
  assign new_n12159_ = ~new_n12156_ & ~new_n12158_;
  assign new_n12160_ = new_n12155_ & new_n12159_;
  assign ys__n17780 = ~new_n12145_ | ~new_n12157_;
  assign new_n12162_ = new_n12143_ & new_n12152_;
  assign new_n12163_ = ~new_n12144_ & ~new_n12162_;
  assign new_n12164_ = ys__n17780 & new_n12163_;
  assign new_n12165_ = new_n12152_ & new_n12157_;
  assign new_n12166_ = new_n12142_ & new_n12157_;
  assign new_n12167_ = ~new_n12165_ & ~new_n12166_;
  assign new_n12168_ = new_n12150_ & new_n12167_;
  assign new_n12169_ = new_n12164_ & new_n12168_;
  assign new_n12170_ = new_n12160_ & new_n12169_;
  assign ys__n574 = ~new_n12151_ & ~new_n12170_;
  assign new_n12172_ = ~ys__n33563 & ~ys__n38922;
  assign new_n12173_ = ys__n38919 & new_n11747_;
  assign new_n12174_ = ~new_n12172_ & new_n12173_;
  assign new_n12175_ = ~ys__n4184 & ~ys__n4810;
  assign new_n12176_ = ~ys__n4192 & new_n12175_;
  assign new_n12177_ = new_n11745_ & ~ys__n17780;
  assign new_n12178_ = new_n12176_ & new_n12177_;
  assign new_n12179_ = new_n12174_ & new_n12178_;
  assign new_n12180_ = new_n11744_ & new_n11747_;
  assign new_n12181_ = ~ys__n4613 & ~ys__n4625;
  assign new_n12182_ = ~ys__n4185 & ~ys__n4810;
  assign new_n12183_ = new_n12181_ & new_n12182_;
  assign new_n12184_ = new_n12165_ & new_n12183_;
  assign new_n12185_ = new_n12180_ & new_n12184_;
  assign new_n12186_ = ys__n47107 & new_n12146_;
  assign new_n12187_ = ys__n30230 & ~ys__n30232;
  assign new_n12188_ = ys__n30232 & ~ys__n33563;
  assign new_n12189_ = ~new_n12187_ & ~new_n12188_;
  assign new_n12190_ = new_n12144_ & new_n12189_;
  assign new_n12191_ = ~new_n12153_ & ~new_n12156_;
  assign new_n12192_ = ~new_n12190_ & new_n12191_;
  assign new_n12193_ = ~new_n12186_ & new_n12192_;
  assign new_n12194_ = ~new_n12185_ & new_n12193_;
  assign new_n12195_ = ~new_n12179_ & new_n12194_;
  assign ys__n576 = ~new_n12170_ & ~new_n12195_;
  assign new_n12197_ = ~ys__n108 & ~ys__n290;
  assign new_n12198_ = ~ys__n110 & ys__n112;
  assign new_n12199_ = ~ys__n1309 & new_n12198_;
  assign new_n12200_ = new_n12197_ & new_n12199_;
  assign new_n12201_ = ~ys__n108 & ~ys__n1309;
  assign new_n12202_ = ~ys__n110 & ~ys__n112;
  assign new_n12203_ = ys__n114 & ~ys__n290;
  assign new_n12204_ = new_n12202_ & new_n12203_;
  assign new_n12205_ = new_n12201_ & new_n12204_;
  assign new_n12206_ = ~new_n12200_ & ~new_n12205_;
  assign new_n12207_ = ~ys__n114 & ys__n118;
  assign new_n12208_ = ~ys__n1309 & new_n12207_;
  assign new_n12209_ = new_n12197_ & new_n12202_;
  assign new_n12210_ = new_n12208_ & new_n12209_;
  assign new_n12211_ = ys__n110 & ~ys__n290;
  assign new_n12212_ = new_n12201_ & new_n12211_;
  assign new_n12213_ = ~ys__n108 & ys__n290;
  assign new_n12214_ = ~ys__n1309 & new_n12213_;
  assign new_n12215_ = ys__n108 & ~ys__n1309;
  assign new_n12216_ = ~ys__n1309 & ~new_n12215_;
  assign new_n12217_ = ~new_n12214_ & new_n12216_;
  assign new_n12218_ = ~new_n12212_ & new_n12217_;
  assign new_n12219_ = ~new_n12210_ & new_n12218_;
  assign new_n12220_ = new_n12206_ & new_n12219_;
  assign new_n12221_ = ys__n112 & new_n12220_;
  assign new_n12222_ = ~ys__n37672 & ys__n37673;
  assign new_n12223_ = ys__n37672 & ~ys__n37673;
  assign new_n12224_ = ~new_n12222_ & ~new_n12223_;
  assign new_n12225_ = ~ys__n18393 & ~new_n12224_;
  assign new_n12226_ = ys__n38861 & ys__n38862;
  assign new_n12227_ = ys__n38863 & ~new_n12226_;
  assign new_n12228_ = ~ys__n33541 & ~ys__n33552;
  assign new_n12229_ = ~ys__n38865 & ~new_n12228_;
  assign new_n12230_ = new_n12227_ & ~new_n12229_;
  assign new_n12231_ = ys__n38864 & ys__n38865;
  assign new_n12232_ = ~ys__n33541 & ys__n38863;
  assign new_n12233_ = ~new_n12227_ & new_n12232_;
  assign new_n12234_ = ~new_n12231_ & ~new_n12233_;
  assign new_n12235_ = ~new_n12230_ & new_n12234_;
  assign new_n12236_ = ~ys__n4750 & ~ys__n4751;
  assign new_n12237_ = ~ys__n4753 & ~ys__n4754;
  assign new_n12238_ = ~ys__n4759 & ~ys__n4761;
  assign new_n12239_ = new_n12237_ & new_n12238_;
  assign new_n12240_ = new_n12236_ & new_n12239_;
  assign new_n12241_ = ~ys__n4756 & ~ys__n4757;
  assign new_n12242_ = ~ys__n4744 & ~ys__n4746;
  assign new_n12243_ = new_n12241_ & new_n12242_;
  assign ys__n4764 = ~new_n12240_ | ~new_n12243_;
  assign new_n12245_ = ~ys__n29117 & ~ys__n4764;
  assign new_n12246_ = ~new_n12235_ & new_n12245_;
  assign ys__n37703 = ys__n24675 | new_n12246_;
  assign new_n12248_ = ys__n33552 & ys__n38865;
  assign new_n12249_ = new_n12227_ & new_n12248_;
  assign new_n12250_ = ~ys__n24675 & ys__n24711;
  assign new_n12251_ = ys__n24675 & ys__n24712;
  assign ys__n18759 = new_n12250_ | new_n12251_;
  assign new_n12253_ = new_n12249_ & ~ys__n18759;
  assign new_n12254_ = ~ys__n38864 & ~new_n12253_;
  assign new_n12255_ = ~ys__n24675 & ~new_n12254_;
  assign new_n12256_ = ys__n37703 & new_n12255_;
  assign ys__n1020 = ys__n4783 | ys__n4784;
  assign new_n12258_ = ~ys__n33545 & ys__n1020;
  assign new_n12259_ = ~ys__n4764 & new_n12258_;
  assign new_n12260_ = ~ys__n844 & ~ys__n3214;
  assign new_n12261_ = ~ys__n18070 & ~ys__n18071;
  assign new_n12262_ = new_n12260_ & new_n12261_;
  assign new_n12263_ = ~new_n12259_ & new_n12262_;
  assign new_n12264_ = ~new_n12256_ & new_n12263_;
  assign new_n12265_ = ys__n18270 & new_n12264_;
  assign new_n12266_ = ~ys__n18270 & ~new_n12264_;
  assign new_n12267_ = ~new_n12265_ & ~new_n12266_;
  assign new_n12268_ = ~ys__n18271 & ~new_n12267_;
  assign new_n12269_ = ys__n18270 & ys__n18271;
  assign ys__n18272 = new_n12268_ | new_n12269_;
  assign new_n12271_ = ~ys__n18393 & ys__n18272;
  assign new_n12272_ = ys__n18271 & ys__n18393;
  assign ys__n27603 = new_n12271_ | new_n12272_;
  assign new_n12274_ = ys__n18393 & ys__n27603;
  assign new_n12275_ = ~new_n12225_ & ~new_n12274_;
  assign new_n12276_ = ~ys__n18208 & ~new_n12275_;
  assign new_n12277_ = ys__n18090 & new_n12276_;
  assign new_n12278_ = ys__n19203 & ~ys__n19215;
  assign new_n12279_ = new_n12215_ & new_n12278_;
  assign new_n12280_ = new_n12277_ & new_n12279_;
  assign new_n12281_ = ys__n18317 & ~new_n12275_;
  assign new_n12282_ = ~ys__n17941 & ~ys__n17943;
  assign new_n12283_ = ys__n18090 & new_n12282_;
  assign new_n12284_ = new_n12210_ & new_n12283_;
  assign new_n12285_ = ~new_n12275_ & new_n12284_;
  assign new_n12286_ = new_n12276_ & new_n12285_;
  assign new_n12287_ = ~new_n12281_ & new_n12286_;
  assign new_n12288_ = ~new_n12280_ & ~new_n12287_;
  assign new_n12289_ = ~new_n12220_ & ~new_n12288_;
  assign ys__n628 = new_n12221_ | new_n12289_;
  assign new_n12291_ = ys__n114 & new_n12220_;
  assign new_n12292_ = ~new_n12220_ & new_n12284_;
  assign new_n12293_ = ~new_n12275_ & new_n12292_;
  assign new_n12294_ = ~new_n12276_ & new_n12293_;
  assign new_n12295_ = ~new_n12281_ & new_n12294_;
  assign ys__n630 = new_n12291_ | new_n12295_;
  assign new_n12297_ = ~ys__n748 & ys__n750;
  assign new_n12298_ = new_n11791_ & new_n12297_;
  assign new_n12299_ = ys__n522 & ys__n524;
  assign new_n12300_ = ys__n526 & ys__n528;
  assign new_n12301_ = new_n12299_ & new_n12300_;
  assign new_n12302_ = ~ys__n512 & ys__n520;
  assign new_n12303_ = ys__n530 & ~ys__n752;
  assign new_n12304_ = new_n12302_ & new_n12303_;
  assign new_n12305_ = new_n12301_ & new_n12304_;
  assign new_n12306_ = ~ys__n23730 & ~ys__n28243;
  assign new_n12307_ = new_n11964_ & new_n12306_;
  assign new_n12308_ = new_n12305_ & new_n12307_;
  assign new_n12309_ = new_n12298_ & new_n12308_;
  assign new_n12310_ = ~ys__n23627 & ~new_n12309_;
  assign new_n12311_ = ys__n22880 & new_n12309_;
  assign new_n12312_ = ~new_n12310_ & ~new_n12311_;
  assign new_n12313_ = ys__n23627 & ys__n23717;
  assign new_n12314_ = ~ys__n23730 & new_n12313_;
  assign new_n12315_ = ~new_n12312_ & ~new_n12314_;
  assign new_n12316_ = ys__n23328 & new_n12314_;
  assign new_n12317_ = ~new_n12315_ & ~new_n12316_;
  assign new_n12318_ = ~ys__n23730 & ys__n28243;
  assign new_n12319_ = new_n11964_ & new_n12318_;
  assign new_n12320_ = new_n11810_ & new_n12319_;
  assign new_n12321_ = ~new_n12317_ & ~new_n12320_;
  assign new_n12322_ = ys__n450 & new_n12320_;
  assign new_n12323_ = ~new_n12321_ & ~new_n12322_;
  assign new_n12324_ = new_n11802_ & new_n12297_;
  assign new_n12325_ = new_n11784_ & new_n12297_;
  assign new_n12326_ = ~new_n12324_ & ~new_n12325_;
  assign new_n12327_ = new_n11766_ & new_n11796_;
  assign new_n12328_ = new_n11796_ & new_n12297_;
  assign new_n12329_ = ~new_n12298_ & ~new_n12328_;
  assign new_n12330_ = ~new_n12327_ & new_n12329_;
  assign new_n12331_ = new_n12326_ & new_n12330_;
  assign new_n12332_ = new_n11766_ & new_n11806_;
  assign new_n12333_ = new_n11775_ & new_n11801_;
  assign new_n12334_ = new_n11766_ & new_n12333_;
  assign new_n12335_ = ~new_n12332_ & ~new_n12334_;
  assign new_n12336_ = new_n11781_ & new_n12335_;
  assign new_n12337_ = new_n11766_ & new_n11802_;
  assign new_n12338_ = new_n11764_ & new_n11778_;
  assign new_n12339_ = new_n12297_ & new_n12338_;
  assign new_n12340_ = ~new_n11785_ & ~new_n12339_;
  assign new_n12341_ = ~new_n12337_ & new_n12340_;
  assign new_n12342_ = new_n12336_ & new_n12341_;
  assign new_n12343_ = new_n12331_ & new_n12342_;
  assign new_n12344_ = ~ys__n4494 & ~ys__n4496;
  assign new_n12345_ = ys__n512 & ~ys__n632;
  assign new_n12346_ = new_n12344_ & new_n12345_;
  assign new_n12347_ = ~ys__n520 & new_n12346_;
  assign new_n12348_ = ~ys__n4478 & ~ys__n4480;
  assign new_n12349_ = ~ys__n514 & ~ys__n2024;
  assign new_n12350_ = new_n12348_ & new_n12349_;
  assign new_n12351_ = ~ys__n516 & new_n12350_;
  assign new_n12352_ = new_n12347_ & new_n12351_;
  assign new_n12353_ = ~ys__n28720 & new_n12352_;
  assign new_n12354_ = ys__n514 & ~ys__n2024;
  assign new_n12355_ = new_n12348_ & new_n12354_;
  assign new_n12356_ = ~ys__n516 & new_n12355_;
  assign new_n12357_ = new_n12347_ & new_n12356_;
  assign new_n12358_ = ys__n28720 & new_n12357_;
  assign new_n12359_ = ~new_n12353_ & ~new_n12358_;
  assign new_n12360_ = new_n12324_ & new_n12359_;
  assign new_n12361_ = new_n12298_ & ~new_n12305_;
  assign new_n12362_ = ys__n516 & new_n12350_;
  assign new_n12363_ = ys__n516 & new_n12355_;
  assign new_n12364_ = ~new_n12362_ & ~new_n12363_;
  assign new_n12365_ = ~new_n12351_ & ~new_n12356_;
  assign new_n12366_ = new_n12364_ & new_n12365_;
  assign new_n12367_ = new_n12327_ & new_n12366_;
  assign new_n12368_ = ~new_n12361_ & ~new_n12367_;
  assign new_n12369_ = ~new_n12360_ & new_n12368_;
  assign new_n12370_ = ~ys__n28719 & new_n12352_;
  assign new_n12371_ = ys__n28719 & new_n12357_;
  assign new_n12372_ = ~new_n12370_ & ~new_n12371_;
  assign new_n12373_ = new_n12325_ & new_n12372_;
  assign new_n12374_ = ~ys__n28718 & new_n12352_;
  assign new_n12375_ = ys__n28718 & new_n12357_;
  assign new_n12376_ = ~new_n12374_ & ~new_n12375_;
  assign new_n12377_ = new_n12328_ & new_n12376_;
  assign new_n12378_ = ~new_n12373_ & ~new_n12377_;
  assign new_n12379_ = new_n12369_ & new_n12378_;
  assign new_n12380_ = ~new_n12343_ & ~new_n12379_;
  assign new_n12381_ = ~new_n12343_ & ~new_n12380_;
  assign new_n12382_ = ~ys__n28243 & ~new_n12381_;
  assign new_n12383_ = ~new_n11767_ & ~new_n11785_;
  assign new_n12384_ = new_n11792_ & new_n12338_;
  assign new_n12385_ = ~new_n11807_ & ~new_n12384_;
  assign new_n12386_ = new_n12383_ & new_n12385_;
  assign new_n12387_ = new_n11781_ & new_n11805_;
  assign new_n12388_ = new_n12386_ & new_n12387_;
  assign new_n12389_ = new_n11800_ & new_n12388_;
  assign new_n12390_ = new_n11767_ & new_n11772_;
  assign new_n12391_ = ~ys__n526 & ~ys__n528;
  assign new_n12392_ = ~ys__n522 & ~ys__n524;
  assign new_n12393_ = new_n12391_ & new_n12392_;
  assign new_n12394_ = ~ys__n530 & new_n12393_;
  assign new_n12395_ = ~ys__n23730 & new_n12394_;
  assign new_n12396_ = new_n12394_ & ~new_n12395_;
  assign new_n12397_ = new_n12384_ & ~new_n12396_;
  assign new_n12398_ = ~new_n12390_ & ~new_n12397_;
  assign new_n12399_ = ~new_n12389_ & ~new_n12398_;
  assign new_n12400_ = ~new_n12389_ & ~new_n12399_;
  assign new_n12401_ = ys__n28243 & ~new_n12400_;
  assign new_n12402_ = ~new_n12382_ & ~new_n12401_;
  assign new_n12403_ = ~ys__n23730 & new_n11964_;
  assign new_n12404_ = ~new_n12402_ & new_n12403_;
  assign new_n12405_ = ~new_n12323_ & ~new_n12404_;
  assign new_n12406_ = ~ys__n23339 & ys__n23548;
  assign new_n12407_ = ys__n23550 & new_n12406_;
  assign new_n12408_ = ~ys__n23339 & ~ys__n23548;
  assign new_n12409_ = ys__n23339 & ys__n23548;
  assign new_n12410_ = ~new_n12408_ & ~new_n12409_;
  assign new_n12411_ = ys__n22464 & ys__n23339;
  assign new_n12412_ = ys__n23550 & new_n12411_;
  assign new_n12413_ = ~new_n12410_ & new_n12412_;
  assign new_n12414_ = ~new_n12407_ & ~new_n12413_;
  assign new_n12415_ = ys__n23552 & ys__n23554;
  assign new_n12416_ = ys__n23556 & ys__n23558;
  assign new_n12417_ = new_n12415_ & new_n12416_;
  assign new_n12418_ = ~new_n12414_ & new_n12417_;
  assign new_n12419_ = ys__n23560 & ys__n23562;
  assign new_n12420_ = ys__n23564 & ys__n23566;
  assign new_n12421_ = new_n12419_ & new_n12420_;
  assign new_n12422_ = ys__n23568 & ys__n23570;
  assign new_n12423_ = ys__n23572 & ys__n23574;
  assign new_n12424_ = new_n12422_ & new_n12423_;
  assign new_n12425_ = new_n12421_ & new_n12424_;
  assign new_n12426_ = new_n12418_ & new_n12425_;
  assign new_n12427_ = ys__n450 & ~new_n12426_;
  assign new_n12428_ = ys__n420 & ys__n442;
  assign new_n12429_ = ys__n440 & ys__n444;
  assign new_n12430_ = new_n12428_ & new_n12429_;
  assign new_n12431_ = ys__n438 & ys__n446;
  assign new_n12432_ = ys__n434 & ys__n436;
  assign new_n12433_ = new_n12431_ & new_n12432_;
  assign new_n12434_ = new_n12430_ & new_n12433_;
  assign new_n12435_ = ys__n432 & ys__n448;
  assign new_n12436_ = ys__n428 & ys__n430;
  assign new_n12437_ = new_n12435_ & new_n12436_;
  assign new_n12438_ = new_n12434_ & new_n12437_;
  assign new_n12439_ = ys__n426 & new_n12438_;
  assign new_n12440_ = ~ys__n450 & new_n12439_;
  assign new_n12441_ = ys__n450 & ~new_n12439_;
  assign new_n12442_ = ~new_n12440_ & ~new_n12441_;
  assign new_n12443_ = new_n12426_ & ~new_n12442_;
  assign ys__n23539 = new_n12427_ | new_n12443_;
  assign new_n12445_ = new_n12404_ & ys__n23539;
  assign new_n12446_ = ~new_n12405_ & ~new_n12445_;
  assign new_n12447_ = ~new_n11785_ & ~new_n12337_;
  assign new_n12448_ = ~ys__n23717 & ~ys__n23730;
  assign new_n12449_ = ~ys__n28243 & new_n12448_;
  assign new_n12450_ = ~new_n12447_ & new_n12449_;
  assign new_n12451_ = ~ys__n23729 & ys__n23730;
  assign new_n12452_ = ~new_n12450_ & ~new_n12451_;
  assign new_n12453_ = ys__n23627 & ~new_n12452_;
  assign new_n12454_ = new_n12339_ & new_n12449_;
  assign new_n12455_ = ys__n23729 & ys__n23730;
  assign new_n12456_ = ~new_n12454_ & ~new_n12455_;
  assign new_n12457_ = ys__n23627 & ~new_n12456_;
  assign new_n12458_ = ~new_n12453_ & ~new_n12457_;
  assign new_n12459_ = ~new_n12446_ & new_n12458_;
  assign new_n12460_ = ys__n450 & ~new_n12458_;
  assign new_n12461_ = ~new_n12459_ & ~new_n12460_;
  assign new_n12462_ = new_n12324_ & ~new_n12359_;
  assign new_n12463_ = new_n12327_ & ~new_n12366_;
  assign new_n12464_ = new_n12336_ & ~new_n12463_;
  assign new_n12465_ = ~new_n12462_ & new_n12464_;
  assign new_n12466_ = new_n12325_ & ~new_n12372_;
  assign new_n12467_ = new_n12328_ & ~new_n12376_;
  assign new_n12468_ = ~new_n12466_ & ~new_n12467_;
  assign new_n12469_ = new_n12465_ & new_n12468_;
  assign new_n12470_ = ~new_n12327_ & ~new_n12328_;
  assign new_n12471_ = new_n12326_ & new_n12470_;
  assign new_n12472_ = new_n12336_ & new_n12471_;
  assign new_n12473_ = ~ys__n28243 & ~new_n12472_;
  assign new_n12474_ = ~new_n12469_ & new_n12473_;
  assign new_n12475_ = ys__n28243 & new_n11790_;
  assign new_n12476_ = ~new_n12474_ & ~new_n12475_;
  assign new_n12477_ = new_n12403_ & ~new_n12476_;
  assign new_n12478_ = ~new_n12461_ & ~new_n12477_;
  assign new_n12479_ = ys__n634 & ~ys__n28243;
  assign new_n12480_ = ~ys__n256 & ~ys__n744;
  assign new_n12481_ = ys__n550 & new_n12480_;
  assign new_n12482_ = ys__n256 & ys__n28641;
  assign new_n12483_ = ~ys__n256 & ys__n744;
  assign new_n12484_ = ys__n4488 & new_n12483_;
  assign new_n12485_ = ~new_n12482_ & ~new_n12484_;
  assign new_n12486_ = ~new_n12481_ & new_n12485_;
  assign new_n12487_ = ~ys__n256 & ~new_n12483_;
  assign new_n12488_ = ~new_n12480_ & new_n12487_;
  assign new_n12489_ = ys__n28243 & ~new_n12488_;
  assign new_n12490_ = ~new_n12486_ & new_n12489_;
  assign new_n12491_ = ~new_n12479_ & ~new_n12490_;
  assign new_n12492_ = ys__n420 & ~new_n12491_;
  assign new_n12493_ = ~ys__n420 & ~new_n12491_;
  assign new_n12494_ = ys__n420 & new_n12491_;
  assign new_n12495_ = ~new_n12493_ & ~new_n12494_;
  assign new_n12496_ = ys__n528 & ~ys__n28243;
  assign new_n12497_ = ys__n526 & new_n12480_;
  assign new_n12498_ = ys__n256 & ys__n526;
  assign new_n12499_ = ys__n526 & new_n12483_;
  assign new_n12500_ = ~new_n12498_ & ~new_n12499_;
  assign new_n12501_ = ~new_n12497_ & new_n12500_;
  assign new_n12502_ = new_n12489_ & ~new_n12501_;
  assign new_n12503_ = ~new_n12496_ & ~new_n12502_;
  assign new_n12504_ = ~ys__n23548 & ~new_n12503_;
  assign new_n12505_ = ys__n23548 & new_n12503_;
  assign new_n12506_ = ~new_n12504_ & ~new_n12505_;
  assign new_n12507_ = ys__n526 & ~ys__n28243;
  assign new_n12508_ = ys__n524 & new_n12480_;
  assign new_n12509_ = ys__n256 & ys__n524;
  assign new_n12510_ = ys__n524 & new_n12483_;
  assign new_n12511_ = ~new_n12509_ & ~new_n12510_;
  assign new_n12512_ = ~new_n12508_ & new_n12511_;
  assign new_n12513_ = new_n12489_ & ~new_n12512_;
  assign new_n12514_ = ~new_n12507_ & ~new_n12513_;
  assign new_n12515_ = ~ys__n23550 & ~new_n12514_;
  assign new_n12516_ = ys__n23550 & new_n12514_;
  assign new_n12517_ = ~new_n12515_ & ~new_n12516_;
  assign new_n12518_ = ys__n528 & new_n12480_;
  assign new_n12519_ = ys__n256 & ys__n528;
  assign new_n12520_ = ys__n528 & new_n12483_;
  assign new_n12521_ = ~new_n12519_ & ~new_n12520_;
  assign new_n12522_ = ~new_n12518_ & new_n12521_;
  assign new_n12523_ = new_n12489_ & ~new_n12522_;
  assign new_n12524_ = ys__n22464 & new_n12523_;
  assign new_n12525_ = ~new_n12517_ & new_n12524_;
  assign new_n12526_ = ~new_n12506_ & new_n12525_;
  assign new_n12527_ = ys__n23550 & ~new_n12514_;
  assign new_n12528_ = ys__n23548 & ~new_n12503_;
  assign new_n12529_ = ~new_n12517_ & new_n12528_;
  assign new_n12530_ = ~new_n12527_ & ~new_n12529_;
  assign new_n12531_ = ~new_n12526_ & new_n12530_;
  assign new_n12532_ = ys__n752 & ~ys__n28243;
  assign new_n12533_ = ys__n736 & new_n12480_;
  assign new_n12534_ = ys__n256 & ys__n28633;
  assign new_n12535_ = ys__n736 & new_n12483_;
  assign new_n12536_ = ~new_n12534_ & ~new_n12535_;
  assign new_n12537_ = ~new_n12533_ & new_n12536_;
  assign new_n12538_ = new_n12489_ & ~new_n12537_;
  assign new_n12539_ = ~new_n12532_ & ~new_n12538_;
  assign new_n12540_ = ~ys__n23558 & ~new_n12539_;
  assign new_n12541_ = ys__n23558 & new_n12539_;
  assign new_n12542_ = ~new_n12540_ & ~new_n12541_;
  assign new_n12543_ = ys__n530 & ~ys__n28243;
  assign new_n12544_ = ys__n752 & new_n12480_;
  assign new_n12545_ = ys__n256 & ys__n28632;
  assign new_n12546_ = ys__n752 & new_n12483_;
  assign new_n12547_ = ~new_n12545_ & ~new_n12546_;
  assign new_n12548_ = ~new_n12544_ & new_n12547_;
  assign new_n12549_ = new_n12489_ & ~new_n12548_;
  assign new_n12550_ = ~new_n12543_ & ~new_n12549_;
  assign new_n12551_ = ~ys__n23556 & ~new_n12550_;
  assign new_n12552_ = ys__n23556 & new_n12550_;
  assign new_n12553_ = ~new_n12551_ & ~new_n12552_;
  assign new_n12554_ = ~new_n12542_ & ~new_n12553_;
  assign new_n12555_ = ys__n522 & ~ys__n28243;
  assign new_n12556_ = ys__n530 & new_n12480_;
  assign new_n12557_ = ys__n256 & ys__n530;
  assign new_n12558_ = ys__n530 & new_n12483_;
  assign new_n12559_ = ~new_n12557_ & ~new_n12558_;
  assign new_n12560_ = ~new_n12556_ & new_n12559_;
  assign new_n12561_ = new_n12489_ & ~new_n12560_;
  assign new_n12562_ = ~new_n12555_ & ~new_n12561_;
  assign new_n12563_ = ~ys__n23554 & ~new_n12562_;
  assign new_n12564_ = ys__n23554 & new_n12562_;
  assign new_n12565_ = ~new_n12563_ & ~new_n12564_;
  assign new_n12566_ = ys__n524 & ~ys__n28243;
  assign new_n12567_ = ys__n522 & new_n12480_;
  assign new_n12568_ = ys__n256 & ys__n522;
  assign new_n12569_ = ys__n522 & new_n12483_;
  assign new_n12570_ = ~new_n12568_ & ~new_n12569_;
  assign new_n12571_ = ~new_n12567_ & new_n12570_;
  assign new_n12572_ = new_n12489_ & ~new_n12571_;
  assign new_n12573_ = ~new_n12566_ & ~new_n12572_;
  assign new_n12574_ = ~ys__n23552 & ~new_n12573_;
  assign new_n12575_ = ys__n23552 & new_n12573_;
  assign new_n12576_ = ~new_n12574_ & ~new_n12575_;
  assign new_n12577_ = ~new_n12565_ & ~new_n12576_;
  assign new_n12578_ = new_n12554_ & new_n12577_;
  assign new_n12579_ = ~new_n12531_ & new_n12578_;
  assign new_n12580_ = ys__n23554 & ~new_n12562_;
  assign new_n12581_ = ys__n23552 & ~new_n12573_;
  assign new_n12582_ = ~new_n12565_ & new_n12581_;
  assign new_n12583_ = ~new_n12580_ & ~new_n12582_;
  assign new_n12584_ = new_n12554_ & ~new_n12583_;
  assign new_n12585_ = ys__n23558 & ~new_n12539_;
  assign new_n12586_ = ys__n23556 & ~new_n12550_;
  assign new_n12587_ = ~new_n12542_ & new_n12586_;
  assign new_n12588_ = ~new_n12585_ & ~new_n12587_;
  assign new_n12589_ = ~new_n12584_ & new_n12588_;
  assign new_n12590_ = ~new_n12579_ & new_n12589_;
  assign new_n12591_ = ys__n636 & ~ys__n28243;
  assign new_n12592_ = ys__n256 & ys__n28640;
  assign new_n12593_ = ~new_n12484_ & ~new_n12592_;
  assign new_n12594_ = ~new_n12481_ & new_n12593_;
  assign new_n12595_ = new_n12489_ & ~new_n12594_;
  assign new_n12596_ = ~new_n12591_ & ~new_n12595_;
  assign new_n12597_ = ~ys__n23574 & ~new_n12596_;
  assign new_n12598_ = ys__n23574 & new_n12596_;
  assign new_n12599_ = ~new_n12597_ & ~new_n12598_;
  assign new_n12600_ = ys__n638 & ~ys__n28243;
  assign new_n12601_ = ys__n256 & ys__n28639;
  assign new_n12602_ = ~new_n12484_ & ~new_n12601_;
  assign new_n12603_ = ~new_n12481_ & new_n12602_;
  assign new_n12604_ = new_n12489_ & ~new_n12603_;
  assign new_n12605_ = ~new_n12600_ & ~new_n12604_;
  assign new_n12606_ = ~ys__n23572 & ~new_n12605_;
  assign new_n12607_ = ys__n23572 & new_n12605_;
  assign new_n12608_ = ~new_n12606_ & ~new_n12607_;
  assign new_n12609_ = ~new_n12599_ & ~new_n12608_;
  assign new_n12610_ = ys__n640 & ~ys__n28243;
  assign new_n12611_ = ys__n256 & ys__n28638;
  assign new_n12612_ = ~new_n12484_ & ~new_n12611_;
  assign new_n12613_ = ~new_n12481_ & new_n12612_;
  assign new_n12614_ = new_n12489_ & ~new_n12613_;
  assign new_n12615_ = ~new_n12610_ & ~new_n12614_;
  assign new_n12616_ = ~ys__n23570 & ~new_n12615_;
  assign new_n12617_ = ys__n23570 & new_n12615_;
  assign new_n12618_ = ~new_n12616_ & ~new_n12617_;
  assign new_n12619_ = ys__n550 & ~ys__n28243;
  assign new_n12620_ = ys__n256 & ys__n28637;
  assign new_n12621_ = ~new_n12484_ & ~new_n12620_;
  assign new_n12622_ = ~new_n12481_ & new_n12621_;
  assign new_n12623_ = new_n12489_ & ~new_n12622_;
  assign new_n12624_ = ~new_n12619_ & ~new_n12623_;
  assign new_n12625_ = ~ys__n23568 & ~new_n12624_;
  assign new_n12626_ = ys__n23568 & new_n12624_;
  assign new_n12627_ = ~new_n12625_ & ~new_n12626_;
  assign new_n12628_ = ~new_n12618_ & ~new_n12627_;
  assign new_n12629_ = new_n12609_ & new_n12628_;
  assign new_n12630_ = ys__n548 & ~ys__n28243;
  assign new_n12631_ = ys__n256 & ys__n47660;
  assign new_n12632_ = ~new_n12484_ & ~new_n12631_;
  assign new_n12633_ = ~new_n12481_ & new_n12632_;
  assign new_n12634_ = new_n12489_ & ~new_n12633_;
  assign new_n12635_ = ~new_n12630_ & ~new_n12634_;
  assign new_n12636_ = ~ys__n23566 & ~new_n12635_;
  assign new_n12637_ = ys__n23566 & new_n12635_;
  assign new_n12638_ = ~new_n12636_ & ~new_n12637_;
  assign new_n12639_ = ys__n518 & ~ys__n28243;
  assign new_n12640_ = ys__n548 & new_n12480_;
  assign new_n12641_ = ys__n256 & ys__n28636;
  assign new_n12642_ = ~new_n12484_ & ~new_n12641_;
  assign new_n12643_ = ~new_n12640_ & new_n12642_;
  assign new_n12644_ = new_n12489_ & ~new_n12643_;
  assign new_n12645_ = ~new_n12639_ & ~new_n12644_;
  assign new_n12646_ = ~ys__n23564 & ~new_n12645_;
  assign new_n12647_ = ys__n23564 & new_n12645_;
  assign new_n12648_ = ~new_n12646_ & ~new_n12647_;
  assign new_n12649_ = ~new_n12638_ & ~new_n12648_;
  assign new_n12650_ = ys__n4488 & ~ys__n28243;
  assign new_n12651_ = ys__n518 & new_n12480_;
  assign new_n12652_ = ys__n256 & ys__n28635;
  assign new_n12653_ = ~new_n12484_ & ~new_n12652_;
  assign new_n12654_ = ~new_n12651_ & new_n12653_;
  assign new_n12655_ = new_n12489_ & ~new_n12654_;
  assign new_n12656_ = ~new_n12650_ & ~new_n12655_;
  assign new_n12657_ = ~ys__n23562 & ~new_n12656_;
  assign new_n12658_ = ys__n23562 & new_n12656_;
  assign new_n12659_ = ~new_n12657_ & ~new_n12658_;
  assign new_n12660_ = ys__n736 & ~ys__n28243;
  assign new_n12661_ = ys__n4488 & new_n12480_;
  assign new_n12662_ = ys__n256 & ys__n28634;
  assign new_n12663_ = ~new_n12484_ & ~new_n12662_;
  assign new_n12664_ = ~new_n12661_ & new_n12663_;
  assign new_n12665_ = new_n12489_ & ~new_n12664_;
  assign new_n12666_ = ~new_n12660_ & ~new_n12665_;
  assign new_n12667_ = ~ys__n23560 & ~new_n12666_;
  assign new_n12668_ = ys__n23560 & new_n12666_;
  assign new_n12669_ = ~new_n12667_ & ~new_n12668_;
  assign new_n12670_ = ~new_n12659_ & ~new_n12669_;
  assign new_n12671_ = new_n12649_ & new_n12670_;
  assign new_n12672_ = new_n12629_ & new_n12671_;
  assign new_n12673_ = ~new_n12590_ & new_n12672_;
  assign new_n12674_ = ys__n23562 & ~new_n12656_;
  assign new_n12675_ = ys__n23560 & ~new_n12666_;
  assign new_n12676_ = ~new_n12659_ & new_n12675_;
  assign new_n12677_ = ~new_n12674_ & ~new_n12676_;
  assign new_n12678_ = new_n12649_ & ~new_n12677_;
  assign new_n12679_ = ys__n23566 & ~new_n12635_;
  assign new_n12680_ = ys__n23564 & ~new_n12645_;
  assign new_n12681_ = ~new_n12638_ & new_n12680_;
  assign new_n12682_ = ~new_n12679_ & ~new_n12681_;
  assign new_n12683_ = ~new_n12678_ & new_n12682_;
  assign new_n12684_ = new_n12629_ & ~new_n12683_;
  assign new_n12685_ = ys__n23570 & ~new_n12615_;
  assign new_n12686_ = ys__n23568 & ~new_n12624_;
  assign new_n12687_ = ~new_n12618_ & new_n12686_;
  assign new_n12688_ = ~new_n12685_ & ~new_n12687_;
  assign new_n12689_ = new_n12609_ & ~new_n12688_;
  assign new_n12690_ = ys__n23574 & ~new_n12596_;
  assign new_n12691_ = ys__n23572 & ~new_n12605_;
  assign new_n12692_ = ~new_n12599_ & new_n12691_;
  assign new_n12693_ = ~new_n12690_ & ~new_n12692_;
  assign new_n12694_ = ~new_n12689_ & new_n12693_;
  assign new_n12695_ = ~new_n12684_ & new_n12694_;
  assign new_n12696_ = ~new_n12673_ & new_n12695_;
  assign new_n12697_ = ~new_n12495_ & ~new_n12696_;
  assign new_n12698_ = ~new_n12492_ & ~new_n12697_;
  assign new_n12699_ = ys__n642 & ~ys__n28243;
  assign new_n12700_ = ~new_n12490_ & ~new_n12699_;
  assign new_n12701_ = new_n12698_ & new_n12700_;
  assign new_n12702_ = ~new_n12698_ & ~new_n12700_;
  assign new_n12703_ = ~new_n12701_ & ~new_n12702_;
  assign new_n12704_ = ys__n450 & ~new_n12703_;
  assign new_n12705_ = ~ys__n440 & ys__n442;
  assign new_n12706_ = ~ys__n440 & ~new_n12705_;
  assign new_n12707_ = ~ys__n438 & ~ys__n444;
  assign new_n12708_ = ~new_n12706_ & new_n12707_;
  assign new_n12709_ = ~ys__n438 & ys__n444;
  assign new_n12710_ = ~ys__n438 & ~new_n12709_;
  assign new_n12711_ = ~new_n12708_ & new_n12710_;
  assign new_n12712_ = ~ys__n432 & ~ys__n436;
  assign new_n12713_ = ~ys__n434 & ~ys__n446;
  assign new_n12714_ = new_n12712_ & new_n12713_;
  assign new_n12715_ = ~new_n12711_ & new_n12714_;
  assign new_n12716_ = ~ys__n434 & ys__n446;
  assign new_n12717_ = ~ys__n434 & ~new_n12716_;
  assign new_n12718_ = new_n12712_ & ~new_n12717_;
  assign new_n12719_ = ~ys__n432 & ys__n436;
  assign new_n12720_ = ~ys__n432 & ~new_n12719_;
  assign new_n12721_ = ~new_n12718_ & new_n12720_;
  assign new_n12722_ = ~new_n12715_ & new_n12721_;
  assign new_n12723_ = ~ys__n426 & ~ys__n430;
  assign new_n12724_ = ~ys__n428 & ~ys__n448;
  assign new_n12725_ = new_n12723_ & new_n12724_;
  assign new_n12726_ = ~new_n12722_ & new_n12725_;
  assign new_n12727_ = ~ys__n428 & ys__n448;
  assign new_n12728_ = ~ys__n428 & ~new_n12727_;
  assign new_n12729_ = new_n12723_ & ~new_n12728_;
  assign new_n12730_ = ~ys__n426 & ys__n430;
  assign new_n12731_ = ~ys__n426 & ~new_n12730_;
  assign new_n12732_ = ~new_n12729_ & new_n12731_;
  assign new_n12733_ = ~new_n12726_ & new_n12732_;
  assign new_n12734_ = ys__n450 & ~new_n12733_;
  assign new_n12735_ = ~ys__n450 & new_n12733_;
  assign new_n12736_ = ~new_n12734_ & ~new_n12735_;
  assign new_n12737_ = new_n12698_ & ~new_n12700_;
  assign new_n12738_ = ~new_n12736_ & new_n12737_;
  assign new_n12739_ = ys__n428 & ys__n448;
  assign new_n12740_ = ys__n426 & ys__n430;
  assign new_n12741_ = new_n12739_ & new_n12740_;
  assign new_n12742_ = ys__n440 & ys__n442;
  assign new_n12743_ = ys__n438 & ys__n444;
  assign new_n12744_ = new_n12742_ & new_n12743_;
  assign new_n12745_ = ys__n434 & ys__n446;
  assign new_n12746_ = ys__n432 & ys__n436;
  assign new_n12747_ = new_n12745_ & new_n12746_;
  assign new_n12748_ = new_n12744_ & new_n12747_;
  assign new_n12749_ = new_n12741_ & new_n12748_;
  assign new_n12750_ = ~ys__n450 & new_n12749_;
  assign new_n12751_ = ys__n450 & ~new_n12749_;
  assign new_n12752_ = ~new_n12750_ & ~new_n12751_;
  assign new_n12753_ = ~new_n12698_ & new_n12700_;
  assign new_n12754_ = ~new_n12752_ & new_n12753_;
  assign new_n12755_ = ~new_n12738_ & ~new_n12754_;
  assign new_n12756_ = ~new_n12704_ & new_n12755_;
  assign new_n12757_ = ~new_n12737_ & ~new_n12753_;
  assign new_n12758_ = new_n12703_ & new_n12757_;
  assign new_n12759_ = new_n12477_ & ~new_n12758_;
  assign new_n12760_ = ~new_n12756_ & new_n12759_;
  assign new_n12761_ = ~new_n12478_ & ~new_n12760_;
  assign new_n12762_ = ys__n23627 & ys__n4566;
  assign new_n12763_ = ~new_n11820_ & ~new_n12762_;
  assign new_n12764_ = ~new_n12761_ & new_n12763_;
  assign new_n12765_ = ~ys__n935 & ys__n28446;
  assign new_n12766_ = ~ys__n935 & ~new_n12765_;
  assign new_n12767_ = new_n12762_ & ~new_n12766_;
  assign new_n12768_ = new_n11820_ & ~new_n12762_;
  assign new_n12769_ = ys__n47690 & new_n12768_;
  assign new_n12770_ = ~new_n12767_ & ~new_n12769_;
  assign new_n12771_ = ~new_n12764_ & new_n12770_;
  assign new_n12772_ = ~new_n12762_ & ~new_n12768_;
  assign new_n12773_ = ~new_n12763_ & new_n12772_;
  assign new_n12774_ = new_n11947_ & ~new_n12773_;
  assign new_n12775_ = ~new_n12771_ & new_n12774_;
  assign new_n12776_ = ~new_n11952_ & ~new_n12762_;
  assign new_n12777_ = ~new_n12761_ & new_n12776_;
  assign new_n12778_ = new_n11952_ & ~new_n12762_;
  assign new_n12779_ = ys__n47690 & new_n12778_;
  assign new_n12780_ = ~new_n12767_ & ~new_n12779_;
  assign new_n12781_ = ~new_n12777_ & new_n12780_;
  assign new_n12782_ = ~new_n12762_ & ~new_n12778_;
  assign new_n12783_ = ~new_n12776_ & new_n12782_;
  assign new_n12784_ = ~new_n11947_ & ~new_n12783_;
  assign new_n12785_ = ~new_n12781_ & new_n12784_;
  assign ys__n714 = new_n12775_ | new_n12785_;
  assign new_n12787_ = ys__n22884 & new_n12309_;
  assign new_n12788_ = ~new_n12310_ & ~new_n12787_;
  assign new_n12789_ = ~new_n12314_ & ~new_n12788_;
  assign new_n12790_ = ys__n23332 & new_n12314_;
  assign new_n12791_ = ~new_n12789_ & ~new_n12790_;
  assign new_n12792_ = ~new_n12320_ & ~new_n12791_;
  assign new_n12793_ = ys__n422 & new_n12320_;
  assign new_n12794_ = ~new_n12792_ & ~new_n12793_;
  assign new_n12795_ = ~new_n12404_ & ~new_n12794_;
  assign new_n12796_ = ys__n422 & ~new_n12426_;
  assign new_n12797_ = ys__n426 & ys__n450;
  assign new_n12798_ = new_n12438_ & new_n12797_;
  assign new_n12799_ = ys__n424 & new_n12798_;
  assign new_n12800_ = ~ys__n422 & new_n12799_;
  assign new_n12801_ = ys__n422 & ~new_n12799_;
  assign new_n12802_ = ~new_n12800_ & ~new_n12801_;
  assign new_n12803_ = new_n12426_ & ~new_n12802_;
  assign ys__n23543 = new_n12796_ | new_n12803_;
  assign new_n12805_ = new_n12404_ & ys__n23543;
  assign new_n12806_ = ~new_n12795_ & ~new_n12805_;
  assign new_n12807_ = new_n12458_ & ~new_n12806_;
  assign new_n12808_ = ys__n422 & ~new_n12458_;
  assign new_n12809_ = ~new_n12807_ & ~new_n12808_;
  assign new_n12810_ = ~new_n12477_ & ~new_n12809_;
  assign new_n12811_ = ys__n422 & ~new_n12703_;
  assign new_n12812_ = ~ys__n424 & ~ys__n450;
  assign new_n12813_ = ~new_n12733_ & new_n12812_;
  assign new_n12814_ = ~ys__n424 & ys__n450;
  assign new_n12815_ = ~ys__n424 & ~new_n12814_;
  assign new_n12816_ = ~new_n12813_ & new_n12815_;
  assign new_n12817_ = ys__n422 & ~new_n12816_;
  assign new_n12818_ = ~ys__n422 & new_n12816_;
  assign new_n12819_ = ~new_n12817_ & ~new_n12818_;
  assign new_n12820_ = new_n12737_ & ~new_n12819_;
  assign new_n12821_ = ys__n424 & ys__n450;
  assign new_n12822_ = new_n12749_ & new_n12821_;
  assign new_n12823_ = ~ys__n422 & new_n12822_;
  assign new_n12824_ = ys__n422 & ~new_n12822_;
  assign new_n12825_ = ~new_n12823_ & ~new_n12824_;
  assign new_n12826_ = new_n12753_ & ~new_n12825_;
  assign new_n12827_ = ~new_n12820_ & ~new_n12826_;
  assign new_n12828_ = ~new_n12811_ & new_n12827_;
  assign new_n12829_ = new_n12759_ & ~new_n12828_;
  assign new_n12830_ = ~new_n12810_ & ~new_n12829_;
  assign new_n12831_ = new_n12763_ & ~new_n12830_;
  assign new_n12832_ = ys__n38311 & new_n12768_;
  assign new_n12833_ = ~new_n12762_ & ~new_n12832_;
  assign new_n12834_ = ~new_n12831_ & new_n12833_;
  assign new_n12835_ = new_n12774_ & ~new_n12834_;
  assign new_n12836_ = new_n12776_ & ~new_n12830_;
  assign new_n12837_ = ys__n38311 & new_n12778_;
  assign new_n12838_ = ~new_n12762_ & ~new_n12837_;
  assign new_n12839_ = ~new_n12836_ & new_n12838_;
  assign new_n12840_ = new_n12784_ & ~new_n12839_;
  assign ys__n716 = new_n12835_ | new_n12840_;
  assign new_n12842_ = ys__n19203 & ys__n38178;
  assign new_n12843_ = ~new_n12212_ & ~new_n12214_;
  assign new_n12844_ = new_n12842_ & ~new_n12843_;
  assign new_n12845_ = ~ys__n1301 & ys__n1309;
  assign new_n12846_ = ~ys__n1301 & ys__n19215;
  assign new_n12847_ = ys__n19203 & new_n12215_;
  assign new_n12848_ = new_n12846_ & new_n12847_;
  assign new_n12849_ = ~new_n12845_ & ~new_n12848_;
  assign new_n12850_ = ~new_n12844_ & new_n12849_;
  assign new_n12851_ = new_n12216_ & new_n12843_;
  assign ys__n732 = ~new_n12850_ & ~new_n12851_;
  assign new_n12853_ = ~ys__n37670 & ys__n37671;
  assign new_n12854_ = ys__n37670 & ~ys__n37671;
  assign new_n12855_ = ~new_n12853_ & ~new_n12854_;
  assign new_n12856_ = ~ys__n18393 & ~new_n12855_;
  assign new_n12857_ = ~ys__n18393 & ~new_n12856_;
  assign new_n12858_ = ~ys__n18393 & ~new_n12857_;
  assign new_n12859_ = ys__n18393 & ys__n27738;
  assign new_n12860_ = ~new_n12858_ & ~new_n12859_;
  assign new_n12861_ = ys__n732 & new_n12860_;
  assign new_n12862_ = ys__n826 & ~new_n12861_;
  assign new_n12863_ = ys__n828 & new_n12861_;
  assign new_n12864_ = ~new_n12862_ & ~new_n12863_;
  assign new_n12865_ = ~ys__n732 & ~new_n12860_;
  assign new_n12866_ = ~new_n12864_ & ~new_n12865_;
  assign new_n12867_ = ys__n824 & new_n12865_;
  assign ys__n730 = new_n12866_ | new_n12867_;
  assign new_n12869_ = ~ys__n889 & ~ys__n4184;
  assign new_n12870_ = ~ys__n4192 & new_n12869_;
  assign new_n12871_ = new_n11747_ & new_n12870_;
  assign ys__n740 = ~new_n11745_ | ~new_n12871_;
  assign new_n12873_ = ys__n23641 & ~ys__n23645;
  assign new_n12874_ = ys__n23645 & ys__n23650;
  assign new_n12875_ = ~new_n12873_ & ~new_n12874_;
  assign ys__n754 = ~ys__n23652 & ~new_n12875_;
  assign new_n12877_ = ys__n23645 & ys__n23647;
  assign ys__n756 = ~ys__n23652 & new_n12877_;
  assign new_n12879_ = ys__n108 & new_n12220_;
  assign new_n12880_ = ~ys__n19203 & new_n12215_;
  assign new_n12881_ = ~new_n12200_ & ~new_n12880_;
  assign new_n12882_ = ~new_n12220_ & ~new_n12881_;
  assign ys__n786 = new_n12879_ | new_n12882_;
  assign new_n12884_ = ys__n1301 & ys__n1309;
  assign new_n12885_ = ys__n1301 & ys__n19203;
  assign new_n12886_ = ys__n19215 & new_n12885_;
  assign new_n12887_ = new_n12215_ & new_n12886_;
  assign new_n12888_ = ~new_n12884_ & ~new_n12887_;
  assign ys__n788 = ~new_n12220_ & ~new_n12888_;
  assign new_n12890_ = ys__n118 & new_n12220_;
  assign new_n12891_ = ~new_n12281_ & ~new_n12283_;
  assign new_n12892_ = ~new_n12281_ & ~new_n12891_;
  assign new_n12893_ = ~new_n12275_ & ~new_n12892_;
  assign new_n12894_ = ~new_n12275_ & ~new_n12893_;
  assign new_n12895_ = new_n12210_ & ~new_n12894_;
  assign new_n12896_ = ~ys__n19215 & ~new_n12277_;
  assign new_n12897_ = ~new_n12846_ & ~new_n12896_;
  assign new_n12898_ = new_n12847_ & ~new_n12897_;
  assign new_n12899_ = new_n12214_ & new_n12842_;
  assign new_n12900_ = ~new_n12845_ & ~new_n12899_;
  assign new_n12901_ = ~new_n12898_ & new_n12900_;
  assign new_n12902_ = ~new_n12895_ & new_n12901_;
  assign new_n12903_ = ~new_n12220_ & ~new_n12902_;
  assign ys__n790 = new_n12890_ | new_n12903_;
  assign new_n12905_ = ys__n290 & new_n12220_;
  assign new_n12906_ = ~ys__n18389 & new_n12205_;
  assign new_n12907_ = new_n12214_ & ~new_n12842_;
  assign new_n12908_ = ~ys__n308 & ~ys__n310;
  assign new_n12909_ = new_n12842_ & new_n12908_;
  assign new_n12910_ = new_n12212_ & new_n12909_;
  assign new_n12911_ = ~new_n12907_ & ~new_n12910_;
  assign new_n12912_ = ~new_n12906_ & new_n12911_;
  assign new_n12913_ = ~new_n12220_ & ~new_n12912_;
  assign ys__n792 = new_n12905_ | new_n12913_;
  assign new_n12915_ = ys__n110 & new_n12220_;
  assign new_n12916_ = new_n12842_ & ~new_n12908_;
  assign new_n12917_ = new_n12842_ & ~new_n12916_;
  assign new_n12918_ = new_n12212_ & ~new_n12917_;
  assign new_n12919_ = ys__n18389 & new_n12205_;
  assign new_n12920_ = ~new_n12918_ & ~new_n12919_;
  assign new_n12921_ = ~new_n12220_ & ~new_n12920_;
  assign ys__n794 = new_n12915_ | new_n12921_;
  assign new_n12923_ = ys__n18283 & new_n12264_;
  assign ys__n37676 = ys__n18070 | new_n12259_;
  assign new_n12925_ = ~ys__n3214 & ys__n37676;
  assign new_n12926_ = ~ys__n3214 & ~new_n12925_;
  assign new_n12927_ = ~ys__n844 & new_n12256_;
  assign new_n12928_ = ~ys__n37678 & ~ys__n37679;
  assign new_n12929_ = ys__n844 & ~new_n12928_;
  assign new_n12930_ = ys__n844 & ys__n37682;
  assign new_n12931_ = ys__n18071 & ~new_n12930_;
  assign new_n12932_ = ~new_n12929_ & new_n12931_;
  assign new_n12933_ = ~new_n12927_ & ~new_n12932_;
  assign new_n12934_ = new_n12926_ & ~new_n12933_;
  assign new_n12935_ = ~new_n12264_ & new_n12934_;
  assign new_n12936_ = ~new_n12923_ & ~new_n12935_;
  assign new_n12937_ = ~ys__n18271 & ~new_n12936_;
  assign new_n12938_ = ys__n18271 & ys__n18283;
  assign ys__n18284 = new_n12937_ | new_n12938_;
  assign new_n12940_ = ys__n18286 & new_n12264_;
  assign new_n12941_ = ys__n844 & new_n12926_;
  assign new_n12942_ = ~new_n12264_ & new_n12941_;
  assign new_n12943_ = ~new_n12934_ & new_n12942_;
  assign new_n12944_ = ~new_n12940_ & ~new_n12943_;
  assign new_n12945_ = ~ys__n18271 & ~new_n12944_;
  assign new_n12946_ = ys__n18271 & ys__n18286;
  assign ys__n18287 = new_n12945_ | new_n12946_;
  assign new_n12948_ = ys__n18984 & ys__n18287;
  assign new_n12949_ = ~ys__n18284 & new_n12948_;
  assign new_n12950_ = ys__n54 & ~ys__n4764;
  assign new_n12951_ = ys__n24667 & ys__n4764;
  assign ys__n18820 = new_n12950_ | new_n12951_;
  assign new_n12953_ = ~ys__n18071 & ys__n18820;
  assign new_n12954_ = ys__n18071 & ys__n18821;
  assign new_n12955_ = ~new_n12953_ & ~new_n12954_;
  assign new_n12956_ = ~new_n12256_ & ~new_n12955_;
  assign new_n12957_ = ys__n24667 & ~ys__n24675;
  assign new_n12958_ = ys__n24675 & ys__n24707;
  assign ys__n18738 = new_n12957_ | new_n12958_;
  assign new_n12960_ = new_n12256_ & ys__n18738;
  assign ys__n18739 = new_n12956_ | new_n12960_;
  assign new_n12962_ = ys__n18284 & ys__n18739;
  assign new_n12963_ = ~new_n12949_ & ~new_n12962_;
  assign new_n12964_ = ys__n18280 & new_n12264_;
  assign new_n12965_ = ~new_n12264_ & new_n12925_;
  assign new_n12966_ = ~new_n12964_ & ~new_n12965_;
  assign new_n12967_ = ~ys__n18271 & ~new_n12966_;
  assign new_n12968_ = ys__n18271 & ys__n18280;
  assign ys__n18281 = new_n12967_ | new_n12968_;
  assign new_n12970_ = ~new_n12963_ & ~ys__n18281;
  assign new_n12971_ = ys__n18636 & ~new_n12259_;
  assign new_n12972_ = ys__n74 & new_n12259_;
  assign ys__n18637 = new_n12971_ | new_n12972_;
  assign new_n12974_ = ys__n18281 & ys__n18637;
  assign new_n12975_ = ~new_n12970_ & ~new_n12974_;
  assign new_n12976_ = ys__n18277 & new_n12264_;
  assign new_n12977_ = ys__n3214 & ~new_n12264_;
  assign new_n12978_ = ~new_n12976_ & ~new_n12977_;
  assign new_n12979_ = ~ys__n18271 & ~new_n12978_;
  assign new_n12980_ = ys__n18271 & ys__n18277;
  assign ys__n18278 = new_n12979_ | new_n12980_;
  assign new_n12982_ = ~new_n12975_ & ~ys__n18278;
  assign new_n12983_ = ys__n18885 & ys__n18278;
  assign ys__n796 = new_n12982_ | new_n12983_;
  assign new_n12985_ = ys__n18983 & ys__n18287;
  assign new_n12986_ = ~ys__n18284 & new_n12985_;
  assign new_n12987_ = ys__n56 & ~ys__n4764;
  assign new_n12988_ = ys__n24666 & ys__n4764;
  assign ys__n18818 = new_n12987_ | new_n12988_;
  assign new_n12990_ = ~ys__n18071 & ys__n18818;
  assign new_n12991_ = ys__n18071 & ys__n18819;
  assign new_n12992_ = ~new_n12990_ & ~new_n12991_;
  assign new_n12993_ = ~new_n12256_ & ~new_n12992_;
  assign new_n12994_ = ys__n24666 & ~ys__n24675;
  assign new_n12995_ = ys__n24675 & ys__n24706;
  assign ys__n18735 = new_n12994_ | new_n12995_;
  assign new_n12997_ = new_n12256_ & ys__n18735;
  assign ys__n18736 = new_n12993_ | new_n12997_;
  assign new_n12999_ = ys__n18284 & ys__n18736;
  assign new_n13000_ = ~new_n12986_ & ~new_n12999_;
  assign new_n13001_ = ~ys__n18281 & ~new_n13000_;
  assign new_n13002_ = ys__n18634 & ~new_n12259_;
  assign new_n13003_ = ys__n76 & new_n12259_;
  assign ys__n18635 = new_n13002_ | new_n13003_;
  assign new_n13005_ = ys__n18281 & ys__n18635;
  assign new_n13006_ = ~new_n13001_ & ~new_n13005_;
  assign new_n13007_ = ~ys__n18278 & ~new_n13006_;
  assign new_n13008_ = ys__n18883 & ys__n18278;
  assign ys__n798 = new_n13007_ | new_n13008_;
  assign new_n13010_ = ys__n18982 & ys__n18287;
  assign new_n13011_ = ~ys__n18284 & new_n13010_;
  assign new_n13012_ = ys__n58 & ~ys__n4764;
  assign new_n13013_ = ys__n24665 & ys__n4764;
  assign ys__n18816 = new_n13012_ | new_n13013_;
  assign new_n13015_ = ~ys__n18071 & ys__n18816;
  assign new_n13016_ = ys__n18071 & ys__n18817;
  assign new_n13017_ = ~new_n13015_ & ~new_n13016_;
  assign new_n13018_ = ~new_n12256_ & ~new_n13017_;
  assign new_n13019_ = ys__n24665 & ~ys__n24675;
  assign new_n13020_ = ys__n24675 & ys__n24705;
  assign ys__n18732 = new_n13019_ | new_n13020_;
  assign new_n13022_ = new_n12256_ & ys__n18732;
  assign ys__n18733 = new_n13018_ | new_n13022_;
  assign new_n13024_ = ys__n18284 & ys__n18733;
  assign new_n13025_ = ~new_n13011_ & ~new_n13024_;
  assign new_n13026_ = ~ys__n18281 & ~new_n13025_;
  assign new_n13027_ = ys__n18632 & ~new_n12259_;
  assign new_n13028_ = ys__n78 & new_n12259_;
  assign ys__n18633 = new_n13027_ | new_n13028_;
  assign new_n13030_ = ys__n18281 & ys__n18633;
  assign new_n13031_ = ~new_n13026_ & ~new_n13030_;
  assign new_n13032_ = ~ys__n18278 & ~new_n13031_;
  assign new_n13033_ = ys__n18881 & ys__n18278;
  assign ys__n800 = new_n13032_ | new_n13033_;
  assign new_n13035_ = ys__n18981 & ys__n18287;
  assign new_n13036_ = ~ys__n18284 & new_n13035_;
  assign new_n13037_ = ys__n60 & ~ys__n4764;
  assign new_n13038_ = ys__n24664 & ys__n4764;
  assign ys__n18814 = new_n13037_ | new_n13038_;
  assign new_n13040_ = ~ys__n18071 & ys__n18814;
  assign new_n13041_ = ys__n18071 & ys__n18815;
  assign new_n13042_ = ~new_n13040_ & ~new_n13041_;
  assign new_n13043_ = ~new_n12256_ & ~new_n13042_;
  assign new_n13044_ = ys__n24664 & ~ys__n24675;
  assign new_n13045_ = ys__n24675 & ys__n24704;
  assign ys__n18729 = new_n13044_ | new_n13045_;
  assign new_n13047_ = new_n12256_ & ys__n18729;
  assign ys__n18730 = new_n13043_ | new_n13047_;
  assign new_n13049_ = ys__n18284 & ys__n18730;
  assign new_n13050_ = ~new_n13036_ & ~new_n13049_;
  assign new_n13051_ = ~ys__n18281 & ~new_n13050_;
  assign new_n13052_ = ys__n18630 & ~new_n12259_;
  assign new_n13053_ = ys__n70 & new_n12259_;
  assign ys__n18631 = new_n13052_ | new_n13053_;
  assign new_n13055_ = ys__n18281 & ys__n18631;
  assign new_n13056_ = ~new_n13051_ & ~new_n13055_;
  assign new_n13057_ = ~ys__n18278 & ~new_n13056_;
  assign new_n13058_ = ys__n18879 & ys__n18278;
  assign ys__n802 = new_n13057_ | new_n13058_;
  assign new_n13060_ = ys__n18980 & ys__n18287;
  assign new_n13061_ = ~ys__n18284 & new_n13060_;
  assign new_n13062_ = ys__n62 & ~ys__n4764;
  assign new_n13063_ = ys__n24663 & ys__n4764;
  assign ys__n18812 = new_n13062_ | new_n13063_;
  assign new_n13065_ = ~ys__n18071 & ys__n18812;
  assign new_n13066_ = ys__n18071 & ys__n18813;
  assign new_n13067_ = ~new_n13065_ & ~new_n13066_;
  assign new_n13068_ = ~new_n12256_ & ~new_n13067_;
  assign new_n13069_ = ys__n24663 & ~ys__n24675;
  assign new_n13070_ = ys__n24675 & ys__n24703;
  assign ys__n18726 = new_n13069_ | new_n13070_;
  assign new_n13072_ = new_n12256_ & ys__n18726;
  assign ys__n18727 = new_n13068_ | new_n13072_;
  assign new_n13074_ = ys__n18284 & ys__n18727;
  assign new_n13075_ = ~new_n13061_ & ~new_n13074_;
  assign new_n13076_ = ~ys__n18281 & ~new_n13075_;
  assign new_n13077_ = ys__n18628 & ~new_n12259_;
  assign new_n13078_ = ys__n72 & new_n12259_;
  assign ys__n18629 = new_n13077_ | new_n13078_;
  assign new_n13080_ = ys__n18281 & ys__n18629;
  assign new_n13081_ = ~new_n13076_ & ~new_n13080_;
  assign new_n13082_ = ~ys__n18278 & ~new_n13081_;
  assign new_n13083_ = ys__n18877 & ys__n18278;
  assign ys__n804 = new_n13082_ | new_n13083_;
  assign new_n13085_ = ys__n18977 & ys__n18287;
  assign new_n13086_ = ~ys__n18284 & new_n13085_;
  assign new_n13087_ = ys__n24657 & ~ys__n4764;
  assign new_n13088_ = ys__n24658 & ys__n4764;
  assign ys__n18806 = new_n13087_ | new_n13088_;
  assign new_n13090_ = ~ys__n18071 & ys__n18806;
  assign new_n13091_ = ys__n18071 & ys__n18807;
  assign new_n13092_ = ~new_n13090_ & ~new_n13091_;
  assign new_n13093_ = ~new_n12256_ & ~new_n13092_;
  assign new_n13094_ = ys__n24658 & ~ys__n24675;
  assign new_n13095_ = ys__n24675 & ys__n24700;
  assign ys__n18717 = new_n13094_ | new_n13095_;
  assign new_n13097_ = new_n12256_ & ys__n18717;
  assign ys__n18718 = new_n13093_ | new_n13097_;
  assign new_n13099_ = ys__n18284 & ys__n18718;
  assign new_n13100_ = ~new_n13086_ & ~new_n13099_;
  assign new_n13101_ = ~ys__n18281 & ~new_n13100_;
  assign new_n13102_ = ys__n18619 & ~new_n12259_;
  assign new_n13103_ = ys__n18620 & new_n12259_;
  assign ys__n18621 = new_n13102_ | new_n13103_;
  assign new_n13105_ = ys__n18281 & ys__n18621;
  assign new_n13106_ = ~new_n13101_ & ~new_n13105_;
  assign new_n13107_ = ~ys__n18278 & ~new_n13106_;
  assign new_n13108_ = ys__n18871 & ys__n18278;
  assign ys__n806 = new_n13107_ | new_n13108_;
  assign new_n13110_ = ys__n18986 & ys__n18287;
  assign new_n13111_ = ~ys__n18284 & new_n13110_;
  assign new_n13112_ = ys__n24670 & ~ys__n4764;
  assign new_n13113_ = ys__n24671 & ys__n4764;
  assign ys__n18824 = new_n13112_ | new_n13113_;
  assign new_n13115_ = ~ys__n18071 & ys__n18824;
  assign new_n13116_ = ys__n18071 & ys__n18825;
  assign new_n13117_ = ~new_n13115_ & ~new_n13116_;
  assign new_n13118_ = ~new_n12256_ & ~new_n13117_;
  assign new_n13119_ = ys__n24671 & ~ys__n24675;
  assign new_n13120_ = ys__n24675 & ys__n24709;
  assign ys__n18744 = new_n13119_ | new_n13120_;
  assign new_n13122_ = new_n12256_ & ys__n18744;
  assign ys__n18745 = new_n13118_ | new_n13122_;
  assign new_n13124_ = ys__n18284 & ys__n18745;
  assign new_n13125_ = ~new_n13111_ & ~new_n13124_;
  assign new_n13126_ = ~ys__n18281 & ~new_n13125_;
  assign new_n13127_ = ys__n18641 & ~new_n12259_;
  assign new_n13128_ = ys__n18642 & new_n12259_;
  assign ys__n18643 = new_n13127_ | new_n13128_;
  assign new_n13130_ = ys__n18281 & ys__n18643;
  assign new_n13131_ = ~new_n13126_ & ~new_n13130_;
  assign new_n13132_ = ~ys__n18278 & ~new_n13131_;
  assign new_n13133_ = ys__n18889 & ys__n18278;
  assign ys__n808 = new_n13132_ | new_n13133_;
  assign new_n13135_ = ys__n18985 & ys__n18287;
  assign new_n13136_ = ~ys__n18284 & new_n13135_;
  assign new_n13137_ = ys__n24668 & ~ys__n4764;
  assign new_n13138_ = ys__n24669 & ys__n4764;
  assign ys__n18822 = new_n13137_ | new_n13138_;
  assign new_n13140_ = ~ys__n18071 & ys__n18822;
  assign new_n13141_ = ys__n18071 & ys__n18823;
  assign new_n13142_ = ~new_n13140_ & ~new_n13141_;
  assign new_n13143_ = ~new_n12256_ & ~new_n13142_;
  assign new_n13144_ = ys__n24669 & ~ys__n24675;
  assign new_n13145_ = ys__n24675 & ys__n24708;
  assign ys__n18741 = new_n13144_ | new_n13145_;
  assign new_n13147_ = new_n12256_ & ys__n18741;
  assign ys__n18742 = new_n13143_ | new_n13147_;
  assign new_n13149_ = ys__n18284 & ys__n18742;
  assign new_n13150_ = ~new_n13136_ & ~new_n13149_;
  assign new_n13151_ = ~ys__n18281 & ~new_n13150_;
  assign new_n13152_ = ys__n18638 & ~new_n12259_;
  assign new_n13153_ = ys__n18639 & new_n12259_;
  assign ys__n18640 = new_n13152_ | new_n13153_;
  assign new_n13155_ = ys__n18281 & ys__n18640;
  assign new_n13156_ = ~new_n13151_ & ~new_n13155_;
  assign new_n13157_ = ~ys__n18278 & ~new_n13156_;
  assign new_n13158_ = ys__n18887 & ys__n18278;
  assign ys__n810 = new_n13157_ | new_n13158_;
  assign new_n13160_ = ys__n18987 & ys__n18287;
  assign new_n13161_ = ~ys__n18284 & new_n13160_;
  assign new_n13162_ = ys__n24672 & ~ys__n4764;
  assign new_n13163_ = ys__n24673 & ys__n4764;
  assign ys__n18826 = new_n13162_ | new_n13163_;
  assign new_n13165_ = ~ys__n18071 & ys__n18826;
  assign new_n13166_ = ys__n18071 & ys__n18827;
  assign new_n13167_ = ~new_n13165_ & ~new_n13166_;
  assign new_n13168_ = ~new_n12256_ & ~new_n13167_;
  assign new_n13169_ = ys__n24673 & ~ys__n24675;
  assign new_n13170_ = ys__n24675 & ys__n24710;
  assign ys__n18747 = new_n13169_ | new_n13170_;
  assign new_n13172_ = new_n12256_ & ys__n18747;
  assign ys__n18748 = new_n13168_ | new_n13172_;
  assign new_n13174_ = ys__n18284 & ys__n18748;
  assign new_n13175_ = ~new_n13161_ & ~new_n13174_;
  assign new_n13176_ = ~ys__n18281 & ~new_n13175_;
  assign new_n13177_ = ys__n18644 & ~new_n12259_;
  assign new_n13178_ = ys__n18645 & new_n12259_;
  assign ys__n18646 = new_n13177_ | new_n13178_;
  assign new_n13180_ = ys__n18281 & ys__n18646;
  assign new_n13181_ = ~new_n13176_ & ~new_n13180_;
  assign new_n13182_ = ~ys__n18278 & ~new_n13181_;
  assign new_n13183_ = ys__n18891 & ys__n18278;
  assign ys__n812 = new_n13182_ | new_n13183_;
  assign new_n13185_ = ys__n20273 & ys__n738;
  assign ys__n814 = ~new_n12020_ & new_n13185_;
  assign new_n13187_ = ys__n29896 & ~new_n11737_;
  assign new_n13188_ = ~new_n11735_ & new_n13187_;
  assign new_n13189_ = ~ys__n23764 & new_n13188_;
  assign new_n13190_ = ys__n29912 & ~new_n11737_;
  assign new_n13191_ = ~new_n11735_ & new_n13190_;
  assign new_n13192_ = ~ys__n22466 & new_n13191_;
  assign new_n13193_ = ys__n22466 & new_n13188_;
  assign new_n13194_ = ~new_n13192_ & ~new_n13193_;
  assign new_n13195_ = ys__n23764 & ~new_n13194_;
  assign new_n13196_ = ~new_n13189_ & ~new_n13195_;
  assign new_n13197_ = ~new_n11993_ & ~new_n13196_;
  assign new_n13198_ = ys__n23764 & ~new_n11998_;
  assign new_n13199_ = ~new_n13197_ & ~new_n13198_;
  assign ys__n25435 = ~new_n11999_ & ~new_n13199_;
  assign new_n13201_ = ~ys__n19256 & ys__n25435;
  assign new_n13202_ = ys__n634 & ys__n19256;
  assign new_n13203_ = ~new_n13201_ & ~new_n13202_;
  assign new_n13204_ = ys__n874 & ~new_n13203_;
  assign ys__n862 = ys__n2 | ~new_n13204_;
  assign new_n13206_ = ys__n37703 & ~new_n12255_;
  assign new_n13207_ = ~ys__n37674 & ys__n37675;
  assign new_n13208_ = ys__n37674 & ~ys__n37675;
  assign new_n13209_ = ~new_n13207_ & ~new_n13208_;
  assign new_n13210_ = ~ys__n18393 & ~new_n13209_;
  assign new_n13211_ = ys__n18393 & new_n12283_;
  assign new_n13212_ = ~new_n12281_ & new_n13211_;
  assign new_n13213_ = ~new_n12281_ & ~new_n13212_;
  assign new_n13214_ = new_n12210_ & ~new_n12275_;
  assign new_n13215_ = ~new_n13213_ & new_n13214_;
  assign new_n13216_ = ys__n18393 & ys__n19203;
  assign new_n13217_ = ~ys__n19215 & new_n13216_;
  assign new_n13218_ = new_n12215_ & new_n13217_;
  assign new_n13219_ = new_n12277_ & new_n13218_;
  assign new_n13220_ = ~ys__n18393 & ~new_n12206_;
  assign new_n13221_ = ~new_n13219_ & ~new_n13220_;
  assign new_n13222_ = ~new_n13215_ & new_n13221_;
  assign new_n13223_ = ~new_n12210_ & ~new_n12215_;
  assign new_n13224_ = new_n12206_ & new_n13223_;
  assign ys__n27605 = ~new_n13222_ & ~new_n13224_;
  assign new_n13226_ = ys__n18393 & ys__n27605;
  assign new_n13227_ = ~new_n13210_ & ~new_n13226_;
  assign new_n13228_ = ys__n33300 & ys__n37692;
  assign new_n13229_ = new_n13227_ & ~new_n13228_;
  assign new_n13230_ = ~ys__n18317 & ~new_n13229_;
  assign new_n13231_ = ~ys__n33300 & ~ys__n37694;
  assign new_n13232_ = ~ys__n37696 & new_n13227_;
  assign new_n13233_ = ~new_n13231_ & ~new_n13232_;
  assign new_n13234_ = ys__n18271 & ys__n37692;
  assign new_n13235_ = ~new_n13233_ & ~new_n13234_;
  assign new_n13236_ = ys__n18317 & ~new_n13235_;
  assign new_n13237_ = ~new_n13230_ & ~new_n13236_;
  assign new_n13238_ = ~ys__n33309 & ~ys__n33311;
  assign new_n13239_ = ~ys__n33313 & new_n13238_;
  assign new_n13240_ = ~new_n13237_ & new_n13239_;
  assign ys__n863 = new_n13206_ & ~new_n13240_;
  assign new_n13242_ = ~new_n13206_ & new_n13240_;
  assign ys__n865 = ys__n863 | new_n13242_;
  assign ys__n866 = ~ys__n2 | new_n13204_;
  assign new_n13245_ = ys__n29895 & ~new_n11737_;
  assign new_n13246_ = ~new_n11735_ & new_n13245_;
  assign new_n13247_ = ~ys__n23764 & new_n13246_;
  assign new_n13248_ = ys__n29911 & ~new_n11737_;
  assign new_n13249_ = ~new_n11735_ & new_n13248_;
  assign new_n13250_ = ~ys__n22466 & new_n13249_;
  assign new_n13251_ = ys__n22466 & new_n13246_;
  assign new_n13252_ = ~new_n13250_ & ~new_n13251_;
  assign new_n13253_ = ys__n23764 & ~new_n13252_;
  assign new_n13254_ = ~new_n13247_ & ~new_n13253_;
  assign new_n13255_ = ~new_n11993_ & ~new_n13254_;
  assign new_n13256_ = ~new_n13198_ & ~new_n13255_;
  assign ys__n25434 = ~new_n11999_ & ~new_n13256_;
  assign new_n13258_ = ~ys__n19256 & ys__n25434;
  assign new_n13259_ = ys__n636 & ys__n19256;
  assign new_n13260_ = ~new_n13258_ & ~new_n13259_;
  assign new_n13261_ = ys__n874 & ~new_n13260_;
  assign ys__n868 = ys__n866 | new_n13261_;
  assign new_n13263_ = ys__n29894 & ~new_n11737_;
  assign new_n13264_ = ~new_n11735_ & new_n13263_;
  assign new_n13265_ = ~ys__n23764 & new_n13264_;
  assign new_n13266_ = ys__n29910 & ~new_n11737_;
  assign new_n13267_ = ~new_n11735_ & new_n13266_;
  assign new_n13268_ = ~ys__n22466 & new_n13267_;
  assign new_n13269_ = ys__n22466 & new_n13264_;
  assign new_n13270_ = ~new_n13268_ & ~new_n13269_;
  assign new_n13271_ = ys__n23764 & ~new_n13270_;
  assign new_n13272_ = ~new_n13265_ & ~new_n13271_;
  assign ys__n25433 = new_n12000_ & ~new_n13272_;
  assign new_n13274_ = ~ys__n19256 & ys__n25433;
  assign new_n13275_ = ys__n638 & ys__n19256;
  assign new_n13276_ = ~new_n13274_ & ~new_n13275_;
  assign new_n13277_ = ys__n874 & ~new_n13276_;
  assign new_n13278_ = new_n13261_ & new_n13277_;
  assign ys__n870 = ys__n862 | ~new_n13278_;
  assign new_n13280_ = ys__n18120 & ~ys__n740;
  assign ys__n871 = ~ys__n874 | new_n13280_;
  assign new_n13282_ = ~ys__n140 & ~ys__n214;
  assign new_n13283_ = ys__n216 & ~ys__n218;
  assign new_n13284_ = new_n13282_ & new_n13283_;
  assign new_n13285_ = ~ys__n216 & ys__n218;
  assign new_n13286_ = new_n13282_ & new_n13285_;
  assign new_n13287_ = ~new_n13284_ & ~new_n13286_;
  assign new_n13288_ = ~ys__n216 & ~ys__n218;
  assign new_n13289_ = ~ys__n140 & ys__n214;
  assign new_n13290_ = new_n13288_ & new_n13289_;
  assign new_n13291_ = new_n13287_ & ~new_n13290_;
  assign ys__n872 = ys__n871 | new_n13291_;
  assign new_n13293_ = ~ys__n140 & ~ys__n210;
  assign new_n13294_ = ys__n66 & ~ys__n212;
  assign new_n13295_ = new_n13293_ & new_n13294_;
  assign new_n13296_ = ~ys__n66 & ys__n212;
  assign new_n13297_ = new_n13293_ & new_n13296_;
  assign new_n13298_ = ~new_n13295_ & ~new_n13297_;
  assign new_n13299_ = ~ys__n66 & ~ys__n212;
  assign new_n13300_ = ~ys__n140 & ys__n210;
  assign new_n13301_ = new_n13299_ & new_n13300_;
  assign new_n13302_ = new_n13298_ & ~new_n13301_;
  assign ys__n873 = ys__n871 | new_n13302_;
  assign new_n13304_ = ~ys__n140 & ~ys__n298;
  assign new_n13305_ = ~ys__n300 & ys__n302;
  assign new_n13306_ = new_n13304_ & new_n13305_;
  assign new_n13307_ = ~ys__n140 & ~ys__n302;
  assign new_n13308_ = ~ys__n298 & ys__n300;
  assign new_n13309_ = new_n13307_ & new_n13308_;
  assign new_n13310_ = ys__n298 & ~ys__n300;
  assign new_n13311_ = new_n13307_ & new_n13310_;
  assign new_n13312_ = ~new_n13309_ & ~new_n13311_;
  assign new_n13313_ = ~new_n13306_ & new_n13312_;
  assign ys__n876 = ys__n874 & ~new_n13313_;
  assign new_n13315_ = ~ys__n140 & ~ys__n580;
  assign new_n13316_ = ~ys__n582 & ys__n584;
  assign new_n13317_ = new_n13315_ & new_n13316_;
  assign new_n13318_ = ~ys__n140 & ~ys__n584;
  assign new_n13319_ = ~ys__n580 & ys__n582;
  assign new_n13320_ = new_n13318_ & new_n13319_;
  assign new_n13321_ = ys__n580 & ~ys__n582;
  assign new_n13322_ = new_n13318_ & new_n13321_;
  assign new_n13323_ = ~new_n13320_ & ~new_n13322_;
  assign new_n13324_ = ~new_n13317_ & new_n13323_;
  assign ys__n878 = ys__n874 & ~new_n13324_;
  assign new_n13326_ = ~ys__n138 & ~ys__n140;
  assign new_n13327_ = ~ys__n120 & ys__n142;
  assign new_n13328_ = new_n13326_ & new_n13327_;
  assign new_n13329_ = ys__n120 & ~ys__n142;
  assign new_n13330_ = new_n13326_ & new_n13329_;
  assign new_n13331_ = ~new_n13328_ & ~new_n13330_;
  assign new_n13332_ = ~ys__n120 & ~ys__n142;
  assign new_n13333_ = ys__n138 & ~ys__n140;
  assign new_n13334_ = new_n13332_ & new_n13333_;
  assign new_n13335_ = new_n13331_ & ~new_n13334_;
  assign ys__n879 = ys__n871 | new_n13335_;
  assign new_n13337_ = ~ys__n140 & ~ys__n392;
  assign new_n13338_ = ~ys__n394 & ys__n396;
  assign new_n13339_ = new_n13337_ & new_n13338_;
  assign new_n13340_ = ~ys__n140 & ~ys__n396;
  assign new_n13341_ = ~ys__n392 & ys__n394;
  assign new_n13342_ = new_n13340_ & new_n13341_;
  assign new_n13343_ = ys__n392 & ~ys__n394;
  assign new_n13344_ = new_n13340_ & new_n13343_;
  assign new_n13345_ = ~new_n13342_ & ~new_n13344_;
  assign new_n13346_ = ~new_n13339_ & new_n13345_;
  assign ys__n881 = ys__n874 & ~new_n13346_;
  assign new_n13348_ = ~ys__n2779 & ~ys__n30816;
  assign new_n13349_ = ys__n30819 & new_n13348_;
  assign new_n13350_ = ys__n30815 & ys__n30816;
  assign new_n13351_ = ~new_n13349_ & ~new_n13350_;
  assign new_n13352_ = ~ys__n562 & ~new_n13351_;
  assign new_n13353_ = ys__n562 & new_n13351_;
  assign ys__n888 = new_n13352_ | new_n13353_;
  assign new_n13355_ = ~ys__n846 & ys__n874;
  assign new_n13356_ = ~ys__n889 & new_n13355_;
  assign new_n13357_ = ~ys__n4184 & ~ys__n4185;
  assign new_n13358_ = new_n12181_ & new_n13357_;
  assign new_n13359_ = ~ys__n4176 & ~ys__n4627;
  assign new_n13360_ = ~ys__n4177 & ~ys__n4698;
  assign new_n13361_ = new_n13359_ & new_n13360_;
  assign new_n13362_ = new_n13358_ & new_n13361_;
  assign ys__n900 = ~new_n13356_ | ~new_n13362_;
  assign ys__n902 = ~ys__n874 | ~new_n13237_;
  assign ys__n904 = ys__n30223 | ~ys__n740;
  assign new_n13366_ = ys__n38305 & ~ys__n738;
  assign ys__n911 = ~ys__n4566 & new_n13366_;
  assign new_n13368_ = ys__n30820 & new_n13348_;
  assign new_n13369_ = ys__n30816 & ys__n30818;
  assign new_n13370_ = ~new_n13368_ & ~new_n13369_;
  assign new_n13371_ = ~ys__n398 & ~new_n13370_;
  assign new_n13372_ = ys__n398 & new_n13370_;
  assign ys__n920 = new_n13371_ | new_n13372_;
  assign new_n13374_ = ys__n172 & ys__n338;
  assign new_n13375_ = ~ys__n172 & ~ys__n338;
  assign new_n13376_ = ~ys__n172 & ys__n338;
  assign new_n13377_ = ~new_n13375_ & ~new_n13376_;
  assign new_n13378_ = ~new_n13374_ & new_n13377_;
  assign new_n13379_ = ys__n22 & ~ys__n316;
  assign new_n13380_ = ~ys__n22 & ~ys__n316;
  assign new_n13381_ = ~new_n13379_ & ~new_n13380_;
  assign new_n13382_ = ~ys__n22 & ys__n316;
  assign new_n13383_ = new_n13381_ & ~new_n13382_;
  assign new_n13384_ = ys__n172 & ~ys__n338;
  assign new_n13385_ = ~new_n13383_ & new_n13384_;
  assign new_n13386_ = new_n13378_ & ~new_n13385_;
  assign new_n13387_ = ~ys__n35047 & ys__n46240;
  assign new_n13388_ = ~ys__n46230 & ys__n46239;
  assign new_n13389_ = ys__n46230 & ~ys__n46239;
  assign new_n13390_ = ~new_n13388_ & ~new_n13389_;
  assign new_n13391_ = ys__n46238 & ~new_n13390_;
  assign ys__n18210 = new_n13387_ | new_n13391_;
  assign new_n13393_ = ~ys__n44 & ys__n6115;
  assign new_n13394_ = ~ys__n44 & ~new_n13393_;
  assign new_n13395_ = ~ys__n18208 & new_n13394_;
  assign new_n13396_ = ys__n18210 & new_n13395_;
  assign new_n13397_ = ~ys__n6120 & ~ys__n6121;
  assign new_n13398_ = ~ys__n6123 & ~ys__n6124;
  assign new_n13399_ = new_n13397_ & new_n13398_;
  assign new_n13400_ = ~ys__n6118 & ~ys__n6119;
  assign new_n13401_ = ys__n46 & ~ys__n340;
  assign new_n13402_ = ys__n18317 & new_n13401_;
  assign new_n13403_ = new_n13400_ & new_n13402_;
  assign new_n13404_ = new_n13399_ & new_n13403_;
  assign new_n13405_ = ys__n40 & ys__n42;
  assign new_n13406_ = ~ys__n6133 & ~ys__n6134;
  assign new_n13407_ = new_n13405_ & new_n13406_;
  assign new_n13408_ = ~ys__n6126 & ~ys__n6127;
  assign new_n13409_ = ~ys__n6129 & ~ys__n6130;
  assign new_n13410_ = new_n13408_ & new_n13409_;
  assign new_n13411_ = new_n13407_ & new_n13410_;
  assign new_n13412_ = ys__n32 & ys__n34;
  assign new_n13413_ = ys__n36 & ys__n38;
  assign new_n13414_ = new_n13412_ & new_n13413_;
  assign new_n13415_ = ys__n24 & ys__n26;
  assign new_n13416_ = ys__n28 & ys__n30;
  assign new_n13417_ = new_n13415_ & new_n13416_;
  assign new_n13418_ = new_n13414_ & new_n13417_;
  assign new_n13419_ = new_n13411_ & new_n13418_;
  assign new_n13420_ = new_n13404_ & new_n13419_;
  assign new_n13421_ = new_n13396_ & new_n13420_;
  assign ys__n923 = new_n13386_ & new_n13421_;
  assign new_n13423_ = ys__n38307 & ~ys__n738;
  assign ys__n927 = ~ys__n4566 & new_n13423_;
  assign new_n13425_ = ys__n754 & ys__n756;
  assign new_n13426_ = ~ys__n738 & new_n13425_;
  assign new_n13427_ = ys__n478 & new_n13426_;
  assign new_n13428_ = ys__n482 & new_n13427_;
  assign ys__n929 = ~ys__n480 & new_n13428_;
  assign ys__n930 = ~ys__n738 & ys__n478;
  assign new_n13431_ = ys__n38220 & ~ys__n4566;
  assign new_n13432_ = ~ys__n935 & ~new_n13431_;
  assign ys__n932 = ~ys__n738 & ~new_n13432_;
  assign new_n13434_ = ys__n38221 & ~ys__n738;
  assign ys__n934 = ~ys__n4566 & new_n13434_;
  assign ys__n936 = ys__n935 & ~ys__n738;
  assign new_n13437_ = ~ys__n38407 & ~ys__n38408;
  assign new_n13438_ = ~ys__n226 & new_n13437_;
  assign new_n13439_ = ys__n478 & new_n13438_;
  assign new_n13440_ = ys__n226 & ys__n478;
  assign new_n13441_ = ~ys__n226 & ~new_n13437_;
  assign new_n13442_ = ys__n478 & new_n13441_;
  assign new_n13443_ = ~new_n13440_ & ~new_n13442_;
  assign new_n13444_ = ~new_n13439_ & new_n13443_;
  assign ys__n942 = ~ys__n738 & ~new_n13444_;
  assign new_n13446_ = ys__n326 & ~ys__n332;
  assign new_n13447_ = ~ys__n328 & ~ys__n330;
  assign new_n13448_ = ~ys__n336 & new_n13447_;
  assign new_n13449_ = new_n13446_ & new_n13448_;
  assign new_n13450_ = ys__n328 & ~ys__n330;
  assign new_n13451_ = ~ys__n336 & new_n13446_;
  assign new_n13452_ = new_n13450_ & new_n13451_;
  assign new_n13453_ = ~new_n13449_ & ~new_n13452_;
  assign new_n13454_ = ~ys__n328 & ys__n330;
  assign new_n13455_ = new_n13451_ & new_n13454_;
  assign new_n13456_ = ys__n328 & ys__n330;
  assign new_n13457_ = new_n13451_ & new_n13456_;
  assign new_n13458_ = ~new_n13455_ & ~new_n13457_;
  assign new_n13459_ = new_n13453_ & new_n13458_;
  assign new_n13460_ = ys__n326 & ys__n332;
  assign new_n13461_ = ys__n336 & new_n13460_;
  assign new_n13462_ = new_n13456_ & new_n13461_;
  assign new_n13463_ = new_n13459_ & ~new_n13462_;
  assign ys__n944 = ys__n602 & ~new_n13463_;
  assign new_n13465_ = ~ys__n4176 & new_n11747_;
  assign new_n13466_ = new_n11743_ & new_n13465_;
  assign new_n13467_ = new_n11742_ & new_n13466_;
  assign ys__n30832 = ys__n4698 | ~new_n13467_;
  assign ys__n948 = ~ys__n4566 & ~ys__n30832;
  assign new_n13470_ = ~ys__n160 & ys__n344;
  assign new_n13471_ = ys__n342 & ys__n350;
  assign new_n13472_ = new_n13470_ & new_n13471_;
  assign new_n13473_ = ys__n348 & ~ys__n2924;
  assign new_n13474_ = ~ys__n162 & ~ys__n346;
  assign new_n13475_ = new_n13473_ & new_n13474_;
  assign new_n13476_ = ys__n352 & new_n13475_;
  assign new_n13477_ = new_n13472_ & new_n13476_;
  assign new_n13478_ = ~ys__n342 & ys__n350;
  assign new_n13479_ = new_n13470_ & new_n13478_;
  assign new_n13480_ = ys__n352 & new_n13479_;
  assign new_n13481_ = new_n13475_ & new_n13480_;
  assign new_n13482_ = ys__n162 & ys__n346;
  assign new_n13483_ = new_n13473_ & new_n13482_;
  assign new_n13484_ = new_n13480_ & new_n13483_;
  assign new_n13485_ = ~new_n13481_ & ~new_n13484_;
  assign new_n13486_ = ~new_n13477_ & new_n13485_;
  assign ys__n949 = ys__n948 & ~new_n13486_;
  assign new_n13488_ = ~new_n13375_ & ~new_n13384_;
  assign new_n13489_ = ~new_n13376_ & new_n13488_;
  assign new_n13490_ = ys__n22 & ys__n316;
  assign new_n13491_ = ~new_n13380_ & ~new_n13382_;
  assign new_n13492_ = ~new_n13490_ & new_n13491_;
  assign new_n13493_ = new_n13374_ & ~new_n13492_;
  assign new_n13494_ = new_n13489_ & ~new_n13493_;
  assign new_n13495_ = ys__n46 & ys__n340;
  assign new_n13496_ = ys__n18317 & new_n13495_;
  assign new_n13497_ = new_n13400_ & new_n13496_;
  assign new_n13498_ = new_n13399_ & new_n13497_;
  assign new_n13499_ = new_n13419_ & new_n13498_;
  assign new_n13500_ = new_n13396_ & new_n13499_;
  assign ys__n970 = new_n13494_ & new_n13500_;
  assign new_n13502_ = ~new_n13379_ & ~new_n13382_;
  assign new_n13503_ = ~new_n13490_ & new_n13502_;
  assign new_n13504_ = new_n13374_ & ~new_n13503_;
  assign new_n13505_ = new_n13489_ & ~new_n13504_;
  assign ys__n972 = new_n13500_ & new_n13505_;
  assign new_n13507_ = new_n13381_ & ~new_n13490_;
  assign new_n13508_ = new_n13374_ & ~new_n13507_;
  assign new_n13509_ = new_n13489_ & ~new_n13508_;
  assign ys__n974 = new_n13500_ & new_n13509_;
  assign new_n13511_ = ~new_n13376_ & ~new_n13384_;
  assign new_n13512_ = ~new_n13374_ & new_n13511_;
  assign new_n13513_ = new_n13375_ & ~new_n13503_;
  assign new_n13514_ = new_n13512_ & ~new_n13513_;
  assign ys__n976 = new_n13500_ & new_n13514_;
  assign new_n13516_ = new_n13375_ & ~new_n13492_;
  assign new_n13517_ = new_n13512_ & ~new_n13516_;
  assign ys__n978 = new_n13500_ & new_n13517_;
  assign new_n13519_ = new_n13374_ & ~new_n13383_;
  assign new_n13520_ = new_n13489_ & ~new_n13519_;
  assign ys__n980 = new_n13500_ & new_n13520_;
  assign new_n13522_ = new_n13384_ & ~new_n13503_;
  assign new_n13523_ = new_n13378_ & ~new_n13522_;
  assign ys__n982 = new_n13500_ & new_n13523_;
  assign new_n13525_ = ~ys__n46 & ys__n340;
  assign new_n13526_ = ys__n18317 & new_n13525_;
  assign new_n13527_ = new_n13400_ & new_n13526_;
  assign new_n13528_ = new_n13399_ & new_n13527_;
  assign new_n13529_ = new_n13419_ & new_n13528_;
  assign new_n13530_ = new_n13396_ & new_n13529_;
  assign new_n13531_ = new_n13375_ & new_n13383_;
  assign ys__n989 = new_n13530_ & new_n13531_;
  assign ys__n991 = new_n13386_ & new_n13500_;
  assign new_n13534_ = new_n13384_ & ~new_n13507_;
  assign new_n13535_ = new_n13378_ & ~new_n13534_;
  assign ys__n993 = new_n13500_ & new_n13535_;
  assign new_n13537_ = new_n13375_ & ~new_n13383_;
  assign new_n13538_ = new_n13512_ & ~new_n13537_;
  assign ys__n995 = new_n13500_ & new_n13538_;
  assign new_n13540_ = new_n13376_ & ~new_n13492_;
  assign new_n13541_ = ~new_n13374_ & new_n13488_;
  assign new_n13542_ = ~new_n13540_ & new_n13541_;
  assign ys__n999 = new_n13500_ & new_n13542_;
  assign new_n13544_ = new_n13376_ & ~new_n13503_;
  assign new_n13545_ = new_n13541_ & ~new_n13544_;
  assign ys__n1001 = new_n13500_ & new_n13545_;
  assign new_n13547_ = new_n13376_ & ~new_n13383_;
  assign new_n13548_ = new_n13541_ & ~new_n13547_;
  assign ys__n1004 = new_n13500_ & new_n13548_;
  assign new_n13550_ = new_n13376_ & ~new_n13507_;
  assign new_n13551_ = new_n13541_ & ~new_n13550_;
  assign ys__n1007 = new_n13500_ & new_n13551_;
  assign new_n13553_ = new_n13375_ & ~new_n13507_;
  assign new_n13554_ = new_n13512_ & ~new_n13553_;
  assign ys__n1009 = new_n13500_ & new_n13554_;
  assign new_n13556_ = new_n13384_ & ~new_n13492_;
  assign new_n13557_ = new_n13378_ & ~new_n13556_;
  assign ys__n1013 = new_n13500_ & new_n13557_;
  assign new_n13559_ = ys__n1020 & new_n13290_;
  assign new_n13560_ = ~ys__n30223 & new_n13286_;
  assign ys__n16191 = new_n13559_ | new_n13560_;
  assign new_n13562_ = ys__n740 & new_n13284_;
  assign new_n13563_ = ~ys__n1020 & ~ys__n740;
  assign new_n13564_ = ~ys__n1020 & new_n13290_;
  assign new_n13565_ = ~new_n13563_ & new_n13564_;
  assign new_n13566_ = ~new_n13562_ & ~new_n13565_;
  assign ys__n1028 = ~ys__n16191 & new_n13566_;
  assign new_n13568_ = ~ys__n18121 & ~ys__n18122;
  assign ys__n1030 = ys__n18124 & ~new_n13568_;
  assign ys__n1031 = ys__n1029 | ys__n1030;
  assign ys__n1032 = ~ys__n874 | ys__n1029;
  assign ys__n1037 = ~ys__n874 | ys__n1036;
  assign new_n13573_ = ~ys__n1029 & ~ys__n1038;
  assign ys__n1040 = ys__n1037 | ~new_n13573_;
  assign ys__n3021 = ys__n874 & ys__n1048;
  assign ys__n1043 = ys__n140 | ~ys__n3021;
  assign new_n13577_ = new_n13376_ & new_n13503_;
  assign ys__n1046 = new_n13530_ & new_n13577_;
  assign ys__n1047 = ys__n140 | ~ys__n874;
  assign ys__n1049 = ys__n1048 | ys__n1047;
  assign new_n13581_ = ys__n1020 & new_n13301_;
  assign new_n13582_ = ~ys__n30223 & new_n13297_;
  assign ys__n16427 = new_n13581_ | new_n13582_;
  assign new_n13584_ = ys__n740 & new_n13295_;
  assign new_n13585_ = ~ys__n1020 & new_n13301_;
  assign new_n13586_ = ~new_n13563_ & new_n13585_;
  assign new_n13587_ = ~new_n13584_ & ~new_n13586_;
  assign ys__n1060 = ~ys__n16427 & new_n13587_;
  assign new_n13589_ = ys__n1020 & new_n13334_;
  assign new_n13590_ = ~ys__n30223 & new_n13330_;
  assign ys__n16721 = new_n13589_ | new_n13590_;
  assign new_n13592_ = ys__n740 & new_n13328_;
  assign new_n13593_ = ~ys__n1020 & new_n13334_;
  assign new_n13594_ = ~new_n13563_ & new_n13593_;
  assign new_n13595_ = ~new_n13592_ & ~new_n13594_;
  assign ys__n1071 = ~ys__n16721 & new_n13595_;
  assign ys__n1074 = ys__n1072 | ys__n1073;
  assign ys__n1075 = ~ys__n874 | ys__n1072;
  assign ys__n1077 = ~ys__n874 | ys__n1076;
  assign ys__n1079 = ys__n1072 | ys__n1078;
  assign ys__n1080 = ys__n1077 | ys__n1079;
  assign ys__n1448 = ys__n874 & ys__n1084;
  assign ys__n1083 = ys__n140 | ~ys__n1448;
  assign ys__n1085 = ys__n1084 | ys__n1047;
  assign ys__n1088 = ys__n1106 & ~ys__n33479;
  assign new_n13606_ = ~ys__n33481 & ys__n33495;
  assign new_n13607_ = ys__n1088 & new_n13606_;
  assign ys__n1087 = ys__n874 & new_n13607_;
  assign new_n13609_ = ~ys__n1098 & ~ys__n1107;
  assign new_n13610_ = ~ys__n1129 & new_n13609_;
  assign new_n13611_ = ~ys__n24463 & new_n13610_;
  assign ys__n1089 = ys__n24519 & ~new_n13611_;
  assign ys__n1090 = ys__n1088 | ys__n1089;
  assign ys__n1091 = ~ys__n874 | ys__n1088;
  assign ys__n1141 = ~ys__n874 | ys__n1094;
  assign ys__n1095 = ~ys__n1106 | ys__n1141;
  assign new_n13617_ = ~ys__n1094 & ~ys__n1106;
  assign new_n13618_ = ys__n874 & ~ys__n1098;
  assign new_n13619_ = ~ys__n1099 & ys__n1107;
  assign new_n13620_ = new_n13618_ & new_n13619_;
  assign ys__n1103 = ~new_n13617_ | ~new_n13620_;
  assign new_n13622_ = ~ys__n1109 & ~ys__n1110;
  assign new_n13623_ = ys__n1129 & new_n13622_;
  assign new_n13624_ = ~ys__n1099 & ~ys__n1107;
  assign new_n13625_ = new_n13618_ & new_n13624_;
  assign new_n13626_ = new_n13617_ & new_n13625_;
  assign ys__n1115 = ~new_n13623_ | ~new_n13626_;
  assign new_n13628_ = ~ys__n1098 & ~ys__n1106;
  assign new_n13629_ = ~ys__n1141 & new_n13628_;
  assign new_n13630_ = ~ys__n1107 & ~ys__n1109;
  assign new_n13631_ = ~ys__n1110 & ~ys__n1129;
  assign new_n13632_ = new_n13630_ & new_n13631_;
  assign new_n13633_ = new_n13629_ & new_n13632_;
  assign new_n13634_ = ~ys__n1119 & ~ys__n1120;
  assign new_n13635_ = ~ys__n1099 & ~ys__n1116;
  assign new_n13636_ = ~ys__n1117 & new_n13635_;
  assign new_n13637_ = new_n13634_ & new_n13636_;
  assign ys__n1125 = ~new_n13633_ | ~new_n13637_;
  assign new_n13639_ = ~ys__n1119 & new_n13635_;
  assign ys__n1128 = ~new_n13633_ | ~new_n13639_;
  assign new_n13641_ = ~ys__n1099 & ~ys__n1119;
  assign ys__n1135 = ~new_n13633_ | ~new_n13641_;
  assign new_n13643_ = ~ys__n1099 & ~ys__n1110;
  assign new_n13644_ = new_n13630_ & new_n13643_;
  assign ys__n1138 = ~new_n13629_ | ~new_n13644_;
  assign ys__n1142 = ~new_n13624_ | ~new_n13629_;
  assign ys__n1143 = ys__n1106 | ys__n1141;
  assign ys__n3118 = ys__n874 & ys__n1147;
  assign ys__n1146 = ys__n140 | ~ys__n3118;
  assign ys__n1148 = ys__n1147 | ys__n1047;
  assign new_n13651_ = ~ys__n1154 & ~ys__n1156;
  assign new_n13652_ = ~ys__n1157 & ys__n24591;
  assign new_n13653_ = new_n13651_ & new_n13652_;
  assign ys__n18137 = ys__n1151 | ys__n1153;
  assign new_n13655_ = ~ys__n1047 & ~ys__n18137;
  assign ys__n1161 = ~new_n13653_ | ~new_n13655_;
  assign ys__n1163 = new_n13421_ & new_n13548_;
  assign ys__n1164 = new_n13421_ & new_n13551_;
  assign ys__n1165 = new_n13421_ & new_n13542_;
  assign new_n13660_ = new_n13375_ & new_n13507_;
  assign ys__n1167 = new_n13530_ & new_n13660_;
  assign new_n13662_ = ~ys__n738 & new_n11954_;
  assign ys__n1170 = new_n12477_ & new_n13662_;
  assign ys__n1171 = ~ys__n874 | new_n13242_;
  assign ys__n1183 = ~ys__n858 | new_n13240_;
  assign ys__n1189 = ~ys__n856 | new_n13240_;
  assign ys__n1195 = ~ys__n854 | new_n13240_;
  assign ys__n1201 = ~ys__n852 | new_n13240_;
  assign ys__n1207 = ~ys__n850 | new_n13240_;
  assign ys__n1213 = ~ys__n848 | new_n13240_;
  assign ys__n1219 = ~ys__n846 | new_n13240_;
  assign ys__n1222 = ~ys__n844 | new_n13240_;
  assign ys__n1228 = ~ys__n842 | new_n13240_;
  assign ys__n1234 = ~ys__n840 | new_n13240_;
  assign ys__n1240 = ~ys__n838 | new_n13240_;
  assign ys__n1246 = ~ys__n836 | new_n13240_;
  assign ys__n1252 = ~ys__n834 | new_n13240_;
  assign ys__n1258 = ~ys__n832 | new_n13240_;
  assign ys__n1261 = ~ys__n830 | new_n13240_;
  assign ys__n1266 = ~ys__n828 | ~new_n12860_;
  assign ys__n1272 = ~ys__n826 | ~new_n12860_;
  assign ys__n1278 = ~ys__n824 | ~new_n12860_;
  assign ys__n1284 = ~ys__n822 | ~new_n12860_;
  assign ys__n1290 = ~ys__n820 | ~new_n12860_;
  assign ys__n1296 = ~ys__n818 | ~new_n12860_;
  assign ys__n1303 = ~ys__n816 | ~new_n12860_;
  assign new_n13687_ = new_n13384_ & new_n13507_;
  assign ys__n1377 = new_n13530_ & new_n13687_;
  assign new_n13689_ = ~ys__n536 & ~ys__n538;
  assign new_n13690_ = ys__n33403 & ~new_n13689_;
  assign new_n13691_ = ~ys__n935 & ys__n30863;
  assign new_n13692_ = ~ys__n33384 & new_n13691_;
  assign new_n13693_ = ~new_n13690_ & new_n13692_;
  assign new_n13694_ = ~ys__n738 & new_n13693_;
  assign ys__n1386 = ys__n4566 & new_n13694_;
  assign new_n13696_ = new_n13383_ & new_n13384_;
  assign ys__n1445 = new_n13530_ & new_n13696_;
  assign new_n13698_ = ~ys__n252 & ~ys__n254;
  assign new_n13699_ = ~ys__n250 & new_n13698_;
  assign new_n13700_ = ~ys__n246 & ~ys__n270;
  assign new_n13701_ = ys__n20273 & ys__n814;
  assign new_n13702_ = ~ys__n278 & new_n13701_;
  assign new_n13703_ = new_n13700_ & new_n13702_;
  assign ys__n1470 = ~new_n13699_ | ~new_n13703_;
  assign ys__n1591 = new_n13421_ & new_n13538_;
  assign ys__n1598 = ys__n44892 & ~ys__n4566;
  assign new_n13707_ = ~ys__n44840 & ~ys__n44842;
  assign new_n13708_ = ~ys__n4566 & ~new_n13707_;
  assign new_n13709_ = ys__n874 & ~ys__n1598;
  assign ys__n1601 = new_n13708_ | ~new_n13709_;
  assign ys__n1616 = new_n13421_ & new_n13523_;
  assign ys__n38453 = ~ys__n564 | ~new_n13689_;
  assign new_n13713_ = ~new_n12124_ & ~ys__n38453;
  assign new_n13714_ = ~new_n12139_ & ~new_n13713_;
  assign new_n13715_ = new_n12140_ & new_n13714_;
  assign new_n13716_ = ~new_n13693_ & new_n13713_;
  assign new_n13717_ = ~ys__n738 & ys__n4566;
  assign new_n13718_ = ~new_n13716_ & new_n13717_;
  assign new_n13719_ = ys__n738 & ~new_n13713_;
  assign new_n13720_ = ~new_n13718_ & ~new_n13719_;
  assign ys__n1790 = ~new_n13715_ & new_n13720_;
  assign new_n13722_ = ys__n33384 & ys__n38451;
  assign new_n13723_ = ~ys__n4177 & ~ys__n33394;
  assign ys__n26555 = ys__n34959 & new_n13723_;
  assign ys__n1802 = new_n13722_ | ys__n26555;
  assign new_n13726_ = ~ys__n348 & ~ys__n2924;
  assign new_n13727_ = ~ys__n162 & ys__n346;
  assign new_n13728_ = new_n13726_ & new_n13727_;
  assign new_n13729_ = ~ys__n342 & ~ys__n350;
  assign new_n13730_ = ys__n160 & ~ys__n344;
  assign new_n13731_ = new_n13729_ & new_n13730_;
  assign new_n13732_ = ys__n352 & new_n13731_;
  assign new_n13733_ = new_n13728_ & new_n13732_;
  assign new_n13734_ = ys__n342 & ~ys__n350;
  assign new_n13735_ = ys__n352 & new_n13730_;
  assign new_n13736_ = new_n13734_ & new_n13735_;
  assign new_n13737_ = new_n13728_ & new_n13736_;
  assign new_n13738_ = ~new_n13733_ & ~new_n13737_;
  assign new_n13739_ = ~ys__n160 & ~ys__n344;
  assign new_n13740_ = new_n13471_ & new_n13739_;
  assign new_n13741_ = ys__n352 & new_n13483_;
  assign new_n13742_ = new_n13740_ & new_n13741_;
  assign ys__n1817 = ~new_n13738_ | new_n13742_;
  assign new_n13744_ = new_n13376_ & new_n13383_;
  assign ys__n1835 = new_n13530_ & new_n13744_;
  assign new_n13746_ = ys__n480 & ~ys__n754;
  assign new_n13747_ = ~ys__n482 & ~ys__n756;
  assign new_n13748_ = new_n13746_ & new_n13747_;
  assign new_n13749_ = ys__n23652 & new_n13748_;
  assign new_n13750_ = new_n12107_ & new_n13748_;
  assign new_n13751_ = ys__n478 & new_n13750_;
  assign new_n13752_ = ~new_n13749_ & new_n13751_;
  assign new_n13753_ = ys__n478 & ~ys__n756;
  assign new_n13754_ = new_n12108_ & new_n13753_;
  assign new_n13755_ = ys__n482 & new_n13754_;
  assign new_n13756_ = new_n13746_ & new_n13755_;
  assign new_n13757_ = ~new_n13750_ & new_n13756_;
  assign new_n13758_ = ~new_n13749_ & new_n13757_;
  assign new_n13759_ = ~new_n13752_ & ~new_n13758_;
  assign new_n13760_ = ys__n478 & new_n13749_;
  assign new_n13761_ = new_n13759_ & ~new_n13760_;
  assign ys__n1837 = ~ys__n738 & ~new_n13761_;
  assign new_n13763_ = ys__n564 & ~new_n13689_;
  assign ys__n2152 = ys__n1386 | new_n13763_;
  assign new_n13765_ = new_n13384_ & new_n13492_;
  assign ys__n2365 = new_n13530_ & new_n13765_;
  assign new_n13767_ = new_n13384_ & new_n13503_;
  assign ys__n2400 = new_n13530_ & new_n13767_;
  assign new_n13769_ = ys__n38304 & ~ys__n4566;
  assign ys__n2423 = ~ys__n738 & new_n13769_;
  assign new_n13771_ = ys__n45046 & ys__n45580;
  assign new_n13772_ = ~ys__n45046 & ~ys__n45580;
  assign new_n13773_ = ~ys__n45622 & ~new_n13772_;
  assign new_n13774_ = ~new_n13771_ & new_n13773_;
  assign new_n13775_ = ys__n45049 & ys__n45582;
  assign new_n13776_ = ~ys__n45049 & ~ys__n45582;
  assign new_n13777_ = ~ys__n45623 & ~new_n13776_;
  assign new_n13778_ = ~new_n13775_ & new_n13777_;
  assign new_n13779_ = ~new_n13774_ & ~new_n13778_;
  assign new_n13780_ = ys__n45052 & ys__n45584;
  assign new_n13781_ = ~ys__n45052 & ~ys__n45584;
  assign new_n13782_ = ~ys__n45624 & ~new_n13781_;
  assign new_n13783_ = ~new_n13780_ & new_n13782_;
  assign new_n13784_ = ys__n45055 & ys__n45586;
  assign new_n13785_ = ~ys__n45055 & ~ys__n45586;
  assign new_n13786_ = ~ys__n45625 & ~new_n13785_;
  assign new_n13787_ = ~new_n13784_ & new_n13786_;
  assign new_n13788_ = ~new_n13783_ & ~new_n13787_;
  assign new_n13789_ = new_n13779_ & new_n13788_;
  assign new_n13790_ = ys__n45034 & ys__n45572;
  assign new_n13791_ = ~ys__n45034 & ~ys__n45572;
  assign new_n13792_ = ~ys__n45618 & ~new_n13791_;
  assign new_n13793_ = ~new_n13790_ & new_n13792_;
  assign new_n13794_ = ys__n45037 & ys__n45574;
  assign new_n13795_ = ~ys__n45037 & ~ys__n45574;
  assign new_n13796_ = ~ys__n45619 & ~new_n13795_;
  assign new_n13797_ = ~new_n13794_ & new_n13796_;
  assign new_n13798_ = ~new_n13793_ & ~new_n13797_;
  assign new_n13799_ = ys__n45040 & ys__n45576;
  assign new_n13800_ = ~ys__n45040 & ~ys__n45576;
  assign new_n13801_ = ~ys__n45620 & ~new_n13800_;
  assign new_n13802_ = ~new_n13799_ & new_n13801_;
  assign new_n13803_ = ys__n45043 & ys__n45578;
  assign new_n13804_ = ~ys__n45043 & ~ys__n45578;
  assign new_n13805_ = ~ys__n45621 & ~new_n13804_;
  assign new_n13806_ = ~new_n13803_ & new_n13805_;
  assign new_n13807_ = ~new_n13802_ & ~new_n13806_;
  assign new_n13808_ = new_n13798_ & new_n13807_;
  assign new_n13809_ = new_n13789_ & new_n13808_;
  assign new_n13810_ = ys__n45070 & ys__n45596;
  assign new_n13811_ = ~ys__n45070 & ~ys__n45596;
  assign new_n13812_ = ~ys__n45630 & ~new_n13811_;
  assign new_n13813_ = ~new_n13810_ & new_n13812_;
  assign new_n13814_ = ys__n45073 & ys__n45598;
  assign new_n13815_ = ~ys__n45073 & ~ys__n45598;
  assign new_n13816_ = ~ys__n45631 & ~new_n13815_;
  assign new_n13817_ = ~new_n13814_ & new_n13816_;
  assign new_n13818_ = ~new_n13813_ & ~new_n13817_;
  assign new_n13819_ = ys__n45076 & ys__n45600;
  assign new_n13820_ = ~ys__n45076 & ~ys__n45600;
  assign new_n13821_ = ~ys__n45632 & ~new_n13820_;
  assign new_n13822_ = ~new_n13819_ & new_n13821_;
  assign new_n13823_ = ys__n45079 & ys__n45602;
  assign new_n13824_ = ~ys__n45079 & ~ys__n45602;
  assign new_n13825_ = ~ys__n45633 & ~new_n13824_;
  assign new_n13826_ = ~new_n13823_ & new_n13825_;
  assign new_n13827_ = ~new_n13822_ & ~new_n13826_;
  assign new_n13828_ = new_n13818_ & new_n13827_;
  assign new_n13829_ = ys__n45058 & ys__n45588;
  assign new_n13830_ = ~ys__n45058 & ~ys__n45588;
  assign new_n13831_ = ~ys__n45626 & ~new_n13830_;
  assign new_n13832_ = ~new_n13829_ & new_n13831_;
  assign new_n13833_ = ys__n45061 & ys__n45590;
  assign new_n13834_ = ~ys__n45061 & ~ys__n45590;
  assign new_n13835_ = ~ys__n45627 & ~new_n13834_;
  assign new_n13836_ = ~new_n13833_ & new_n13835_;
  assign new_n13837_ = ~new_n13832_ & ~new_n13836_;
  assign new_n13838_ = ys__n45064 & ys__n45592;
  assign new_n13839_ = ~ys__n45064 & ~ys__n45592;
  assign new_n13840_ = ~ys__n45628 & ~new_n13839_;
  assign new_n13841_ = ~new_n13838_ & new_n13840_;
  assign new_n13842_ = ys__n45067 & ys__n45594;
  assign new_n13843_ = ~ys__n45067 & ~ys__n45594;
  assign new_n13844_ = ~ys__n45629 & ~new_n13843_;
  assign new_n13845_ = ~new_n13842_ & new_n13844_;
  assign new_n13846_ = ~new_n13841_ & ~new_n13845_;
  assign new_n13847_ = new_n13837_ & new_n13846_;
  assign new_n13848_ = new_n13828_ & new_n13847_;
  assign new_n13849_ = new_n13809_ & new_n13848_;
  assign new_n13850_ = ys__n44992 & ys__n45544;
  assign new_n13851_ = ~ys__n44992 & ~ys__n45544;
  assign new_n13852_ = ~ys__n45604 & ~new_n13851_;
  assign new_n13853_ = ~new_n13850_ & new_n13852_;
  assign new_n13854_ = ys__n44995 & ys__n45546;
  assign new_n13855_ = ~ys__n44995 & ~ys__n45546;
  assign new_n13856_ = ~ys__n45605 & ~new_n13855_;
  assign new_n13857_ = ~new_n13854_ & new_n13856_;
  assign new_n13858_ = ~new_n13853_ & ~new_n13857_;
  assign new_n13859_ = ys__n44998 & ys__n45548;
  assign new_n13860_ = ~ys__n44998 & ~ys__n45548;
  assign new_n13861_ = ~ys__n45606 & ~new_n13860_;
  assign new_n13862_ = ~new_n13859_ & new_n13861_;
  assign new_n13863_ = ys__n45001 & ys__n45550;
  assign new_n13864_ = ~ys__n45001 & ~ys__n45550;
  assign new_n13865_ = ~ys__n45607 & ~new_n13864_;
  assign new_n13866_ = ~new_n13863_ & new_n13865_;
  assign new_n13867_ = ~new_n13862_ & ~new_n13866_;
  assign new_n13868_ = ys__n45004 & ys__n45552;
  assign new_n13869_ = ~ys__n45004 & ~ys__n45552;
  assign new_n13870_ = ~ys__n45608 & ~new_n13869_;
  assign new_n13871_ = ~new_n13868_ & new_n13870_;
  assign new_n13872_ = ys__n45007 & ys__n45554;
  assign new_n13873_ = ~ys__n45007 & ~ys__n45554;
  assign new_n13874_ = ~ys__n45609 & ~new_n13873_;
  assign new_n13875_ = ~new_n13872_ & new_n13874_;
  assign new_n13876_ = ~new_n13871_ & ~new_n13875_;
  assign new_n13877_ = new_n13867_ & new_n13876_;
  assign new_n13878_ = new_n13858_ & new_n13877_;
  assign new_n13879_ = ys__n45022 & ys__n45564;
  assign new_n13880_ = ~ys__n45022 & ~ys__n45564;
  assign new_n13881_ = ~ys__n45614 & ~new_n13880_;
  assign new_n13882_ = ~new_n13879_ & new_n13881_;
  assign new_n13883_ = ys__n45025 & ys__n45566;
  assign new_n13884_ = ~ys__n45025 & ~ys__n45566;
  assign new_n13885_ = ~ys__n45615 & ~new_n13884_;
  assign new_n13886_ = ~new_n13883_ & new_n13885_;
  assign new_n13887_ = ~new_n13882_ & ~new_n13886_;
  assign new_n13888_ = ys__n45028 & ys__n45568;
  assign new_n13889_ = ~ys__n45028 & ~ys__n45568;
  assign new_n13890_ = ~ys__n45616 & ~new_n13889_;
  assign new_n13891_ = ~new_n13888_ & new_n13890_;
  assign new_n13892_ = ys__n45031 & ys__n45570;
  assign new_n13893_ = ~ys__n45031 & ~ys__n45570;
  assign new_n13894_ = ~ys__n45617 & ~new_n13893_;
  assign new_n13895_ = ~new_n13892_ & new_n13894_;
  assign new_n13896_ = ~new_n13891_ & ~new_n13895_;
  assign new_n13897_ = new_n13887_ & new_n13896_;
  assign new_n13898_ = ys__n45010 & ys__n45556;
  assign new_n13899_ = ~ys__n45010 & ~ys__n45556;
  assign new_n13900_ = ~ys__n45610 & ~new_n13899_;
  assign new_n13901_ = ~new_n13898_ & new_n13900_;
  assign new_n13902_ = ys__n45013 & ys__n45558;
  assign new_n13903_ = ~ys__n45013 & ~ys__n45558;
  assign new_n13904_ = ~ys__n45611 & ~new_n13903_;
  assign new_n13905_ = ~new_n13902_ & new_n13904_;
  assign new_n13906_ = ~new_n13901_ & ~new_n13905_;
  assign new_n13907_ = ys__n45016 & ys__n45560;
  assign new_n13908_ = ~ys__n45016 & ~ys__n45560;
  assign new_n13909_ = ~ys__n45612 & ~new_n13908_;
  assign new_n13910_ = ~new_n13907_ & new_n13909_;
  assign new_n13911_ = ys__n45019 & ys__n45562;
  assign new_n13912_ = ~ys__n45019 & ~ys__n45562;
  assign new_n13913_ = ~ys__n45613 & ~new_n13912_;
  assign new_n13914_ = ~new_n13911_ & new_n13913_;
  assign new_n13915_ = ~new_n13910_ & ~new_n13914_;
  assign new_n13916_ = new_n13906_ & new_n13915_;
  assign new_n13917_ = new_n13897_ & new_n13916_;
  assign new_n13918_ = new_n13878_ & new_n13917_;
  assign new_n13919_ = new_n13849_ & new_n13918_;
  assign new_n13920_ = ys__n45172 & ys__n45674;
  assign new_n13921_ = ~ys__n45172 & ~ys__n45674;
  assign new_n13922_ = ~ys__n45700 & ~new_n13921_;
  assign new_n13923_ = ~new_n13920_ & new_n13922_;
  assign new_n13924_ = ys__n45175 & ys__n45676;
  assign new_n13925_ = ~ys__n45175 & ~ys__n45676;
  assign new_n13926_ = ~ys__n45700 & ~new_n13925_;
  assign new_n13927_ = ~new_n13924_ & new_n13926_;
  assign new_n13928_ = ~new_n13923_ & ~new_n13927_;
  assign new_n13929_ = ys__n45178 & ys__n45678;
  assign new_n13930_ = ~ys__n45178 & ~ys__n45678;
  assign new_n13931_ = ~ys__n45700 & ~new_n13930_;
  assign new_n13932_ = ~new_n13929_ & new_n13931_;
  assign new_n13933_ = ys__n45181 & ys__n45680;
  assign new_n13934_ = ~ys__n45181 & ~ys__n45680;
  assign new_n13935_ = ~ys__n45700 & ~new_n13934_;
  assign new_n13936_ = ~new_n13933_ & new_n13935_;
  assign new_n13937_ = ~new_n13932_ & ~new_n13936_;
  assign new_n13938_ = new_n13928_ & new_n13937_;
  assign new_n13939_ = ys__n45160 & ys__n45666;
  assign new_n13940_ = ~ys__n45160 & ~ys__n45666;
  assign new_n13941_ = ~ys__n45700 & ~new_n13940_;
  assign new_n13942_ = ~new_n13939_ & new_n13941_;
  assign new_n13943_ = ys__n45163 & ys__n45668;
  assign new_n13944_ = ~ys__n45163 & ~ys__n45668;
  assign new_n13945_ = ~ys__n45700 & ~new_n13944_;
  assign new_n13946_ = ~new_n13943_ & new_n13945_;
  assign new_n13947_ = ~new_n13942_ & ~new_n13946_;
  assign new_n13948_ = ys__n45166 & ys__n45670;
  assign new_n13949_ = ~ys__n45166 & ~ys__n45670;
  assign new_n13950_ = ~ys__n45700 & ~new_n13949_;
  assign new_n13951_ = ~new_n13948_ & new_n13950_;
  assign new_n13952_ = ys__n45169 & ys__n45672;
  assign new_n13953_ = ~ys__n45169 & ~ys__n45672;
  assign new_n13954_ = ~ys__n45700 & ~new_n13953_;
  assign new_n13955_ = ~new_n13952_ & new_n13954_;
  assign new_n13956_ = ~new_n13951_ & ~new_n13955_;
  assign new_n13957_ = new_n13947_ & new_n13956_;
  assign new_n13958_ = new_n13938_ & new_n13957_;
  assign new_n13959_ = ys__n45196 & ys__n45690;
  assign new_n13960_ = ~ys__n45196 & ~ys__n45690;
  assign new_n13961_ = ~ys__n45701 & ~new_n13960_;
  assign new_n13962_ = ~new_n13959_ & new_n13961_;
  assign new_n13963_ = ys__n45199 & ys__n45692;
  assign new_n13964_ = ~ys__n45199 & ~ys__n45692;
  assign new_n13965_ = ~ys__n45701 & ~new_n13964_;
  assign new_n13966_ = ~new_n13963_ & new_n13965_;
  assign new_n13967_ = ~new_n13962_ & ~new_n13966_;
  assign new_n13968_ = ys__n45202 & ys__n45694;
  assign new_n13969_ = ~ys__n45202 & ~ys__n45694;
  assign new_n13970_ = ~ys__n45701 & ~new_n13969_;
  assign new_n13971_ = ~new_n13968_ & new_n13970_;
  assign new_n13972_ = ys__n45205 & ys__n45696;
  assign new_n13973_ = ~ys__n45205 & ~ys__n45696;
  assign new_n13974_ = ~ys__n45701 & ~new_n13973_;
  assign new_n13975_ = ~new_n13972_ & new_n13974_;
  assign new_n13976_ = ~new_n13971_ & ~new_n13975_;
  assign new_n13977_ = new_n13967_ & new_n13976_;
  assign new_n13978_ = ys__n45184 & ys__n45682;
  assign new_n13979_ = ~ys__n45184 & ~ys__n45682;
  assign new_n13980_ = ~ys__n45701 & ~new_n13979_;
  assign new_n13981_ = ~new_n13978_ & new_n13980_;
  assign new_n13982_ = ys__n45187 & ys__n45684;
  assign new_n13983_ = ~ys__n45187 & ~ys__n45684;
  assign new_n13984_ = ~ys__n45701 & ~new_n13983_;
  assign new_n13985_ = ~new_n13982_ & new_n13984_;
  assign new_n13986_ = ~new_n13981_ & ~new_n13985_;
  assign new_n13987_ = ys__n45190 & ys__n45686;
  assign new_n13988_ = ~ys__n45190 & ~ys__n45686;
  assign new_n13989_ = ~ys__n45701 & ~new_n13988_;
  assign new_n13990_ = ~new_n13987_ & new_n13989_;
  assign new_n13991_ = ys__n45193 & ys__n45688;
  assign new_n13992_ = ~ys__n45193 & ~ys__n45688;
  assign new_n13993_ = ~ys__n45701 & ~new_n13992_;
  assign new_n13994_ = ~new_n13991_ & new_n13993_;
  assign new_n13995_ = ~new_n13990_ & ~new_n13994_;
  assign new_n13996_ = new_n13986_ & new_n13995_;
  assign new_n13997_ = new_n13977_ & new_n13996_;
  assign new_n13998_ = new_n13958_ & new_n13997_;
  assign new_n13999_ = ys__n45124 & ys__n45642;
  assign new_n14000_ = ~ys__n45124 & ~ys__n45642;
  assign new_n14001_ = ~ys__n45698 & ~new_n14000_;
  assign new_n14002_ = ~new_n13999_ & new_n14001_;
  assign new_n14003_ = ys__n45127 & ys__n45644;
  assign new_n14004_ = ~ys__n45127 & ~ys__n45644;
  assign new_n14005_ = ~ys__n45698 & ~new_n14004_;
  assign new_n14006_ = ~new_n14003_ & new_n14005_;
  assign new_n14007_ = ~new_n14002_ & ~new_n14006_;
  assign new_n14008_ = ys__n45130 & ys__n45646;
  assign new_n14009_ = ~ys__n45130 & ~ys__n45646;
  assign new_n14010_ = ~ys__n45698 & ~new_n14009_;
  assign new_n14011_ = ~new_n14008_ & new_n14010_;
  assign new_n14012_ = ys__n45133 & ys__n45648;
  assign new_n14013_ = ~ys__n45133 & ~ys__n45648;
  assign new_n14014_ = ~ys__n45698 & ~new_n14013_;
  assign new_n14015_ = ~new_n14012_ & new_n14014_;
  assign new_n14016_ = ~new_n14011_ & ~new_n14015_;
  assign new_n14017_ = new_n14007_ & new_n14016_;
  assign new_n14018_ = ys__n45112 & ys__n45634;
  assign new_n14019_ = ~ys__n45112 & ~ys__n45634;
  assign new_n14020_ = ~ys__n45698 & ~new_n14019_;
  assign new_n14021_ = ~new_n14018_ & new_n14020_;
  assign new_n14022_ = ys__n45115 & ys__n45636;
  assign new_n14023_ = ~ys__n45115 & ~ys__n45636;
  assign new_n14024_ = ~ys__n45698 & ~new_n14023_;
  assign new_n14025_ = ~new_n14022_ & new_n14024_;
  assign new_n14026_ = ~new_n14021_ & ~new_n14025_;
  assign new_n14027_ = ys__n45118 & ys__n45638;
  assign new_n14028_ = ~ys__n45118 & ~ys__n45638;
  assign new_n14029_ = ~ys__n45698 & ~new_n14028_;
  assign new_n14030_ = ~new_n14027_ & new_n14029_;
  assign new_n14031_ = ys__n45121 & ys__n45640;
  assign new_n14032_ = ~ys__n45121 & ~ys__n45640;
  assign new_n14033_ = ~ys__n45698 & ~new_n14032_;
  assign new_n14034_ = ~new_n14031_ & new_n14033_;
  assign new_n14035_ = ~new_n14030_ & ~new_n14034_;
  assign new_n14036_ = new_n14026_ & new_n14035_;
  assign new_n14037_ = new_n14017_ & new_n14036_;
  assign new_n14038_ = ys__n45148 & ys__n45658;
  assign new_n14039_ = ~ys__n45148 & ~ys__n45658;
  assign new_n14040_ = ~ys__n45699 & ~new_n14039_;
  assign new_n14041_ = ~new_n14038_ & new_n14040_;
  assign new_n14042_ = ys__n45151 & ys__n45660;
  assign new_n14043_ = ~ys__n45151 & ~ys__n45660;
  assign new_n14044_ = ~ys__n45699 & ~new_n14043_;
  assign new_n14045_ = ~new_n14042_ & new_n14044_;
  assign new_n14046_ = ~new_n14041_ & ~new_n14045_;
  assign new_n14047_ = ys__n45154 & ys__n45662;
  assign new_n14048_ = ~ys__n45154 & ~ys__n45662;
  assign new_n14049_ = ~ys__n45699 & ~new_n14048_;
  assign new_n14050_ = ~new_n14047_ & new_n14049_;
  assign new_n14051_ = ys__n45157 & ys__n45664;
  assign new_n14052_ = ~ys__n45157 & ~ys__n45664;
  assign new_n14053_ = ~ys__n45699 & ~new_n14052_;
  assign new_n14054_ = ~new_n14051_ & new_n14053_;
  assign new_n14055_ = ~new_n14050_ & ~new_n14054_;
  assign new_n14056_ = new_n14046_ & new_n14055_;
  assign new_n14057_ = ys__n45136 & ys__n45650;
  assign new_n14058_ = ~ys__n45136 & ~ys__n45650;
  assign new_n14059_ = ~ys__n45699 & ~new_n14058_;
  assign new_n14060_ = ~new_n14057_ & new_n14059_;
  assign new_n14061_ = ys__n45139 & ys__n45652;
  assign new_n14062_ = ~ys__n45139 & ~ys__n45652;
  assign new_n14063_ = ~ys__n45699 & ~new_n14062_;
  assign new_n14064_ = ~new_n14061_ & new_n14063_;
  assign new_n14065_ = ~new_n14060_ & ~new_n14064_;
  assign new_n14066_ = ys__n45142 & ys__n45654;
  assign new_n14067_ = ~ys__n45142 & ~ys__n45654;
  assign new_n14068_ = ~ys__n45699 & ~new_n14067_;
  assign new_n14069_ = ~new_n14066_ & new_n14068_;
  assign new_n14070_ = ys__n45145 & ys__n45656;
  assign new_n14071_ = ~ys__n45145 & ~ys__n45656;
  assign new_n14072_ = ~ys__n45699 & ~new_n14071_;
  assign new_n14073_ = ~new_n14070_ & new_n14072_;
  assign new_n14074_ = ~new_n14069_ & ~new_n14073_;
  assign new_n14075_ = new_n14065_ & new_n14074_;
  assign new_n14076_ = new_n14056_ & new_n14075_;
  assign new_n14077_ = new_n14037_ & new_n14076_;
  assign new_n14078_ = new_n13998_ & new_n14077_;
  assign new_n14079_ = new_n13919_ & new_n14078_;
  assign new_n14080_ = ys__n45702 & new_n14079_;
  assign new_n14081_ = ys__n45046 & ys__n45416;
  assign new_n14082_ = ~ys__n45046 & ~ys__n45416;
  assign new_n14083_ = ~ys__n45458 & ~new_n14082_;
  assign new_n14084_ = ~new_n14081_ & new_n14083_;
  assign new_n14085_ = ys__n45049 & ys__n45418;
  assign new_n14086_ = ~ys__n45049 & ~ys__n45418;
  assign new_n14087_ = ~ys__n45459 & ~new_n14086_;
  assign new_n14088_ = ~new_n14085_ & new_n14087_;
  assign new_n14089_ = ~new_n14084_ & ~new_n14088_;
  assign new_n14090_ = ys__n45052 & ys__n45420;
  assign new_n14091_ = ~ys__n45052 & ~ys__n45420;
  assign new_n14092_ = ~ys__n45460 & ~new_n14091_;
  assign new_n14093_ = ~new_n14090_ & new_n14092_;
  assign new_n14094_ = ys__n45055 & ys__n45422;
  assign new_n14095_ = ~ys__n45055 & ~ys__n45422;
  assign new_n14096_ = ~ys__n45461 & ~new_n14095_;
  assign new_n14097_ = ~new_n14094_ & new_n14096_;
  assign new_n14098_ = ~new_n14093_ & ~new_n14097_;
  assign new_n14099_ = new_n14089_ & new_n14098_;
  assign new_n14100_ = ys__n45034 & ys__n45408;
  assign new_n14101_ = ~ys__n45034 & ~ys__n45408;
  assign new_n14102_ = ~ys__n45454 & ~new_n14101_;
  assign new_n14103_ = ~new_n14100_ & new_n14102_;
  assign new_n14104_ = ys__n45037 & ys__n45410;
  assign new_n14105_ = ~ys__n45037 & ~ys__n45410;
  assign new_n14106_ = ~ys__n45455 & ~new_n14105_;
  assign new_n14107_ = ~new_n14104_ & new_n14106_;
  assign new_n14108_ = ~new_n14103_ & ~new_n14107_;
  assign new_n14109_ = ys__n45040 & ys__n45412;
  assign new_n14110_ = ~ys__n45040 & ~ys__n45412;
  assign new_n14111_ = ~ys__n45456 & ~new_n14110_;
  assign new_n14112_ = ~new_n14109_ & new_n14111_;
  assign new_n14113_ = ys__n45043 & ys__n45414;
  assign new_n14114_ = ~ys__n45043 & ~ys__n45414;
  assign new_n14115_ = ~ys__n45457 & ~new_n14114_;
  assign new_n14116_ = ~new_n14113_ & new_n14115_;
  assign new_n14117_ = ~new_n14112_ & ~new_n14116_;
  assign new_n14118_ = new_n14108_ & new_n14117_;
  assign new_n14119_ = new_n14099_ & new_n14118_;
  assign new_n14120_ = ys__n45070 & ys__n45432;
  assign new_n14121_ = ~ys__n45070 & ~ys__n45432;
  assign new_n14122_ = ~ys__n45466 & ~new_n14121_;
  assign new_n14123_ = ~new_n14120_ & new_n14122_;
  assign new_n14124_ = ys__n45073 & ys__n45434;
  assign new_n14125_ = ~ys__n45073 & ~ys__n45434;
  assign new_n14126_ = ~ys__n45467 & ~new_n14125_;
  assign new_n14127_ = ~new_n14124_ & new_n14126_;
  assign new_n14128_ = ~new_n14123_ & ~new_n14127_;
  assign new_n14129_ = ys__n45076 & ys__n45436;
  assign new_n14130_ = ~ys__n45076 & ~ys__n45436;
  assign new_n14131_ = ~ys__n45468 & ~new_n14130_;
  assign new_n14132_ = ~new_n14129_ & new_n14131_;
  assign new_n14133_ = ys__n45079 & ys__n45438;
  assign new_n14134_ = ~ys__n45079 & ~ys__n45438;
  assign new_n14135_ = ~ys__n45469 & ~new_n14134_;
  assign new_n14136_ = ~new_n14133_ & new_n14135_;
  assign new_n14137_ = ~new_n14132_ & ~new_n14136_;
  assign new_n14138_ = new_n14128_ & new_n14137_;
  assign new_n14139_ = ys__n45058 & ys__n45424;
  assign new_n14140_ = ~ys__n45058 & ~ys__n45424;
  assign new_n14141_ = ~ys__n45462 & ~new_n14140_;
  assign new_n14142_ = ~new_n14139_ & new_n14141_;
  assign new_n14143_ = ys__n45061 & ys__n45426;
  assign new_n14144_ = ~ys__n45061 & ~ys__n45426;
  assign new_n14145_ = ~ys__n45463 & ~new_n14144_;
  assign new_n14146_ = ~new_n14143_ & new_n14145_;
  assign new_n14147_ = ~new_n14142_ & ~new_n14146_;
  assign new_n14148_ = ys__n45064 & ys__n45428;
  assign new_n14149_ = ~ys__n45064 & ~ys__n45428;
  assign new_n14150_ = ~ys__n45464 & ~new_n14149_;
  assign new_n14151_ = ~new_n14148_ & new_n14150_;
  assign new_n14152_ = ys__n45067 & ys__n45430;
  assign new_n14153_ = ~ys__n45067 & ~ys__n45430;
  assign new_n14154_ = ~ys__n45465 & ~new_n14153_;
  assign new_n14155_ = ~new_n14152_ & new_n14154_;
  assign new_n14156_ = ~new_n14151_ & ~new_n14155_;
  assign new_n14157_ = new_n14147_ & new_n14156_;
  assign new_n14158_ = new_n14138_ & new_n14157_;
  assign new_n14159_ = new_n14119_ & new_n14158_;
  assign new_n14160_ = ys__n44992 & ys__n45380;
  assign new_n14161_ = ~ys__n44992 & ~ys__n45380;
  assign new_n14162_ = ~ys__n45440 & ~new_n14161_;
  assign new_n14163_ = ~new_n14160_ & new_n14162_;
  assign new_n14164_ = ys__n44995 & ys__n45382;
  assign new_n14165_ = ~ys__n44995 & ~ys__n45382;
  assign new_n14166_ = ~ys__n45441 & ~new_n14165_;
  assign new_n14167_ = ~new_n14164_ & new_n14166_;
  assign new_n14168_ = ~new_n14163_ & ~new_n14167_;
  assign new_n14169_ = ys__n44998 & ys__n45384;
  assign new_n14170_ = ~ys__n44998 & ~ys__n45384;
  assign new_n14171_ = ~ys__n45442 & ~new_n14170_;
  assign new_n14172_ = ~new_n14169_ & new_n14171_;
  assign new_n14173_ = ys__n45001 & ys__n45386;
  assign new_n14174_ = ~ys__n45001 & ~ys__n45386;
  assign new_n14175_ = ~ys__n45443 & ~new_n14174_;
  assign new_n14176_ = ~new_n14173_ & new_n14175_;
  assign new_n14177_ = ~new_n14172_ & ~new_n14176_;
  assign new_n14178_ = ys__n45004 & ys__n45388;
  assign new_n14179_ = ~ys__n45004 & ~ys__n45388;
  assign new_n14180_ = ~ys__n45444 & ~new_n14179_;
  assign new_n14181_ = ~new_n14178_ & new_n14180_;
  assign new_n14182_ = ys__n45007 & ys__n45390;
  assign new_n14183_ = ~ys__n45007 & ~ys__n45390;
  assign new_n14184_ = ~ys__n45445 & ~new_n14183_;
  assign new_n14185_ = ~new_n14182_ & new_n14184_;
  assign new_n14186_ = ~new_n14181_ & ~new_n14185_;
  assign new_n14187_ = new_n14177_ & new_n14186_;
  assign new_n14188_ = new_n14168_ & new_n14187_;
  assign new_n14189_ = ys__n45022 & ys__n45400;
  assign new_n14190_ = ~ys__n45022 & ~ys__n45400;
  assign new_n14191_ = ~ys__n45450 & ~new_n14190_;
  assign new_n14192_ = ~new_n14189_ & new_n14191_;
  assign new_n14193_ = ys__n45025 & ys__n45402;
  assign new_n14194_ = ~ys__n45025 & ~ys__n45402;
  assign new_n14195_ = ~ys__n45451 & ~new_n14194_;
  assign new_n14196_ = ~new_n14193_ & new_n14195_;
  assign new_n14197_ = ~new_n14192_ & ~new_n14196_;
  assign new_n14198_ = ys__n45028 & ys__n45404;
  assign new_n14199_ = ~ys__n45028 & ~ys__n45404;
  assign new_n14200_ = ~ys__n45452 & ~new_n14199_;
  assign new_n14201_ = ~new_n14198_ & new_n14200_;
  assign new_n14202_ = ys__n45031 & ys__n45406;
  assign new_n14203_ = ~ys__n45031 & ~ys__n45406;
  assign new_n14204_ = ~ys__n45453 & ~new_n14203_;
  assign new_n14205_ = ~new_n14202_ & new_n14204_;
  assign new_n14206_ = ~new_n14201_ & ~new_n14205_;
  assign new_n14207_ = new_n14197_ & new_n14206_;
  assign new_n14208_ = ys__n45010 & ys__n45392;
  assign new_n14209_ = ~ys__n45010 & ~ys__n45392;
  assign new_n14210_ = ~ys__n45446 & ~new_n14209_;
  assign new_n14211_ = ~new_n14208_ & new_n14210_;
  assign new_n14212_ = ys__n45013 & ys__n45394;
  assign new_n14213_ = ~ys__n45013 & ~ys__n45394;
  assign new_n14214_ = ~ys__n45447 & ~new_n14213_;
  assign new_n14215_ = ~new_n14212_ & new_n14214_;
  assign new_n14216_ = ~new_n14211_ & ~new_n14215_;
  assign new_n14217_ = ys__n45016 & ys__n45396;
  assign new_n14218_ = ~ys__n45016 & ~ys__n45396;
  assign new_n14219_ = ~ys__n45448 & ~new_n14218_;
  assign new_n14220_ = ~new_n14217_ & new_n14219_;
  assign new_n14221_ = ys__n45019 & ys__n45398;
  assign new_n14222_ = ~ys__n45019 & ~ys__n45398;
  assign new_n14223_ = ~ys__n45449 & ~new_n14222_;
  assign new_n14224_ = ~new_n14221_ & new_n14223_;
  assign new_n14225_ = ~new_n14220_ & ~new_n14224_;
  assign new_n14226_ = new_n14216_ & new_n14225_;
  assign new_n14227_ = new_n14207_ & new_n14226_;
  assign new_n14228_ = new_n14188_ & new_n14227_;
  assign new_n14229_ = new_n14159_ & new_n14228_;
  assign new_n14230_ = ys__n45172 & ys__n45510;
  assign new_n14231_ = ~ys__n45172 & ~ys__n45510;
  assign new_n14232_ = ~ys__n45536 & ~new_n14231_;
  assign new_n14233_ = ~new_n14230_ & new_n14232_;
  assign new_n14234_ = ys__n45175 & ys__n45512;
  assign new_n14235_ = ~ys__n45175 & ~ys__n45512;
  assign new_n14236_ = ~ys__n45536 & ~new_n14235_;
  assign new_n14237_ = ~new_n14234_ & new_n14236_;
  assign new_n14238_ = ~new_n14233_ & ~new_n14237_;
  assign new_n14239_ = ys__n45178 & ys__n45514;
  assign new_n14240_ = ~ys__n45178 & ~ys__n45514;
  assign new_n14241_ = ~ys__n45536 & ~new_n14240_;
  assign new_n14242_ = ~new_n14239_ & new_n14241_;
  assign new_n14243_ = ys__n45181 & ys__n45516;
  assign new_n14244_ = ~ys__n45181 & ~ys__n45516;
  assign new_n14245_ = ~ys__n45536 & ~new_n14244_;
  assign new_n14246_ = ~new_n14243_ & new_n14245_;
  assign new_n14247_ = ~new_n14242_ & ~new_n14246_;
  assign new_n14248_ = new_n14238_ & new_n14247_;
  assign new_n14249_ = ys__n45160 & ys__n45502;
  assign new_n14250_ = ~ys__n45160 & ~ys__n45502;
  assign new_n14251_ = ~ys__n45536 & ~new_n14250_;
  assign new_n14252_ = ~new_n14249_ & new_n14251_;
  assign new_n14253_ = ys__n45163 & ys__n45504;
  assign new_n14254_ = ~ys__n45163 & ~ys__n45504;
  assign new_n14255_ = ~ys__n45536 & ~new_n14254_;
  assign new_n14256_ = ~new_n14253_ & new_n14255_;
  assign new_n14257_ = ~new_n14252_ & ~new_n14256_;
  assign new_n14258_ = ys__n45166 & ys__n45506;
  assign new_n14259_ = ~ys__n45166 & ~ys__n45506;
  assign new_n14260_ = ~ys__n45536 & ~new_n14259_;
  assign new_n14261_ = ~new_n14258_ & new_n14260_;
  assign new_n14262_ = ys__n45169 & ys__n45508;
  assign new_n14263_ = ~ys__n45169 & ~ys__n45508;
  assign new_n14264_ = ~ys__n45536 & ~new_n14263_;
  assign new_n14265_ = ~new_n14262_ & new_n14264_;
  assign new_n14266_ = ~new_n14261_ & ~new_n14265_;
  assign new_n14267_ = new_n14257_ & new_n14266_;
  assign new_n14268_ = new_n14248_ & new_n14267_;
  assign new_n14269_ = ys__n45196 & ys__n45526;
  assign new_n14270_ = ~ys__n45196 & ~ys__n45526;
  assign new_n14271_ = ~ys__n45537 & ~new_n14270_;
  assign new_n14272_ = ~new_n14269_ & new_n14271_;
  assign new_n14273_ = ys__n45199 & ys__n45528;
  assign new_n14274_ = ~ys__n45199 & ~ys__n45528;
  assign new_n14275_ = ~ys__n45537 & ~new_n14274_;
  assign new_n14276_ = ~new_n14273_ & new_n14275_;
  assign new_n14277_ = ~new_n14272_ & ~new_n14276_;
  assign new_n14278_ = ys__n45202 & ys__n45530;
  assign new_n14279_ = ~ys__n45202 & ~ys__n45530;
  assign new_n14280_ = ~ys__n45537 & ~new_n14279_;
  assign new_n14281_ = ~new_n14278_ & new_n14280_;
  assign new_n14282_ = ys__n45205 & ys__n45532;
  assign new_n14283_ = ~ys__n45205 & ~ys__n45532;
  assign new_n14284_ = ~ys__n45537 & ~new_n14283_;
  assign new_n14285_ = ~new_n14282_ & new_n14284_;
  assign new_n14286_ = ~new_n14281_ & ~new_n14285_;
  assign new_n14287_ = new_n14277_ & new_n14286_;
  assign new_n14288_ = ys__n45184 & ys__n45518;
  assign new_n14289_ = ~ys__n45184 & ~ys__n45518;
  assign new_n14290_ = ~ys__n45537 & ~new_n14289_;
  assign new_n14291_ = ~new_n14288_ & new_n14290_;
  assign new_n14292_ = ys__n45187 & ys__n45520;
  assign new_n14293_ = ~ys__n45187 & ~ys__n45520;
  assign new_n14294_ = ~ys__n45537 & ~new_n14293_;
  assign new_n14295_ = ~new_n14292_ & new_n14294_;
  assign new_n14296_ = ~new_n14291_ & ~new_n14295_;
  assign new_n14297_ = ys__n45190 & ys__n45522;
  assign new_n14298_ = ~ys__n45190 & ~ys__n45522;
  assign new_n14299_ = ~ys__n45537 & ~new_n14298_;
  assign new_n14300_ = ~new_n14297_ & new_n14299_;
  assign new_n14301_ = ys__n45193 & ys__n45524;
  assign new_n14302_ = ~ys__n45193 & ~ys__n45524;
  assign new_n14303_ = ~ys__n45537 & ~new_n14302_;
  assign new_n14304_ = ~new_n14301_ & new_n14303_;
  assign new_n14305_ = ~new_n14300_ & ~new_n14304_;
  assign new_n14306_ = new_n14296_ & new_n14305_;
  assign new_n14307_ = new_n14287_ & new_n14306_;
  assign new_n14308_ = new_n14268_ & new_n14307_;
  assign new_n14309_ = ys__n45124 & ys__n45478;
  assign new_n14310_ = ~ys__n45124 & ~ys__n45478;
  assign new_n14311_ = ~ys__n45534 & ~new_n14310_;
  assign new_n14312_ = ~new_n14309_ & new_n14311_;
  assign new_n14313_ = ys__n45127 & ys__n45480;
  assign new_n14314_ = ~ys__n45127 & ~ys__n45480;
  assign new_n14315_ = ~ys__n45534 & ~new_n14314_;
  assign new_n14316_ = ~new_n14313_ & new_n14315_;
  assign new_n14317_ = ~new_n14312_ & ~new_n14316_;
  assign new_n14318_ = ys__n45130 & ys__n45482;
  assign new_n14319_ = ~ys__n45130 & ~ys__n45482;
  assign new_n14320_ = ~ys__n45534 & ~new_n14319_;
  assign new_n14321_ = ~new_n14318_ & new_n14320_;
  assign new_n14322_ = ys__n45133 & ys__n45484;
  assign new_n14323_ = ~ys__n45133 & ~ys__n45484;
  assign new_n14324_ = ~ys__n45534 & ~new_n14323_;
  assign new_n14325_ = ~new_n14322_ & new_n14324_;
  assign new_n14326_ = ~new_n14321_ & ~new_n14325_;
  assign new_n14327_ = new_n14317_ & new_n14326_;
  assign new_n14328_ = ys__n45112 & ys__n45470;
  assign new_n14329_ = ~ys__n45112 & ~ys__n45470;
  assign new_n14330_ = ~ys__n45534 & ~new_n14329_;
  assign new_n14331_ = ~new_n14328_ & new_n14330_;
  assign new_n14332_ = ys__n45115 & ys__n45472;
  assign new_n14333_ = ~ys__n45115 & ~ys__n45472;
  assign new_n14334_ = ~ys__n45534 & ~new_n14333_;
  assign new_n14335_ = ~new_n14332_ & new_n14334_;
  assign new_n14336_ = ~new_n14331_ & ~new_n14335_;
  assign new_n14337_ = ys__n45118 & ys__n45474;
  assign new_n14338_ = ~ys__n45118 & ~ys__n45474;
  assign new_n14339_ = ~ys__n45534 & ~new_n14338_;
  assign new_n14340_ = ~new_n14337_ & new_n14339_;
  assign new_n14341_ = ys__n45121 & ys__n45476;
  assign new_n14342_ = ~ys__n45121 & ~ys__n45476;
  assign new_n14343_ = ~ys__n45534 & ~new_n14342_;
  assign new_n14344_ = ~new_n14341_ & new_n14343_;
  assign new_n14345_ = ~new_n14340_ & ~new_n14344_;
  assign new_n14346_ = new_n14336_ & new_n14345_;
  assign new_n14347_ = new_n14327_ & new_n14346_;
  assign new_n14348_ = ys__n45148 & ys__n45494;
  assign new_n14349_ = ~ys__n45148 & ~ys__n45494;
  assign new_n14350_ = ~ys__n45535 & ~new_n14349_;
  assign new_n14351_ = ~new_n14348_ & new_n14350_;
  assign new_n14352_ = ys__n45151 & ys__n45496;
  assign new_n14353_ = ~ys__n45151 & ~ys__n45496;
  assign new_n14354_ = ~ys__n45535 & ~new_n14353_;
  assign new_n14355_ = ~new_n14352_ & new_n14354_;
  assign new_n14356_ = ~new_n14351_ & ~new_n14355_;
  assign new_n14357_ = ys__n45154 & ys__n45498;
  assign new_n14358_ = ~ys__n45154 & ~ys__n45498;
  assign new_n14359_ = ~ys__n45535 & ~new_n14358_;
  assign new_n14360_ = ~new_n14357_ & new_n14359_;
  assign new_n14361_ = ys__n45157 & ys__n45500;
  assign new_n14362_ = ~ys__n45157 & ~ys__n45500;
  assign new_n14363_ = ~ys__n45535 & ~new_n14362_;
  assign new_n14364_ = ~new_n14361_ & new_n14363_;
  assign new_n14365_ = ~new_n14360_ & ~new_n14364_;
  assign new_n14366_ = new_n14356_ & new_n14365_;
  assign new_n14367_ = ys__n45136 & ys__n45486;
  assign new_n14368_ = ~ys__n45136 & ~ys__n45486;
  assign new_n14369_ = ~ys__n45535 & ~new_n14368_;
  assign new_n14370_ = ~new_n14367_ & new_n14369_;
  assign new_n14371_ = ys__n45139 & ys__n45488;
  assign new_n14372_ = ~ys__n45139 & ~ys__n45488;
  assign new_n14373_ = ~ys__n45535 & ~new_n14372_;
  assign new_n14374_ = ~new_n14371_ & new_n14373_;
  assign new_n14375_ = ~new_n14370_ & ~new_n14374_;
  assign new_n14376_ = ys__n45142 & ys__n45490;
  assign new_n14377_ = ~ys__n45142 & ~ys__n45490;
  assign new_n14378_ = ~ys__n45535 & ~new_n14377_;
  assign new_n14379_ = ~new_n14376_ & new_n14378_;
  assign new_n14380_ = ys__n45145 & ys__n45492;
  assign new_n14381_ = ~ys__n45145 & ~ys__n45492;
  assign new_n14382_ = ~ys__n45535 & ~new_n14381_;
  assign new_n14383_ = ~new_n14380_ & new_n14382_;
  assign new_n14384_ = ~new_n14379_ & ~new_n14383_;
  assign new_n14385_ = new_n14375_ & new_n14384_;
  assign new_n14386_ = new_n14366_ & new_n14385_;
  assign new_n14387_ = new_n14347_ & new_n14386_;
  assign new_n14388_ = new_n14308_ & new_n14387_;
  assign new_n14389_ = new_n14229_ & new_n14388_;
  assign new_n14390_ = ys__n45538 & new_n14389_;
  assign new_n14391_ = ~new_n14080_ & ~new_n14390_;
  assign new_n14392_ = ys__n45046 & ys__n45252;
  assign new_n14393_ = ~ys__n45046 & ~ys__n45252;
  assign new_n14394_ = ~ys__n45294 & ~new_n14393_;
  assign new_n14395_ = ~new_n14392_ & new_n14394_;
  assign new_n14396_ = ys__n45049 & ys__n45254;
  assign new_n14397_ = ~ys__n45049 & ~ys__n45254;
  assign new_n14398_ = ~ys__n45295 & ~new_n14397_;
  assign new_n14399_ = ~new_n14396_ & new_n14398_;
  assign new_n14400_ = ~new_n14395_ & ~new_n14399_;
  assign new_n14401_ = ys__n45052 & ys__n45256;
  assign new_n14402_ = ~ys__n45052 & ~ys__n45256;
  assign new_n14403_ = ~ys__n45296 & ~new_n14402_;
  assign new_n14404_ = ~new_n14401_ & new_n14403_;
  assign new_n14405_ = ys__n45055 & ys__n45258;
  assign new_n14406_ = ~ys__n45055 & ~ys__n45258;
  assign new_n14407_ = ~ys__n45297 & ~new_n14406_;
  assign new_n14408_ = ~new_n14405_ & new_n14407_;
  assign new_n14409_ = ~new_n14404_ & ~new_n14408_;
  assign new_n14410_ = new_n14400_ & new_n14409_;
  assign new_n14411_ = ys__n45034 & ys__n45244;
  assign new_n14412_ = ~ys__n45034 & ~ys__n45244;
  assign new_n14413_ = ~ys__n45290 & ~new_n14412_;
  assign new_n14414_ = ~new_n14411_ & new_n14413_;
  assign new_n14415_ = ys__n45037 & ys__n45246;
  assign new_n14416_ = ~ys__n45037 & ~ys__n45246;
  assign new_n14417_ = ~ys__n45291 & ~new_n14416_;
  assign new_n14418_ = ~new_n14415_ & new_n14417_;
  assign new_n14419_ = ~new_n14414_ & ~new_n14418_;
  assign new_n14420_ = ys__n45040 & ys__n45248;
  assign new_n14421_ = ~ys__n45040 & ~ys__n45248;
  assign new_n14422_ = ~ys__n45292 & ~new_n14421_;
  assign new_n14423_ = ~new_n14420_ & new_n14422_;
  assign new_n14424_ = ys__n45043 & ys__n45250;
  assign new_n14425_ = ~ys__n45043 & ~ys__n45250;
  assign new_n14426_ = ~ys__n45293 & ~new_n14425_;
  assign new_n14427_ = ~new_n14424_ & new_n14426_;
  assign new_n14428_ = ~new_n14423_ & ~new_n14427_;
  assign new_n14429_ = new_n14419_ & new_n14428_;
  assign new_n14430_ = new_n14410_ & new_n14429_;
  assign new_n14431_ = ys__n45070 & ys__n45268;
  assign new_n14432_ = ~ys__n45070 & ~ys__n45268;
  assign new_n14433_ = ~ys__n45302 & ~new_n14432_;
  assign new_n14434_ = ~new_n14431_ & new_n14433_;
  assign new_n14435_ = ys__n45073 & ys__n45270;
  assign new_n14436_ = ~ys__n45073 & ~ys__n45270;
  assign new_n14437_ = ~ys__n45303 & ~new_n14436_;
  assign new_n14438_ = ~new_n14435_ & new_n14437_;
  assign new_n14439_ = ~new_n14434_ & ~new_n14438_;
  assign new_n14440_ = ys__n45076 & ys__n45272;
  assign new_n14441_ = ~ys__n45076 & ~ys__n45272;
  assign new_n14442_ = ~ys__n45304 & ~new_n14441_;
  assign new_n14443_ = ~new_n14440_ & new_n14442_;
  assign new_n14444_ = ys__n45079 & ys__n45274;
  assign new_n14445_ = ~ys__n45079 & ~ys__n45274;
  assign new_n14446_ = ~ys__n45305 & ~new_n14445_;
  assign new_n14447_ = ~new_n14444_ & new_n14446_;
  assign new_n14448_ = ~new_n14443_ & ~new_n14447_;
  assign new_n14449_ = new_n14439_ & new_n14448_;
  assign new_n14450_ = ys__n45058 & ys__n45260;
  assign new_n14451_ = ~ys__n45058 & ~ys__n45260;
  assign new_n14452_ = ~ys__n45298 & ~new_n14451_;
  assign new_n14453_ = ~new_n14450_ & new_n14452_;
  assign new_n14454_ = ys__n45061 & ys__n45262;
  assign new_n14455_ = ~ys__n45061 & ~ys__n45262;
  assign new_n14456_ = ~ys__n45299 & ~new_n14455_;
  assign new_n14457_ = ~new_n14454_ & new_n14456_;
  assign new_n14458_ = ~new_n14453_ & ~new_n14457_;
  assign new_n14459_ = ys__n45064 & ys__n45264;
  assign new_n14460_ = ~ys__n45064 & ~ys__n45264;
  assign new_n14461_ = ~ys__n45300 & ~new_n14460_;
  assign new_n14462_ = ~new_n14459_ & new_n14461_;
  assign new_n14463_ = ys__n45067 & ys__n45266;
  assign new_n14464_ = ~ys__n45067 & ~ys__n45266;
  assign new_n14465_ = ~ys__n45301 & ~new_n14464_;
  assign new_n14466_ = ~new_n14463_ & new_n14465_;
  assign new_n14467_ = ~new_n14462_ & ~new_n14466_;
  assign new_n14468_ = new_n14458_ & new_n14467_;
  assign new_n14469_ = new_n14449_ & new_n14468_;
  assign new_n14470_ = new_n14430_ & new_n14469_;
  assign new_n14471_ = ys__n44992 & ys__n45216;
  assign new_n14472_ = ~ys__n44992 & ~ys__n45216;
  assign new_n14473_ = ~ys__n45276 & ~new_n14472_;
  assign new_n14474_ = ~new_n14471_ & new_n14473_;
  assign new_n14475_ = ys__n44995 & ys__n45218;
  assign new_n14476_ = ~ys__n44995 & ~ys__n45218;
  assign new_n14477_ = ~ys__n45277 & ~new_n14476_;
  assign new_n14478_ = ~new_n14475_ & new_n14477_;
  assign new_n14479_ = ~new_n14474_ & ~new_n14478_;
  assign new_n14480_ = ys__n44998 & ys__n45220;
  assign new_n14481_ = ~ys__n44998 & ~ys__n45220;
  assign new_n14482_ = ~ys__n45278 & ~new_n14481_;
  assign new_n14483_ = ~new_n14480_ & new_n14482_;
  assign new_n14484_ = ys__n45001 & ys__n45222;
  assign new_n14485_ = ~ys__n45001 & ~ys__n45222;
  assign new_n14486_ = ~ys__n45279 & ~new_n14485_;
  assign new_n14487_ = ~new_n14484_ & new_n14486_;
  assign new_n14488_ = ~new_n14483_ & ~new_n14487_;
  assign new_n14489_ = ys__n45004 & ys__n45224;
  assign new_n14490_ = ~ys__n45004 & ~ys__n45224;
  assign new_n14491_ = ~ys__n45280 & ~new_n14490_;
  assign new_n14492_ = ~new_n14489_ & new_n14491_;
  assign new_n14493_ = ys__n45007 & ys__n45226;
  assign new_n14494_ = ~ys__n45007 & ~ys__n45226;
  assign new_n14495_ = ~ys__n45281 & ~new_n14494_;
  assign new_n14496_ = ~new_n14493_ & new_n14495_;
  assign new_n14497_ = ~new_n14492_ & ~new_n14496_;
  assign new_n14498_ = new_n14488_ & new_n14497_;
  assign new_n14499_ = new_n14479_ & new_n14498_;
  assign new_n14500_ = ys__n45022 & ys__n45236;
  assign new_n14501_ = ~ys__n45022 & ~ys__n45236;
  assign new_n14502_ = ~ys__n45286 & ~new_n14501_;
  assign new_n14503_ = ~new_n14500_ & new_n14502_;
  assign new_n14504_ = ys__n45025 & ys__n45238;
  assign new_n14505_ = ~ys__n45025 & ~ys__n45238;
  assign new_n14506_ = ~ys__n45287 & ~new_n14505_;
  assign new_n14507_ = ~new_n14504_ & new_n14506_;
  assign new_n14508_ = ~new_n14503_ & ~new_n14507_;
  assign new_n14509_ = ys__n45028 & ys__n45240;
  assign new_n14510_ = ~ys__n45028 & ~ys__n45240;
  assign new_n14511_ = ~ys__n45288 & ~new_n14510_;
  assign new_n14512_ = ~new_n14509_ & new_n14511_;
  assign new_n14513_ = ys__n45031 & ys__n45242;
  assign new_n14514_ = ~ys__n45031 & ~ys__n45242;
  assign new_n14515_ = ~ys__n45289 & ~new_n14514_;
  assign new_n14516_ = ~new_n14513_ & new_n14515_;
  assign new_n14517_ = ~new_n14512_ & ~new_n14516_;
  assign new_n14518_ = new_n14508_ & new_n14517_;
  assign new_n14519_ = ys__n45010 & ys__n45228;
  assign new_n14520_ = ~ys__n45010 & ~ys__n45228;
  assign new_n14521_ = ~ys__n45282 & ~new_n14520_;
  assign new_n14522_ = ~new_n14519_ & new_n14521_;
  assign new_n14523_ = ys__n45013 & ys__n45230;
  assign new_n14524_ = ~ys__n45013 & ~ys__n45230;
  assign new_n14525_ = ~ys__n45283 & ~new_n14524_;
  assign new_n14526_ = ~new_n14523_ & new_n14525_;
  assign new_n14527_ = ~new_n14522_ & ~new_n14526_;
  assign new_n14528_ = ys__n45016 & ys__n45232;
  assign new_n14529_ = ~ys__n45016 & ~ys__n45232;
  assign new_n14530_ = ~ys__n45284 & ~new_n14529_;
  assign new_n14531_ = ~new_n14528_ & new_n14530_;
  assign new_n14532_ = ys__n45019 & ys__n45234;
  assign new_n14533_ = ~ys__n45019 & ~ys__n45234;
  assign new_n14534_ = ~ys__n45285 & ~new_n14533_;
  assign new_n14535_ = ~new_n14532_ & new_n14534_;
  assign new_n14536_ = ~new_n14531_ & ~new_n14535_;
  assign new_n14537_ = new_n14527_ & new_n14536_;
  assign new_n14538_ = new_n14518_ & new_n14537_;
  assign new_n14539_ = new_n14499_ & new_n14538_;
  assign new_n14540_ = new_n14470_ & new_n14539_;
  assign new_n14541_ = ys__n45172 & ys__n45346;
  assign new_n14542_ = ~ys__n45172 & ~ys__n45346;
  assign new_n14543_ = ~ys__n45372 & ~new_n14542_;
  assign new_n14544_ = ~new_n14541_ & new_n14543_;
  assign new_n14545_ = ys__n45175 & ys__n45348;
  assign new_n14546_ = ~ys__n45175 & ~ys__n45348;
  assign new_n14547_ = ~ys__n45372 & ~new_n14546_;
  assign new_n14548_ = ~new_n14545_ & new_n14547_;
  assign new_n14549_ = ~new_n14544_ & ~new_n14548_;
  assign new_n14550_ = ys__n45178 & ys__n45350;
  assign new_n14551_ = ~ys__n45178 & ~ys__n45350;
  assign new_n14552_ = ~ys__n45372 & ~new_n14551_;
  assign new_n14553_ = ~new_n14550_ & new_n14552_;
  assign new_n14554_ = ys__n45181 & ys__n45352;
  assign new_n14555_ = ~ys__n45181 & ~ys__n45352;
  assign new_n14556_ = ~ys__n45372 & ~new_n14555_;
  assign new_n14557_ = ~new_n14554_ & new_n14556_;
  assign new_n14558_ = ~new_n14553_ & ~new_n14557_;
  assign new_n14559_ = new_n14549_ & new_n14558_;
  assign new_n14560_ = ys__n45160 & ys__n45338;
  assign new_n14561_ = ~ys__n45160 & ~ys__n45338;
  assign new_n14562_ = ~ys__n45372 & ~new_n14561_;
  assign new_n14563_ = ~new_n14560_ & new_n14562_;
  assign new_n14564_ = ys__n45163 & ys__n45340;
  assign new_n14565_ = ~ys__n45163 & ~ys__n45340;
  assign new_n14566_ = ~ys__n45372 & ~new_n14565_;
  assign new_n14567_ = ~new_n14564_ & new_n14566_;
  assign new_n14568_ = ~new_n14563_ & ~new_n14567_;
  assign new_n14569_ = ys__n45166 & ys__n45342;
  assign new_n14570_ = ~ys__n45166 & ~ys__n45342;
  assign new_n14571_ = ~ys__n45372 & ~new_n14570_;
  assign new_n14572_ = ~new_n14569_ & new_n14571_;
  assign new_n14573_ = ys__n45169 & ys__n45344;
  assign new_n14574_ = ~ys__n45169 & ~ys__n45344;
  assign new_n14575_ = ~ys__n45372 & ~new_n14574_;
  assign new_n14576_ = ~new_n14573_ & new_n14575_;
  assign new_n14577_ = ~new_n14572_ & ~new_n14576_;
  assign new_n14578_ = new_n14568_ & new_n14577_;
  assign new_n14579_ = new_n14559_ & new_n14578_;
  assign new_n14580_ = ys__n45196 & ys__n45362;
  assign new_n14581_ = ~ys__n45196 & ~ys__n45362;
  assign new_n14582_ = ~ys__n45373 & ~new_n14581_;
  assign new_n14583_ = ~new_n14580_ & new_n14582_;
  assign new_n14584_ = ys__n45199 & ys__n45364;
  assign new_n14585_ = ~ys__n45199 & ~ys__n45364;
  assign new_n14586_ = ~ys__n45373 & ~new_n14585_;
  assign new_n14587_ = ~new_n14584_ & new_n14586_;
  assign new_n14588_ = ~new_n14583_ & ~new_n14587_;
  assign new_n14589_ = ys__n45202 & ys__n45366;
  assign new_n14590_ = ~ys__n45202 & ~ys__n45366;
  assign new_n14591_ = ~ys__n45373 & ~new_n14590_;
  assign new_n14592_ = ~new_n14589_ & new_n14591_;
  assign new_n14593_ = ys__n45205 & ys__n45368;
  assign new_n14594_ = ~ys__n45205 & ~ys__n45368;
  assign new_n14595_ = ~ys__n45373 & ~new_n14594_;
  assign new_n14596_ = ~new_n14593_ & new_n14595_;
  assign new_n14597_ = ~new_n14592_ & ~new_n14596_;
  assign new_n14598_ = new_n14588_ & new_n14597_;
  assign new_n14599_ = ys__n45184 & ys__n45354;
  assign new_n14600_ = ~ys__n45184 & ~ys__n45354;
  assign new_n14601_ = ~ys__n45373 & ~new_n14600_;
  assign new_n14602_ = ~new_n14599_ & new_n14601_;
  assign new_n14603_ = ys__n45187 & ys__n45356;
  assign new_n14604_ = ~ys__n45187 & ~ys__n45356;
  assign new_n14605_ = ~ys__n45373 & ~new_n14604_;
  assign new_n14606_ = ~new_n14603_ & new_n14605_;
  assign new_n14607_ = ~new_n14602_ & ~new_n14606_;
  assign new_n14608_ = ys__n45190 & ys__n45358;
  assign new_n14609_ = ~ys__n45190 & ~ys__n45358;
  assign new_n14610_ = ~ys__n45373 & ~new_n14609_;
  assign new_n14611_ = ~new_n14608_ & new_n14610_;
  assign new_n14612_ = ys__n45193 & ys__n45360;
  assign new_n14613_ = ~ys__n45193 & ~ys__n45360;
  assign new_n14614_ = ~ys__n45373 & ~new_n14613_;
  assign new_n14615_ = ~new_n14612_ & new_n14614_;
  assign new_n14616_ = ~new_n14611_ & ~new_n14615_;
  assign new_n14617_ = new_n14607_ & new_n14616_;
  assign new_n14618_ = new_n14598_ & new_n14617_;
  assign new_n14619_ = new_n14579_ & new_n14618_;
  assign new_n14620_ = ys__n45124 & ys__n45314;
  assign new_n14621_ = ~ys__n45124 & ~ys__n45314;
  assign new_n14622_ = ~ys__n45370 & ~new_n14621_;
  assign new_n14623_ = ~new_n14620_ & new_n14622_;
  assign new_n14624_ = ys__n45127 & ys__n45316;
  assign new_n14625_ = ~ys__n45127 & ~ys__n45316;
  assign new_n14626_ = ~ys__n45370 & ~new_n14625_;
  assign new_n14627_ = ~new_n14624_ & new_n14626_;
  assign new_n14628_ = ~new_n14623_ & ~new_n14627_;
  assign new_n14629_ = ys__n45130 & ys__n45318;
  assign new_n14630_ = ~ys__n45130 & ~ys__n45318;
  assign new_n14631_ = ~ys__n45370 & ~new_n14630_;
  assign new_n14632_ = ~new_n14629_ & new_n14631_;
  assign new_n14633_ = ys__n45133 & ys__n45320;
  assign new_n14634_ = ~ys__n45133 & ~ys__n45320;
  assign new_n14635_ = ~ys__n45370 & ~new_n14634_;
  assign new_n14636_ = ~new_n14633_ & new_n14635_;
  assign new_n14637_ = ~new_n14632_ & ~new_n14636_;
  assign new_n14638_ = new_n14628_ & new_n14637_;
  assign new_n14639_ = ys__n45112 & ys__n45306;
  assign new_n14640_ = ~ys__n45112 & ~ys__n45306;
  assign new_n14641_ = ~ys__n45370 & ~new_n14640_;
  assign new_n14642_ = ~new_n14639_ & new_n14641_;
  assign new_n14643_ = ys__n45115 & ys__n45308;
  assign new_n14644_ = ~ys__n45115 & ~ys__n45308;
  assign new_n14645_ = ~ys__n45370 & ~new_n14644_;
  assign new_n14646_ = ~new_n14643_ & new_n14645_;
  assign new_n14647_ = ~new_n14642_ & ~new_n14646_;
  assign new_n14648_ = ys__n45118 & ys__n45310;
  assign new_n14649_ = ~ys__n45118 & ~ys__n45310;
  assign new_n14650_ = ~ys__n45370 & ~new_n14649_;
  assign new_n14651_ = ~new_n14648_ & new_n14650_;
  assign new_n14652_ = ys__n45121 & ys__n45312;
  assign new_n14653_ = ~ys__n45121 & ~ys__n45312;
  assign new_n14654_ = ~ys__n45370 & ~new_n14653_;
  assign new_n14655_ = ~new_n14652_ & new_n14654_;
  assign new_n14656_ = ~new_n14651_ & ~new_n14655_;
  assign new_n14657_ = new_n14647_ & new_n14656_;
  assign new_n14658_ = new_n14638_ & new_n14657_;
  assign new_n14659_ = ys__n45148 & ys__n45330;
  assign new_n14660_ = ~ys__n45148 & ~ys__n45330;
  assign new_n14661_ = ~ys__n45371 & ~new_n14660_;
  assign new_n14662_ = ~new_n14659_ & new_n14661_;
  assign new_n14663_ = ys__n45151 & ys__n45332;
  assign new_n14664_ = ~ys__n45151 & ~ys__n45332;
  assign new_n14665_ = ~ys__n45371 & ~new_n14664_;
  assign new_n14666_ = ~new_n14663_ & new_n14665_;
  assign new_n14667_ = ~new_n14662_ & ~new_n14666_;
  assign new_n14668_ = ys__n45154 & ys__n45334;
  assign new_n14669_ = ~ys__n45154 & ~ys__n45334;
  assign new_n14670_ = ~ys__n45371 & ~new_n14669_;
  assign new_n14671_ = ~new_n14668_ & new_n14670_;
  assign new_n14672_ = ys__n45157 & ys__n45336;
  assign new_n14673_ = ~ys__n45157 & ~ys__n45336;
  assign new_n14674_ = ~ys__n45371 & ~new_n14673_;
  assign new_n14675_ = ~new_n14672_ & new_n14674_;
  assign new_n14676_ = ~new_n14671_ & ~new_n14675_;
  assign new_n14677_ = new_n14667_ & new_n14676_;
  assign new_n14678_ = ys__n45136 & ys__n45322;
  assign new_n14679_ = ~ys__n45136 & ~ys__n45322;
  assign new_n14680_ = ~ys__n45371 & ~new_n14679_;
  assign new_n14681_ = ~new_n14678_ & new_n14680_;
  assign new_n14682_ = ys__n45139 & ys__n45324;
  assign new_n14683_ = ~ys__n45139 & ~ys__n45324;
  assign new_n14684_ = ~ys__n45371 & ~new_n14683_;
  assign new_n14685_ = ~new_n14682_ & new_n14684_;
  assign new_n14686_ = ~new_n14681_ & ~new_n14685_;
  assign new_n14687_ = ys__n45142 & ys__n45326;
  assign new_n14688_ = ~ys__n45142 & ~ys__n45326;
  assign new_n14689_ = ~ys__n45371 & ~new_n14688_;
  assign new_n14690_ = ~new_n14687_ & new_n14689_;
  assign new_n14691_ = ys__n45145 & ys__n45328;
  assign new_n14692_ = ~ys__n45145 & ~ys__n45328;
  assign new_n14693_ = ~ys__n45371 & ~new_n14692_;
  assign new_n14694_ = ~new_n14691_ & new_n14693_;
  assign new_n14695_ = ~new_n14690_ & ~new_n14694_;
  assign new_n14696_ = new_n14686_ & new_n14695_;
  assign new_n14697_ = new_n14677_ & new_n14696_;
  assign new_n14698_ = new_n14658_ & new_n14697_;
  assign new_n14699_ = new_n14619_ & new_n14698_;
  assign new_n14700_ = new_n14540_ & new_n14699_;
  assign new_n14701_ = ys__n45374 & new_n14700_;
  assign new_n14702_ = ys__n45046 & ys__n45047;
  assign new_n14703_ = ~ys__n45046 & ~ys__n45047;
  assign new_n14704_ = ~ys__n45100 & ~new_n14703_;
  assign new_n14705_ = ~new_n14702_ & new_n14704_;
  assign new_n14706_ = ys__n45049 & ys__n45050;
  assign new_n14707_ = ~ys__n45049 & ~ys__n45050;
  assign new_n14708_ = ~ys__n45101 & ~new_n14707_;
  assign new_n14709_ = ~new_n14706_ & new_n14708_;
  assign new_n14710_ = ~new_n14705_ & ~new_n14709_;
  assign new_n14711_ = ys__n45052 & ys__n45053;
  assign new_n14712_ = ~ys__n45052 & ~ys__n45053;
  assign new_n14713_ = ~ys__n45102 & ~new_n14712_;
  assign new_n14714_ = ~new_n14711_ & new_n14713_;
  assign new_n14715_ = ys__n45055 & ys__n45056;
  assign new_n14716_ = ~ys__n45055 & ~ys__n45056;
  assign new_n14717_ = ~ys__n45103 & ~new_n14716_;
  assign new_n14718_ = ~new_n14715_ & new_n14717_;
  assign new_n14719_ = ~new_n14714_ & ~new_n14718_;
  assign new_n14720_ = new_n14710_ & new_n14719_;
  assign new_n14721_ = ys__n45034 & ys__n45035;
  assign new_n14722_ = ~ys__n45034 & ~ys__n45035;
  assign new_n14723_ = ~ys__n45096 & ~new_n14722_;
  assign new_n14724_ = ~new_n14721_ & new_n14723_;
  assign new_n14725_ = ys__n45037 & ys__n45038;
  assign new_n14726_ = ~ys__n45037 & ~ys__n45038;
  assign new_n14727_ = ~ys__n45097 & ~new_n14726_;
  assign new_n14728_ = ~new_n14725_ & new_n14727_;
  assign new_n14729_ = ~new_n14724_ & ~new_n14728_;
  assign new_n14730_ = ys__n45040 & ys__n45041;
  assign new_n14731_ = ~ys__n45040 & ~ys__n45041;
  assign new_n14732_ = ~ys__n45098 & ~new_n14731_;
  assign new_n14733_ = ~new_n14730_ & new_n14732_;
  assign new_n14734_ = ys__n45043 & ys__n45044;
  assign new_n14735_ = ~ys__n45043 & ~ys__n45044;
  assign new_n14736_ = ~ys__n45099 & ~new_n14735_;
  assign new_n14737_ = ~new_n14734_ & new_n14736_;
  assign new_n14738_ = ~new_n14733_ & ~new_n14737_;
  assign new_n14739_ = new_n14729_ & new_n14738_;
  assign new_n14740_ = new_n14720_ & new_n14739_;
  assign new_n14741_ = ys__n45070 & ys__n45071;
  assign new_n14742_ = ~ys__n45070 & ~ys__n45071;
  assign new_n14743_ = ~ys__n45108 & ~new_n14742_;
  assign new_n14744_ = ~new_n14741_ & new_n14743_;
  assign new_n14745_ = ys__n45073 & ys__n45074;
  assign new_n14746_ = ~ys__n45073 & ~ys__n45074;
  assign new_n14747_ = ~ys__n45109 & ~new_n14746_;
  assign new_n14748_ = ~new_n14745_ & new_n14747_;
  assign new_n14749_ = ~new_n14744_ & ~new_n14748_;
  assign new_n14750_ = ys__n45076 & ys__n45077;
  assign new_n14751_ = ~ys__n45076 & ~ys__n45077;
  assign new_n14752_ = ~ys__n45110 & ~new_n14751_;
  assign new_n14753_ = ~new_n14750_ & new_n14752_;
  assign new_n14754_ = ys__n45079 & ys__n45080;
  assign new_n14755_ = ~ys__n45079 & ~ys__n45080;
  assign new_n14756_ = ~ys__n45111 & ~new_n14755_;
  assign new_n14757_ = ~new_n14754_ & new_n14756_;
  assign new_n14758_ = ~new_n14753_ & ~new_n14757_;
  assign new_n14759_ = new_n14749_ & new_n14758_;
  assign new_n14760_ = ys__n45058 & ys__n45059;
  assign new_n14761_ = ~ys__n45058 & ~ys__n45059;
  assign new_n14762_ = ~ys__n45104 & ~new_n14761_;
  assign new_n14763_ = ~new_n14760_ & new_n14762_;
  assign new_n14764_ = ys__n45061 & ys__n45062;
  assign new_n14765_ = ~ys__n45061 & ~ys__n45062;
  assign new_n14766_ = ~ys__n45105 & ~new_n14765_;
  assign new_n14767_ = ~new_n14764_ & new_n14766_;
  assign new_n14768_ = ~new_n14763_ & ~new_n14767_;
  assign new_n14769_ = ys__n45064 & ys__n45065;
  assign new_n14770_ = ~ys__n45064 & ~ys__n45065;
  assign new_n14771_ = ~ys__n45106 & ~new_n14770_;
  assign new_n14772_ = ~new_n14769_ & new_n14771_;
  assign new_n14773_ = ys__n45067 & ys__n45068;
  assign new_n14774_ = ~ys__n45067 & ~ys__n45068;
  assign new_n14775_ = ~ys__n45107 & ~new_n14774_;
  assign new_n14776_ = ~new_n14773_ & new_n14775_;
  assign new_n14777_ = ~new_n14772_ & ~new_n14776_;
  assign new_n14778_ = new_n14768_ & new_n14777_;
  assign new_n14779_ = new_n14759_ & new_n14778_;
  assign new_n14780_ = new_n14740_ & new_n14779_;
  assign new_n14781_ = ys__n44992 & ys__n44993;
  assign new_n14782_ = ~ys__n44992 & ~ys__n44993;
  assign new_n14783_ = ~ys__n45082 & ~new_n14782_;
  assign new_n14784_ = ~new_n14781_ & new_n14783_;
  assign new_n14785_ = ys__n44995 & ys__n44996;
  assign new_n14786_ = ~ys__n44995 & ~ys__n44996;
  assign new_n14787_ = ~ys__n45083 & ~new_n14786_;
  assign new_n14788_ = ~new_n14785_ & new_n14787_;
  assign new_n14789_ = ~new_n14784_ & ~new_n14788_;
  assign new_n14790_ = ys__n44998 & ys__n44999;
  assign new_n14791_ = ~ys__n44998 & ~ys__n44999;
  assign new_n14792_ = ~ys__n45084 & ~new_n14791_;
  assign new_n14793_ = ~new_n14790_ & new_n14792_;
  assign new_n14794_ = ys__n45001 & ys__n45002;
  assign new_n14795_ = ~ys__n45001 & ~ys__n45002;
  assign new_n14796_ = ~ys__n45085 & ~new_n14795_;
  assign new_n14797_ = ~new_n14794_ & new_n14796_;
  assign new_n14798_ = ~new_n14793_ & ~new_n14797_;
  assign new_n14799_ = ys__n45004 & ys__n45005;
  assign new_n14800_ = ~ys__n45004 & ~ys__n45005;
  assign new_n14801_ = ~ys__n45086 & ~new_n14800_;
  assign new_n14802_ = ~new_n14799_ & new_n14801_;
  assign new_n14803_ = ys__n45007 & ys__n45008;
  assign new_n14804_ = ~ys__n45007 & ~ys__n45008;
  assign new_n14805_ = ~ys__n45087 & ~new_n14804_;
  assign new_n14806_ = ~new_n14803_ & new_n14805_;
  assign new_n14807_ = ~new_n14802_ & ~new_n14806_;
  assign new_n14808_ = new_n14798_ & new_n14807_;
  assign new_n14809_ = new_n14789_ & new_n14808_;
  assign new_n14810_ = ys__n45022 & ys__n45023;
  assign new_n14811_ = ~ys__n45022 & ~ys__n45023;
  assign new_n14812_ = ~ys__n45092 & ~new_n14811_;
  assign new_n14813_ = ~new_n14810_ & new_n14812_;
  assign new_n14814_ = ys__n45025 & ys__n45026;
  assign new_n14815_ = ~ys__n45025 & ~ys__n45026;
  assign new_n14816_ = ~ys__n45093 & ~new_n14815_;
  assign new_n14817_ = ~new_n14814_ & new_n14816_;
  assign new_n14818_ = ~new_n14813_ & ~new_n14817_;
  assign new_n14819_ = ys__n45028 & ys__n45029;
  assign new_n14820_ = ~ys__n45028 & ~ys__n45029;
  assign new_n14821_ = ~ys__n45094 & ~new_n14820_;
  assign new_n14822_ = ~new_n14819_ & new_n14821_;
  assign new_n14823_ = ys__n45031 & ys__n45032;
  assign new_n14824_ = ~ys__n45031 & ~ys__n45032;
  assign new_n14825_ = ~ys__n45095 & ~new_n14824_;
  assign new_n14826_ = ~new_n14823_ & new_n14825_;
  assign new_n14827_ = ~new_n14822_ & ~new_n14826_;
  assign new_n14828_ = new_n14818_ & new_n14827_;
  assign new_n14829_ = ys__n45010 & ys__n45011;
  assign new_n14830_ = ~ys__n45010 & ~ys__n45011;
  assign new_n14831_ = ~ys__n45088 & ~new_n14830_;
  assign new_n14832_ = ~new_n14829_ & new_n14831_;
  assign new_n14833_ = ys__n45013 & ys__n45014;
  assign new_n14834_ = ~ys__n45013 & ~ys__n45014;
  assign new_n14835_ = ~ys__n45089 & ~new_n14834_;
  assign new_n14836_ = ~new_n14833_ & new_n14835_;
  assign new_n14837_ = ~new_n14832_ & ~new_n14836_;
  assign new_n14838_ = ys__n45016 & ys__n45017;
  assign new_n14839_ = ~ys__n45016 & ~ys__n45017;
  assign new_n14840_ = ~ys__n45090 & ~new_n14839_;
  assign new_n14841_ = ~new_n14838_ & new_n14840_;
  assign new_n14842_ = ys__n45019 & ys__n45020;
  assign new_n14843_ = ~ys__n45019 & ~ys__n45020;
  assign new_n14844_ = ~ys__n45091 & ~new_n14843_;
  assign new_n14845_ = ~new_n14842_ & new_n14844_;
  assign new_n14846_ = ~new_n14841_ & ~new_n14845_;
  assign new_n14847_ = new_n14837_ & new_n14846_;
  assign new_n14848_ = new_n14828_ & new_n14847_;
  assign new_n14849_ = new_n14809_ & new_n14848_;
  assign new_n14850_ = new_n14780_ & new_n14849_;
  assign new_n14851_ = ys__n45172 & ys__n45173;
  assign new_n14852_ = ~ys__n45172 & ~ys__n45173;
  assign new_n14853_ = ~ys__n45210 & ~new_n14852_;
  assign new_n14854_ = ~new_n14851_ & new_n14853_;
  assign new_n14855_ = ys__n45175 & ys__n45176;
  assign new_n14856_ = ~ys__n45175 & ~ys__n45176;
  assign new_n14857_ = ~ys__n45210 & ~new_n14856_;
  assign new_n14858_ = ~new_n14855_ & new_n14857_;
  assign new_n14859_ = ~new_n14854_ & ~new_n14858_;
  assign new_n14860_ = ys__n45178 & ys__n45179;
  assign new_n14861_ = ~ys__n45178 & ~ys__n45179;
  assign new_n14862_ = ~ys__n45210 & ~new_n14861_;
  assign new_n14863_ = ~new_n14860_ & new_n14862_;
  assign new_n14864_ = ys__n45181 & ys__n45182;
  assign new_n14865_ = ~ys__n45181 & ~ys__n45182;
  assign new_n14866_ = ~ys__n45210 & ~new_n14865_;
  assign new_n14867_ = ~new_n14864_ & new_n14866_;
  assign new_n14868_ = ~new_n14863_ & ~new_n14867_;
  assign new_n14869_ = new_n14859_ & new_n14868_;
  assign new_n14870_ = ys__n45160 & ys__n45161;
  assign new_n14871_ = ~ys__n45160 & ~ys__n45161;
  assign new_n14872_ = ~ys__n45210 & ~new_n14871_;
  assign new_n14873_ = ~new_n14870_ & new_n14872_;
  assign new_n14874_ = ys__n45163 & ys__n45164;
  assign new_n14875_ = ~ys__n45163 & ~ys__n45164;
  assign new_n14876_ = ~ys__n45210 & ~new_n14875_;
  assign new_n14877_ = ~new_n14874_ & new_n14876_;
  assign new_n14878_ = ~new_n14873_ & ~new_n14877_;
  assign new_n14879_ = ys__n45166 & ys__n45167;
  assign new_n14880_ = ~ys__n45166 & ~ys__n45167;
  assign new_n14881_ = ~ys__n45210 & ~new_n14880_;
  assign new_n14882_ = ~new_n14879_ & new_n14881_;
  assign new_n14883_ = ys__n45169 & ys__n45170;
  assign new_n14884_ = ~ys__n45169 & ~ys__n45170;
  assign new_n14885_ = ~ys__n45210 & ~new_n14884_;
  assign new_n14886_ = ~new_n14883_ & new_n14885_;
  assign new_n14887_ = ~new_n14882_ & ~new_n14886_;
  assign new_n14888_ = new_n14878_ & new_n14887_;
  assign new_n14889_ = new_n14869_ & new_n14888_;
  assign new_n14890_ = ys__n45196 & ys__n45197;
  assign new_n14891_ = ~ys__n45196 & ~ys__n45197;
  assign new_n14892_ = ~ys__n45211 & ~new_n14891_;
  assign new_n14893_ = ~new_n14890_ & new_n14892_;
  assign new_n14894_ = ys__n45199 & ys__n45200;
  assign new_n14895_ = ~ys__n45199 & ~ys__n45200;
  assign new_n14896_ = ~ys__n45211 & ~new_n14895_;
  assign new_n14897_ = ~new_n14894_ & new_n14896_;
  assign new_n14898_ = ~new_n14893_ & ~new_n14897_;
  assign new_n14899_ = ys__n45202 & ys__n45203;
  assign new_n14900_ = ~ys__n45202 & ~ys__n45203;
  assign new_n14901_ = ~ys__n45211 & ~new_n14900_;
  assign new_n14902_ = ~new_n14899_ & new_n14901_;
  assign new_n14903_ = ys__n45205 & ys__n45206;
  assign new_n14904_ = ~ys__n45205 & ~ys__n45206;
  assign new_n14905_ = ~ys__n45211 & ~new_n14904_;
  assign new_n14906_ = ~new_n14903_ & new_n14905_;
  assign new_n14907_ = ~new_n14902_ & ~new_n14906_;
  assign new_n14908_ = new_n14898_ & new_n14907_;
  assign new_n14909_ = ys__n45184 & ys__n45185;
  assign new_n14910_ = ~ys__n45184 & ~ys__n45185;
  assign new_n14911_ = ~ys__n45211 & ~new_n14910_;
  assign new_n14912_ = ~new_n14909_ & new_n14911_;
  assign new_n14913_ = ys__n45187 & ys__n45188;
  assign new_n14914_ = ~ys__n45187 & ~ys__n45188;
  assign new_n14915_ = ~ys__n45211 & ~new_n14914_;
  assign new_n14916_ = ~new_n14913_ & new_n14915_;
  assign new_n14917_ = ~new_n14912_ & ~new_n14916_;
  assign new_n14918_ = ys__n45190 & ys__n45191;
  assign new_n14919_ = ~ys__n45190 & ~ys__n45191;
  assign new_n14920_ = ~ys__n45211 & ~new_n14919_;
  assign new_n14921_ = ~new_n14918_ & new_n14920_;
  assign new_n14922_ = ys__n45193 & ys__n45194;
  assign new_n14923_ = ~ys__n45193 & ~ys__n45194;
  assign new_n14924_ = ~ys__n45211 & ~new_n14923_;
  assign new_n14925_ = ~new_n14922_ & new_n14924_;
  assign new_n14926_ = ~new_n14921_ & ~new_n14925_;
  assign new_n14927_ = new_n14917_ & new_n14926_;
  assign new_n14928_ = new_n14908_ & new_n14927_;
  assign new_n14929_ = new_n14889_ & new_n14928_;
  assign new_n14930_ = ys__n45124 & ys__n45125;
  assign new_n14931_ = ~ys__n45124 & ~ys__n45125;
  assign new_n14932_ = ~ys__n45208 & ~new_n14931_;
  assign new_n14933_ = ~new_n14930_ & new_n14932_;
  assign new_n14934_ = ys__n45127 & ys__n45128;
  assign new_n14935_ = ~ys__n45127 & ~ys__n45128;
  assign new_n14936_ = ~ys__n45208 & ~new_n14935_;
  assign new_n14937_ = ~new_n14934_ & new_n14936_;
  assign new_n14938_ = ~new_n14933_ & ~new_n14937_;
  assign new_n14939_ = ys__n45130 & ys__n45131;
  assign new_n14940_ = ~ys__n45130 & ~ys__n45131;
  assign new_n14941_ = ~ys__n45208 & ~new_n14940_;
  assign new_n14942_ = ~new_n14939_ & new_n14941_;
  assign new_n14943_ = ys__n45133 & ys__n45134;
  assign new_n14944_ = ~ys__n45133 & ~ys__n45134;
  assign new_n14945_ = ~ys__n45208 & ~new_n14944_;
  assign new_n14946_ = ~new_n14943_ & new_n14945_;
  assign new_n14947_ = ~new_n14942_ & ~new_n14946_;
  assign new_n14948_ = new_n14938_ & new_n14947_;
  assign new_n14949_ = ys__n45112 & ys__n45113;
  assign new_n14950_ = ~ys__n45112 & ~ys__n45113;
  assign new_n14951_ = ~ys__n45208 & ~new_n14950_;
  assign new_n14952_ = ~new_n14949_ & new_n14951_;
  assign new_n14953_ = ys__n45115 & ys__n45116;
  assign new_n14954_ = ~ys__n45115 & ~ys__n45116;
  assign new_n14955_ = ~ys__n45208 & ~new_n14954_;
  assign new_n14956_ = ~new_n14953_ & new_n14955_;
  assign new_n14957_ = ~new_n14952_ & ~new_n14956_;
  assign new_n14958_ = ys__n45118 & ys__n45119;
  assign new_n14959_ = ~ys__n45118 & ~ys__n45119;
  assign new_n14960_ = ~ys__n45208 & ~new_n14959_;
  assign new_n14961_ = ~new_n14958_ & new_n14960_;
  assign new_n14962_ = ys__n45121 & ys__n45122;
  assign new_n14963_ = ~ys__n45121 & ~ys__n45122;
  assign new_n14964_ = ~ys__n45208 & ~new_n14963_;
  assign new_n14965_ = ~new_n14962_ & new_n14964_;
  assign new_n14966_ = ~new_n14961_ & ~new_n14965_;
  assign new_n14967_ = new_n14957_ & new_n14966_;
  assign new_n14968_ = new_n14948_ & new_n14967_;
  assign new_n14969_ = ys__n45148 & ys__n45149;
  assign new_n14970_ = ~ys__n45148 & ~ys__n45149;
  assign new_n14971_ = ~ys__n45209 & ~new_n14970_;
  assign new_n14972_ = ~new_n14969_ & new_n14971_;
  assign new_n14973_ = ys__n45151 & ys__n45152;
  assign new_n14974_ = ~ys__n45151 & ~ys__n45152;
  assign new_n14975_ = ~ys__n45209 & ~new_n14974_;
  assign new_n14976_ = ~new_n14973_ & new_n14975_;
  assign new_n14977_ = ~new_n14972_ & ~new_n14976_;
  assign new_n14978_ = ys__n45154 & ys__n45155;
  assign new_n14979_ = ~ys__n45154 & ~ys__n45155;
  assign new_n14980_ = ~ys__n45209 & ~new_n14979_;
  assign new_n14981_ = ~new_n14978_ & new_n14980_;
  assign new_n14982_ = ys__n45157 & ys__n45158;
  assign new_n14983_ = ~ys__n45157 & ~ys__n45158;
  assign new_n14984_ = ~ys__n45209 & ~new_n14983_;
  assign new_n14985_ = ~new_n14982_ & new_n14984_;
  assign new_n14986_ = ~new_n14981_ & ~new_n14985_;
  assign new_n14987_ = new_n14977_ & new_n14986_;
  assign new_n14988_ = ys__n45136 & ys__n45137;
  assign new_n14989_ = ~ys__n45136 & ~ys__n45137;
  assign new_n14990_ = ~ys__n45209 & ~new_n14989_;
  assign new_n14991_ = ~new_n14988_ & new_n14990_;
  assign new_n14992_ = ys__n45139 & ys__n45140;
  assign new_n14993_ = ~ys__n45139 & ~ys__n45140;
  assign new_n14994_ = ~ys__n45209 & ~new_n14993_;
  assign new_n14995_ = ~new_n14992_ & new_n14994_;
  assign new_n14996_ = ~new_n14991_ & ~new_n14995_;
  assign new_n14997_ = ys__n45142 & ys__n45143;
  assign new_n14998_ = ~ys__n45142 & ~ys__n45143;
  assign new_n14999_ = ~ys__n45209 & ~new_n14998_;
  assign new_n15000_ = ~new_n14997_ & new_n14999_;
  assign new_n15001_ = ys__n45145 & ys__n45146;
  assign new_n15002_ = ~ys__n45145 & ~ys__n45146;
  assign new_n15003_ = ~ys__n45209 & ~new_n15002_;
  assign new_n15004_ = ~new_n15001_ & new_n15003_;
  assign new_n15005_ = ~new_n15000_ & ~new_n15004_;
  assign new_n15006_ = new_n14996_ & new_n15005_;
  assign new_n15007_ = new_n14987_ & new_n15006_;
  assign new_n15008_ = new_n14968_ & new_n15007_;
  assign new_n15009_ = new_n14929_ & new_n15008_;
  assign new_n15010_ = new_n14850_ & new_n15009_;
  assign new_n15011_ = ys__n45212 & new_n15010_;
  assign new_n15012_ = ~new_n14701_ & ~new_n15011_;
  assign new_n15013_ = new_n14391_ & new_n15012_;
  assign new_n15014_ = ~ys__n23850 & ~ys__n30214;
  assign new_n15015_ = ys__n38906 & new_n15014_;
  assign new_n15016_ = ~ys__n38902 & ~ys__n38904;
  assign new_n15017_ = ~new_n15015_ & new_n15016_;
  assign new_n15018_ = ~new_n15013_ & ~new_n15017_;
  assign new_n15019_ = ~ys__n262 & ~ys__n18101;
  assign new_n15020_ = ~ys__n18106 & new_n15019_;
  assign new_n15021_ = ~ys__n4566 & new_n15020_;
  assign new_n15022_ = ~ys__n22799 & ys__n38272;
  assign new_n15023_ = ys__n22794 & ~ys__n33359;
  assign new_n15024_ = ~ys__n33375 & ~ys__n33389;
  assign new_n15025_ = new_n15023_ & new_n15024_;
  assign ys__n33357 = ~new_n15022_ & new_n15025_;
  assign new_n15027_ = ~ys__n33375 & ~ys__n33357;
  assign new_n15028_ = ~ys__n33350 & ~ys__n33352;
  assign new_n15029_ = new_n15027_ & new_n15028_;
  assign new_n15030_ = ys__n38259 & new_n15029_;
  assign new_n15031_ = new_n15029_ & ~new_n15030_;
  assign new_n15032_ = ys__n38257 & new_n15031_;
  assign new_n15033_ = ~ys__n38278 & ~ys__n38279;
  assign new_n15034_ = ~ys__n38277 & new_n15033_;
  assign new_n15035_ = new_n15031_ & ~new_n15034_;
  assign new_n15036_ = ~new_n15032_ & new_n15035_;
  assign new_n15037_ = ys__n33350 & new_n15027_;
  assign new_n15038_ = ys__n33352 & new_n15027_;
  assign new_n15039_ = ~ys__n33357 & ~new_n15038_;
  assign new_n15040_ = ~new_n15037_ & new_n15039_;
  assign new_n15041_ = ~new_n15030_ & new_n15040_;
  assign new_n15042_ = ~new_n15032_ & new_n15041_;
  assign new_n15043_ = ~new_n15036_ & new_n15042_;
  assign new_n15044_ = new_n15021_ & ~new_n15043_;
  assign new_n15045_ = ~ys__n738 & new_n15044_;
  assign new_n15046_ = ~new_n15018_ & new_n15045_;
  assign new_n15047_ = ys__n38236 & new_n15027_;
  assign new_n15048_ = ys__n38237 & new_n15027_;
  assign new_n15049_ = ~new_n15047_ & ~new_n15048_;
  assign new_n15050_ = new_n15040_ & new_n15049_;
  assign new_n15051_ = new_n15021_ & ~new_n15050_;
  assign new_n15052_ = ~ys__n738 & new_n15051_;
  assign new_n15053_ = new_n15018_ & new_n15052_;
  assign new_n15054_ = ~new_n15046_ & ~new_n15053_;
  assign new_n15055_ = ys__n874 & ~ys__n738;
  assign new_n15056_ = new_n15030_ & new_n15055_;
  assign new_n15057_ = ~new_n15018_ & new_n15056_;
  assign ys__n2491 = ~new_n15054_ & new_n15057_;
  assign ys__n2535 = ys__n196 & ~ys__n4566;
  assign ys__n2536 = ys__n874 & ys__n2535;
  assign new_n15061_ = ~ys__n768 & ~ys__n776;
  assign new_n15062_ = ~ys__n778 & ~ys__n4168;
  assign new_n15063_ = new_n15061_ & new_n15062_;
  assign new_n15064_ = ~ys__n600 & ~ys__n602;
  assign new_n15065_ = ~ys__n604 & ~ys__n698;
  assign new_n15066_ = new_n15064_ & new_n15065_;
  assign new_n15067_ = ~ys__n598 & ~ys__n774;
  assign new_n15068_ = ~ys__n770 & ~ys__n784;
  assign new_n15069_ = new_n15067_ & ~new_n15068_;
  assign new_n15070_ = new_n15066_ & new_n15069_;
  assign ys__n2582 = new_n15063_ & new_n15070_;
  assign new_n15072_ = new_n13376_ & new_n13492_;
  assign ys__n2635 = new_n13530_ & new_n15072_;
  assign new_n15074_ = ~ys__n4832 & ~ys__n4833;
  assign new_n15075_ = ys__n164 & ~ys__n4826;
  assign new_n15076_ = ys__n354 & new_n15075_;
  assign ys__n2651 = new_n15074_ & new_n15076_;
  assign ys__n2653 = ys__n2652 | ys__n2651;
  assign new_n15079_ = new_n13375_ & new_n13492_;
  assign ys__n2655 = new_n13530_ & new_n15079_;
  assign new_n15081_ = new_n13375_ & new_n13503_;
  assign ys__n2674 = new_n13530_ & new_n15081_;
  assign ys__n2684 = new_n13421_ & new_n13545_;
  assign new_n15084_ = ~ys__n738 & new_n15027_;
  assign new_n15085_ = new_n15021_ & new_n15084_;
  assign ys__n2733 = ~ys__n874 | new_n15085_;
  assign ys__n2776 = new_n13421_ & new_n13509_;
  assign new_n15088_ = ys__n38219 & ~ys__n738;
  assign ys__n2778 = ~ys__n4566 & new_n15088_;
  assign ys__n2780 = ys__n874 & ys__n2779;
  assign ys__n2782 = ~ys__n740 | new_n13344_;
  assign new_n15092_ = ~ys__n738 & ~new_n15049_;
  assign new_n15093_ = ~new_n15054_ & new_n15092_;
  assign new_n15094_ = ~new_n15037_ & ~new_n15038_;
  assign new_n15095_ = ~ys__n738 & ~new_n15094_;
  assign new_n15096_ = ~new_n15054_ & new_n15095_;
  assign ys__n2804 = new_n15093_ | new_n15096_;
  assign new_n15098_ = ys__n874 & ~ys__n34959;
  assign ys__n2806 = ys__n740 & new_n15098_;
  assign new_n15100_ = ~new_n12205_ & ~new_n12212_;
  assign new_n15101_ = new_n12212_ & ~new_n12842_;
  assign ys__n2845 = ~new_n15100_ & ~new_n15101_;
  assign new_n15103_ = ys__n828 & ~new_n12861_;
  assign new_n15104_ = ~new_n12861_ & ~new_n15103_;
  assign new_n15105_ = ~new_n12865_ & ~new_n15104_;
  assign new_n15106_ = ys__n826 & new_n12865_;
  assign ys__n4603 = new_n15105_ | new_n15106_;
  assign new_n15108_ = ~new_n12860_ & ~ys__n4603;
  assign new_n15109_ = new_n12861_ & ys__n730;
  assign new_n15110_ = ~ys__n732 & new_n12860_;
  assign new_n15111_ = ~new_n15109_ & ~new_n15110_;
  assign ys__n2855 = ~new_n15108_ & new_n15111_;
  assign ys__n3024 = new_n13421_ & new_n13517_;
  assign ys__n3035 = ~ys__n740 | new_n13311_;
  assign new_n15115_ = ~ys__n452 & ys__n24427;
  assign new_n15116_ = ys__n452 & ~ys__n24427;
  assign new_n15117_ = ~new_n15115_ & ~new_n15116_;
  assign new_n15118_ = ~ys__n35426 & ys__n38695;
  assign new_n15119_ = ys__n35426 & ~ys__n38695;
  assign new_n15120_ = ~new_n15118_ & ~new_n15119_;
  assign new_n15121_ = new_n15117_ & new_n15120_;
  assign new_n15122_ = ys__n1098 & ys__n24519;
  assign new_n15123_ = new_n15121_ & new_n15122_;
  assign new_n15124_ = ys__n24463 & ys__n24519;
  assign new_n15125_ = ~ys__n1110 & ~ys__n1120;
  assign new_n15126_ = ~new_n15124_ & new_n15125_;
  assign ys__n3039 = new_n15123_ | ~new_n15126_;
  assign ys__n3040 = ~ys__n740 | ys__n3039;
  assign ys__n3051 = new_n13421_ & new_n13514_;
  assign ys__n3061 = new_n13421_ & new_n13535_;
  assign ys__n3068 = new_n12861_ | new_n12865_;
  assign ys__n3083 = new_n13421_ & new_n13557_;
  assign new_n15133_ = ~ys__n164 & ~ys__n354;
  assign new_n15134_ = ~ys__n4826 & new_n15133_;
  assign new_n15135_ = new_n15074_ & new_n15134_;
  assign new_n15136_ = ~ys__n402 & new_n15135_;
  assign new_n15137_ = ys__n402 & ~ys__n408;
  assign new_n15138_ = ~ys__n404 & new_n15137_;
  assign ys__n3085 = new_n15136_ | ~new_n15138_;
  assign new_n15140_ = new_n13376_ & new_n13507_;
  assign ys__n3097 = new_n13530_ & new_n15140_;
  assign ys__n3106 = new_n13421_ & new_n13520_;
  assign ys__n3114 = new_n13421_ & new_n13494_;
  assign ys__n3115 = new_n13421_ & new_n13554_;
  assign ys__n3121 = new_n13421_ & new_n13505_;
  assign new_n15146_ = ~ys__n46 & ~ys__n340;
  assign new_n15147_ = new_n13400_ & new_n15146_;
  assign new_n15148_ = new_n13399_ & new_n15147_;
  assign new_n15149_ = ~ys__n44 & ~ys__n6115;
  assign new_n15150_ = new_n13380_ & new_n15149_;
  assign new_n15151_ = ~ys__n6112 & ~ys__n6113;
  assign new_n15152_ = ys__n18317 & new_n13375_;
  assign new_n15153_ = new_n15151_ & new_n15152_;
  assign new_n15154_ = new_n15150_ & new_n15153_;
  assign new_n15155_ = new_n15148_ & new_n15154_;
  assign new_n15156_ = new_n13419_ & new_n15155_;
  assign ys__n3195 = ~ys__n874 | new_n15156_;
  assign new_n15158_ = ~ys__n18821 & ~ys__n38090;
  assign new_n15159_ = ys__n18821 & ys__n38090;
  assign new_n15160_ = ~new_n15158_ & ~new_n15159_;
  assign new_n15161_ = ~ys__n18823 & ~ys__n38091;
  assign new_n15162_ = ys__n18823 & ys__n38091;
  assign new_n15163_ = ~new_n15161_ & ~new_n15162_;
  assign new_n15164_ = ~new_n15160_ & ~new_n15163_;
  assign new_n15165_ = ~ys__n18825 & ~ys__n38092;
  assign new_n15166_ = ys__n18825 & ys__n38092;
  assign new_n15167_ = ~new_n15165_ & ~new_n15166_;
  assign new_n15168_ = ~ys__n18827 & ~ys__n38093;
  assign new_n15169_ = ys__n18827 & ys__n38093;
  assign new_n15170_ = ~new_n15168_ & ~new_n15169_;
  assign new_n15171_ = ~new_n15167_ & ~new_n15170_;
  assign new_n15172_ = new_n15164_ & new_n15171_;
  assign new_n15173_ = ~ys__n18813 & ~ys__n38086;
  assign new_n15174_ = ys__n18813 & ys__n38086;
  assign new_n15175_ = ~new_n15173_ & ~new_n15174_;
  assign new_n15176_ = ~ys__n18815 & ~ys__n38087;
  assign new_n15177_ = ys__n18815 & ys__n38087;
  assign new_n15178_ = ~new_n15176_ & ~new_n15177_;
  assign new_n15179_ = ~new_n15175_ & ~new_n15178_;
  assign new_n15180_ = ~ys__n18817 & ~ys__n38088;
  assign new_n15181_ = ys__n18817 & ys__n38088;
  assign new_n15182_ = ~new_n15180_ & ~new_n15181_;
  assign new_n15183_ = ~ys__n18819 & ~ys__n38089;
  assign new_n15184_ = ys__n18819 & ys__n38089;
  assign new_n15185_ = ~new_n15183_ & ~new_n15184_;
  assign new_n15186_ = ~new_n15182_ & ~new_n15185_;
  assign new_n15187_ = new_n15179_ & new_n15186_;
  assign new_n15188_ = ~ys__n18805 & ~ys__n38082;
  assign new_n15189_ = ys__n18805 & ys__n38082;
  assign new_n15190_ = ~new_n15188_ & ~new_n15189_;
  assign new_n15191_ = ~ys__n18807 & ~ys__n38083;
  assign new_n15192_ = ys__n18807 & ys__n38083;
  assign new_n15193_ = ~new_n15191_ & ~new_n15192_;
  assign new_n15194_ = ~new_n15190_ & ~new_n15193_;
  assign new_n15195_ = ~ys__n18809 & ~ys__n38084;
  assign new_n15196_ = ys__n18809 & ys__n38084;
  assign new_n15197_ = ~new_n15195_ & ~new_n15196_;
  assign new_n15198_ = ~ys__n18811 & ~ys__n38085;
  assign new_n15199_ = ys__n18811 & ys__n38085;
  assign new_n15200_ = ~new_n15198_ & ~new_n15199_;
  assign new_n15201_ = ~new_n15197_ & ~new_n15200_;
  assign new_n15202_ = new_n15194_ & new_n15201_;
  assign new_n15203_ = new_n15187_ & new_n15202_;
  assign new_n15204_ = new_n15172_ & new_n15203_;
  assign new_n15205_ = ~ys__n18781 & ~ys__n38070;
  assign new_n15206_ = ys__n18781 & ys__n38070;
  assign new_n15207_ = ~new_n15205_ & ~new_n15206_;
  assign new_n15208_ = ~ys__n18783 & ~ys__n38071;
  assign new_n15209_ = ys__n18783 & ys__n38071;
  assign new_n15210_ = ~new_n15208_ & ~new_n15209_;
  assign new_n15211_ = ~new_n15207_ & ~new_n15210_;
  assign new_n15212_ = ~ys__n18785 & ~ys__n38072;
  assign new_n15213_ = ys__n18785 & ys__n38072;
  assign new_n15214_ = ~new_n15212_ & ~new_n15213_;
  assign new_n15215_ = ~ys__n18787 & ~ys__n38073;
  assign new_n15216_ = ys__n18787 & ys__n38073;
  assign new_n15217_ = ~new_n15215_ & ~new_n15216_;
  assign new_n15218_ = ~new_n15214_ & ~new_n15217_;
  assign new_n15219_ = new_n15211_ & new_n15218_;
  assign new_n15220_ = ~ys__n18773 & ~ys__n38066;
  assign new_n15221_ = ys__n18773 & ys__n38066;
  assign new_n15222_ = ~new_n15220_ & ~new_n15221_;
  assign new_n15223_ = ~ys__n18775 & ~ys__n38067;
  assign new_n15224_ = ys__n18775 & ys__n38067;
  assign new_n15225_ = ~new_n15223_ & ~new_n15224_;
  assign new_n15226_ = ~new_n15222_ & ~new_n15225_;
  assign new_n15227_ = ~ys__n18777 & ~ys__n38068;
  assign new_n15228_ = ys__n18777 & ys__n38068;
  assign new_n15229_ = ~new_n15227_ & ~new_n15228_;
  assign new_n15230_ = ~ys__n18779 & ~ys__n38069;
  assign new_n15231_ = ys__n18779 & ys__n38069;
  assign new_n15232_ = ~new_n15230_ & ~new_n15231_;
  assign new_n15233_ = ~new_n15229_ & ~new_n15232_;
  assign new_n15234_ = new_n15226_ & new_n15233_;
  assign new_n15235_ = new_n15219_ & new_n15234_;
  assign new_n15236_ = ~ys__n18797 & ~ys__n38078;
  assign new_n15237_ = ys__n18797 & ys__n38078;
  assign new_n15238_ = ~new_n15236_ & ~new_n15237_;
  assign new_n15239_ = ~ys__n18799 & ~ys__n38079;
  assign new_n15240_ = ys__n18799 & ys__n38079;
  assign new_n15241_ = ~new_n15239_ & ~new_n15240_;
  assign new_n15242_ = ~new_n15238_ & ~new_n15241_;
  assign new_n15243_ = ~ys__n18801 & ~ys__n38080;
  assign new_n15244_ = ys__n18801 & ys__n38080;
  assign new_n15245_ = ~new_n15243_ & ~new_n15244_;
  assign new_n15246_ = ~ys__n18803 & ~ys__n38081;
  assign new_n15247_ = ys__n18803 & ys__n38081;
  assign new_n15248_ = ~new_n15246_ & ~new_n15247_;
  assign new_n15249_ = ~new_n15245_ & ~new_n15248_;
  assign new_n15250_ = new_n15242_ & new_n15249_;
  assign new_n15251_ = ~ys__n18789 & ~ys__n38074;
  assign new_n15252_ = ys__n18789 & ys__n38074;
  assign new_n15253_ = ~new_n15251_ & ~new_n15252_;
  assign new_n15254_ = ~ys__n18791 & ~ys__n38075;
  assign new_n15255_ = ys__n18791 & ys__n38075;
  assign new_n15256_ = ~new_n15254_ & ~new_n15255_;
  assign new_n15257_ = ~new_n15253_ & ~new_n15256_;
  assign new_n15258_ = ~ys__n18793 & ~ys__n38076;
  assign new_n15259_ = ys__n18793 & ys__n38076;
  assign new_n15260_ = ~new_n15258_ & ~new_n15259_;
  assign new_n15261_ = ~ys__n18795 & ~ys__n38077;
  assign new_n15262_ = ys__n18795 & ys__n38077;
  assign new_n15263_ = ~new_n15261_ & ~new_n15262_;
  assign new_n15264_ = ~new_n15260_ & ~new_n15263_;
  assign new_n15265_ = new_n15257_ & new_n15264_;
  assign new_n15266_ = new_n15250_ & new_n15265_;
  assign new_n15267_ = new_n15235_ & new_n15266_;
  assign new_n15268_ = new_n15204_ & new_n15267_;
  assign new_n15269_ = ~ys__n37746 & ~new_n15268_;
  assign new_n15270_ = ys__n836 & ~new_n15269_;
  assign new_n15271_ = ~ys__n18821 & ~ys__n38062;
  assign new_n15272_ = ys__n18821 & ys__n38062;
  assign new_n15273_ = ~new_n15271_ & ~new_n15272_;
  assign new_n15274_ = ~ys__n18823 & ~ys__n38063;
  assign new_n15275_ = ys__n18823 & ys__n38063;
  assign new_n15276_ = ~new_n15274_ & ~new_n15275_;
  assign new_n15277_ = ~new_n15273_ & ~new_n15276_;
  assign new_n15278_ = ~ys__n18825 & ~ys__n38064;
  assign new_n15279_ = ys__n18825 & ys__n38064;
  assign new_n15280_ = ~new_n15278_ & ~new_n15279_;
  assign new_n15281_ = ~ys__n18827 & ~ys__n38065;
  assign new_n15282_ = ys__n18827 & ys__n38065;
  assign new_n15283_ = ~new_n15281_ & ~new_n15282_;
  assign new_n15284_ = ~new_n15280_ & ~new_n15283_;
  assign new_n15285_ = new_n15277_ & new_n15284_;
  assign new_n15286_ = ~ys__n18813 & ~ys__n38058;
  assign new_n15287_ = ys__n18813 & ys__n38058;
  assign new_n15288_ = ~new_n15286_ & ~new_n15287_;
  assign new_n15289_ = ~ys__n18815 & ~ys__n38059;
  assign new_n15290_ = ys__n18815 & ys__n38059;
  assign new_n15291_ = ~new_n15289_ & ~new_n15290_;
  assign new_n15292_ = ~new_n15288_ & ~new_n15291_;
  assign new_n15293_ = ~ys__n18817 & ~ys__n38060;
  assign new_n15294_ = ys__n18817 & ys__n38060;
  assign new_n15295_ = ~new_n15293_ & ~new_n15294_;
  assign new_n15296_ = ~ys__n18819 & ~ys__n38061;
  assign new_n15297_ = ys__n18819 & ys__n38061;
  assign new_n15298_ = ~new_n15296_ & ~new_n15297_;
  assign new_n15299_ = ~new_n15295_ & ~new_n15298_;
  assign new_n15300_ = new_n15292_ & new_n15299_;
  assign new_n15301_ = ~ys__n18805 & ~ys__n38054;
  assign new_n15302_ = ys__n18805 & ys__n38054;
  assign new_n15303_ = ~new_n15301_ & ~new_n15302_;
  assign new_n15304_ = ~ys__n18807 & ~ys__n38055;
  assign new_n15305_ = ys__n18807 & ys__n38055;
  assign new_n15306_ = ~new_n15304_ & ~new_n15305_;
  assign new_n15307_ = ~new_n15303_ & ~new_n15306_;
  assign new_n15308_ = ~ys__n18809 & ~ys__n38056;
  assign new_n15309_ = ys__n18809 & ys__n38056;
  assign new_n15310_ = ~new_n15308_ & ~new_n15309_;
  assign new_n15311_ = ~ys__n18811 & ~ys__n38057;
  assign new_n15312_ = ys__n18811 & ys__n38057;
  assign new_n15313_ = ~new_n15311_ & ~new_n15312_;
  assign new_n15314_ = ~new_n15310_ & ~new_n15313_;
  assign new_n15315_ = new_n15307_ & new_n15314_;
  assign new_n15316_ = new_n15300_ & new_n15315_;
  assign new_n15317_ = new_n15285_ & new_n15316_;
  assign new_n15318_ = ~ys__n18781 & ~ys__n38042;
  assign new_n15319_ = ys__n18781 & ys__n38042;
  assign new_n15320_ = ~new_n15318_ & ~new_n15319_;
  assign new_n15321_ = ~ys__n18783 & ~ys__n38043;
  assign new_n15322_ = ys__n18783 & ys__n38043;
  assign new_n15323_ = ~new_n15321_ & ~new_n15322_;
  assign new_n15324_ = ~new_n15320_ & ~new_n15323_;
  assign new_n15325_ = ~ys__n18785 & ~ys__n38044;
  assign new_n15326_ = ys__n18785 & ys__n38044;
  assign new_n15327_ = ~new_n15325_ & ~new_n15326_;
  assign new_n15328_ = ~ys__n18787 & ~ys__n38045;
  assign new_n15329_ = ys__n18787 & ys__n38045;
  assign new_n15330_ = ~new_n15328_ & ~new_n15329_;
  assign new_n15331_ = ~new_n15327_ & ~new_n15330_;
  assign new_n15332_ = new_n15324_ & new_n15331_;
  assign new_n15333_ = ~ys__n18773 & ~ys__n38038;
  assign new_n15334_ = ys__n18773 & ys__n38038;
  assign new_n15335_ = ~new_n15333_ & ~new_n15334_;
  assign new_n15336_ = ~ys__n18775 & ~ys__n38039;
  assign new_n15337_ = ys__n18775 & ys__n38039;
  assign new_n15338_ = ~new_n15336_ & ~new_n15337_;
  assign new_n15339_ = ~new_n15335_ & ~new_n15338_;
  assign new_n15340_ = ~ys__n18777 & ~ys__n38040;
  assign new_n15341_ = ys__n18777 & ys__n38040;
  assign new_n15342_ = ~new_n15340_ & ~new_n15341_;
  assign new_n15343_ = ~ys__n18779 & ~ys__n38041;
  assign new_n15344_ = ys__n18779 & ys__n38041;
  assign new_n15345_ = ~new_n15343_ & ~new_n15344_;
  assign new_n15346_ = ~new_n15342_ & ~new_n15345_;
  assign new_n15347_ = new_n15339_ & new_n15346_;
  assign new_n15348_ = new_n15332_ & new_n15347_;
  assign new_n15349_ = ~ys__n18797 & ~ys__n38050;
  assign new_n15350_ = ys__n18797 & ys__n38050;
  assign new_n15351_ = ~new_n15349_ & ~new_n15350_;
  assign new_n15352_ = ~ys__n18799 & ~ys__n38051;
  assign new_n15353_ = ys__n18799 & ys__n38051;
  assign new_n15354_ = ~new_n15352_ & ~new_n15353_;
  assign new_n15355_ = ~new_n15351_ & ~new_n15354_;
  assign new_n15356_ = ~ys__n18801 & ~ys__n38052;
  assign new_n15357_ = ys__n18801 & ys__n38052;
  assign new_n15358_ = ~new_n15356_ & ~new_n15357_;
  assign new_n15359_ = ~ys__n18803 & ~ys__n38053;
  assign new_n15360_ = ys__n18803 & ys__n38053;
  assign new_n15361_ = ~new_n15359_ & ~new_n15360_;
  assign new_n15362_ = ~new_n15358_ & ~new_n15361_;
  assign new_n15363_ = new_n15355_ & new_n15362_;
  assign new_n15364_ = ~ys__n18789 & ~ys__n38046;
  assign new_n15365_ = ys__n18789 & ys__n38046;
  assign new_n15366_ = ~new_n15364_ & ~new_n15365_;
  assign new_n15367_ = ~ys__n18791 & ~ys__n38047;
  assign new_n15368_ = ys__n18791 & ys__n38047;
  assign new_n15369_ = ~new_n15367_ & ~new_n15368_;
  assign new_n15370_ = ~new_n15366_ & ~new_n15369_;
  assign new_n15371_ = ~ys__n18793 & ~ys__n38048;
  assign new_n15372_ = ys__n18793 & ys__n38048;
  assign new_n15373_ = ~new_n15371_ & ~new_n15372_;
  assign new_n15374_ = ~ys__n18795 & ~ys__n38049;
  assign new_n15375_ = ys__n18795 & ys__n38049;
  assign new_n15376_ = ~new_n15374_ & ~new_n15375_;
  assign new_n15377_ = ~new_n15373_ & ~new_n15376_;
  assign new_n15378_ = new_n15370_ & new_n15377_;
  assign new_n15379_ = new_n15363_ & new_n15378_;
  assign new_n15380_ = new_n15348_ & new_n15379_;
  assign new_n15381_ = new_n15317_ & new_n15380_;
  assign new_n15382_ = ~ys__n37747 & ~new_n15381_;
  assign new_n15383_ = ys__n834 & ~new_n15382_;
  assign new_n15384_ = ~new_n15270_ & ~new_n15383_;
  assign new_n15385_ = ~ys__n18821 & ~ys__n38034;
  assign new_n15386_ = ys__n18821 & ys__n38034;
  assign new_n15387_ = ~new_n15385_ & ~new_n15386_;
  assign new_n15388_ = ~ys__n18823 & ~ys__n38035;
  assign new_n15389_ = ys__n18823 & ys__n38035;
  assign new_n15390_ = ~new_n15388_ & ~new_n15389_;
  assign new_n15391_ = ~new_n15387_ & ~new_n15390_;
  assign new_n15392_ = ~ys__n18825 & ~ys__n38036;
  assign new_n15393_ = ys__n18825 & ys__n38036;
  assign new_n15394_ = ~new_n15392_ & ~new_n15393_;
  assign new_n15395_ = ~ys__n18827 & ~ys__n38037;
  assign new_n15396_ = ys__n18827 & ys__n38037;
  assign new_n15397_ = ~new_n15395_ & ~new_n15396_;
  assign new_n15398_ = ~new_n15394_ & ~new_n15397_;
  assign new_n15399_ = new_n15391_ & new_n15398_;
  assign new_n15400_ = ~ys__n18813 & ~ys__n38030;
  assign new_n15401_ = ys__n18813 & ys__n38030;
  assign new_n15402_ = ~new_n15400_ & ~new_n15401_;
  assign new_n15403_ = ~ys__n18815 & ~ys__n38031;
  assign new_n15404_ = ys__n18815 & ys__n38031;
  assign new_n15405_ = ~new_n15403_ & ~new_n15404_;
  assign new_n15406_ = ~new_n15402_ & ~new_n15405_;
  assign new_n15407_ = ~ys__n18817 & ~ys__n38032;
  assign new_n15408_ = ys__n18817 & ys__n38032;
  assign new_n15409_ = ~new_n15407_ & ~new_n15408_;
  assign new_n15410_ = ~ys__n18819 & ~ys__n38033;
  assign new_n15411_ = ys__n18819 & ys__n38033;
  assign new_n15412_ = ~new_n15410_ & ~new_n15411_;
  assign new_n15413_ = ~new_n15409_ & ~new_n15412_;
  assign new_n15414_ = new_n15406_ & new_n15413_;
  assign new_n15415_ = ~ys__n18805 & ~ys__n38026;
  assign new_n15416_ = ys__n18805 & ys__n38026;
  assign new_n15417_ = ~new_n15415_ & ~new_n15416_;
  assign new_n15418_ = ~ys__n18807 & ~ys__n38027;
  assign new_n15419_ = ys__n18807 & ys__n38027;
  assign new_n15420_ = ~new_n15418_ & ~new_n15419_;
  assign new_n15421_ = ~new_n15417_ & ~new_n15420_;
  assign new_n15422_ = ~ys__n18809 & ~ys__n38028;
  assign new_n15423_ = ys__n18809 & ys__n38028;
  assign new_n15424_ = ~new_n15422_ & ~new_n15423_;
  assign new_n15425_ = ~ys__n18811 & ~ys__n38029;
  assign new_n15426_ = ys__n18811 & ys__n38029;
  assign new_n15427_ = ~new_n15425_ & ~new_n15426_;
  assign new_n15428_ = ~new_n15424_ & ~new_n15427_;
  assign new_n15429_ = new_n15421_ & new_n15428_;
  assign new_n15430_ = new_n15414_ & new_n15429_;
  assign new_n15431_ = new_n15399_ & new_n15430_;
  assign new_n15432_ = ~ys__n18781 & ~ys__n38014;
  assign new_n15433_ = ys__n18781 & ys__n38014;
  assign new_n15434_ = ~new_n15432_ & ~new_n15433_;
  assign new_n15435_ = ~ys__n18783 & ~ys__n38015;
  assign new_n15436_ = ys__n18783 & ys__n38015;
  assign new_n15437_ = ~new_n15435_ & ~new_n15436_;
  assign new_n15438_ = ~new_n15434_ & ~new_n15437_;
  assign new_n15439_ = ~ys__n18785 & ~ys__n38016;
  assign new_n15440_ = ys__n18785 & ys__n38016;
  assign new_n15441_ = ~new_n15439_ & ~new_n15440_;
  assign new_n15442_ = ~ys__n18787 & ~ys__n38017;
  assign new_n15443_ = ys__n18787 & ys__n38017;
  assign new_n15444_ = ~new_n15442_ & ~new_n15443_;
  assign new_n15445_ = ~new_n15441_ & ~new_n15444_;
  assign new_n15446_ = new_n15438_ & new_n15445_;
  assign new_n15447_ = ~ys__n18773 & ~ys__n38010;
  assign new_n15448_ = ys__n18773 & ys__n38010;
  assign new_n15449_ = ~new_n15447_ & ~new_n15448_;
  assign new_n15450_ = ~ys__n18775 & ~ys__n38011;
  assign new_n15451_ = ys__n18775 & ys__n38011;
  assign new_n15452_ = ~new_n15450_ & ~new_n15451_;
  assign new_n15453_ = ~new_n15449_ & ~new_n15452_;
  assign new_n15454_ = ~ys__n18777 & ~ys__n38012;
  assign new_n15455_ = ys__n18777 & ys__n38012;
  assign new_n15456_ = ~new_n15454_ & ~new_n15455_;
  assign new_n15457_ = ~ys__n18779 & ~ys__n38013;
  assign new_n15458_ = ys__n18779 & ys__n38013;
  assign new_n15459_ = ~new_n15457_ & ~new_n15458_;
  assign new_n15460_ = ~new_n15456_ & ~new_n15459_;
  assign new_n15461_ = new_n15453_ & new_n15460_;
  assign new_n15462_ = new_n15446_ & new_n15461_;
  assign new_n15463_ = ~ys__n18797 & ~ys__n38022;
  assign new_n15464_ = ys__n18797 & ys__n38022;
  assign new_n15465_ = ~new_n15463_ & ~new_n15464_;
  assign new_n15466_ = ~ys__n18799 & ~ys__n38023;
  assign new_n15467_ = ys__n18799 & ys__n38023;
  assign new_n15468_ = ~new_n15466_ & ~new_n15467_;
  assign new_n15469_ = ~new_n15465_ & ~new_n15468_;
  assign new_n15470_ = ~ys__n18801 & ~ys__n38024;
  assign new_n15471_ = ys__n18801 & ys__n38024;
  assign new_n15472_ = ~new_n15470_ & ~new_n15471_;
  assign new_n15473_ = ~ys__n18803 & ~ys__n38025;
  assign new_n15474_ = ys__n18803 & ys__n38025;
  assign new_n15475_ = ~new_n15473_ & ~new_n15474_;
  assign new_n15476_ = ~new_n15472_ & ~new_n15475_;
  assign new_n15477_ = new_n15469_ & new_n15476_;
  assign new_n15478_ = ~ys__n18789 & ~ys__n38018;
  assign new_n15479_ = ys__n18789 & ys__n38018;
  assign new_n15480_ = ~new_n15478_ & ~new_n15479_;
  assign new_n15481_ = ~ys__n18791 & ~ys__n38019;
  assign new_n15482_ = ys__n18791 & ys__n38019;
  assign new_n15483_ = ~new_n15481_ & ~new_n15482_;
  assign new_n15484_ = ~new_n15480_ & ~new_n15483_;
  assign new_n15485_ = ~ys__n18793 & ~ys__n38020;
  assign new_n15486_ = ys__n18793 & ys__n38020;
  assign new_n15487_ = ~new_n15485_ & ~new_n15486_;
  assign new_n15488_ = ~ys__n18795 & ~ys__n38021;
  assign new_n15489_ = ys__n18795 & ys__n38021;
  assign new_n15490_ = ~new_n15488_ & ~new_n15489_;
  assign new_n15491_ = ~new_n15487_ & ~new_n15490_;
  assign new_n15492_ = new_n15484_ & new_n15491_;
  assign new_n15493_ = new_n15477_ & new_n15492_;
  assign new_n15494_ = new_n15462_ & new_n15493_;
  assign new_n15495_ = new_n15431_ & new_n15494_;
  assign new_n15496_ = ~ys__n37748 & ~new_n15495_;
  assign new_n15497_ = ys__n832 & ~new_n15496_;
  assign new_n15498_ = ~ys__n18821 & ~ys__n38006;
  assign new_n15499_ = ys__n18821 & ys__n38006;
  assign new_n15500_ = ~new_n15498_ & ~new_n15499_;
  assign new_n15501_ = ~ys__n18823 & ~ys__n38007;
  assign new_n15502_ = ys__n18823 & ys__n38007;
  assign new_n15503_ = ~new_n15501_ & ~new_n15502_;
  assign new_n15504_ = ~new_n15500_ & ~new_n15503_;
  assign new_n15505_ = ~ys__n18825 & ~ys__n38008;
  assign new_n15506_ = ys__n18825 & ys__n38008;
  assign new_n15507_ = ~new_n15505_ & ~new_n15506_;
  assign new_n15508_ = ~ys__n18827 & ~ys__n38009;
  assign new_n15509_ = ys__n18827 & ys__n38009;
  assign new_n15510_ = ~new_n15508_ & ~new_n15509_;
  assign new_n15511_ = ~new_n15507_ & ~new_n15510_;
  assign new_n15512_ = new_n15504_ & new_n15511_;
  assign new_n15513_ = ~ys__n18813 & ~ys__n38002;
  assign new_n15514_ = ys__n18813 & ys__n38002;
  assign new_n15515_ = ~new_n15513_ & ~new_n15514_;
  assign new_n15516_ = ~ys__n18815 & ~ys__n38003;
  assign new_n15517_ = ys__n18815 & ys__n38003;
  assign new_n15518_ = ~new_n15516_ & ~new_n15517_;
  assign new_n15519_ = ~new_n15515_ & ~new_n15518_;
  assign new_n15520_ = ~ys__n18817 & ~ys__n38004;
  assign new_n15521_ = ys__n18817 & ys__n38004;
  assign new_n15522_ = ~new_n15520_ & ~new_n15521_;
  assign new_n15523_ = ~ys__n18819 & ~ys__n38005;
  assign new_n15524_ = ys__n18819 & ys__n38005;
  assign new_n15525_ = ~new_n15523_ & ~new_n15524_;
  assign new_n15526_ = ~new_n15522_ & ~new_n15525_;
  assign new_n15527_ = new_n15519_ & new_n15526_;
  assign new_n15528_ = ~ys__n18805 & ~ys__n37998;
  assign new_n15529_ = ys__n18805 & ys__n37998;
  assign new_n15530_ = ~new_n15528_ & ~new_n15529_;
  assign new_n15531_ = ~ys__n18807 & ~ys__n37999;
  assign new_n15532_ = ys__n18807 & ys__n37999;
  assign new_n15533_ = ~new_n15531_ & ~new_n15532_;
  assign new_n15534_ = ~new_n15530_ & ~new_n15533_;
  assign new_n15535_ = ~ys__n18809 & ~ys__n38000;
  assign new_n15536_ = ys__n18809 & ys__n38000;
  assign new_n15537_ = ~new_n15535_ & ~new_n15536_;
  assign new_n15538_ = ~ys__n18811 & ~ys__n38001;
  assign new_n15539_ = ys__n18811 & ys__n38001;
  assign new_n15540_ = ~new_n15538_ & ~new_n15539_;
  assign new_n15541_ = ~new_n15537_ & ~new_n15540_;
  assign new_n15542_ = new_n15534_ & new_n15541_;
  assign new_n15543_ = new_n15527_ & new_n15542_;
  assign new_n15544_ = new_n15512_ & new_n15543_;
  assign new_n15545_ = ~ys__n18781 & ~ys__n37986;
  assign new_n15546_ = ys__n18781 & ys__n37986;
  assign new_n15547_ = ~new_n15545_ & ~new_n15546_;
  assign new_n15548_ = ~ys__n18783 & ~ys__n37987;
  assign new_n15549_ = ys__n18783 & ys__n37987;
  assign new_n15550_ = ~new_n15548_ & ~new_n15549_;
  assign new_n15551_ = ~new_n15547_ & ~new_n15550_;
  assign new_n15552_ = ~ys__n18785 & ~ys__n37988;
  assign new_n15553_ = ys__n18785 & ys__n37988;
  assign new_n15554_ = ~new_n15552_ & ~new_n15553_;
  assign new_n15555_ = ~ys__n18787 & ~ys__n37989;
  assign new_n15556_ = ys__n18787 & ys__n37989;
  assign new_n15557_ = ~new_n15555_ & ~new_n15556_;
  assign new_n15558_ = ~new_n15554_ & ~new_n15557_;
  assign new_n15559_ = new_n15551_ & new_n15558_;
  assign new_n15560_ = ~ys__n18773 & ~ys__n37982;
  assign new_n15561_ = ys__n18773 & ys__n37982;
  assign new_n15562_ = ~new_n15560_ & ~new_n15561_;
  assign new_n15563_ = ~ys__n18775 & ~ys__n37983;
  assign new_n15564_ = ys__n18775 & ys__n37983;
  assign new_n15565_ = ~new_n15563_ & ~new_n15564_;
  assign new_n15566_ = ~new_n15562_ & ~new_n15565_;
  assign new_n15567_ = ~ys__n18777 & ~ys__n37984;
  assign new_n15568_ = ys__n18777 & ys__n37984;
  assign new_n15569_ = ~new_n15567_ & ~new_n15568_;
  assign new_n15570_ = ~ys__n18779 & ~ys__n37985;
  assign new_n15571_ = ys__n18779 & ys__n37985;
  assign new_n15572_ = ~new_n15570_ & ~new_n15571_;
  assign new_n15573_ = ~new_n15569_ & ~new_n15572_;
  assign new_n15574_ = new_n15566_ & new_n15573_;
  assign new_n15575_ = new_n15559_ & new_n15574_;
  assign new_n15576_ = ~ys__n18797 & ~ys__n37994;
  assign new_n15577_ = ys__n18797 & ys__n37994;
  assign new_n15578_ = ~new_n15576_ & ~new_n15577_;
  assign new_n15579_ = ~ys__n18799 & ~ys__n37995;
  assign new_n15580_ = ys__n18799 & ys__n37995;
  assign new_n15581_ = ~new_n15579_ & ~new_n15580_;
  assign new_n15582_ = ~new_n15578_ & ~new_n15581_;
  assign new_n15583_ = ~ys__n18801 & ~ys__n37996;
  assign new_n15584_ = ys__n18801 & ys__n37996;
  assign new_n15585_ = ~new_n15583_ & ~new_n15584_;
  assign new_n15586_ = ~ys__n18803 & ~ys__n37997;
  assign new_n15587_ = ys__n18803 & ys__n37997;
  assign new_n15588_ = ~new_n15586_ & ~new_n15587_;
  assign new_n15589_ = ~new_n15585_ & ~new_n15588_;
  assign new_n15590_ = new_n15582_ & new_n15589_;
  assign new_n15591_ = ~ys__n18789 & ~ys__n37990;
  assign new_n15592_ = ys__n18789 & ys__n37990;
  assign new_n15593_ = ~new_n15591_ & ~new_n15592_;
  assign new_n15594_ = ~ys__n18791 & ~ys__n37991;
  assign new_n15595_ = ys__n18791 & ys__n37991;
  assign new_n15596_ = ~new_n15594_ & ~new_n15595_;
  assign new_n15597_ = ~new_n15593_ & ~new_n15596_;
  assign new_n15598_ = ~ys__n18793 & ~ys__n37992;
  assign new_n15599_ = ys__n18793 & ys__n37992;
  assign new_n15600_ = ~new_n15598_ & ~new_n15599_;
  assign new_n15601_ = ~ys__n18795 & ~ys__n37993;
  assign new_n15602_ = ys__n18795 & ys__n37993;
  assign new_n15603_ = ~new_n15601_ & ~new_n15602_;
  assign new_n15604_ = ~new_n15600_ & ~new_n15603_;
  assign new_n15605_ = new_n15597_ & new_n15604_;
  assign new_n15606_ = new_n15590_ & new_n15605_;
  assign new_n15607_ = new_n15575_ & new_n15606_;
  assign new_n15608_ = new_n15544_ & new_n15607_;
  assign new_n15609_ = ~ys__n37749 & ~new_n15608_;
  assign new_n15610_ = ys__n830 & ~new_n15609_;
  assign new_n15611_ = ~new_n15497_ & ~new_n15610_;
  assign new_n15612_ = new_n15384_ & new_n15611_;
  assign new_n15613_ = ~ys__n18821 & ~ys__n18984;
  assign new_n15614_ = ys__n18821 & ys__n18984;
  assign new_n15615_ = ~new_n15613_ & ~new_n15614_;
  assign new_n15616_ = ~ys__n18823 & ~ys__n18985;
  assign new_n15617_ = ys__n18823 & ys__n18985;
  assign new_n15618_ = ~new_n15616_ & ~new_n15617_;
  assign new_n15619_ = ~new_n15615_ & ~new_n15618_;
  assign new_n15620_ = ~ys__n18825 & ~ys__n18986;
  assign new_n15621_ = ys__n18825 & ys__n18986;
  assign new_n15622_ = ~new_n15620_ & ~new_n15621_;
  assign new_n15623_ = ~ys__n18827 & ~ys__n18987;
  assign new_n15624_ = ys__n18827 & ys__n18987;
  assign new_n15625_ = ~new_n15623_ & ~new_n15624_;
  assign new_n15626_ = ~new_n15622_ & ~new_n15625_;
  assign new_n15627_ = new_n15619_ & new_n15626_;
  assign new_n15628_ = ~ys__n18813 & ~ys__n18980;
  assign new_n15629_ = ys__n18813 & ys__n18980;
  assign new_n15630_ = ~new_n15628_ & ~new_n15629_;
  assign new_n15631_ = ~ys__n18815 & ~ys__n18981;
  assign new_n15632_ = ys__n18815 & ys__n18981;
  assign new_n15633_ = ~new_n15631_ & ~new_n15632_;
  assign new_n15634_ = ~new_n15630_ & ~new_n15633_;
  assign new_n15635_ = ~ys__n18817 & ~ys__n18982;
  assign new_n15636_ = ys__n18817 & ys__n18982;
  assign new_n15637_ = ~new_n15635_ & ~new_n15636_;
  assign new_n15638_ = ~ys__n18819 & ~ys__n18983;
  assign new_n15639_ = ys__n18819 & ys__n18983;
  assign new_n15640_ = ~new_n15638_ & ~new_n15639_;
  assign new_n15641_ = ~new_n15637_ & ~new_n15640_;
  assign new_n15642_ = new_n15634_ & new_n15641_;
  assign new_n15643_ = ~ys__n18805 & ~ys__n18976;
  assign new_n15644_ = ys__n18805 & ys__n18976;
  assign new_n15645_ = ~new_n15643_ & ~new_n15644_;
  assign new_n15646_ = ~ys__n18807 & ~ys__n18977;
  assign new_n15647_ = ys__n18807 & ys__n18977;
  assign new_n15648_ = ~new_n15646_ & ~new_n15647_;
  assign new_n15649_ = ~new_n15645_ & ~new_n15648_;
  assign new_n15650_ = ~ys__n18809 & ~ys__n18978;
  assign new_n15651_ = ys__n18809 & ys__n18978;
  assign new_n15652_ = ~new_n15650_ & ~new_n15651_;
  assign new_n15653_ = ~ys__n18811 & ~ys__n18979;
  assign new_n15654_ = ys__n18811 & ys__n18979;
  assign new_n15655_ = ~new_n15653_ & ~new_n15654_;
  assign new_n15656_ = ~new_n15652_ & ~new_n15655_;
  assign new_n15657_ = new_n15649_ & new_n15656_;
  assign new_n15658_ = new_n15642_ & new_n15657_;
  assign new_n15659_ = new_n15627_ & new_n15658_;
  assign new_n15660_ = ~ys__n18781 & ~ys__n18964;
  assign new_n15661_ = ys__n18781 & ys__n18964;
  assign new_n15662_ = ~new_n15660_ & ~new_n15661_;
  assign new_n15663_ = ~ys__n18783 & ~ys__n18965;
  assign new_n15664_ = ys__n18783 & ys__n18965;
  assign new_n15665_ = ~new_n15663_ & ~new_n15664_;
  assign new_n15666_ = ~new_n15662_ & ~new_n15665_;
  assign new_n15667_ = ~ys__n18785 & ~ys__n18966;
  assign new_n15668_ = ys__n18785 & ys__n18966;
  assign new_n15669_ = ~new_n15667_ & ~new_n15668_;
  assign new_n15670_ = ~ys__n18787 & ~ys__n18967;
  assign new_n15671_ = ys__n18787 & ys__n18967;
  assign new_n15672_ = ~new_n15670_ & ~new_n15671_;
  assign new_n15673_ = ~new_n15669_ & ~new_n15672_;
  assign new_n15674_ = new_n15666_ & new_n15673_;
  assign new_n15675_ = ~ys__n18773 & ~ys__n18960;
  assign new_n15676_ = ys__n18773 & ys__n18960;
  assign new_n15677_ = ~new_n15675_ & ~new_n15676_;
  assign new_n15678_ = ~ys__n18775 & ~ys__n18961;
  assign new_n15679_ = ys__n18775 & ys__n18961;
  assign new_n15680_ = ~new_n15678_ & ~new_n15679_;
  assign new_n15681_ = ~new_n15677_ & ~new_n15680_;
  assign new_n15682_ = ~ys__n18777 & ~ys__n18962;
  assign new_n15683_ = ys__n18777 & ys__n18962;
  assign new_n15684_ = ~new_n15682_ & ~new_n15683_;
  assign new_n15685_ = ~ys__n18779 & ~ys__n18963;
  assign new_n15686_ = ys__n18779 & ys__n18963;
  assign new_n15687_ = ~new_n15685_ & ~new_n15686_;
  assign new_n15688_ = ~new_n15684_ & ~new_n15687_;
  assign new_n15689_ = new_n15681_ & new_n15688_;
  assign new_n15690_ = new_n15674_ & new_n15689_;
  assign new_n15691_ = ~ys__n18797 & ~ys__n18972;
  assign new_n15692_ = ys__n18797 & ys__n18972;
  assign new_n15693_ = ~new_n15691_ & ~new_n15692_;
  assign new_n15694_ = ~ys__n18799 & ~ys__n18973;
  assign new_n15695_ = ys__n18799 & ys__n18973;
  assign new_n15696_ = ~new_n15694_ & ~new_n15695_;
  assign new_n15697_ = ~new_n15693_ & ~new_n15696_;
  assign new_n15698_ = ~ys__n18801 & ~ys__n18974;
  assign new_n15699_ = ys__n18801 & ys__n18974;
  assign new_n15700_ = ~new_n15698_ & ~new_n15699_;
  assign new_n15701_ = ~ys__n18803 & ~ys__n18975;
  assign new_n15702_ = ys__n18803 & ys__n18975;
  assign new_n15703_ = ~new_n15701_ & ~new_n15702_;
  assign new_n15704_ = ~new_n15700_ & ~new_n15703_;
  assign new_n15705_ = new_n15697_ & new_n15704_;
  assign new_n15706_ = ~ys__n18789 & ~ys__n18968;
  assign new_n15707_ = ys__n18789 & ys__n18968;
  assign new_n15708_ = ~new_n15706_ & ~new_n15707_;
  assign new_n15709_ = ~ys__n18791 & ~ys__n18969;
  assign new_n15710_ = ys__n18791 & ys__n18969;
  assign new_n15711_ = ~new_n15709_ & ~new_n15710_;
  assign new_n15712_ = ~new_n15708_ & ~new_n15711_;
  assign new_n15713_ = ~ys__n18793 & ~ys__n18970;
  assign new_n15714_ = ys__n18793 & ys__n18970;
  assign new_n15715_ = ~new_n15713_ & ~new_n15714_;
  assign new_n15716_ = ~ys__n18795 & ~ys__n18971;
  assign new_n15717_ = ys__n18795 & ys__n18971;
  assign new_n15718_ = ~new_n15716_ & ~new_n15717_;
  assign new_n15719_ = ~new_n15715_ & ~new_n15718_;
  assign new_n15720_ = new_n15712_ & new_n15719_;
  assign new_n15721_ = new_n15705_ & new_n15720_;
  assign new_n15722_ = new_n15690_ & new_n15721_;
  assign new_n15723_ = new_n15659_ & new_n15722_;
  assign new_n15724_ = ~ys__n19166 & ~new_n15723_;
  assign new_n15725_ = ys__n844 & ~new_n15724_;
  assign new_n15726_ = ~ys__n18821 & ~ys__n38174;
  assign new_n15727_ = ys__n18821 & ys__n38174;
  assign new_n15728_ = ~new_n15726_ & ~new_n15727_;
  assign new_n15729_ = ~ys__n18823 & ~ys__n38175;
  assign new_n15730_ = ys__n18823 & ys__n38175;
  assign new_n15731_ = ~new_n15729_ & ~new_n15730_;
  assign new_n15732_ = ~new_n15728_ & ~new_n15731_;
  assign new_n15733_ = ~ys__n18825 & ~ys__n38176;
  assign new_n15734_ = ys__n18825 & ys__n38176;
  assign new_n15735_ = ~new_n15733_ & ~new_n15734_;
  assign new_n15736_ = ~ys__n18827 & ~ys__n38177;
  assign new_n15737_ = ys__n18827 & ys__n38177;
  assign new_n15738_ = ~new_n15736_ & ~new_n15737_;
  assign new_n15739_ = ~new_n15735_ & ~new_n15738_;
  assign new_n15740_ = new_n15732_ & new_n15739_;
  assign new_n15741_ = ~ys__n18813 & ~ys__n38170;
  assign new_n15742_ = ys__n18813 & ys__n38170;
  assign new_n15743_ = ~new_n15741_ & ~new_n15742_;
  assign new_n15744_ = ~ys__n18815 & ~ys__n38171;
  assign new_n15745_ = ys__n18815 & ys__n38171;
  assign new_n15746_ = ~new_n15744_ & ~new_n15745_;
  assign new_n15747_ = ~new_n15743_ & ~new_n15746_;
  assign new_n15748_ = ~ys__n18817 & ~ys__n38172;
  assign new_n15749_ = ys__n18817 & ys__n38172;
  assign new_n15750_ = ~new_n15748_ & ~new_n15749_;
  assign new_n15751_ = ~ys__n18819 & ~ys__n38173;
  assign new_n15752_ = ys__n18819 & ys__n38173;
  assign new_n15753_ = ~new_n15751_ & ~new_n15752_;
  assign new_n15754_ = ~new_n15750_ & ~new_n15753_;
  assign new_n15755_ = new_n15747_ & new_n15754_;
  assign new_n15756_ = ~ys__n18805 & ~ys__n38166;
  assign new_n15757_ = ys__n18805 & ys__n38166;
  assign new_n15758_ = ~new_n15756_ & ~new_n15757_;
  assign new_n15759_ = ~ys__n18807 & ~ys__n38167;
  assign new_n15760_ = ys__n18807 & ys__n38167;
  assign new_n15761_ = ~new_n15759_ & ~new_n15760_;
  assign new_n15762_ = ~new_n15758_ & ~new_n15761_;
  assign new_n15763_ = ~ys__n18809 & ~ys__n38168;
  assign new_n15764_ = ys__n18809 & ys__n38168;
  assign new_n15765_ = ~new_n15763_ & ~new_n15764_;
  assign new_n15766_ = ~ys__n18811 & ~ys__n38169;
  assign new_n15767_ = ys__n18811 & ys__n38169;
  assign new_n15768_ = ~new_n15766_ & ~new_n15767_;
  assign new_n15769_ = ~new_n15765_ & ~new_n15768_;
  assign new_n15770_ = new_n15762_ & new_n15769_;
  assign new_n15771_ = new_n15755_ & new_n15770_;
  assign new_n15772_ = new_n15740_ & new_n15771_;
  assign new_n15773_ = ~ys__n18781 & ~ys__n38154;
  assign new_n15774_ = ys__n18781 & ys__n38154;
  assign new_n15775_ = ~new_n15773_ & ~new_n15774_;
  assign new_n15776_ = ~ys__n18783 & ~ys__n38155;
  assign new_n15777_ = ys__n18783 & ys__n38155;
  assign new_n15778_ = ~new_n15776_ & ~new_n15777_;
  assign new_n15779_ = ~new_n15775_ & ~new_n15778_;
  assign new_n15780_ = ~ys__n18785 & ~ys__n38156;
  assign new_n15781_ = ys__n18785 & ys__n38156;
  assign new_n15782_ = ~new_n15780_ & ~new_n15781_;
  assign new_n15783_ = ~ys__n18787 & ~ys__n38157;
  assign new_n15784_ = ys__n18787 & ys__n38157;
  assign new_n15785_ = ~new_n15783_ & ~new_n15784_;
  assign new_n15786_ = ~new_n15782_ & ~new_n15785_;
  assign new_n15787_ = new_n15779_ & new_n15786_;
  assign new_n15788_ = ~ys__n18773 & ~ys__n38150;
  assign new_n15789_ = ys__n18773 & ys__n38150;
  assign new_n15790_ = ~new_n15788_ & ~new_n15789_;
  assign new_n15791_ = ~ys__n18775 & ~ys__n38151;
  assign new_n15792_ = ys__n18775 & ys__n38151;
  assign new_n15793_ = ~new_n15791_ & ~new_n15792_;
  assign new_n15794_ = ~new_n15790_ & ~new_n15793_;
  assign new_n15795_ = ~ys__n18777 & ~ys__n38152;
  assign new_n15796_ = ys__n18777 & ys__n38152;
  assign new_n15797_ = ~new_n15795_ & ~new_n15796_;
  assign new_n15798_ = ~ys__n18779 & ~ys__n38153;
  assign new_n15799_ = ys__n18779 & ys__n38153;
  assign new_n15800_ = ~new_n15798_ & ~new_n15799_;
  assign new_n15801_ = ~new_n15797_ & ~new_n15800_;
  assign new_n15802_ = new_n15794_ & new_n15801_;
  assign new_n15803_ = new_n15787_ & new_n15802_;
  assign new_n15804_ = ~ys__n18797 & ~ys__n38162;
  assign new_n15805_ = ys__n18797 & ys__n38162;
  assign new_n15806_ = ~new_n15804_ & ~new_n15805_;
  assign new_n15807_ = ~ys__n18799 & ~ys__n38163;
  assign new_n15808_ = ys__n18799 & ys__n38163;
  assign new_n15809_ = ~new_n15807_ & ~new_n15808_;
  assign new_n15810_ = ~new_n15806_ & ~new_n15809_;
  assign new_n15811_ = ~ys__n18801 & ~ys__n38164;
  assign new_n15812_ = ys__n18801 & ys__n38164;
  assign new_n15813_ = ~new_n15811_ & ~new_n15812_;
  assign new_n15814_ = ~ys__n18803 & ~ys__n38165;
  assign new_n15815_ = ys__n18803 & ys__n38165;
  assign new_n15816_ = ~new_n15814_ & ~new_n15815_;
  assign new_n15817_ = ~new_n15813_ & ~new_n15816_;
  assign new_n15818_ = new_n15810_ & new_n15817_;
  assign new_n15819_ = ~ys__n18789 & ~ys__n38158;
  assign new_n15820_ = ys__n18789 & ys__n38158;
  assign new_n15821_ = ~new_n15819_ & ~new_n15820_;
  assign new_n15822_ = ~ys__n18791 & ~ys__n38159;
  assign new_n15823_ = ys__n18791 & ys__n38159;
  assign new_n15824_ = ~new_n15822_ & ~new_n15823_;
  assign new_n15825_ = ~new_n15821_ & ~new_n15824_;
  assign new_n15826_ = ~ys__n18793 & ~ys__n38160;
  assign new_n15827_ = ys__n18793 & ys__n38160;
  assign new_n15828_ = ~new_n15826_ & ~new_n15827_;
  assign new_n15829_ = ~ys__n18795 & ~ys__n38161;
  assign new_n15830_ = ys__n18795 & ys__n38161;
  assign new_n15831_ = ~new_n15829_ & ~new_n15830_;
  assign new_n15832_ = ~new_n15828_ & ~new_n15831_;
  assign new_n15833_ = new_n15825_ & new_n15832_;
  assign new_n15834_ = new_n15818_ & new_n15833_;
  assign new_n15835_ = new_n15803_ & new_n15834_;
  assign new_n15836_ = new_n15772_ & new_n15835_;
  assign new_n15837_ = ~ys__n37743 & ~new_n15836_;
  assign new_n15838_ = ys__n842 & ~new_n15837_;
  assign new_n15839_ = ~new_n15725_ & ~new_n15838_;
  assign new_n15840_ = ~ys__n18821 & ~ys__n38146;
  assign new_n15841_ = ys__n18821 & ys__n38146;
  assign new_n15842_ = ~new_n15840_ & ~new_n15841_;
  assign new_n15843_ = ~ys__n18823 & ~ys__n38147;
  assign new_n15844_ = ys__n18823 & ys__n38147;
  assign new_n15845_ = ~new_n15843_ & ~new_n15844_;
  assign new_n15846_ = ~new_n15842_ & ~new_n15845_;
  assign new_n15847_ = ~ys__n18825 & ~ys__n38148;
  assign new_n15848_ = ys__n18825 & ys__n38148;
  assign new_n15849_ = ~new_n15847_ & ~new_n15848_;
  assign new_n15850_ = ~ys__n18827 & ~ys__n38149;
  assign new_n15851_ = ys__n18827 & ys__n38149;
  assign new_n15852_ = ~new_n15850_ & ~new_n15851_;
  assign new_n15853_ = ~new_n15849_ & ~new_n15852_;
  assign new_n15854_ = new_n15846_ & new_n15853_;
  assign new_n15855_ = ~ys__n18813 & ~ys__n38142;
  assign new_n15856_ = ys__n18813 & ys__n38142;
  assign new_n15857_ = ~new_n15855_ & ~new_n15856_;
  assign new_n15858_ = ~ys__n18815 & ~ys__n38143;
  assign new_n15859_ = ys__n18815 & ys__n38143;
  assign new_n15860_ = ~new_n15858_ & ~new_n15859_;
  assign new_n15861_ = ~new_n15857_ & ~new_n15860_;
  assign new_n15862_ = ~ys__n18817 & ~ys__n38144;
  assign new_n15863_ = ys__n18817 & ys__n38144;
  assign new_n15864_ = ~new_n15862_ & ~new_n15863_;
  assign new_n15865_ = ~ys__n18819 & ~ys__n38145;
  assign new_n15866_ = ys__n18819 & ys__n38145;
  assign new_n15867_ = ~new_n15865_ & ~new_n15866_;
  assign new_n15868_ = ~new_n15864_ & ~new_n15867_;
  assign new_n15869_ = new_n15861_ & new_n15868_;
  assign new_n15870_ = ~ys__n18805 & ~ys__n38138;
  assign new_n15871_ = ys__n18805 & ys__n38138;
  assign new_n15872_ = ~new_n15870_ & ~new_n15871_;
  assign new_n15873_ = ~ys__n18807 & ~ys__n38139;
  assign new_n15874_ = ys__n18807 & ys__n38139;
  assign new_n15875_ = ~new_n15873_ & ~new_n15874_;
  assign new_n15876_ = ~new_n15872_ & ~new_n15875_;
  assign new_n15877_ = ~ys__n18809 & ~ys__n38140;
  assign new_n15878_ = ys__n18809 & ys__n38140;
  assign new_n15879_ = ~new_n15877_ & ~new_n15878_;
  assign new_n15880_ = ~ys__n18811 & ~ys__n38141;
  assign new_n15881_ = ys__n18811 & ys__n38141;
  assign new_n15882_ = ~new_n15880_ & ~new_n15881_;
  assign new_n15883_ = ~new_n15879_ & ~new_n15882_;
  assign new_n15884_ = new_n15876_ & new_n15883_;
  assign new_n15885_ = new_n15869_ & new_n15884_;
  assign new_n15886_ = new_n15854_ & new_n15885_;
  assign new_n15887_ = ~ys__n18781 & ~ys__n38126;
  assign new_n15888_ = ys__n18781 & ys__n38126;
  assign new_n15889_ = ~new_n15887_ & ~new_n15888_;
  assign new_n15890_ = ~ys__n18783 & ~ys__n38127;
  assign new_n15891_ = ys__n18783 & ys__n38127;
  assign new_n15892_ = ~new_n15890_ & ~new_n15891_;
  assign new_n15893_ = ~new_n15889_ & ~new_n15892_;
  assign new_n15894_ = ~ys__n18785 & ~ys__n38128;
  assign new_n15895_ = ys__n18785 & ys__n38128;
  assign new_n15896_ = ~new_n15894_ & ~new_n15895_;
  assign new_n15897_ = ~ys__n18787 & ~ys__n38129;
  assign new_n15898_ = ys__n18787 & ys__n38129;
  assign new_n15899_ = ~new_n15897_ & ~new_n15898_;
  assign new_n15900_ = ~new_n15896_ & ~new_n15899_;
  assign new_n15901_ = new_n15893_ & new_n15900_;
  assign new_n15902_ = ~ys__n18773 & ~ys__n38122;
  assign new_n15903_ = ys__n18773 & ys__n38122;
  assign new_n15904_ = ~new_n15902_ & ~new_n15903_;
  assign new_n15905_ = ~ys__n18775 & ~ys__n38123;
  assign new_n15906_ = ys__n18775 & ys__n38123;
  assign new_n15907_ = ~new_n15905_ & ~new_n15906_;
  assign new_n15908_ = ~new_n15904_ & ~new_n15907_;
  assign new_n15909_ = ~ys__n18777 & ~ys__n38124;
  assign new_n15910_ = ys__n18777 & ys__n38124;
  assign new_n15911_ = ~new_n15909_ & ~new_n15910_;
  assign new_n15912_ = ~ys__n18779 & ~ys__n38125;
  assign new_n15913_ = ys__n18779 & ys__n38125;
  assign new_n15914_ = ~new_n15912_ & ~new_n15913_;
  assign new_n15915_ = ~new_n15911_ & ~new_n15914_;
  assign new_n15916_ = new_n15908_ & new_n15915_;
  assign new_n15917_ = new_n15901_ & new_n15916_;
  assign new_n15918_ = ~ys__n18797 & ~ys__n38134;
  assign new_n15919_ = ys__n18797 & ys__n38134;
  assign new_n15920_ = ~new_n15918_ & ~new_n15919_;
  assign new_n15921_ = ~ys__n18799 & ~ys__n38135;
  assign new_n15922_ = ys__n18799 & ys__n38135;
  assign new_n15923_ = ~new_n15921_ & ~new_n15922_;
  assign new_n15924_ = ~new_n15920_ & ~new_n15923_;
  assign new_n15925_ = ~ys__n18801 & ~ys__n38136;
  assign new_n15926_ = ys__n18801 & ys__n38136;
  assign new_n15927_ = ~new_n15925_ & ~new_n15926_;
  assign new_n15928_ = ~ys__n18803 & ~ys__n38137;
  assign new_n15929_ = ys__n18803 & ys__n38137;
  assign new_n15930_ = ~new_n15928_ & ~new_n15929_;
  assign new_n15931_ = ~new_n15927_ & ~new_n15930_;
  assign new_n15932_ = new_n15924_ & new_n15931_;
  assign new_n15933_ = ~ys__n18789 & ~ys__n38130;
  assign new_n15934_ = ys__n18789 & ys__n38130;
  assign new_n15935_ = ~new_n15933_ & ~new_n15934_;
  assign new_n15936_ = ~ys__n18791 & ~ys__n38131;
  assign new_n15937_ = ys__n18791 & ys__n38131;
  assign new_n15938_ = ~new_n15936_ & ~new_n15937_;
  assign new_n15939_ = ~new_n15935_ & ~new_n15938_;
  assign new_n15940_ = ~ys__n18793 & ~ys__n38132;
  assign new_n15941_ = ys__n18793 & ys__n38132;
  assign new_n15942_ = ~new_n15940_ & ~new_n15941_;
  assign new_n15943_ = ~ys__n18795 & ~ys__n38133;
  assign new_n15944_ = ys__n18795 & ys__n38133;
  assign new_n15945_ = ~new_n15943_ & ~new_n15944_;
  assign new_n15946_ = ~new_n15942_ & ~new_n15945_;
  assign new_n15947_ = new_n15939_ & new_n15946_;
  assign new_n15948_ = new_n15932_ & new_n15947_;
  assign new_n15949_ = new_n15917_ & new_n15948_;
  assign new_n15950_ = new_n15886_ & new_n15949_;
  assign new_n15951_ = ~ys__n37744 & ~new_n15950_;
  assign new_n15952_ = ys__n840 & ~new_n15951_;
  assign new_n15953_ = ~ys__n18821 & ~ys__n38118;
  assign new_n15954_ = ys__n18821 & ys__n38118;
  assign new_n15955_ = ~new_n15953_ & ~new_n15954_;
  assign new_n15956_ = ~ys__n18823 & ~ys__n38119;
  assign new_n15957_ = ys__n18823 & ys__n38119;
  assign new_n15958_ = ~new_n15956_ & ~new_n15957_;
  assign new_n15959_ = ~new_n15955_ & ~new_n15958_;
  assign new_n15960_ = ~ys__n18825 & ~ys__n38120;
  assign new_n15961_ = ys__n18825 & ys__n38120;
  assign new_n15962_ = ~new_n15960_ & ~new_n15961_;
  assign new_n15963_ = ~ys__n18827 & ~ys__n38121;
  assign new_n15964_ = ys__n18827 & ys__n38121;
  assign new_n15965_ = ~new_n15963_ & ~new_n15964_;
  assign new_n15966_ = ~new_n15962_ & ~new_n15965_;
  assign new_n15967_ = new_n15959_ & new_n15966_;
  assign new_n15968_ = ~ys__n18813 & ~ys__n38114;
  assign new_n15969_ = ys__n18813 & ys__n38114;
  assign new_n15970_ = ~new_n15968_ & ~new_n15969_;
  assign new_n15971_ = ~ys__n18815 & ~ys__n38115;
  assign new_n15972_ = ys__n18815 & ys__n38115;
  assign new_n15973_ = ~new_n15971_ & ~new_n15972_;
  assign new_n15974_ = ~new_n15970_ & ~new_n15973_;
  assign new_n15975_ = ~ys__n18817 & ~ys__n38116;
  assign new_n15976_ = ys__n18817 & ys__n38116;
  assign new_n15977_ = ~new_n15975_ & ~new_n15976_;
  assign new_n15978_ = ~ys__n18819 & ~ys__n38117;
  assign new_n15979_ = ys__n18819 & ys__n38117;
  assign new_n15980_ = ~new_n15978_ & ~new_n15979_;
  assign new_n15981_ = ~new_n15977_ & ~new_n15980_;
  assign new_n15982_ = new_n15974_ & new_n15981_;
  assign new_n15983_ = ~ys__n18805 & ~ys__n38110;
  assign new_n15984_ = ys__n18805 & ys__n38110;
  assign new_n15985_ = ~new_n15983_ & ~new_n15984_;
  assign new_n15986_ = ~ys__n18807 & ~ys__n38111;
  assign new_n15987_ = ys__n18807 & ys__n38111;
  assign new_n15988_ = ~new_n15986_ & ~new_n15987_;
  assign new_n15989_ = ~new_n15985_ & ~new_n15988_;
  assign new_n15990_ = ~ys__n18809 & ~ys__n38112;
  assign new_n15991_ = ys__n18809 & ys__n38112;
  assign new_n15992_ = ~new_n15990_ & ~new_n15991_;
  assign new_n15993_ = ~ys__n18811 & ~ys__n38113;
  assign new_n15994_ = ys__n18811 & ys__n38113;
  assign new_n15995_ = ~new_n15993_ & ~new_n15994_;
  assign new_n15996_ = ~new_n15992_ & ~new_n15995_;
  assign new_n15997_ = new_n15989_ & new_n15996_;
  assign new_n15998_ = new_n15982_ & new_n15997_;
  assign new_n15999_ = new_n15967_ & new_n15998_;
  assign new_n16000_ = ~ys__n18781 & ~ys__n38098;
  assign new_n16001_ = ys__n18781 & ys__n38098;
  assign new_n16002_ = ~new_n16000_ & ~new_n16001_;
  assign new_n16003_ = ~ys__n18783 & ~ys__n38099;
  assign new_n16004_ = ys__n18783 & ys__n38099;
  assign new_n16005_ = ~new_n16003_ & ~new_n16004_;
  assign new_n16006_ = ~new_n16002_ & ~new_n16005_;
  assign new_n16007_ = ~ys__n18785 & ~ys__n38100;
  assign new_n16008_ = ys__n18785 & ys__n38100;
  assign new_n16009_ = ~new_n16007_ & ~new_n16008_;
  assign new_n16010_ = ~ys__n18787 & ~ys__n38101;
  assign new_n16011_ = ys__n18787 & ys__n38101;
  assign new_n16012_ = ~new_n16010_ & ~new_n16011_;
  assign new_n16013_ = ~new_n16009_ & ~new_n16012_;
  assign new_n16014_ = new_n16006_ & new_n16013_;
  assign new_n16015_ = ~ys__n18773 & ~ys__n38094;
  assign new_n16016_ = ys__n18773 & ys__n38094;
  assign new_n16017_ = ~new_n16015_ & ~new_n16016_;
  assign new_n16018_ = ~ys__n18775 & ~ys__n38095;
  assign new_n16019_ = ys__n18775 & ys__n38095;
  assign new_n16020_ = ~new_n16018_ & ~new_n16019_;
  assign new_n16021_ = ~new_n16017_ & ~new_n16020_;
  assign new_n16022_ = ~ys__n18777 & ~ys__n38096;
  assign new_n16023_ = ys__n18777 & ys__n38096;
  assign new_n16024_ = ~new_n16022_ & ~new_n16023_;
  assign new_n16025_ = ~ys__n18779 & ~ys__n38097;
  assign new_n16026_ = ys__n18779 & ys__n38097;
  assign new_n16027_ = ~new_n16025_ & ~new_n16026_;
  assign new_n16028_ = ~new_n16024_ & ~new_n16027_;
  assign new_n16029_ = new_n16021_ & new_n16028_;
  assign new_n16030_ = new_n16014_ & new_n16029_;
  assign new_n16031_ = ~ys__n18797 & ~ys__n38106;
  assign new_n16032_ = ys__n18797 & ys__n38106;
  assign new_n16033_ = ~new_n16031_ & ~new_n16032_;
  assign new_n16034_ = ~ys__n18799 & ~ys__n38107;
  assign new_n16035_ = ys__n18799 & ys__n38107;
  assign new_n16036_ = ~new_n16034_ & ~new_n16035_;
  assign new_n16037_ = ~new_n16033_ & ~new_n16036_;
  assign new_n16038_ = ~ys__n18801 & ~ys__n38108;
  assign new_n16039_ = ys__n18801 & ys__n38108;
  assign new_n16040_ = ~new_n16038_ & ~new_n16039_;
  assign new_n16041_ = ~ys__n18803 & ~ys__n38109;
  assign new_n16042_ = ys__n18803 & ys__n38109;
  assign new_n16043_ = ~new_n16041_ & ~new_n16042_;
  assign new_n16044_ = ~new_n16040_ & ~new_n16043_;
  assign new_n16045_ = new_n16037_ & new_n16044_;
  assign new_n16046_ = ~ys__n18789 & ~ys__n38102;
  assign new_n16047_ = ys__n18789 & ys__n38102;
  assign new_n16048_ = ~new_n16046_ & ~new_n16047_;
  assign new_n16049_ = ~ys__n18791 & ~ys__n38103;
  assign new_n16050_ = ys__n18791 & ys__n38103;
  assign new_n16051_ = ~new_n16049_ & ~new_n16050_;
  assign new_n16052_ = ~new_n16048_ & ~new_n16051_;
  assign new_n16053_ = ~ys__n18793 & ~ys__n38104;
  assign new_n16054_ = ys__n18793 & ys__n38104;
  assign new_n16055_ = ~new_n16053_ & ~new_n16054_;
  assign new_n16056_ = ~ys__n18795 & ~ys__n38105;
  assign new_n16057_ = ys__n18795 & ys__n38105;
  assign new_n16058_ = ~new_n16056_ & ~new_n16057_;
  assign new_n16059_ = ~new_n16055_ & ~new_n16058_;
  assign new_n16060_ = new_n16052_ & new_n16059_;
  assign new_n16061_ = new_n16045_ & new_n16060_;
  assign new_n16062_ = new_n16030_ & new_n16061_;
  assign new_n16063_ = new_n15999_ & new_n16062_;
  assign new_n16064_ = ~ys__n37745 & ~new_n16063_;
  assign new_n16065_ = ys__n838 & ~new_n16064_;
  assign new_n16066_ = ~new_n15952_ & ~new_n16065_;
  assign new_n16067_ = new_n15839_ & new_n16066_;
  assign new_n16068_ = new_n15612_ & new_n16067_;
  assign new_n16069_ = ~ys__n18821 & ~ys__n37866;
  assign new_n16070_ = ys__n18821 & ys__n37866;
  assign new_n16071_ = ~new_n16069_ & ~new_n16070_;
  assign new_n16072_ = ~ys__n18823 & ~ys__n37867;
  assign new_n16073_ = ys__n18823 & ys__n37867;
  assign new_n16074_ = ~new_n16072_ & ~new_n16073_;
  assign new_n16075_ = ~new_n16071_ & ~new_n16074_;
  assign new_n16076_ = ~ys__n18825 & ~ys__n37868;
  assign new_n16077_ = ys__n18825 & ys__n37868;
  assign new_n16078_ = ~new_n16076_ & ~new_n16077_;
  assign new_n16079_ = ~ys__n18827 & ~ys__n37869;
  assign new_n16080_ = ys__n18827 & ys__n37869;
  assign new_n16081_ = ~new_n16079_ & ~new_n16080_;
  assign new_n16082_ = ~new_n16078_ & ~new_n16081_;
  assign new_n16083_ = new_n16075_ & new_n16082_;
  assign new_n16084_ = ~ys__n18813 & ~ys__n37862;
  assign new_n16085_ = ys__n18813 & ys__n37862;
  assign new_n16086_ = ~new_n16084_ & ~new_n16085_;
  assign new_n16087_ = ~ys__n18815 & ~ys__n37863;
  assign new_n16088_ = ys__n18815 & ys__n37863;
  assign new_n16089_ = ~new_n16087_ & ~new_n16088_;
  assign new_n16090_ = ~new_n16086_ & ~new_n16089_;
  assign new_n16091_ = ~ys__n18817 & ~ys__n37864;
  assign new_n16092_ = ys__n18817 & ys__n37864;
  assign new_n16093_ = ~new_n16091_ & ~new_n16092_;
  assign new_n16094_ = ~ys__n18819 & ~ys__n37865;
  assign new_n16095_ = ys__n18819 & ys__n37865;
  assign new_n16096_ = ~new_n16094_ & ~new_n16095_;
  assign new_n16097_ = ~new_n16093_ & ~new_n16096_;
  assign new_n16098_ = new_n16090_ & new_n16097_;
  assign new_n16099_ = ~ys__n18805 & ~ys__n37858;
  assign new_n16100_ = ys__n18805 & ys__n37858;
  assign new_n16101_ = ~new_n16099_ & ~new_n16100_;
  assign new_n16102_ = ~ys__n18807 & ~ys__n37859;
  assign new_n16103_ = ys__n18807 & ys__n37859;
  assign new_n16104_ = ~new_n16102_ & ~new_n16103_;
  assign new_n16105_ = ~new_n16101_ & ~new_n16104_;
  assign new_n16106_ = ~ys__n18809 & ~ys__n37860;
  assign new_n16107_ = ys__n18809 & ys__n37860;
  assign new_n16108_ = ~new_n16106_ & ~new_n16107_;
  assign new_n16109_ = ~ys__n18811 & ~ys__n37861;
  assign new_n16110_ = ys__n18811 & ys__n37861;
  assign new_n16111_ = ~new_n16109_ & ~new_n16110_;
  assign new_n16112_ = ~new_n16108_ & ~new_n16111_;
  assign new_n16113_ = new_n16105_ & new_n16112_;
  assign new_n16114_ = new_n16098_ & new_n16113_;
  assign new_n16115_ = new_n16083_ & new_n16114_;
  assign new_n16116_ = ~ys__n18781 & ~ys__n37846;
  assign new_n16117_ = ys__n18781 & ys__n37846;
  assign new_n16118_ = ~new_n16116_ & ~new_n16117_;
  assign new_n16119_ = ~ys__n18783 & ~ys__n37847;
  assign new_n16120_ = ys__n18783 & ys__n37847;
  assign new_n16121_ = ~new_n16119_ & ~new_n16120_;
  assign new_n16122_ = ~new_n16118_ & ~new_n16121_;
  assign new_n16123_ = ~ys__n18785 & ~ys__n37848;
  assign new_n16124_ = ys__n18785 & ys__n37848;
  assign new_n16125_ = ~new_n16123_ & ~new_n16124_;
  assign new_n16126_ = ~ys__n18787 & ~ys__n37849;
  assign new_n16127_ = ys__n18787 & ys__n37849;
  assign new_n16128_ = ~new_n16126_ & ~new_n16127_;
  assign new_n16129_ = ~new_n16125_ & ~new_n16128_;
  assign new_n16130_ = new_n16122_ & new_n16129_;
  assign new_n16131_ = ~ys__n18773 & ~ys__n37842;
  assign new_n16132_ = ys__n18773 & ys__n37842;
  assign new_n16133_ = ~new_n16131_ & ~new_n16132_;
  assign new_n16134_ = ~ys__n18775 & ~ys__n37843;
  assign new_n16135_ = ys__n18775 & ys__n37843;
  assign new_n16136_ = ~new_n16134_ & ~new_n16135_;
  assign new_n16137_ = ~new_n16133_ & ~new_n16136_;
  assign new_n16138_ = ~ys__n18777 & ~ys__n37844;
  assign new_n16139_ = ys__n18777 & ys__n37844;
  assign new_n16140_ = ~new_n16138_ & ~new_n16139_;
  assign new_n16141_ = ~ys__n18779 & ~ys__n37845;
  assign new_n16142_ = ys__n18779 & ys__n37845;
  assign new_n16143_ = ~new_n16141_ & ~new_n16142_;
  assign new_n16144_ = ~new_n16140_ & ~new_n16143_;
  assign new_n16145_ = new_n16137_ & new_n16144_;
  assign new_n16146_ = new_n16130_ & new_n16145_;
  assign new_n16147_ = ~ys__n18797 & ~ys__n37854;
  assign new_n16148_ = ys__n18797 & ys__n37854;
  assign new_n16149_ = ~new_n16147_ & ~new_n16148_;
  assign new_n16150_ = ~ys__n18799 & ~ys__n37855;
  assign new_n16151_ = ys__n18799 & ys__n37855;
  assign new_n16152_ = ~new_n16150_ & ~new_n16151_;
  assign new_n16153_ = ~new_n16149_ & ~new_n16152_;
  assign new_n16154_ = ~ys__n18801 & ~ys__n37856;
  assign new_n16155_ = ys__n18801 & ys__n37856;
  assign new_n16156_ = ~new_n16154_ & ~new_n16155_;
  assign new_n16157_ = ~ys__n18803 & ~ys__n37857;
  assign new_n16158_ = ys__n18803 & ys__n37857;
  assign new_n16159_ = ~new_n16157_ & ~new_n16158_;
  assign new_n16160_ = ~new_n16156_ & ~new_n16159_;
  assign new_n16161_ = new_n16153_ & new_n16160_;
  assign new_n16162_ = ~ys__n18789 & ~ys__n37850;
  assign new_n16163_ = ys__n18789 & ys__n37850;
  assign new_n16164_ = ~new_n16162_ & ~new_n16163_;
  assign new_n16165_ = ~ys__n18791 & ~ys__n37851;
  assign new_n16166_ = ys__n18791 & ys__n37851;
  assign new_n16167_ = ~new_n16165_ & ~new_n16166_;
  assign new_n16168_ = ~new_n16164_ & ~new_n16167_;
  assign new_n16169_ = ~ys__n18793 & ~ys__n37852;
  assign new_n16170_ = ys__n18793 & ys__n37852;
  assign new_n16171_ = ~new_n16169_ & ~new_n16170_;
  assign new_n16172_ = ~ys__n18795 & ~ys__n37853;
  assign new_n16173_ = ys__n18795 & ys__n37853;
  assign new_n16174_ = ~new_n16172_ & ~new_n16173_;
  assign new_n16175_ = ~new_n16171_ & ~new_n16174_;
  assign new_n16176_ = new_n16168_ & new_n16175_;
  assign new_n16177_ = new_n16161_ & new_n16176_;
  assign new_n16178_ = new_n16146_ & new_n16177_;
  assign new_n16179_ = new_n16115_ & new_n16178_;
  assign new_n16180_ = ~ys__n37754 & ~new_n16179_;
  assign new_n16181_ = ys__n850 & ~new_n16180_;
  assign new_n16182_ = ~ys__n18821 & ~ys__n37838;
  assign new_n16183_ = ys__n18821 & ys__n37838;
  assign new_n16184_ = ~new_n16182_ & ~new_n16183_;
  assign new_n16185_ = ~ys__n18823 & ~ys__n37839;
  assign new_n16186_ = ys__n18823 & ys__n37839;
  assign new_n16187_ = ~new_n16185_ & ~new_n16186_;
  assign new_n16188_ = ~new_n16184_ & ~new_n16187_;
  assign new_n16189_ = ~ys__n18825 & ~ys__n37840;
  assign new_n16190_ = ys__n18825 & ys__n37840;
  assign new_n16191_ = ~new_n16189_ & ~new_n16190_;
  assign new_n16192_ = ~ys__n18827 & ~ys__n37841;
  assign new_n16193_ = ys__n18827 & ys__n37841;
  assign new_n16194_ = ~new_n16192_ & ~new_n16193_;
  assign new_n16195_ = ~new_n16191_ & ~new_n16194_;
  assign new_n16196_ = new_n16188_ & new_n16195_;
  assign new_n16197_ = ~ys__n18813 & ~ys__n37834;
  assign new_n16198_ = ys__n18813 & ys__n37834;
  assign new_n16199_ = ~new_n16197_ & ~new_n16198_;
  assign new_n16200_ = ~ys__n18815 & ~ys__n37835;
  assign new_n16201_ = ys__n18815 & ys__n37835;
  assign new_n16202_ = ~new_n16200_ & ~new_n16201_;
  assign new_n16203_ = ~new_n16199_ & ~new_n16202_;
  assign new_n16204_ = ~ys__n18817 & ~ys__n37836;
  assign new_n16205_ = ys__n18817 & ys__n37836;
  assign new_n16206_ = ~new_n16204_ & ~new_n16205_;
  assign new_n16207_ = ~ys__n18819 & ~ys__n37837;
  assign new_n16208_ = ys__n18819 & ys__n37837;
  assign new_n16209_ = ~new_n16207_ & ~new_n16208_;
  assign new_n16210_ = ~new_n16206_ & ~new_n16209_;
  assign new_n16211_ = new_n16203_ & new_n16210_;
  assign new_n16212_ = ~ys__n18805 & ~ys__n37830;
  assign new_n16213_ = ys__n18805 & ys__n37830;
  assign new_n16214_ = ~new_n16212_ & ~new_n16213_;
  assign new_n16215_ = ~ys__n18807 & ~ys__n37831;
  assign new_n16216_ = ys__n18807 & ys__n37831;
  assign new_n16217_ = ~new_n16215_ & ~new_n16216_;
  assign new_n16218_ = ~new_n16214_ & ~new_n16217_;
  assign new_n16219_ = ~ys__n18809 & ~ys__n37832;
  assign new_n16220_ = ys__n18809 & ys__n37832;
  assign new_n16221_ = ~new_n16219_ & ~new_n16220_;
  assign new_n16222_ = ~ys__n18811 & ~ys__n37833;
  assign new_n16223_ = ys__n18811 & ys__n37833;
  assign new_n16224_ = ~new_n16222_ & ~new_n16223_;
  assign new_n16225_ = ~new_n16221_ & ~new_n16224_;
  assign new_n16226_ = new_n16218_ & new_n16225_;
  assign new_n16227_ = new_n16211_ & new_n16226_;
  assign new_n16228_ = new_n16196_ & new_n16227_;
  assign new_n16229_ = ~ys__n18781 & ~ys__n37818;
  assign new_n16230_ = ys__n18781 & ys__n37818;
  assign new_n16231_ = ~new_n16229_ & ~new_n16230_;
  assign new_n16232_ = ~ys__n18783 & ~ys__n37819;
  assign new_n16233_ = ys__n18783 & ys__n37819;
  assign new_n16234_ = ~new_n16232_ & ~new_n16233_;
  assign new_n16235_ = ~new_n16231_ & ~new_n16234_;
  assign new_n16236_ = ~ys__n18785 & ~ys__n37820;
  assign new_n16237_ = ys__n18785 & ys__n37820;
  assign new_n16238_ = ~new_n16236_ & ~new_n16237_;
  assign new_n16239_ = ~ys__n18787 & ~ys__n37821;
  assign new_n16240_ = ys__n18787 & ys__n37821;
  assign new_n16241_ = ~new_n16239_ & ~new_n16240_;
  assign new_n16242_ = ~new_n16238_ & ~new_n16241_;
  assign new_n16243_ = new_n16235_ & new_n16242_;
  assign new_n16244_ = ~ys__n18773 & ~ys__n37814;
  assign new_n16245_ = ys__n18773 & ys__n37814;
  assign new_n16246_ = ~new_n16244_ & ~new_n16245_;
  assign new_n16247_ = ~ys__n18775 & ~ys__n37815;
  assign new_n16248_ = ys__n18775 & ys__n37815;
  assign new_n16249_ = ~new_n16247_ & ~new_n16248_;
  assign new_n16250_ = ~new_n16246_ & ~new_n16249_;
  assign new_n16251_ = ~ys__n18777 & ~ys__n37816;
  assign new_n16252_ = ys__n18777 & ys__n37816;
  assign new_n16253_ = ~new_n16251_ & ~new_n16252_;
  assign new_n16254_ = ~ys__n18779 & ~ys__n37817;
  assign new_n16255_ = ys__n18779 & ys__n37817;
  assign new_n16256_ = ~new_n16254_ & ~new_n16255_;
  assign new_n16257_ = ~new_n16253_ & ~new_n16256_;
  assign new_n16258_ = new_n16250_ & new_n16257_;
  assign new_n16259_ = new_n16243_ & new_n16258_;
  assign new_n16260_ = ~ys__n18797 & ~ys__n37826;
  assign new_n16261_ = ys__n18797 & ys__n37826;
  assign new_n16262_ = ~new_n16260_ & ~new_n16261_;
  assign new_n16263_ = ~ys__n18799 & ~ys__n37827;
  assign new_n16264_ = ys__n18799 & ys__n37827;
  assign new_n16265_ = ~new_n16263_ & ~new_n16264_;
  assign new_n16266_ = ~new_n16262_ & ~new_n16265_;
  assign new_n16267_ = ~ys__n18801 & ~ys__n37828;
  assign new_n16268_ = ys__n18801 & ys__n37828;
  assign new_n16269_ = ~new_n16267_ & ~new_n16268_;
  assign new_n16270_ = ~ys__n18803 & ~ys__n37829;
  assign new_n16271_ = ys__n18803 & ys__n37829;
  assign new_n16272_ = ~new_n16270_ & ~new_n16271_;
  assign new_n16273_ = ~new_n16269_ & ~new_n16272_;
  assign new_n16274_ = new_n16266_ & new_n16273_;
  assign new_n16275_ = ~ys__n18789 & ~ys__n37822;
  assign new_n16276_ = ys__n18789 & ys__n37822;
  assign new_n16277_ = ~new_n16275_ & ~new_n16276_;
  assign new_n16278_ = ~ys__n18791 & ~ys__n37823;
  assign new_n16279_ = ys__n18791 & ys__n37823;
  assign new_n16280_ = ~new_n16278_ & ~new_n16279_;
  assign new_n16281_ = ~new_n16277_ & ~new_n16280_;
  assign new_n16282_ = ~ys__n18793 & ~ys__n37824;
  assign new_n16283_ = ys__n18793 & ys__n37824;
  assign new_n16284_ = ~new_n16282_ & ~new_n16283_;
  assign new_n16285_ = ~ys__n18795 & ~ys__n37825;
  assign new_n16286_ = ys__n18795 & ys__n37825;
  assign new_n16287_ = ~new_n16285_ & ~new_n16286_;
  assign new_n16288_ = ~new_n16284_ & ~new_n16287_;
  assign new_n16289_ = new_n16281_ & new_n16288_;
  assign new_n16290_ = new_n16274_ & new_n16289_;
  assign new_n16291_ = new_n16259_ & new_n16290_;
  assign new_n16292_ = new_n16228_ & new_n16291_;
  assign new_n16293_ = ~ys__n37755 & ~new_n16292_;
  assign new_n16294_ = ys__n848 & ~new_n16293_;
  assign new_n16295_ = ~new_n16181_ & ~new_n16294_;
  assign new_n16296_ = ~ys__n18821 & ~ys__n37810;
  assign new_n16297_ = ys__n18821 & ys__n37810;
  assign new_n16298_ = ~new_n16296_ & ~new_n16297_;
  assign new_n16299_ = ~ys__n18823 & ~ys__n37811;
  assign new_n16300_ = ys__n18823 & ys__n37811;
  assign new_n16301_ = ~new_n16299_ & ~new_n16300_;
  assign new_n16302_ = ~new_n16298_ & ~new_n16301_;
  assign new_n16303_ = ~ys__n18825 & ~ys__n37812;
  assign new_n16304_ = ys__n18825 & ys__n37812;
  assign new_n16305_ = ~new_n16303_ & ~new_n16304_;
  assign new_n16306_ = ~ys__n18827 & ~ys__n37813;
  assign new_n16307_ = ys__n18827 & ys__n37813;
  assign new_n16308_ = ~new_n16306_ & ~new_n16307_;
  assign new_n16309_ = ~new_n16305_ & ~new_n16308_;
  assign new_n16310_ = new_n16302_ & new_n16309_;
  assign new_n16311_ = ~ys__n18813 & ~ys__n37806;
  assign new_n16312_ = ys__n18813 & ys__n37806;
  assign new_n16313_ = ~new_n16311_ & ~new_n16312_;
  assign new_n16314_ = ~ys__n18815 & ~ys__n37807;
  assign new_n16315_ = ys__n18815 & ys__n37807;
  assign new_n16316_ = ~new_n16314_ & ~new_n16315_;
  assign new_n16317_ = ~new_n16313_ & ~new_n16316_;
  assign new_n16318_ = ~ys__n18817 & ~ys__n37808;
  assign new_n16319_ = ys__n18817 & ys__n37808;
  assign new_n16320_ = ~new_n16318_ & ~new_n16319_;
  assign new_n16321_ = ~ys__n18819 & ~ys__n37809;
  assign new_n16322_ = ys__n18819 & ys__n37809;
  assign new_n16323_ = ~new_n16321_ & ~new_n16322_;
  assign new_n16324_ = ~new_n16320_ & ~new_n16323_;
  assign new_n16325_ = new_n16317_ & new_n16324_;
  assign new_n16326_ = ~ys__n18805 & ~ys__n37802;
  assign new_n16327_ = ys__n18805 & ys__n37802;
  assign new_n16328_ = ~new_n16326_ & ~new_n16327_;
  assign new_n16329_ = ~ys__n18807 & ~ys__n37803;
  assign new_n16330_ = ys__n18807 & ys__n37803;
  assign new_n16331_ = ~new_n16329_ & ~new_n16330_;
  assign new_n16332_ = ~new_n16328_ & ~new_n16331_;
  assign new_n16333_ = ~ys__n18809 & ~ys__n37804;
  assign new_n16334_ = ys__n18809 & ys__n37804;
  assign new_n16335_ = ~new_n16333_ & ~new_n16334_;
  assign new_n16336_ = ~ys__n18811 & ~ys__n37805;
  assign new_n16337_ = ys__n18811 & ys__n37805;
  assign new_n16338_ = ~new_n16336_ & ~new_n16337_;
  assign new_n16339_ = ~new_n16335_ & ~new_n16338_;
  assign new_n16340_ = new_n16332_ & new_n16339_;
  assign new_n16341_ = new_n16325_ & new_n16340_;
  assign new_n16342_ = new_n16310_ & new_n16341_;
  assign new_n16343_ = ~ys__n18781 & ~ys__n37790;
  assign new_n16344_ = ys__n18781 & ys__n37790;
  assign new_n16345_ = ~new_n16343_ & ~new_n16344_;
  assign new_n16346_ = ~ys__n18783 & ~ys__n37791;
  assign new_n16347_ = ys__n18783 & ys__n37791;
  assign new_n16348_ = ~new_n16346_ & ~new_n16347_;
  assign new_n16349_ = ~new_n16345_ & ~new_n16348_;
  assign new_n16350_ = ~ys__n18785 & ~ys__n37792;
  assign new_n16351_ = ys__n18785 & ys__n37792;
  assign new_n16352_ = ~new_n16350_ & ~new_n16351_;
  assign new_n16353_ = ~ys__n18787 & ~ys__n37793;
  assign new_n16354_ = ys__n18787 & ys__n37793;
  assign new_n16355_ = ~new_n16353_ & ~new_n16354_;
  assign new_n16356_ = ~new_n16352_ & ~new_n16355_;
  assign new_n16357_ = new_n16349_ & new_n16356_;
  assign new_n16358_ = ~ys__n18773 & ~ys__n37786;
  assign new_n16359_ = ys__n18773 & ys__n37786;
  assign new_n16360_ = ~new_n16358_ & ~new_n16359_;
  assign new_n16361_ = ~ys__n18775 & ~ys__n37787;
  assign new_n16362_ = ys__n18775 & ys__n37787;
  assign new_n16363_ = ~new_n16361_ & ~new_n16362_;
  assign new_n16364_ = ~new_n16360_ & ~new_n16363_;
  assign new_n16365_ = ~ys__n18777 & ~ys__n37788;
  assign new_n16366_ = ys__n18777 & ys__n37788;
  assign new_n16367_ = ~new_n16365_ & ~new_n16366_;
  assign new_n16368_ = ~ys__n18779 & ~ys__n37789;
  assign new_n16369_ = ys__n18779 & ys__n37789;
  assign new_n16370_ = ~new_n16368_ & ~new_n16369_;
  assign new_n16371_ = ~new_n16367_ & ~new_n16370_;
  assign new_n16372_ = new_n16364_ & new_n16371_;
  assign new_n16373_ = new_n16357_ & new_n16372_;
  assign new_n16374_ = ~ys__n18797 & ~ys__n37798;
  assign new_n16375_ = ys__n18797 & ys__n37798;
  assign new_n16376_ = ~new_n16374_ & ~new_n16375_;
  assign new_n16377_ = ~ys__n18799 & ~ys__n37799;
  assign new_n16378_ = ys__n18799 & ys__n37799;
  assign new_n16379_ = ~new_n16377_ & ~new_n16378_;
  assign new_n16380_ = ~new_n16376_ & ~new_n16379_;
  assign new_n16381_ = ~ys__n18801 & ~ys__n37800;
  assign new_n16382_ = ys__n18801 & ys__n37800;
  assign new_n16383_ = ~new_n16381_ & ~new_n16382_;
  assign new_n16384_ = ~ys__n18803 & ~ys__n37801;
  assign new_n16385_ = ys__n18803 & ys__n37801;
  assign new_n16386_ = ~new_n16384_ & ~new_n16385_;
  assign new_n16387_ = ~new_n16383_ & ~new_n16386_;
  assign new_n16388_ = new_n16380_ & new_n16387_;
  assign new_n16389_ = ~ys__n18789 & ~ys__n37794;
  assign new_n16390_ = ys__n18789 & ys__n37794;
  assign new_n16391_ = ~new_n16389_ & ~new_n16390_;
  assign new_n16392_ = ~ys__n18791 & ~ys__n37795;
  assign new_n16393_ = ys__n18791 & ys__n37795;
  assign new_n16394_ = ~new_n16392_ & ~new_n16393_;
  assign new_n16395_ = ~new_n16391_ & ~new_n16394_;
  assign new_n16396_ = ~ys__n18793 & ~ys__n37796;
  assign new_n16397_ = ys__n18793 & ys__n37796;
  assign new_n16398_ = ~new_n16396_ & ~new_n16397_;
  assign new_n16399_ = ~ys__n18795 & ~ys__n37797;
  assign new_n16400_ = ys__n18795 & ys__n37797;
  assign new_n16401_ = ~new_n16399_ & ~new_n16400_;
  assign new_n16402_ = ~new_n16398_ & ~new_n16401_;
  assign new_n16403_ = new_n16395_ & new_n16402_;
  assign new_n16404_ = new_n16388_ & new_n16403_;
  assign new_n16405_ = new_n16373_ & new_n16404_;
  assign new_n16406_ = new_n16342_ & new_n16405_;
  assign new_n16407_ = ~ys__n37756 & ~new_n16406_;
  assign new_n16408_ = ys__n846 & ~new_n16407_;
  assign new_n16409_ = ~ys__n18821 & ~ys__n37782;
  assign new_n16410_ = ys__n18821 & ys__n37782;
  assign new_n16411_ = ~new_n16409_ & ~new_n16410_;
  assign new_n16412_ = ~ys__n18823 & ~ys__n37783;
  assign new_n16413_ = ys__n18823 & ys__n37783;
  assign new_n16414_ = ~new_n16412_ & ~new_n16413_;
  assign new_n16415_ = ~new_n16411_ & ~new_n16414_;
  assign new_n16416_ = ~ys__n18825 & ~ys__n37784;
  assign new_n16417_ = ys__n18825 & ys__n37784;
  assign new_n16418_ = ~new_n16416_ & ~new_n16417_;
  assign new_n16419_ = ~ys__n18827 & ~ys__n37785;
  assign new_n16420_ = ys__n18827 & ys__n37785;
  assign new_n16421_ = ~new_n16419_ & ~new_n16420_;
  assign new_n16422_ = ~new_n16418_ & ~new_n16421_;
  assign new_n16423_ = new_n16415_ & new_n16422_;
  assign new_n16424_ = ~ys__n18813 & ~ys__n37778;
  assign new_n16425_ = ys__n18813 & ys__n37778;
  assign new_n16426_ = ~new_n16424_ & ~new_n16425_;
  assign new_n16427_ = ~ys__n18815 & ~ys__n37779;
  assign new_n16428_ = ys__n18815 & ys__n37779;
  assign new_n16429_ = ~new_n16427_ & ~new_n16428_;
  assign new_n16430_ = ~new_n16426_ & ~new_n16429_;
  assign new_n16431_ = ~ys__n18817 & ~ys__n37780;
  assign new_n16432_ = ys__n18817 & ys__n37780;
  assign new_n16433_ = ~new_n16431_ & ~new_n16432_;
  assign new_n16434_ = ~ys__n18819 & ~ys__n37781;
  assign new_n16435_ = ys__n18819 & ys__n37781;
  assign new_n16436_ = ~new_n16434_ & ~new_n16435_;
  assign new_n16437_ = ~new_n16433_ & ~new_n16436_;
  assign new_n16438_ = new_n16430_ & new_n16437_;
  assign new_n16439_ = ~ys__n18805 & ~ys__n37774;
  assign new_n16440_ = ys__n18805 & ys__n37774;
  assign new_n16441_ = ~new_n16439_ & ~new_n16440_;
  assign new_n16442_ = ~ys__n18807 & ~ys__n37775;
  assign new_n16443_ = ys__n18807 & ys__n37775;
  assign new_n16444_ = ~new_n16442_ & ~new_n16443_;
  assign new_n16445_ = ~new_n16441_ & ~new_n16444_;
  assign new_n16446_ = ~ys__n18809 & ~ys__n37776;
  assign new_n16447_ = ys__n18809 & ys__n37776;
  assign new_n16448_ = ~new_n16446_ & ~new_n16447_;
  assign new_n16449_ = ~ys__n18811 & ~ys__n37777;
  assign new_n16450_ = ys__n18811 & ys__n37777;
  assign new_n16451_ = ~new_n16449_ & ~new_n16450_;
  assign new_n16452_ = ~new_n16448_ & ~new_n16451_;
  assign new_n16453_ = new_n16445_ & new_n16452_;
  assign new_n16454_ = new_n16438_ & new_n16453_;
  assign new_n16455_ = new_n16423_ & new_n16454_;
  assign new_n16456_ = ~ys__n18781 & ~ys__n37762;
  assign new_n16457_ = ys__n18781 & ys__n37762;
  assign new_n16458_ = ~new_n16456_ & ~new_n16457_;
  assign new_n16459_ = ~ys__n18783 & ~ys__n37763;
  assign new_n16460_ = ys__n18783 & ys__n37763;
  assign new_n16461_ = ~new_n16459_ & ~new_n16460_;
  assign new_n16462_ = ~new_n16458_ & ~new_n16461_;
  assign new_n16463_ = ~ys__n18785 & ~ys__n37764;
  assign new_n16464_ = ys__n18785 & ys__n37764;
  assign new_n16465_ = ~new_n16463_ & ~new_n16464_;
  assign new_n16466_ = ~ys__n18787 & ~ys__n37765;
  assign new_n16467_ = ys__n18787 & ys__n37765;
  assign new_n16468_ = ~new_n16466_ & ~new_n16467_;
  assign new_n16469_ = ~new_n16465_ & ~new_n16468_;
  assign new_n16470_ = new_n16462_ & new_n16469_;
  assign new_n16471_ = ~ys__n18773 & ~ys__n37758;
  assign new_n16472_ = ys__n18773 & ys__n37758;
  assign new_n16473_ = ~new_n16471_ & ~new_n16472_;
  assign new_n16474_ = ~ys__n18775 & ~ys__n37759;
  assign new_n16475_ = ys__n18775 & ys__n37759;
  assign new_n16476_ = ~new_n16474_ & ~new_n16475_;
  assign new_n16477_ = ~new_n16473_ & ~new_n16476_;
  assign new_n16478_ = ~ys__n18777 & ~ys__n37760;
  assign new_n16479_ = ys__n18777 & ys__n37760;
  assign new_n16480_ = ~new_n16478_ & ~new_n16479_;
  assign new_n16481_ = ~ys__n18779 & ~ys__n37761;
  assign new_n16482_ = ys__n18779 & ys__n37761;
  assign new_n16483_ = ~new_n16481_ & ~new_n16482_;
  assign new_n16484_ = ~new_n16480_ & ~new_n16483_;
  assign new_n16485_ = new_n16477_ & new_n16484_;
  assign new_n16486_ = new_n16470_ & new_n16485_;
  assign new_n16487_ = ~ys__n18797 & ~ys__n37770;
  assign new_n16488_ = ys__n18797 & ys__n37770;
  assign new_n16489_ = ~new_n16487_ & ~new_n16488_;
  assign new_n16490_ = ~ys__n18799 & ~ys__n37771;
  assign new_n16491_ = ys__n18799 & ys__n37771;
  assign new_n16492_ = ~new_n16490_ & ~new_n16491_;
  assign new_n16493_ = ~new_n16489_ & ~new_n16492_;
  assign new_n16494_ = ~ys__n18801 & ~ys__n37772;
  assign new_n16495_ = ys__n18801 & ys__n37772;
  assign new_n16496_ = ~new_n16494_ & ~new_n16495_;
  assign new_n16497_ = ~ys__n18803 & ~ys__n37773;
  assign new_n16498_ = ys__n18803 & ys__n37773;
  assign new_n16499_ = ~new_n16497_ & ~new_n16498_;
  assign new_n16500_ = ~new_n16496_ & ~new_n16499_;
  assign new_n16501_ = new_n16493_ & new_n16500_;
  assign new_n16502_ = ~ys__n18789 & ~ys__n37766;
  assign new_n16503_ = ys__n18789 & ys__n37766;
  assign new_n16504_ = ~new_n16502_ & ~new_n16503_;
  assign new_n16505_ = ~ys__n18791 & ~ys__n37767;
  assign new_n16506_ = ys__n18791 & ys__n37767;
  assign new_n16507_ = ~new_n16505_ & ~new_n16506_;
  assign new_n16508_ = ~new_n16504_ & ~new_n16507_;
  assign new_n16509_ = ~ys__n18793 & ~ys__n37768;
  assign new_n16510_ = ys__n18793 & ys__n37768;
  assign new_n16511_ = ~new_n16509_ & ~new_n16510_;
  assign new_n16512_ = ~ys__n18795 & ~ys__n37769;
  assign new_n16513_ = ys__n18795 & ys__n37769;
  assign new_n16514_ = ~new_n16512_ & ~new_n16513_;
  assign new_n16515_ = ~new_n16511_ & ~new_n16514_;
  assign new_n16516_ = new_n16508_ & new_n16515_;
  assign new_n16517_ = new_n16501_ & new_n16516_;
  assign new_n16518_ = new_n16486_ & new_n16517_;
  assign new_n16519_ = new_n16455_ & new_n16518_;
  assign new_n16520_ = ~ys__n37757 & ~new_n16519_;
  assign new_n16521_ = ys__n116 & ~new_n16520_;
  assign new_n16522_ = ~new_n16408_ & ~new_n16521_;
  assign new_n16523_ = new_n16295_ & new_n16522_;
  assign new_n16524_ = ~ys__n18821 & ~ys__n37978;
  assign new_n16525_ = ys__n18821 & ys__n37978;
  assign new_n16526_ = ~new_n16524_ & ~new_n16525_;
  assign new_n16527_ = ~ys__n18823 & ~ys__n37979;
  assign new_n16528_ = ys__n18823 & ys__n37979;
  assign new_n16529_ = ~new_n16527_ & ~new_n16528_;
  assign new_n16530_ = ~new_n16526_ & ~new_n16529_;
  assign new_n16531_ = ~ys__n18825 & ~ys__n37980;
  assign new_n16532_ = ys__n18825 & ys__n37980;
  assign new_n16533_ = ~new_n16531_ & ~new_n16532_;
  assign new_n16534_ = ~ys__n18827 & ~ys__n37981;
  assign new_n16535_ = ys__n18827 & ys__n37981;
  assign new_n16536_ = ~new_n16534_ & ~new_n16535_;
  assign new_n16537_ = ~new_n16533_ & ~new_n16536_;
  assign new_n16538_ = new_n16530_ & new_n16537_;
  assign new_n16539_ = ~ys__n18813 & ~ys__n37974;
  assign new_n16540_ = ys__n18813 & ys__n37974;
  assign new_n16541_ = ~new_n16539_ & ~new_n16540_;
  assign new_n16542_ = ~ys__n18815 & ~ys__n37975;
  assign new_n16543_ = ys__n18815 & ys__n37975;
  assign new_n16544_ = ~new_n16542_ & ~new_n16543_;
  assign new_n16545_ = ~new_n16541_ & ~new_n16544_;
  assign new_n16546_ = ~ys__n18817 & ~ys__n37976;
  assign new_n16547_ = ys__n18817 & ys__n37976;
  assign new_n16548_ = ~new_n16546_ & ~new_n16547_;
  assign new_n16549_ = ~ys__n18819 & ~ys__n37977;
  assign new_n16550_ = ys__n18819 & ys__n37977;
  assign new_n16551_ = ~new_n16549_ & ~new_n16550_;
  assign new_n16552_ = ~new_n16548_ & ~new_n16551_;
  assign new_n16553_ = new_n16545_ & new_n16552_;
  assign new_n16554_ = ~ys__n18805 & ~ys__n37970;
  assign new_n16555_ = ys__n18805 & ys__n37970;
  assign new_n16556_ = ~new_n16554_ & ~new_n16555_;
  assign new_n16557_ = ~ys__n18807 & ~ys__n37971;
  assign new_n16558_ = ys__n18807 & ys__n37971;
  assign new_n16559_ = ~new_n16557_ & ~new_n16558_;
  assign new_n16560_ = ~new_n16556_ & ~new_n16559_;
  assign new_n16561_ = ~ys__n18809 & ~ys__n37972;
  assign new_n16562_ = ys__n18809 & ys__n37972;
  assign new_n16563_ = ~new_n16561_ & ~new_n16562_;
  assign new_n16564_ = ~ys__n18811 & ~ys__n37973;
  assign new_n16565_ = ys__n18811 & ys__n37973;
  assign new_n16566_ = ~new_n16564_ & ~new_n16565_;
  assign new_n16567_ = ~new_n16563_ & ~new_n16566_;
  assign new_n16568_ = new_n16560_ & new_n16567_;
  assign new_n16569_ = new_n16553_ & new_n16568_;
  assign new_n16570_ = new_n16538_ & new_n16569_;
  assign new_n16571_ = ~ys__n18781 & ~ys__n37958;
  assign new_n16572_ = ys__n18781 & ys__n37958;
  assign new_n16573_ = ~new_n16571_ & ~new_n16572_;
  assign new_n16574_ = ~ys__n18783 & ~ys__n37959;
  assign new_n16575_ = ys__n18783 & ys__n37959;
  assign new_n16576_ = ~new_n16574_ & ~new_n16575_;
  assign new_n16577_ = ~new_n16573_ & ~new_n16576_;
  assign new_n16578_ = ~ys__n18785 & ~ys__n37960;
  assign new_n16579_ = ys__n18785 & ys__n37960;
  assign new_n16580_ = ~new_n16578_ & ~new_n16579_;
  assign new_n16581_ = ~ys__n18787 & ~ys__n37961;
  assign new_n16582_ = ys__n18787 & ys__n37961;
  assign new_n16583_ = ~new_n16581_ & ~new_n16582_;
  assign new_n16584_ = ~new_n16580_ & ~new_n16583_;
  assign new_n16585_ = new_n16577_ & new_n16584_;
  assign new_n16586_ = ~ys__n18773 & ~ys__n37954;
  assign new_n16587_ = ys__n18773 & ys__n37954;
  assign new_n16588_ = ~new_n16586_ & ~new_n16587_;
  assign new_n16589_ = ~ys__n18775 & ~ys__n37955;
  assign new_n16590_ = ys__n18775 & ys__n37955;
  assign new_n16591_ = ~new_n16589_ & ~new_n16590_;
  assign new_n16592_ = ~new_n16588_ & ~new_n16591_;
  assign new_n16593_ = ~ys__n18777 & ~ys__n37956;
  assign new_n16594_ = ys__n18777 & ys__n37956;
  assign new_n16595_ = ~new_n16593_ & ~new_n16594_;
  assign new_n16596_ = ~ys__n18779 & ~ys__n37957;
  assign new_n16597_ = ys__n18779 & ys__n37957;
  assign new_n16598_ = ~new_n16596_ & ~new_n16597_;
  assign new_n16599_ = ~new_n16595_ & ~new_n16598_;
  assign new_n16600_ = new_n16592_ & new_n16599_;
  assign new_n16601_ = new_n16585_ & new_n16600_;
  assign new_n16602_ = ~ys__n18797 & ~ys__n37966;
  assign new_n16603_ = ys__n18797 & ys__n37966;
  assign new_n16604_ = ~new_n16602_ & ~new_n16603_;
  assign new_n16605_ = ~ys__n18799 & ~ys__n37967;
  assign new_n16606_ = ys__n18799 & ys__n37967;
  assign new_n16607_ = ~new_n16605_ & ~new_n16606_;
  assign new_n16608_ = ~new_n16604_ & ~new_n16607_;
  assign new_n16609_ = ~ys__n18801 & ~ys__n37968;
  assign new_n16610_ = ys__n18801 & ys__n37968;
  assign new_n16611_ = ~new_n16609_ & ~new_n16610_;
  assign new_n16612_ = ~ys__n18803 & ~ys__n37969;
  assign new_n16613_ = ys__n18803 & ys__n37969;
  assign new_n16614_ = ~new_n16612_ & ~new_n16613_;
  assign new_n16615_ = ~new_n16611_ & ~new_n16614_;
  assign new_n16616_ = new_n16608_ & new_n16615_;
  assign new_n16617_ = ~ys__n18789 & ~ys__n37962;
  assign new_n16618_ = ys__n18789 & ys__n37962;
  assign new_n16619_ = ~new_n16617_ & ~new_n16618_;
  assign new_n16620_ = ~ys__n18791 & ~ys__n37963;
  assign new_n16621_ = ys__n18791 & ys__n37963;
  assign new_n16622_ = ~new_n16620_ & ~new_n16621_;
  assign new_n16623_ = ~new_n16619_ & ~new_n16622_;
  assign new_n16624_ = ~ys__n18793 & ~ys__n37964;
  assign new_n16625_ = ys__n18793 & ys__n37964;
  assign new_n16626_ = ~new_n16624_ & ~new_n16625_;
  assign new_n16627_ = ~ys__n18795 & ~ys__n37965;
  assign new_n16628_ = ys__n18795 & ys__n37965;
  assign new_n16629_ = ~new_n16627_ & ~new_n16628_;
  assign new_n16630_ = ~new_n16626_ & ~new_n16629_;
  assign new_n16631_ = new_n16623_ & new_n16630_;
  assign new_n16632_ = new_n16616_ & new_n16631_;
  assign new_n16633_ = new_n16601_ & new_n16632_;
  assign new_n16634_ = new_n16570_ & new_n16633_;
  assign new_n16635_ = ~ys__n37750 & ~new_n16634_;
  assign new_n16636_ = ys__n858 & ~new_n16635_;
  assign new_n16637_ = ~ys__n18821 & ~ys__n37950;
  assign new_n16638_ = ys__n18821 & ys__n37950;
  assign new_n16639_ = ~new_n16637_ & ~new_n16638_;
  assign new_n16640_ = ~ys__n18823 & ~ys__n37951;
  assign new_n16641_ = ys__n18823 & ys__n37951;
  assign new_n16642_ = ~new_n16640_ & ~new_n16641_;
  assign new_n16643_ = ~new_n16639_ & ~new_n16642_;
  assign new_n16644_ = ~ys__n18825 & ~ys__n37952;
  assign new_n16645_ = ys__n18825 & ys__n37952;
  assign new_n16646_ = ~new_n16644_ & ~new_n16645_;
  assign new_n16647_ = ~ys__n18827 & ~ys__n37953;
  assign new_n16648_ = ys__n18827 & ys__n37953;
  assign new_n16649_ = ~new_n16647_ & ~new_n16648_;
  assign new_n16650_ = ~new_n16646_ & ~new_n16649_;
  assign new_n16651_ = new_n16643_ & new_n16650_;
  assign new_n16652_ = ~ys__n18813 & ~ys__n37946;
  assign new_n16653_ = ys__n18813 & ys__n37946;
  assign new_n16654_ = ~new_n16652_ & ~new_n16653_;
  assign new_n16655_ = ~ys__n18815 & ~ys__n37947;
  assign new_n16656_ = ys__n18815 & ys__n37947;
  assign new_n16657_ = ~new_n16655_ & ~new_n16656_;
  assign new_n16658_ = ~new_n16654_ & ~new_n16657_;
  assign new_n16659_ = ~ys__n18817 & ~ys__n37948;
  assign new_n16660_ = ys__n18817 & ys__n37948;
  assign new_n16661_ = ~new_n16659_ & ~new_n16660_;
  assign new_n16662_ = ~ys__n18819 & ~ys__n37949;
  assign new_n16663_ = ys__n18819 & ys__n37949;
  assign new_n16664_ = ~new_n16662_ & ~new_n16663_;
  assign new_n16665_ = ~new_n16661_ & ~new_n16664_;
  assign new_n16666_ = new_n16658_ & new_n16665_;
  assign new_n16667_ = ~ys__n18805 & ~ys__n37942;
  assign new_n16668_ = ys__n18805 & ys__n37942;
  assign new_n16669_ = ~new_n16667_ & ~new_n16668_;
  assign new_n16670_ = ~ys__n18807 & ~ys__n37943;
  assign new_n16671_ = ys__n18807 & ys__n37943;
  assign new_n16672_ = ~new_n16670_ & ~new_n16671_;
  assign new_n16673_ = ~new_n16669_ & ~new_n16672_;
  assign new_n16674_ = ~ys__n18809 & ~ys__n37944;
  assign new_n16675_ = ys__n18809 & ys__n37944;
  assign new_n16676_ = ~new_n16674_ & ~new_n16675_;
  assign new_n16677_ = ~ys__n18811 & ~ys__n37945;
  assign new_n16678_ = ys__n18811 & ys__n37945;
  assign new_n16679_ = ~new_n16677_ & ~new_n16678_;
  assign new_n16680_ = ~new_n16676_ & ~new_n16679_;
  assign new_n16681_ = new_n16673_ & new_n16680_;
  assign new_n16682_ = new_n16666_ & new_n16681_;
  assign new_n16683_ = new_n16651_ & new_n16682_;
  assign new_n16684_ = ~ys__n18781 & ~ys__n37930;
  assign new_n16685_ = ys__n18781 & ys__n37930;
  assign new_n16686_ = ~new_n16684_ & ~new_n16685_;
  assign new_n16687_ = ~ys__n18783 & ~ys__n37931;
  assign new_n16688_ = ys__n18783 & ys__n37931;
  assign new_n16689_ = ~new_n16687_ & ~new_n16688_;
  assign new_n16690_ = ~new_n16686_ & ~new_n16689_;
  assign new_n16691_ = ~ys__n18785 & ~ys__n37932;
  assign new_n16692_ = ys__n18785 & ys__n37932;
  assign new_n16693_ = ~new_n16691_ & ~new_n16692_;
  assign new_n16694_ = ~ys__n18787 & ~ys__n37933;
  assign new_n16695_ = ys__n18787 & ys__n37933;
  assign new_n16696_ = ~new_n16694_ & ~new_n16695_;
  assign new_n16697_ = ~new_n16693_ & ~new_n16696_;
  assign new_n16698_ = new_n16690_ & new_n16697_;
  assign new_n16699_ = ~ys__n18773 & ~ys__n37926;
  assign new_n16700_ = ys__n18773 & ys__n37926;
  assign new_n16701_ = ~new_n16699_ & ~new_n16700_;
  assign new_n16702_ = ~ys__n18775 & ~ys__n37927;
  assign new_n16703_ = ys__n18775 & ys__n37927;
  assign new_n16704_ = ~new_n16702_ & ~new_n16703_;
  assign new_n16705_ = ~new_n16701_ & ~new_n16704_;
  assign new_n16706_ = ~ys__n18777 & ~ys__n37928;
  assign new_n16707_ = ys__n18777 & ys__n37928;
  assign new_n16708_ = ~new_n16706_ & ~new_n16707_;
  assign new_n16709_ = ~ys__n18779 & ~ys__n37929;
  assign new_n16710_ = ys__n18779 & ys__n37929;
  assign new_n16711_ = ~new_n16709_ & ~new_n16710_;
  assign new_n16712_ = ~new_n16708_ & ~new_n16711_;
  assign new_n16713_ = new_n16705_ & new_n16712_;
  assign new_n16714_ = new_n16698_ & new_n16713_;
  assign new_n16715_ = ~ys__n18797 & ~ys__n37938;
  assign new_n16716_ = ys__n18797 & ys__n37938;
  assign new_n16717_ = ~new_n16715_ & ~new_n16716_;
  assign new_n16718_ = ~ys__n18799 & ~ys__n37939;
  assign new_n16719_ = ys__n18799 & ys__n37939;
  assign new_n16720_ = ~new_n16718_ & ~new_n16719_;
  assign new_n16721_ = ~new_n16717_ & ~new_n16720_;
  assign new_n16722_ = ~ys__n18801 & ~ys__n37940;
  assign new_n16723_ = ys__n18801 & ys__n37940;
  assign new_n16724_ = ~new_n16722_ & ~new_n16723_;
  assign new_n16725_ = ~ys__n18803 & ~ys__n37941;
  assign new_n16726_ = ys__n18803 & ys__n37941;
  assign new_n16727_ = ~new_n16725_ & ~new_n16726_;
  assign new_n16728_ = ~new_n16724_ & ~new_n16727_;
  assign new_n16729_ = new_n16721_ & new_n16728_;
  assign new_n16730_ = ~ys__n18789 & ~ys__n37934;
  assign new_n16731_ = ys__n18789 & ys__n37934;
  assign new_n16732_ = ~new_n16730_ & ~new_n16731_;
  assign new_n16733_ = ~ys__n18791 & ~ys__n37935;
  assign new_n16734_ = ys__n18791 & ys__n37935;
  assign new_n16735_ = ~new_n16733_ & ~new_n16734_;
  assign new_n16736_ = ~new_n16732_ & ~new_n16735_;
  assign new_n16737_ = ~ys__n18793 & ~ys__n37936;
  assign new_n16738_ = ys__n18793 & ys__n37936;
  assign new_n16739_ = ~new_n16737_ & ~new_n16738_;
  assign new_n16740_ = ~ys__n18795 & ~ys__n37937;
  assign new_n16741_ = ys__n18795 & ys__n37937;
  assign new_n16742_ = ~new_n16740_ & ~new_n16741_;
  assign new_n16743_ = ~new_n16739_ & ~new_n16742_;
  assign new_n16744_ = new_n16736_ & new_n16743_;
  assign new_n16745_ = new_n16729_ & new_n16744_;
  assign new_n16746_ = new_n16714_ & new_n16745_;
  assign new_n16747_ = new_n16683_ & new_n16746_;
  assign new_n16748_ = ~ys__n37751 & ~new_n16747_;
  assign new_n16749_ = ys__n856 & ~new_n16748_;
  assign new_n16750_ = ~new_n16636_ & ~new_n16749_;
  assign new_n16751_ = ~ys__n18821 & ~ys__n37922;
  assign new_n16752_ = ys__n18821 & ys__n37922;
  assign new_n16753_ = ~new_n16751_ & ~new_n16752_;
  assign new_n16754_ = ~ys__n18823 & ~ys__n37923;
  assign new_n16755_ = ys__n18823 & ys__n37923;
  assign new_n16756_ = ~new_n16754_ & ~new_n16755_;
  assign new_n16757_ = ~new_n16753_ & ~new_n16756_;
  assign new_n16758_ = ~ys__n18825 & ~ys__n37924;
  assign new_n16759_ = ys__n18825 & ys__n37924;
  assign new_n16760_ = ~new_n16758_ & ~new_n16759_;
  assign new_n16761_ = ~ys__n18827 & ~ys__n37925;
  assign new_n16762_ = ys__n18827 & ys__n37925;
  assign new_n16763_ = ~new_n16761_ & ~new_n16762_;
  assign new_n16764_ = ~new_n16760_ & ~new_n16763_;
  assign new_n16765_ = new_n16757_ & new_n16764_;
  assign new_n16766_ = ~ys__n18813 & ~ys__n37918;
  assign new_n16767_ = ys__n18813 & ys__n37918;
  assign new_n16768_ = ~new_n16766_ & ~new_n16767_;
  assign new_n16769_ = ~ys__n18815 & ~ys__n37919;
  assign new_n16770_ = ys__n18815 & ys__n37919;
  assign new_n16771_ = ~new_n16769_ & ~new_n16770_;
  assign new_n16772_ = ~new_n16768_ & ~new_n16771_;
  assign new_n16773_ = ~ys__n18817 & ~ys__n37920;
  assign new_n16774_ = ys__n18817 & ys__n37920;
  assign new_n16775_ = ~new_n16773_ & ~new_n16774_;
  assign new_n16776_ = ~ys__n18819 & ~ys__n37921;
  assign new_n16777_ = ys__n18819 & ys__n37921;
  assign new_n16778_ = ~new_n16776_ & ~new_n16777_;
  assign new_n16779_ = ~new_n16775_ & ~new_n16778_;
  assign new_n16780_ = new_n16772_ & new_n16779_;
  assign new_n16781_ = ~ys__n18805 & ~ys__n37914;
  assign new_n16782_ = ys__n18805 & ys__n37914;
  assign new_n16783_ = ~new_n16781_ & ~new_n16782_;
  assign new_n16784_ = ~ys__n18807 & ~ys__n37915;
  assign new_n16785_ = ys__n18807 & ys__n37915;
  assign new_n16786_ = ~new_n16784_ & ~new_n16785_;
  assign new_n16787_ = ~new_n16783_ & ~new_n16786_;
  assign new_n16788_ = ~ys__n18809 & ~ys__n37916;
  assign new_n16789_ = ys__n18809 & ys__n37916;
  assign new_n16790_ = ~new_n16788_ & ~new_n16789_;
  assign new_n16791_ = ~ys__n18811 & ~ys__n37917;
  assign new_n16792_ = ys__n18811 & ys__n37917;
  assign new_n16793_ = ~new_n16791_ & ~new_n16792_;
  assign new_n16794_ = ~new_n16790_ & ~new_n16793_;
  assign new_n16795_ = new_n16787_ & new_n16794_;
  assign new_n16796_ = new_n16780_ & new_n16795_;
  assign new_n16797_ = new_n16765_ & new_n16796_;
  assign new_n16798_ = ~ys__n18781 & ~ys__n37902;
  assign new_n16799_ = ys__n18781 & ys__n37902;
  assign new_n16800_ = ~new_n16798_ & ~new_n16799_;
  assign new_n16801_ = ~ys__n18783 & ~ys__n37903;
  assign new_n16802_ = ys__n18783 & ys__n37903;
  assign new_n16803_ = ~new_n16801_ & ~new_n16802_;
  assign new_n16804_ = ~new_n16800_ & ~new_n16803_;
  assign new_n16805_ = ~ys__n18785 & ~ys__n37904;
  assign new_n16806_ = ys__n18785 & ys__n37904;
  assign new_n16807_ = ~new_n16805_ & ~new_n16806_;
  assign new_n16808_ = ~ys__n18787 & ~ys__n37905;
  assign new_n16809_ = ys__n18787 & ys__n37905;
  assign new_n16810_ = ~new_n16808_ & ~new_n16809_;
  assign new_n16811_ = ~new_n16807_ & ~new_n16810_;
  assign new_n16812_ = new_n16804_ & new_n16811_;
  assign new_n16813_ = ~ys__n18773 & ~ys__n37898;
  assign new_n16814_ = ys__n18773 & ys__n37898;
  assign new_n16815_ = ~new_n16813_ & ~new_n16814_;
  assign new_n16816_ = ~ys__n18775 & ~ys__n37899;
  assign new_n16817_ = ys__n18775 & ys__n37899;
  assign new_n16818_ = ~new_n16816_ & ~new_n16817_;
  assign new_n16819_ = ~new_n16815_ & ~new_n16818_;
  assign new_n16820_ = ~ys__n18777 & ~ys__n37900;
  assign new_n16821_ = ys__n18777 & ys__n37900;
  assign new_n16822_ = ~new_n16820_ & ~new_n16821_;
  assign new_n16823_ = ~ys__n18779 & ~ys__n37901;
  assign new_n16824_ = ys__n18779 & ys__n37901;
  assign new_n16825_ = ~new_n16823_ & ~new_n16824_;
  assign new_n16826_ = ~new_n16822_ & ~new_n16825_;
  assign new_n16827_ = new_n16819_ & new_n16826_;
  assign new_n16828_ = new_n16812_ & new_n16827_;
  assign new_n16829_ = ~ys__n18797 & ~ys__n37910;
  assign new_n16830_ = ys__n18797 & ys__n37910;
  assign new_n16831_ = ~new_n16829_ & ~new_n16830_;
  assign new_n16832_ = ~ys__n18799 & ~ys__n37911;
  assign new_n16833_ = ys__n18799 & ys__n37911;
  assign new_n16834_ = ~new_n16832_ & ~new_n16833_;
  assign new_n16835_ = ~new_n16831_ & ~new_n16834_;
  assign new_n16836_ = ~ys__n18801 & ~ys__n37912;
  assign new_n16837_ = ys__n18801 & ys__n37912;
  assign new_n16838_ = ~new_n16836_ & ~new_n16837_;
  assign new_n16839_ = ~ys__n18803 & ~ys__n37913;
  assign new_n16840_ = ys__n18803 & ys__n37913;
  assign new_n16841_ = ~new_n16839_ & ~new_n16840_;
  assign new_n16842_ = ~new_n16838_ & ~new_n16841_;
  assign new_n16843_ = new_n16835_ & new_n16842_;
  assign new_n16844_ = ~ys__n18789 & ~ys__n37906;
  assign new_n16845_ = ys__n18789 & ys__n37906;
  assign new_n16846_ = ~new_n16844_ & ~new_n16845_;
  assign new_n16847_ = ~ys__n18791 & ~ys__n37907;
  assign new_n16848_ = ys__n18791 & ys__n37907;
  assign new_n16849_ = ~new_n16847_ & ~new_n16848_;
  assign new_n16850_ = ~new_n16846_ & ~new_n16849_;
  assign new_n16851_ = ~ys__n18793 & ~ys__n37908;
  assign new_n16852_ = ys__n18793 & ys__n37908;
  assign new_n16853_ = ~new_n16851_ & ~new_n16852_;
  assign new_n16854_ = ~ys__n18795 & ~ys__n37909;
  assign new_n16855_ = ys__n18795 & ys__n37909;
  assign new_n16856_ = ~new_n16854_ & ~new_n16855_;
  assign new_n16857_ = ~new_n16853_ & ~new_n16856_;
  assign new_n16858_ = new_n16850_ & new_n16857_;
  assign new_n16859_ = new_n16843_ & new_n16858_;
  assign new_n16860_ = new_n16828_ & new_n16859_;
  assign new_n16861_ = new_n16797_ & new_n16860_;
  assign new_n16862_ = ~ys__n37752 & ~new_n16861_;
  assign new_n16863_ = ys__n854 & ~new_n16862_;
  assign new_n16864_ = ~ys__n18821 & ~ys__n37894;
  assign new_n16865_ = ys__n18821 & ys__n37894;
  assign new_n16866_ = ~new_n16864_ & ~new_n16865_;
  assign new_n16867_ = ~ys__n18823 & ~ys__n37895;
  assign new_n16868_ = ys__n18823 & ys__n37895;
  assign new_n16869_ = ~new_n16867_ & ~new_n16868_;
  assign new_n16870_ = ~new_n16866_ & ~new_n16869_;
  assign new_n16871_ = ~ys__n18825 & ~ys__n37896;
  assign new_n16872_ = ys__n18825 & ys__n37896;
  assign new_n16873_ = ~new_n16871_ & ~new_n16872_;
  assign new_n16874_ = ~ys__n18827 & ~ys__n37897;
  assign new_n16875_ = ys__n18827 & ys__n37897;
  assign new_n16876_ = ~new_n16874_ & ~new_n16875_;
  assign new_n16877_ = ~new_n16873_ & ~new_n16876_;
  assign new_n16878_ = new_n16870_ & new_n16877_;
  assign new_n16879_ = ~ys__n18813 & ~ys__n37890;
  assign new_n16880_ = ys__n18813 & ys__n37890;
  assign new_n16881_ = ~new_n16879_ & ~new_n16880_;
  assign new_n16882_ = ~ys__n18815 & ~ys__n37891;
  assign new_n16883_ = ys__n18815 & ys__n37891;
  assign new_n16884_ = ~new_n16882_ & ~new_n16883_;
  assign new_n16885_ = ~new_n16881_ & ~new_n16884_;
  assign new_n16886_ = ~ys__n18817 & ~ys__n37892;
  assign new_n16887_ = ys__n18817 & ys__n37892;
  assign new_n16888_ = ~new_n16886_ & ~new_n16887_;
  assign new_n16889_ = ~ys__n18819 & ~ys__n37893;
  assign new_n16890_ = ys__n18819 & ys__n37893;
  assign new_n16891_ = ~new_n16889_ & ~new_n16890_;
  assign new_n16892_ = ~new_n16888_ & ~new_n16891_;
  assign new_n16893_ = new_n16885_ & new_n16892_;
  assign new_n16894_ = ~ys__n18805 & ~ys__n37886;
  assign new_n16895_ = ys__n18805 & ys__n37886;
  assign new_n16896_ = ~new_n16894_ & ~new_n16895_;
  assign new_n16897_ = ~ys__n18807 & ~ys__n37887;
  assign new_n16898_ = ys__n18807 & ys__n37887;
  assign new_n16899_ = ~new_n16897_ & ~new_n16898_;
  assign new_n16900_ = ~new_n16896_ & ~new_n16899_;
  assign new_n16901_ = ~ys__n18809 & ~ys__n37888;
  assign new_n16902_ = ys__n18809 & ys__n37888;
  assign new_n16903_ = ~new_n16901_ & ~new_n16902_;
  assign new_n16904_ = ~ys__n18811 & ~ys__n37889;
  assign new_n16905_ = ys__n18811 & ys__n37889;
  assign new_n16906_ = ~new_n16904_ & ~new_n16905_;
  assign new_n16907_ = ~new_n16903_ & ~new_n16906_;
  assign new_n16908_ = new_n16900_ & new_n16907_;
  assign new_n16909_ = new_n16893_ & new_n16908_;
  assign new_n16910_ = new_n16878_ & new_n16909_;
  assign new_n16911_ = ~ys__n18781 & ~ys__n37874;
  assign new_n16912_ = ys__n18781 & ys__n37874;
  assign new_n16913_ = ~new_n16911_ & ~new_n16912_;
  assign new_n16914_ = ~ys__n18783 & ~ys__n37875;
  assign new_n16915_ = ys__n18783 & ys__n37875;
  assign new_n16916_ = ~new_n16914_ & ~new_n16915_;
  assign new_n16917_ = ~new_n16913_ & ~new_n16916_;
  assign new_n16918_ = ~ys__n18785 & ~ys__n37876;
  assign new_n16919_ = ys__n18785 & ys__n37876;
  assign new_n16920_ = ~new_n16918_ & ~new_n16919_;
  assign new_n16921_ = ~ys__n18787 & ~ys__n37877;
  assign new_n16922_ = ys__n18787 & ys__n37877;
  assign new_n16923_ = ~new_n16921_ & ~new_n16922_;
  assign new_n16924_ = ~new_n16920_ & ~new_n16923_;
  assign new_n16925_ = new_n16917_ & new_n16924_;
  assign new_n16926_ = ~ys__n18773 & ~ys__n37870;
  assign new_n16927_ = ys__n18773 & ys__n37870;
  assign new_n16928_ = ~new_n16926_ & ~new_n16927_;
  assign new_n16929_ = ~ys__n18775 & ~ys__n37871;
  assign new_n16930_ = ys__n18775 & ys__n37871;
  assign new_n16931_ = ~new_n16929_ & ~new_n16930_;
  assign new_n16932_ = ~new_n16928_ & ~new_n16931_;
  assign new_n16933_ = ~ys__n18777 & ~ys__n37872;
  assign new_n16934_ = ys__n18777 & ys__n37872;
  assign new_n16935_ = ~new_n16933_ & ~new_n16934_;
  assign new_n16936_ = ~ys__n18779 & ~ys__n37873;
  assign new_n16937_ = ys__n18779 & ys__n37873;
  assign new_n16938_ = ~new_n16936_ & ~new_n16937_;
  assign new_n16939_ = ~new_n16935_ & ~new_n16938_;
  assign new_n16940_ = new_n16932_ & new_n16939_;
  assign new_n16941_ = new_n16925_ & new_n16940_;
  assign new_n16942_ = ~ys__n18797 & ~ys__n37882;
  assign new_n16943_ = ys__n18797 & ys__n37882;
  assign new_n16944_ = ~new_n16942_ & ~new_n16943_;
  assign new_n16945_ = ~ys__n18799 & ~ys__n37883;
  assign new_n16946_ = ys__n18799 & ys__n37883;
  assign new_n16947_ = ~new_n16945_ & ~new_n16946_;
  assign new_n16948_ = ~new_n16944_ & ~new_n16947_;
  assign new_n16949_ = ~ys__n18801 & ~ys__n37884;
  assign new_n16950_ = ys__n18801 & ys__n37884;
  assign new_n16951_ = ~new_n16949_ & ~new_n16950_;
  assign new_n16952_ = ~ys__n18803 & ~ys__n37885;
  assign new_n16953_ = ys__n18803 & ys__n37885;
  assign new_n16954_ = ~new_n16952_ & ~new_n16953_;
  assign new_n16955_ = ~new_n16951_ & ~new_n16954_;
  assign new_n16956_ = new_n16948_ & new_n16955_;
  assign new_n16957_ = ~ys__n18789 & ~ys__n37878;
  assign new_n16958_ = ys__n18789 & ys__n37878;
  assign new_n16959_ = ~new_n16957_ & ~new_n16958_;
  assign new_n16960_ = ~ys__n18791 & ~ys__n37879;
  assign new_n16961_ = ys__n18791 & ys__n37879;
  assign new_n16962_ = ~new_n16960_ & ~new_n16961_;
  assign new_n16963_ = ~new_n16959_ & ~new_n16962_;
  assign new_n16964_ = ~ys__n18793 & ~ys__n37880;
  assign new_n16965_ = ys__n18793 & ys__n37880;
  assign new_n16966_ = ~new_n16964_ & ~new_n16965_;
  assign new_n16967_ = ~ys__n18795 & ~ys__n37881;
  assign new_n16968_ = ys__n18795 & ys__n37881;
  assign new_n16969_ = ~new_n16967_ & ~new_n16968_;
  assign new_n16970_ = ~new_n16966_ & ~new_n16969_;
  assign new_n16971_ = new_n16963_ & new_n16970_;
  assign new_n16972_ = new_n16956_ & new_n16971_;
  assign new_n16973_ = new_n16941_ & new_n16972_;
  assign new_n16974_ = new_n16910_ & new_n16973_;
  assign new_n16975_ = ~ys__n37753 & ~new_n16974_;
  assign new_n16976_ = ys__n852 & ~new_n16975_;
  assign new_n16977_ = ~new_n16863_ & ~new_n16976_;
  assign new_n16978_ = new_n16750_ & new_n16977_;
  assign new_n16979_ = new_n16523_ & new_n16978_;
  assign ys__n3249 = ~new_n16068_ | ~new_n16979_;
  assign new_n16981_ = ys__n18978 & ys__n18287;
  assign new_n16982_ = ~ys__n18284 & new_n16981_;
  assign new_n16983_ = ys__n24659 & ~ys__n4764;
  assign new_n16984_ = ys__n24660 & ys__n4764;
  assign ys__n18808 = new_n16983_ | new_n16984_;
  assign new_n16986_ = ~ys__n18071 & ys__n18808;
  assign new_n16987_ = ys__n18071 & ys__n18809;
  assign new_n16988_ = ~new_n16986_ & ~new_n16987_;
  assign new_n16989_ = ~new_n12256_ & ~new_n16988_;
  assign new_n16990_ = ys__n24660 & ~ys__n24675;
  assign new_n16991_ = ys__n24675 & ys__n24701;
  assign ys__n18720 = new_n16990_ | new_n16991_;
  assign new_n16993_ = new_n12256_ & ys__n18720;
  assign ys__n18721 = new_n16989_ | new_n16993_;
  assign new_n16995_ = ys__n18284 & ys__n18721;
  assign new_n16996_ = ~new_n16982_ & ~new_n16995_;
  assign new_n16997_ = ~ys__n18281 & ~new_n16996_;
  assign new_n16998_ = ys__n18622 & ~new_n12259_;
  assign new_n16999_ = ys__n18623 & new_n12259_;
  assign ys__n18624 = new_n16998_ | new_n16999_;
  assign new_n17001_ = ys__n18281 & ys__n18624;
  assign new_n17002_ = ~new_n16997_ & ~new_n17001_;
  assign new_n17003_ = ~ys__n18278 & ~new_n17002_;
  assign new_n17004_ = ys__n18873 & ys__n18278;
  assign ys__n3250 = new_n17003_ | new_n17004_;
  assign new_n17006_ = ys__n18979 & ys__n18287;
  assign new_n17007_ = ~ys__n18284 & new_n17006_;
  assign new_n17008_ = ys__n24661 & ~ys__n4764;
  assign new_n17009_ = ys__n24662 & ys__n4764;
  assign ys__n18810 = new_n17008_ | new_n17009_;
  assign new_n17011_ = ~ys__n18071 & ys__n18810;
  assign new_n17012_ = ys__n18071 & ys__n18811;
  assign new_n17013_ = ~new_n17011_ & ~new_n17012_;
  assign new_n17014_ = ~new_n12256_ & ~new_n17013_;
  assign new_n17015_ = ys__n24662 & ~ys__n24675;
  assign new_n17016_ = ys__n24675 & ys__n24702;
  assign ys__n18723 = new_n17015_ | new_n17016_;
  assign new_n17018_ = new_n12256_ & ys__n18723;
  assign ys__n18724 = new_n17014_ | new_n17018_;
  assign new_n17020_ = ys__n18284 & ys__n18724;
  assign new_n17021_ = ~new_n17007_ & ~new_n17020_;
  assign new_n17022_ = ~ys__n18281 & ~new_n17021_;
  assign new_n17023_ = ys__n18625 & ~new_n12259_;
  assign new_n17024_ = ys__n18626 & new_n12259_;
  assign ys__n18627 = new_n17023_ | new_n17024_;
  assign new_n17026_ = ys__n18281 & ys__n18627;
  assign new_n17027_ = ~new_n17022_ & ~new_n17026_;
  assign new_n17028_ = ~ys__n18278 & ~new_n17027_;
  assign new_n17029_ = ys__n18875 & ys__n18278;
  assign ys__n3252 = new_n17028_ | new_n17029_;
  assign new_n17031_ = ~ys__n846 & new_n12181_;
  assign new_n17032_ = new_n13357_ & new_n17031_;
  assign ys__n4189 = ~new_n13361_ | ~new_n17032_;
  assign new_n17034_ = ~ys__n776 & ~ys__n4168;
  assign new_n17035_ = ~ys__n604 & ~ys__n778;
  assign new_n17036_ = new_n17034_ & new_n17035_;
  assign new_n17037_ = ~ys__n698 & ~ys__n768;
  assign new_n17038_ = new_n15064_ & new_n17037_;
  assign new_n17039_ = new_n17036_ & new_n17038_;
  assign new_n17040_ = new_n15067_ & new_n15068_;
  assign new_n17041_ = ys__n772 & new_n17040_;
  assign new_n17042_ = new_n17039_ & new_n17041_;
  assign new_n17043_ = ~ys__n598 & ys__n774;
  assign new_n17044_ = new_n17039_ & new_n17043_;
  assign new_n17045_ = ys__n770 & ~ys__n784;
  assign new_n17046_ = new_n15067_ & new_n17045_;
  assign new_n17047_ = new_n17039_ & new_n17046_;
  assign new_n17048_ = ~new_n17044_ & ~new_n17047_;
  assign new_n17049_ = ~new_n17042_ & new_n17048_;
  assign new_n17050_ = ~ys__n772 & ~ys__n780;
  assign new_n17051_ = ys__n782 & new_n17050_;
  assign new_n17052_ = new_n17040_ & new_n17051_;
  assign new_n17053_ = new_n17039_ & new_n17052_;
  assign new_n17054_ = ~ys__n772 & ys__n780;
  assign new_n17055_ = new_n17040_ & new_n17054_;
  assign new_n17056_ = new_n17039_ & new_n17055_;
  assign new_n17057_ = ~new_n17053_ & ~new_n17056_;
  assign new_n17058_ = ~ys__n782 & ~ys__n2644;
  assign new_n17059_ = new_n17050_ & new_n17058_;
  assign new_n17060_ = new_n17040_ & new_n17059_;
  assign new_n17061_ = new_n17039_ & new_n17060_;
  assign new_n17062_ = ys__n598 & new_n17039_;
  assign new_n17063_ = ~new_n17061_ & ~new_n17062_;
  assign new_n17064_ = new_n17057_ & new_n17063_;
  assign new_n17065_ = ys__n602 & new_n17036_;
  assign new_n17066_ = ys__n698 & new_n15064_;
  assign new_n17067_ = new_n17036_ & new_n17066_;
  assign new_n17068_ = ~new_n17065_ & ~new_n17067_;
  assign new_n17069_ = ys__n600 & ~ys__n602;
  assign new_n17070_ = new_n17036_ & new_n17069_;
  assign new_n17071_ = ~ys__n698 & ys__n768;
  assign new_n17072_ = new_n15064_ & new_n17071_;
  assign new_n17073_ = new_n17036_ & new_n17072_;
  assign new_n17074_ = ~new_n17070_ & ~new_n17073_;
  assign new_n17075_ = new_n17068_ & new_n17074_;
  assign new_n17076_ = ys__n784 & new_n15067_;
  assign new_n17077_ = new_n17039_ & new_n17076_;
  assign new_n17078_ = ys__n604 & new_n17034_;
  assign new_n17079_ = ~ys__n604 & ys__n778;
  assign new_n17080_ = new_n17034_ & new_n17079_;
  assign new_n17081_ = ys__n776 & ~ys__n4168;
  assign new_n17082_ = ~new_n17080_ & ~new_n17081_;
  assign new_n17083_ = ~new_n17078_ & new_n17082_;
  assign new_n17084_ = ~new_n17077_ & new_n17083_;
  assign new_n17085_ = new_n17075_ & new_n17084_;
  assign new_n17086_ = new_n17064_ & new_n17085_;
  assign ys__n4320 = new_n17049_ & new_n17086_;
  assign ys__n4414 = ~ys__n18271 & ~new_n12264_;
  assign ys__n4521 = ~ys__n740 | new_n13322_;
  assign new_n17090_ = new_n12327_ & ~new_n12364_;
  assign new_n17091_ = ~new_n12337_ & ~new_n12339_;
  assign new_n17092_ = ~ys__n530 & ~ys__n752;
  assign new_n17093_ = ~ys__n526 & ys__n528;
  assign new_n17094_ = ys__n522 & ~ys__n524;
  assign new_n17095_ = new_n17093_ & new_n17094_;
  assign new_n17096_ = new_n17092_ & new_n17095_;
  assign new_n17097_ = new_n11766_ & new_n11791_;
  assign new_n17098_ = new_n17096_ & new_n17097_;
  assign new_n17099_ = new_n17091_ & ~new_n17098_;
  assign new_n17100_ = ~new_n17090_ & new_n17099_;
  assign new_n17101_ = ~new_n12327_ & ~new_n17097_;
  assign new_n17102_ = new_n17091_ & new_n17101_;
  assign new_n17103_ = ~ys__n28243 & ~new_n17102_;
  assign new_n17104_ = ~new_n17100_ & new_n17103_;
  assign new_n17105_ = new_n12384_ & new_n12394_;
  assign new_n17106_ = ys__n736 & ~ys__n752;
  assign new_n17107_ = ~ys__n4488 & ~ys__n23730;
  assign new_n17108_ = new_n17106_ & new_n17107_;
  assign new_n17109_ = new_n17105_ & new_n17108_;
  assign new_n17110_ = ~ys__n23730 & ~new_n17109_;
  assign new_n17111_ = ys__n28243 & ~new_n17110_;
  assign new_n17112_ = ~new_n17104_ & ~new_n17111_;
  assign ys__n4588 = ~ys__n738 & ~new_n17112_;
  assign new_n17114_ = ~ys__n23627 & ys__n23629;
  assign new_n17115_ = ~new_n12309_ & new_n17114_;
  assign new_n17116_ = ys__n22882 & new_n12309_;
  assign new_n17117_ = ~new_n17115_ & ~new_n17116_;
  assign new_n17118_ = ~new_n12314_ & ~new_n17117_;
  assign new_n17119_ = ys__n23330 & new_n12314_;
  assign new_n17120_ = ~new_n17118_ & ~new_n17119_;
  assign new_n17121_ = ~new_n12320_ & ~new_n17120_;
  assign new_n17122_ = ys__n424 & new_n12320_;
  assign new_n17123_ = ~new_n17121_ & ~new_n17122_;
  assign new_n17124_ = ~new_n12404_ & ~new_n17123_;
  assign new_n17125_ = ys__n424 & ~new_n12426_;
  assign new_n17126_ = ~ys__n424 & new_n12798_;
  assign new_n17127_ = ys__n424 & ~new_n12798_;
  assign new_n17128_ = ~new_n17126_ & ~new_n17127_;
  assign new_n17129_ = new_n12426_ & ~new_n17128_;
  assign ys__n23541 = new_n17125_ | new_n17129_;
  assign new_n17131_ = new_n12404_ & ys__n23541;
  assign new_n17132_ = ~new_n17124_ & ~new_n17131_;
  assign new_n17133_ = new_n12458_ & ~new_n17132_;
  assign new_n17134_ = ys__n424 & ~new_n12458_;
  assign new_n17135_ = ~new_n17133_ & ~new_n17134_;
  assign new_n17136_ = ~new_n12477_ & ~new_n17135_;
  assign new_n17137_ = ys__n424 & ~new_n12703_;
  assign new_n17138_ = ~ys__n450 & ~new_n12733_;
  assign new_n17139_ = ~ys__n450 & ~new_n17138_;
  assign new_n17140_ = ys__n424 & ~new_n17139_;
  assign new_n17141_ = ~ys__n424 & new_n17139_;
  assign new_n17142_ = ~new_n17140_ & ~new_n17141_;
  assign new_n17143_ = new_n12737_ & ~new_n17142_;
  assign new_n17144_ = ys__n450 & new_n12749_;
  assign new_n17145_ = ~ys__n424 & new_n17144_;
  assign new_n17146_ = ys__n424 & ~new_n17144_;
  assign new_n17147_ = ~new_n17145_ & ~new_n17146_;
  assign new_n17148_ = new_n12753_ & ~new_n17147_;
  assign new_n17149_ = ~new_n17143_ & ~new_n17148_;
  assign new_n17150_ = ~new_n17137_ & new_n17149_;
  assign new_n17151_ = new_n12759_ & ~new_n17150_;
  assign new_n17152_ = ~new_n17136_ & ~new_n17151_;
  assign new_n17153_ = new_n12763_ & ~new_n17152_;
  assign new_n17154_ = ys__n935 & ys__n23629;
  assign new_n17155_ = new_n12762_ & new_n17154_;
  assign new_n17156_ = ys__n47691 & new_n12768_;
  assign new_n17157_ = ~new_n17155_ & ~new_n17156_;
  assign new_n17158_ = ~new_n17153_ & new_n17157_;
  assign new_n17159_ = new_n12774_ & ~new_n17158_;
  assign new_n17160_ = new_n12776_ & ~new_n17152_;
  assign new_n17161_ = ys__n47691 & new_n12778_;
  assign new_n17162_ = ~new_n17155_ & ~new_n17161_;
  assign new_n17163_ = ~new_n17160_ & new_n17162_;
  assign new_n17164_ = new_n12784_ & ~new_n17163_;
  assign ys__n4615 = new_n17159_ | new_n17164_;
  assign new_n17166_ = ~ys__n35098 & ~ys__n35423;
  assign new_n17167_ = ys__n35098 & ys__n35423;
  assign new_n17168_ = ~new_n17166_ & ~new_n17167_;
  assign new_n17169_ = ~ys__n35096 & ~ys__n35421;
  assign new_n17170_ = ys__n35096 & ys__n35421;
  assign new_n17171_ = ~new_n17169_ & ~new_n17170_;
  assign new_n17172_ = ~new_n17168_ & ~new_n17171_;
  assign new_n17173_ = ~ys__n35094 & ~ys__n35419;
  assign new_n17174_ = ys__n35094 & ys__n35419;
  assign new_n17175_ = ~new_n17173_ & ~new_n17174_;
  assign new_n17176_ = ~ys__n35092 & ~ys__n35417;
  assign new_n17177_ = ys__n35092 & ys__n35417;
  assign new_n17178_ = ~new_n17176_ & ~new_n17177_;
  assign new_n17179_ = ~new_n17175_ & ~new_n17178_;
  assign new_n17180_ = new_n17172_ & new_n17179_;
  assign new_n17181_ = ~ys__n35090 & ~ys__n35415;
  assign new_n17182_ = ys__n35090 & ys__n35415;
  assign new_n17183_ = ~new_n17181_ & ~new_n17182_;
  assign new_n17184_ = ~ys__n35088 & ~ys__n35413;
  assign new_n17185_ = ys__n35088 & ys__n35413;
  assign new_n17186_ = ~new_n17184_ & ~new_n17185_;
  assign new_n17187_ = ~new_n17183_ & ~new_n17186_;
  assign new_n17188_ = ~ys__n35086 & ~ys__n48335;
  assign new_n17189_ = ys__n35086 & ys__n48335;
  assign new_n17190_ = ~new_n17188_ & ~new_n17189_;
  assign new_n17191_ = ~ys__n35084 & ~ys__n48334;
  assign new_n17192_ = ys__n35084 & ys__n48334;
  assign new_n17193_ = ~new_n17191_ & ~new_n17192_;
  assign new_n17194_ = ~new_n17190_ & ~new_n17193_;
  assign new_n17195_ = new_n17187_ & new_n17194_;
  assign new_n17196_ = ~ys__n35082 & ~ys__n48333;
  assign new_n17197_ = ys__n35082 & ys__n48333;
  assign new_n17198_ = ~new_n17196_ & ~new_n17197_;
  assign new_n17199_ = ~ys__n35080 & ~ys__n48332;
  assign new_n17200_ = ys__n35080 & ys__n48332;
  assign new_n17201_ = ~new_n17199_ & ~new_n17200_;
  assign new_n17202_ = ~new_n17198_ & ~new_n17201_;
  assign new_n17203_ = ~ys__n35078 & ys__n48331;
  assign new_n17204_ = ~ys__n35078 & ~ys__n48331;
  assign new_n17205_ = ys__n35078 & ys__n48331;
  assign new_n17206_ = ~new_n17204_ & ~new_n17205_;
  assign new_n17207_ = ~ys__n35076 & ys__n48330;
  assign new_n17208_ = ~ys__n35076 & ~ys__n48330;
  assign new_n17209_ = ys__n35076 & ys__n48330;
  assign new_n17210_ = ~new_n17208_ & ~new_n17209_;
  assign new_n17211_ = ~new_n17207_ & new_n17210_;
  assign new_n17212_ = ~new_n17206_ & ~new_n17211_;
  assign new_n17213_ = ~new_n17203_ & ~new_n17212_;
  assign new_n17214_ = new_n17202_ & ~new_n17213_;
  assign new_n17215_ = ~ys__n35082 & ys__n48333;
  assign new_n17216_ = ~ys__n35080 & ys__n48332;
  assign new_n17217_ = ~new_n17198_ & new_n17216_;
  assign new_n17218_ = ~new_n17215_ & ~new_n17217_;
  assign new_n17219_ = ~new_n17214_ & new_n17218_;
  assign new_n17220_ = new_n17195_ & ~new_n17219_;
  assign new_n17221_ = ~ys__n35086 & ys__n48335;
  assign new_n17222_ = ~ys__n35084 & ys__n48334;
  assign new_n17223_ = ~new_n17190_ & new_n17222_;
  assign new_n17224_ = ~new_n17221_ & ~new_n17223_;
  assign new_n17225_ = new_n17187_ & ~new_n17224_;
  assign new_n17226_ = ~ys__n35090 & ys__n35415;
  assign new_n17227_ = ~ys__n35088 & ys__n35413;
  assign new_n17228_ = ~new_n17183_ & new_n17227_;
  assign new_n17229_ = ~new_n17226_ & ~new_n17228_;
  assign new_n17230_ = ~new_n17225_ & new_n17229_;
  assign new_n17231_ = ~new_n17220_ & new_n17230_;
  assign new_n17232_ = new_n17180_ & ~new_n17231_;
  assign new_n17233_ = ~ys__n35094 & ys__n35419;
  assign new_n17234_ = ~ys__n35092 & ys__n35417;
  assign new_n17235_ = ~new_n17175_ & new_n17234_;
  assign new_n17236_ = ~new_n17233_ & ~new_n17235_;
  assign new_n17237_ = new_n17172_ & ~new_n17236_;
  assign new_n17238_ = ~ys__n35098 & ys__n35423;
  assign new_n17239_ = ~ys__n35096 & ys__n35421;
  assign new_n17240_ = ~new_n17168_ & new_n17239_;
  assign new_n17241_ = ~new_n17238_ & ~new_n17240_;
  assign new_n17242_ = ~new_n17237_ & new_n17241_;
  assign new_n17243_ = ~new_n17232_ & new_n17242_;
  assign new_n17244_ = ~new_n17206_ & ~new_n17210_;
  assign new_n17245_ = new_n17202_ & new_n17244_;
  assign new_n17246_ = new_n17180_ & new_n17245_;
  assign new_n17247_ = new_n17195_ & new_n17246_;
  assign new_n17248_ = ~new_n17243_ & ~new_n17247_;
  assign new_n17249_ = ~ys__n33218 & ~ys__n35419;
  assign new_n17250_ = ys__n33218 & ys__n35419;
  assign new_n17251_ = ~new_n17249_ & ~new_n17250_;
  assign new_n17252_ = ~ys__n33216 & ~ys__n35417;
  assign new_n17253_ = ys__n33216 & ys__n35417;
  assign new_n17254_ = ~new_n17252_ & ~new_n17253_;
  assign new_n17255_ = ~new_n17251_ & ~new_n17254_;
  assign new_n17256_ = ~ys__n33222 & ~ys__n35423;
  assign new_n17257_ = ys__n33222 & ys__n35423;
  assign new_n17258_ = ~new_n17256_ & ~new_n17257_;
  assign new_n17259_ = ~ys__n33220 & ~ys__n35421;
  assign new_n17260_ = ys__n33220 & ys__n35421;
  assign new_n17261_ = ~new_n17259_ & ~new_n17260_;
  assign new_n17262_ = ~new_n17258_ & ~new_n17261_;
  assign new_n17263_ = ~ys__n33214 & ~ys__n35415;
  assign new_n17264_ = ys__n33214 & ys__n35415;
  assign new_n17265_ = ~new_n17263_ & ~new_n17264_;
  assign new_n17266_ = ~ys__n33212 & ~ys__n35413;
  assign new_n17267_ = ys__n33212 & ys__n35413;
  assign new_n17268_ = ~new_n17266_ & ~new_n17267_;
  assign new_n17269_ = ~new_n17265_ & ~new_n17268_;
  assign new_n17270_ = new_n17262_ & new_n17269_;
  assign new_n17271_ = new_n17255_ & new_n17270_;
  assign new_n17272_ = ~ys__n33214 & ys__n35415;
  assign new_n17273_ = ~ys__n33212 & ys__n35413;
  assign new_n17274_ = new_n17268_ & ~new_n17273_;
  assign new_n17275_ = ~new_n17265_ & ~new_n17274_;
  assign new_n17276_ = ~new_n17272_ & ~new_n17275_;
  assign new_n17277_ = new_n17255_ & ~new_n17276_;
  assign new_n17278_ = ~ys__n33218 & ys__n35419;
  assign new_n17279_ = ~ys__n33216 & ys__n35417;
  assign new_n17280_ = ~new_n17251_ & new_n17279_;
  assign new_n17281_ = ~new_n17278_ & ~new_n17280_;
  assign new_n17282_ = ~new_n17277_ & new_n17281_;
  assign new_n17283_ = new_n17262_ & ~new_n17282_;
  assign new_n17284_ = ~ys__n33222 & ys__n35423;
  assign new_n17285_ = ~ys__n33220 & ys__n35421;
  assign new_n17286_ = ~new_n17258_ & new_n17285_;
  assign new_n17287_ = ~new_n17284_ & ~new_n17286_;
  assign new_n17288_ = ~new_n17283_ & new_n17287_;
  assign new_n17289_ = ~new_n17271_ & ~new_n17288_;
  assign new_n17290_ = ~new_n17271_ & ~new_n17289_;
  assign new_n17291_ = ~ys__n38847 & ys__n38848;
  assign new_n17292_ = ys__n38847 & ~ys__n38848;
  assign new_n17293_ = ~new_n17291_ & ~new_n17292_;
  assign new_n17294_ = ~ys__n38849 & ys__n38850;
  assign new_n17295_ = ys__n38849 & ~ys__n38850;
  assign new_n17296_ = ~new_n17294_ & ~new_n17295_;
  assign new_n17297_ = new_n17293_ & new_n17296_;
  assign new_n17298_ = ~ys__n38843 & ys__n38844;
  assign new_n17299_ = ys__n38843 & ~ys__n38844;
  assign new_n17300_ = ~new_n17298_ & ~new_n17299_;
  assign new_n17301_ = ~ys__n38845 & ys__n38846;
  assign new_n17302_ = ys__n38845 & ~ys__n38846;
  assign new_n17303_ = ~new_n17301_ & ~new_n17302_;
  assign new_n17304_ = new_n17300_ & new_n17303_;
  assign new_n17305_ = new_n17297_ & new_n17304_;
  assign new_n17306_ = ~ys__n38855 & ys__n38856;
  assign new_n17307_ = ys__n38855 & ~ys__n38856;
  assign new_n17308_ = ~new_n17306_ & ~new_n17307_;
  assign new_n17309_ = ~ys__n38857 & ys__n38858;
  assign new_n17310_ = ys__n38857 & ~ys__n38858;
  assign new_n17311_ = ~new_n17309_ & ~new_n17310_;
  assign new_n17312_ = new_n17308_ & new_n17311_;
  assign new_n17313_ = ~ys__n38851 & ys__n38852;
  assign new_n17314_ = ys__n38851 & ~ys__n38852;
  assign new_n17315_ = ~new_n17313_ & ~new_n17314_;
  assign new_n17316_ = ~ys__n38853 & ys__n38854;
  assign new_n17317_ = ys__n38853 & ~ys__n38854;
  assign new_n17318_ = ~new_n17316_ & ~new_n17317_;
  assign new_n17319_ = new_n17315_ & new_n17318_;
  assign new_n17320_ = new_n17312_ & new_n17319_;
  assign new_n17321_ = new_n17305_ & new_n17320_;
  assign new_n17322_ = ~ys__n38831 & ys__n38832;
  assign new_n17323_ = ys__n38831 & ~ys__n38832;
  assign new_n17324_ = ~new_n17322_ & ~new_n17323_;
  assign new_n17325_ = ~ys__n38833 & ys__n38834;
  assign new_n17326_ = ys__n38833 & ~ys__n38834;
  assign new_n17327_ = ~new_n17325_ & ~new_n17326_;
  assign new_n17328_ = new_n17324_ & new_n17327_;
  assign new_n17329_ = ~ys__n38827 & ys__n38828;
  assign new_n17330_ = ys__n38827 & ~ys__n38828;
  assign new_n17331_ = ~new_n17329_ & ~new_n17330_;
  assign new_n17332_ = ~ys__n38829 & ys__n38830;
  assign new_n17333_ = ys__n38829 & ~ys__n38830;
  assign new_n17334_ = ~new_n17332_ & ~new_n17333_;
  assign new_n17335_ = new_n17331_ & new_n17334_;
  assign new_n17336_ = new_n17328_ & new_n17335_;
  assign new_n17337_ = ~ys__n38839 & ys__n38840;
  assign new_n17338_ = ys__n38839 & ~ys__n38840;
  assign new_n17339_ = ~new_n17337_ & ~new_n17338_;
  assign new_n17340_ = ~ys__n38841 & ys__n38842;
  assign new_n17341_ = ys__n38841 & ~ys__n38842;
  assign new_n17342_ = ~new_n17340_ & ~new_n17341_;
  assign new_n17343_ = new_n17339_ & new_n17342_;
  assign new_n17344_ = ~ys__n38835 & ys__n38836;
  assign new_n17345_ = ys__n38835 & ~ys__n38836;
  assign new_n17346_ = ~new_n17344_ & ~new_n17345_;
  assign new_n17347_ = ~ys__n38837 & ys__n38838;
  assign new_n17348_ = ys__n38837 & ~ys__n38838;
  assign new_n17349_ = ~new_n17347_ & ~new_n17348_;
  assign new_n17350_ = new_n17346_ & new_n17349_;
  assign new_n17351_ = new_n17343_ & new_n17350_;
  assign new_n17352_ = new_n17336_ & new_n17351_;
  assign new_n17353_ = new_n17321_ & new_n17352_;
  assign new_n17354_ = ~new_n17290_ & new_n17353_;
  assign new_n17355_ = ~new_n17248_ & new_n17354_;
  assign new_n17356_ = ~ys__n18149 & ~ys__n18150;
  assign new_n17357_ = ys__n18137 & ~new_n17356_;
  assign ys__n4696 = new_n17355_ & new_n17357_;
  assign new_n17359_ = new_n12144_ & ~new_n12189_;
  assign new_n17360_ = new_n12155_ & new_n12167_;
  assign new_n17361_ = ~new_n17359_ & new_n17360_;
  assign ys__n4791 = ~new_n12170_ & ~new_n17361_;
  assign ys__n4793 = ~new_n12160_ & ~new_n12170_;
  assign new_n17364_ = ~ys__n574 & ~ys__n4791;
  assign new_n17365_ = ~ys__n4793 & new_n17364_;
  assign ys__n4798 = ys__n576 | ~new_n17365_;
  assign ys__n18166 = ys__n402 & ~ys__n4566;
  assign new_n17368_ = ~ys__n164 & ~ys__n398;
  assign new_n17369_ = ~new_n15135_ & new_n17368_;
  assign new_n17370_ = ~ys__n18166 & new_n17369_;
  assign ys__n4817 = ys__n18166 | new_n17370_;
  assign new_n17372_ = ~ys__n164 & ys__n4826;
  assign new_n17373_ = ~new_n15075_ & ~new_n17372_;
  assign new_n17374_ = ~ys__n398 & ~new_n17373_;
  assign new_n17375_ = ~new_n15135_ & new_n17374_;
  assign ys__n4818 = ~ys__n18166 & new_n17375_;
  assign new_n17377_ = ys__n164 & ys__n4826;
  assign new_n17378_ = ~ys__n4832 & new_n17377_;
  assign new_n17379_ = ys__n4832 & ~new_n17377_;
  assign new_n17380_ = ~new_n17378_ & ~new_n17379_;
  assign new_n17381_ = ~ys__n398 & ~new_n15135_;
  assign new_n17382_ = ~new_n17380_ & new_n17381_;
  assign ys__n4820 = ~ys__n18166 & new_n17382_;
  assign new_n17384_ = ys__n4832 & new_n17377_;
  assign new_n17385_ = ~ys__n4833 & new_n17384_;
  assign new_n17386_ = ys__n4833 & ~new_n17384_;
  assign new_n17387_ = ~new_n17385_ & ~new_n17386_;
  assign new_n17388_ = new_n17381_ & ~new_n17387_;
  assign ys__n4821 = ~ys__n18166 & new_n17388_;
  assign new_n17390_ = ys__n4832 & ys__n4833;
  assign new_n17391_ = new_n17377_ & new_n17390_;
  assign new_n17392_ = ~ys__n354 & new_n17391_;
  assign new_n17393_ = ys__n354 & ~new_n17391_;
  assign new_n17394_ = ~new_n17392_ & ~new_n17393_;
  assign new_n17395_ = new_n17381_ & ~new_n17394_;
  assign ys__n4824 = ~ys__n18166 & new_n17395_;
  assign new_n17397_ = ~ys__n4818 & ~ys__n4820;
  assign new_n17398_ = ~ys__n4821 & ~ys__n4824;
  assign new_n17399_ = new_n17397_ & new_n17398_;
  assign ys__n4825 = ys__n4817 | ~new_n17399_;
  assign new_n17401_ = ~new_n13477_ & ~new_n13481_;
  assign new_n17402_ = ~new_n13484_ & new_n17401_;
  assign ys__n4839 = ys__n4836 & new_n17402_;
  assign ys__n4840 = ys__n4837 & new_n17402_;
  assign new_n17405_ = ys__n47661 & ~new_n11954_;
  assign new_n17406_ = ys__n23269 & ~new_n12314_;
  assign new_n17407_ = new_n11954_ & new_n17406_;
  assign ys__n12455 = new_n17405_ | new_n17407_;
  assign new_n17409_ = ys__n47662 & ~new_n11954_;
  assign new_n17410_ = ys__n23271 & ~new_n12314_;
  assign new_n17411_ = ys__n23272 & new_n12314_;
  assign new_n17412_ = ~new_n17410_ & ~new_n17411_;
  assign new_n17413_ = new_n11954_ & ~new_n17412_;
  assign ys__n12458 = new_n17409_ | new_n17413_;
  assign new_n17415_ = ys__n47663 & ~new_n11954_;
  assign new_n17416_ = ys__n23203 & ~new_n12314_;
  assign new_n17417_ = ys__n23274 & new_n12314_;
  assign new_n17418_ = ~new_n17416_ & ~new_n17417_;
  assign new_n17419_ = new_n11954_ & ~new_n17418_;
  assign ys__n12461 = new_n17415_ | new_n17419_;
  assign new_n17421_ = ys__n47664 & ~new_n11954_;
  assign new_n17422_ = ys__n23205 & ~new_n12314_;
  assign new_n17423_ = ys__n23276 & new_n12314_;
  assign new_n17424_ = ~new_n17422_ & ~new_n17423_;
  assign new_n17425_ = new_n11954_ & ~new_n17424_;
  assign ys__n12464 = new_n17421_ | new_n17425_;
  assign new_n17427_ = ys__n47665 & ~new_n11954_;
  assign new_n17428_ = ys__n23207 & ~new_n12314_;
  assign new_n17429_ = ys__n23278 & new_n12314_;
  assign new_n17430_ = ~new_n17428_ & ~new_n17429_;
  assign new_n17431_ = new_n11954_ & ~new_n17430_;
  assign ys__n12467 = new_n17427_ | new_n17431_;
  assign new_n17433_ = ys__n47666 & ~new_n11954_;
  assign new_n17434_ = ys__n23209 & ~new_n12314_;
  assign new_n17435_ = ys__n23280 & new_n12314_;
  assign new_n17436_ = ~new_n17434_ & ~new_n17435_;
  assign new_n17437_ = new_n11954_ & ~new_n17436_;
  assign ys__n12470 = new_n17433_ | new_n17437_;
  assign new_n17439_ = ys__n47667 & ~new_n11954_;
  assign new_n17440_ = ys__n23211 & ~new_n12314_;
  assign new_n17441_ = ys__n23282 & new_n12314_;
  assign new_n17442_ = ~new_n17440_ & ~new_n17441_;
  assign new_n17443_ = new_n11954_ & ~new_n17442_;
  assign ys__n12473 = new_n17439_ | new_n17443_;
  assign new_n17445_ = ys__n47668 & ~new_n11954_;
  assign new_n17446_ = ys__n23213 & ~new_n12314_;
  assign new_n17447_ = ys__n23284 & new_n12314_;
  assign new_n17448_ = ~new_n17446_ & ~new_n17447_;
  assign new_n17449_ = new_n11954_ & ~new_n17448_;
  assign ys__n12476 = new_n17445_ | new_n17449_;
  assign new_n17451_ = ys__n47669 & ~new_n11954_;
  assign new_n17452_ = ys__n23215 & ~new_n12314_;
  assign new_n17453_ = ys__n23286 & new_n12314_;
  assign new_n17454_ = ~new_n17452_ & ~new_n17453_;
  assign new_n17455_ = new_n11954_ & ~new_n17454_;
  assign ys__n12479 = new_n17451_ | new_n17455_;
  assign new_n17457_ = ys__n47670 & ~new_n11954_;
  assign new_n17458_ = ys__n23217 & ~new_n12314_;
  assign new_n17459_ = ys__n23288 & new_n12314_;
  assign new_n17460_ = ~new_n17458_ & ~new_n17459_;
  assign new_n17461_ = new_n11954_ & ~new_n17460_;
  assign ys__n12482 = new_n17457_ | new_n17461_;
  assign new_n17463_ = ys__n47671 & ~new_n11954_;
  assign new_n17464_ = ys__n23219 & ~new_n12314_;
  assign new_n17465_ = ys__n23290 & new_n12314_;
  assign new_n17466_ = ~new_n17464_ & ~new_n17465_;
  assign new_n17467_ = new_n11954_ & ~new_n17466_;
  assign ys__n12485 = new_n17463_ | new_n17467_;
  assign new_n17469_ = ys__n47672 & ~new_n11954_;
  assign new_n17470_ = ys__n23221 & ~new_n12314_;
  assign new_n17471_ = ys__n23292 & new_n12314_;
  assign new_n17472_ = ~new_n17470_ & ~new_n17471_;
  assign new_n17473_ = new_n11954_ & ~new_n17472_;
  assign ys__n12488 = new_n17469_ | new_n17473_;
  assign new_n17475_ = ys__n47673 & ~new_n11954_;
  assign new_n17476_ = ys__n23223 & ~new_n12314_;
  assign new_n17477_ = ys__n23294 & new_n12314_;
  assign new_n17478_ = ~new_n17476_ & ~new_n17477_;
  assign new_n17479_ = new_n11954_ & ~new_n17478_;
  assign ys__n12491 = new_n17475_ | new_n17479_;
  assign new_n17481_ = ys__n47674 & ~new_n11954_;
  assign new_n17482_ = ys__n23225 & ~new_n12314_;
  assign new_n17483_ = ys__n23296 & new_n12314_;
  assign new_n17484_ = ~new_n17482_ & ~new_n17483_;
  assign new_n17485_ = new_n11954_ & ~new_n17484_;
  assign ys__n12494 = new_n17481_ | new_n17485_;
  assign new_n17487_ = ys__n47675 & ~new_n11954_;
  assign new_n17488_ = ys__n23227 & ~new_n12314_;
  assign new_n17489_ = ys__n23298 & new_n12314_;
  assign new_n17490_ = ~new_n17488_ & ~new_n17489_;
  assign new_n17491_ = new_n11954_ & ~new_n17490_;
  assign ys__n12497 = new_n17487_ | new_n17491_;
  assign new_n17493_ = ys__n47676 & ~new_n11954_;
  assign new_n17494_ = ys__n23229 & ~new_n12314_;
  assign new_n17495_ = ys__n23300 & new_n12314_;
  assign new_n17496_ = ~new_n17494_ & ~new_n17495_;
  assign new_n17497_ = new_n11954_ & ~new_n17496_;
  assign ys__n12500 = new_n17493_ | new_n17497_;
  assign new_n17499_ = ys__n47677 & ~new_n11954_;
  assign new_n17500_ = ys__n23231 & ~new_n12314_;
  assign new_n17501_ = ys__n23302 & new_n12314_;
  assign new_n17502_ = ~new_n17500_ & ~new_n17501_;
  assign new_n17503_ = new_n11954_ & ~new_n17502_;
  assign ys__n12503 = new_n17499_ | new_n17503_;
  assign new_n17505_ = ys__n47678 & ~new_n11954_;
  assign new_n17506_ = ys__n23233 & ~new_n12314_;
  assign new_n17507_ = ys__n23304 & new_n12314_;
  assign new_n17508_ = ~new_n17506_ & ~new_n17507_;
  assign new_n17509_ = new_n11954_ & ~new_n17508_;
  assign ys__n12506 = new_n17505_ | new_n17509_;
  assign new_n17511_ = ys__n47679 & ~new_n11954_;
  assign new_n17512_ = ys__n23235 & ~new_n12314_;
  assign new_n17513_ = ys__n23306 & new_n12314_;
  assign new_n17514_ = ~new_n17512_ & ~new_n17513_;
  assign new_n17515_ = new_n11954_ & ~new_n17514_;
  assign ys__n12509 = new_n17511_ | new_n17515_;
  assign new_n17517_ = ys__n47680 & ~new_n11954_;
  assign new_n17518_ = ys__n23237 & ~new_n12314_;
  assign new_n17519_ = ys__n23308 & new_n12314_;
  assign new_n17520_ = ~new_n17518_ & ~new_n17519_;
  assign new_n17521_ = new_n11954_ & ~new_n17520_;
  assign ys__n12512 = new_n17517_ | new_n17521_;
  assign new_n17523_ = ys__n47681 & ~new_n11954_;
  assign new_n17524_ = ys__n23239 & ~new_n12314_;
  assign new_n17525_ = ys__n23310 & new_n12314_;
  assign new_n17526_ = ~new_n17524_ & ~new_n17525_;
  assign new_n17527_ = new_n11954_ & ~new_n17526_;
  assign ys__n12515 = new_n17523_ | new_n17527_;
  assign new_n17529_ = ys__n47682 & ~new_n11954_;
  assign new_n17530_ = ys__n23241 & ~new_n12314_;
  assign new_n17531_ = ys__n23312 & new_n12314_;
  assign new_n17532_ = ~new_n17530_ & ~new_n17531_;
  assign new_n17533_ = new_n11954_ & ~new_n17532_;
  assign ys__n12518 = new_n17529_ | new_n17533_;
  assign new_n17535_ = ys__n47683 & ~new_n11954_;
  assign new_n17536_ = ys__n23243 & ~new_n12314_;
  assign new_n17537_ = ys__n23314 & new_n12314_;
  assign new_n17538_ = ~new_n17536_ & ~new_n17537_;
  assign new_n17539_ = new_n11954_ & ~new_n17538_;
  assign ys__n12521 = new_n17535_ | new_n17539_;
  assign new_n17541_ = ys__n47684 & ~new_n11954_;
  assign new_n17542_ = ys__n23245 & ~new_n12314_;
  assign new_n17543_ = ys__n23316 & new_n12314_;
  assign new_n17544_ = ~new_n17542_ & ~new_n17543_;
  assign new_n17545_ = new_n11954_ & ~new_n17544_;
  assign ys__n12524 = new_n17541_ | new_n17545_;
  assign new_n17547_ = ys__n47685 & ~new_n11954_;
  assign new_n17548_ = ys__n23247 & ~new_n12314_;
  assign new_n17549_ = ys__n23318 & new_n12314_;
  assign new_n17550_ = ~new_n17548_ & ~new_n17549_;
  assign new_n17551_ = new_n11954_ & ~new_n17550_;
  assign ys__n12527 = new_n17547_ | new_n17551_;
  assign new_n17553_ = ys__n47686 & ~new_n11954_;
  assign new_n17554_ = ys__n23249 & ~new_n12314_;
  assign new_n17555_ = ys__n23320 & new_n12314_;
  assign new_n17556_ = ~new_n17554_ & ~new_n17555_;
  assign new_n17557_ = new_n11954_ & ~new_n17556_;
  assign ys__n12530 = new_n17553_ | new_n17557_;
  assign new_n17559_ = ys__n47687 & ~new_n11954_;
  assign new_n17560_ = ys__n23251 & ~new_n12314_;
  assign new_n17561_ = ys__n23322 & new_n12314_;
  assign new_n17562_ = ~new_n17560_ & ~new_n17561_;
  assign new_n17563_ = new_n11954_ & ~new_n17562_;
  assign ys__n12533 = new_n17559_ | new_n17563_;
  assign new_n17565_ = ys__n47688 & ~new_n11954_;
  assign new_n17566_ = ys__n23253 & ~new_n12314_;
  assign new_n17567_ = ys__n23324 & new_n12314_;
  assign new_n17568_ = ~new_n17566_ & ~new_n17567_;
  assign new_n17569_ = new_n11954_ & ~new_n17568_;
  assign ys__n12536 = new_n17565_ | new_n17569_;
  assign new_n17571_ = ys__n47689 & ~new_n11954_;
  assign new_n17572_ = ys__n23255 & ~new_n12314_;
  assign new_n17573_ = ys__n23326 & new_n12314_;
  assign new_n17574_ = ~new_n17572_ & ~new_n17573_;
  assign new_n17575_ = new_n11954_ & ~new_n17574_;
  assign ys__n12539 = new_n17571_ | new_n17575_;
  assign new_n17577_ = ys__n47690 & ~new_n11954_;
  assign new_n17578_ = ys__n23257 & ~new_n12314_;
  assign new_n17579_ = ~new_n12316_ & ~new_n17578_;
  assign new_n17580_ = new_n11954_ & ~new_n17579_;
  assign ys__n12542 = new_n17577_ | new_n17580_;
  assign new_n17582_ = ys__n47691 & ~new_n11954_;
  assign new_n17583_ = ys__n23259 & ~new_n12314_;
  assign new_n17584_ = ~new_n17119_ & ~new_n17583_;
  assign new_n17585_ = new_n11954_ & ~new_n17584_;
  assign ys__n12545 = new_n17582_ | new_n17585_;
  assign new_n17587_ = ys__n38311 & ~new_n11954_;
  assign new_n17588_ = ys__n23261 & ~new_n12314_;
  assign new_n17589_ = ~new_n12790_ & ~new_n17588_;
  assign new_n17590_ = new_n11954_ & ~new_n17589_;
  assign ys__n12548 = new_n17587_ | new_n17590_;
  assign new_n17592_ = ys__n30223 & new_n13286_;
  assign ys__n16188 = new_n13562_ | new_n17592_;
  assign new_n17594_ = ys__n740 & new_n13320_;
  assign new_n17595_ = new_n13322_ & ys__n3039;
  assign ys__n16412 = new_n17594_ | new_n17595_;
  assign new_n17597_ = new_n13322_ & ~ys__n3039;
  assign new_n17598_ = ys__n23850 & new_n13317_;
  assign ys__n16415 = new_n17597_ | new_n17598_;
  assign new_n17600_ = ys__n30223 & new_n13297_;
  assign ys__n16424 = new_n13584_ | new_n17600_;
  assign new_n17602_ = ys__n740 & new_n13309_;
  assign new_n17603_ = new_n13311_ & ys__n3039;
  assign ys__n16706 = new_n17602_ | new_n17603_;
  assign new_n17605_ = new_n13311_ & ~ys__n3039;
  assign new_n17606_ = ys__n23850 & new_n13306_;
  assign ys__n16709 = new_n17605_ | new_n17606_;
  assign new_n17608_ = ys__n30223 & new_n13330_;
  assign ys__n16718 = new_n13592_ | new_n17608_;
  assign new_n17610_ = ys__n740 & new_n13342_;
  assign new_n17611_ = new_n13344_ & ys__n3039;
  assign ys__n17692 = new_n17610_ | new_n17611_;
  assign new_n17613_ = new_n13344_ & ~ys__n3039;
  assign new_n17614_ = ys__n23850 & new_n13339_;
  assign ys__n17697 = new_n17613_ | new_n17614_;
  assign new_n17616_ = ys__n414 & ys__n728;
  assign new_n17617_ = ys__n724 & ys__n726;
  assign new_n17618_ = new_n17616_ & new_n17617_;
  assign new_n17619_ = ys__n718 & ys__n720;
  assign new_n17620_ = ys__n722 & new_n17619_;
  assign ys__n18007 = new_n17618_ & new_n17620_;
  assign new_n17622_ = ys__n714 & ys__n716;
  assign ys__n18009 = ~ys__n4615 & new_n17622_;
  assign new_n17624_ = ys__n312 & ys__n622;
  assign new_n17625_ = ys__n618 & ys__n620;
  assign new_n17626_ = new_n17624_ & new_n17625_;
  assign new_n17627_ = ys__n612 & ys__n614;
  assign new_n17628_ = ys__n616 & new_n17627_;
  assign ys__n18015 = new_n17626_ & new_n17628_;
  assign new_n17630_ = ys__n456 & ys__n710;
  assign new_n17631_ = ys__n706 & ys__n708;
  assign new_n17632_ = new_n17630_ & new_n17631_;
  assign new_n17633_ = ys__n700 & ys__n702;
  assign new_n17634_ = ys__n704 & new_n17633_;
  assign ys__n18019 = new_n17632_ & new_n17634_;
  assign new_n17636_ = ys__n574 & ~ys__n4791;
  assign new_n17637_ = ~ys__n4793 & new_n17636_;
  assign ys__n18028 = ys__n576 & new_n17637_;
  assign new_n17639_ = ~ys__n628 & ~ys__n794;
  assign new_n17640_ = ~ys__n786 & ~ys__n792;
  assign new_n17641_ = ~ys__n788 & new_n17640_;
  assign new_n17642_ = ys__n630 & new_n17641_;
  assign new_n17643_ = new_n17639_ & new_n17642_;
  assign new_n17644_ = ~ys__n790 & new_n17643_;
  assign new_n17645_ = ~ys__n630 & ~ys__n790;
  assign new_n17646_ = ~ys__n794 & new_n17641_;
  assign new_n17647_ = ys__n628 & new_n17646_;
  assign new_n17648_ = new_n17645_ & new_n17647_;
  assign ys__n18078 = new_n17644_ | new_n17648_;
  assign new_n17650_ = ys__n1301 & ~new_n12861_;
  assign new_n17651_ = ys__n816 & new_n12861_;
  assign new_n17652_ = ~new_n17650_ & ~new_n17651_;
  assign ys__n18080 = ~new_n12865_ & ~new_n17652_;
  assign new_n17654_ = new_n17639_ & new_n17645_;
  assign new_n17655_ = ~ys__n786 & ~ys__n788;
  assign new_n17656_ = ys__n792 & new_n17655_;
  assign new_n17657_ = new_n17654_ & new_n17656_;
  assign new_n17658_ = ys__n18080 & new_n17657_;
  assign new_n17659_ = ys__n794 & new_n17641_;
  assign new_n17660_ = ~ys__n628 & new_n17659_;
  assign new_n17661_ = new_n17645_ & new_n17660_;
  assign new_n17662_ = ~ys__n18078 & ~new_n17661_;
  assign ys__n18082 = new_n17658_ | ~new_n17662_;
  assign new_n17664_ = ~new_n17644_ & ~new_n17661_;
  assign new_n17665_ = ~new_n17657_ & new_n17664_;
  assign new_n17666_ = ~ys__n18080 & ~new_n17665_;
  assign new_n17667_ = ys__n786 & ~ys__n788;
  assign new_n17668_ = ~ys__n792 & new_n17667_;
  assign new_n17669_ = new_n17654_ & new_n17668_;
  assign ys__n18089 = new_n17648_ | new_n17669_;
  assign ys__n18087 = new_n17666_ | ys__n18089;
  assign new_n17672_ = ~ys__n630 & new_n17641_;
  assign new_n17673_ = new_n17639_ & new_n17672_;
  assign new_n17674_ = ys__n790 & new_n17673_;
  assign new_n17675_ = ys__n788 & new_n17640_;
  assign new_n17676_ = new_n17654_ & new_n17675_;
  assign ys__n18088 = ~new_n17674_ & ~new_n17676_;
  assign ys__n18125 = ys__n1094 | ys__n1088;
  assign ys__n24256 = ys__n30219 & ~ys__n4566;
  assign new_n17680_ = ~ys__n846 & new_n11743_;
  assign new_n17681_ = new_n13360_ & new_n17680_;
  assign new_n17682_ = new_n12176_ & new_n17681_;
  assign ys__n18227 = ys__n4176 | ~new_n17682_;
  assign new_n17684_ = ys__n24256 & ~ys__n18227;
  assign new_n17685_ = ys__n18149 & ~ys__n4566;
  assign new_n17686_ = ys__n18227 & new_n17685_;
  assign ys__n18128 = new_n17684_ | new_n17686_;
  assign new_n17688_ = ~ys__n4566 & new_n17682_;
  assign new_n17689_ = ys__n4696 & new_n17688_;
  assign new_n17690_ = ~ys__n33509 & ~ys__n4566;
  assign new_n17691_ = ys__n18150 & ys__n18137;
  assign new_n17692_ = new_n17682_ & new_n17691_;
  assign new_n17693_ = ys__n38776 & ys__n38777;
  assign new_n17694_ = new_n17692_ & new_n17693_;
  assign new_n17695_ = new_n17690_ & new_n17694_;
  assign new_n17696_ = new_n17689_ & new_n17695_;
  assign new_n17697_ = new_n17692_ & ~new_n17693_;
  assign new_n17698_ = ~ys__n33511 & new_n17690_;
  assign new_n17699_ = new_n17697_ & new_n17698_;
  assign new_n17700_ = new_n17689_ & new_n17699_;
  assign ys__n33515 = ~new_n17696_ & ~new_n17700_;
  assign new_n17702_ = ~ys__n1156 & ys__n1157;
  assign new_n17703_ = ~ys__n1156 & ~new_n17702_;
  assign new_n17704_ = ~ys__n1154 & ~new_n17703_;
  assign new_n17705_ = ys__n1154 & new_n17682_;
  assign new_n17706_ = ~new_n17704_ & ~new_n17705_;
  assign new_n17707_ = ~ys__n1153 & ~new_n17706_;
  assign new_n17708_ = ~ys__n18149 & ~ys__n33532;
  assign new_n17709_ = ~ys__n4566 & new_n17708_;
  assign new_n17710_ = new_n17689_ & new_n17709_;
  assign new_n17711_ = ys__n1153 & ~new_n17710_;
  assign new_n17712_ = ~new_n17707_ & ~new_n17711_;
  assign new_n17713_ = ~ys__n1151 & ~new_n17712_;
  assign new_n17714_ = ys__n18150 & new_n17689_;
  assign new_n17715_ = ~ys__n4566 & new_n17714_;
  assign new_n17716_ = new_n12176_ & new_n12180_;
  assign new_n17717_ = ys__n1119 & ~new_n17716_;
  assign new_n17718_ = ~ys__n33491 & ys__n33493;
  assign new_n17719_ = ys__n1088 & new_n17718_;
  assign new_n17720_ = new_n17716_ & new_n17719_;
  assign new_n17721_ = ~ys__n4566 & new_n17720_;
  assign new_n17722_ = ~ys__n4696 & new_n17721_;
  assign new_n17723_ = ~new_n17717_ & ~new_n17722_;
  assign new_n17724_ = ys__n24464 & ~new_n17716_;
  assign new_n17725_ = ys__n4696 & new_n17721_;
  assign new_n17726_ = ~new_n17724_ & ~new_n17725_;
  assign new_n17727_ = ys__n24590 & new_n17356_;
  assign new_n17728_ = ys__n1151 & ~new_n17727_;
  assign new_n17729_ = new_n17726_ & new_n17728_;
  assign new_n17730_ = new_n17723_ & new_n17729_;
  assign new_n17731_ = ~new_n17715_ & new_n17730_;
  assign new_n17732_ = ~new_n17713_ & ~new_n17731_;
  assign new_n17733_ = ~ys__n140 & ~new_n17732_;
  assign ys__n18133 = ys__n140 | new_n17733_;
  assign new_n17735_ = ~ys__n1151 & ys__n1153;
  assign new_n17736_ = ~ys__n33532 & new_n17735_;
  assign new_n17737_ = ~ys__n4566 & new_n17736_;
  assign new_n17738_ = new_n17714_ & new_n17737_;
  assign new_n17739_ = ys__n1151 & new_n17715_;
  assign new_n17740_ = ~new_n17738_ & ~new_n17739_;
  assign ys__n18134 = ~ys__n140 & ~new_n17740_;
  assign new_n17742_ = ~ys__n18133 & ~ys__n18134;
  assign new_n17743_ = ys__n23335 & ys__n27855;
  assign new_n17744_ = new_n11904_ & new_n17743_;
  assign new_n17745_ = ~new_n11904_ & ~new_n17743_;
  assign new_n17746_ = ~new_n17744_ & ~new_n17745_;
  assign new_n17747_ = ~new_n11901_ & new_n17746_;
  assign new_n17748_ = new_n11901_ & new_n17746_;
  assign new_n17749_ = ~new_n17747_ & ~new_n17748_;
  assign new_n17750_ = ~new_n11901_ & ~new_n17746_;
  assign new_n17751_ = new_n11901_ & ~new_n17746_;
  assign new_n17752_ = ~new_n17750_ & ~new_n17751_;
  assign new_n17753_ = new_n17749_ & new_n17752_;
  assign new_n17754_ = ~ys__n1509 & ys__n1511;
  assign new_n17755_ = ~new_n17753_ & new_n17754_;
  assign new_n17756_ = ys__n1509 & ~new_n17749_;
  assign new_n17757_ = ~new_n17753_ & new_n17756_;
  assign new_n17758_ = ~new_n17755_ & ~new_n17757_;
  assign new_n17759_ = ~ys__n1508 & ~new_n17758_;
  assign new_n17760_ = ys__n1508 & new_n17748_;
  assign new_n17761_ = ~new_n17753_ & new_n17760_;
  assign ys__n20045 = new_n17759_ | new_n17761_;
  assign new_n17763_ = ys__n1509 & ~new_n17752_;
  assign new_n17764_ = ~new_n17753_ & new_n17763_;
  assign new_n17765_ = ~new_n17755_ & ~new_n17764_;
  assign new_n17766_ = ~ys__n1508 & ~new_n17765_;
  assign new_n17767_ = ys__n1508 & new_n17751_;
  assign new_n17768_ = ~new_n17753_ & new_n17767_;
  assign ys__n20040 = new_n17766_ | new_n17768_;
  assign ys__n33521 = ~ys__n20045 | ~ys__n20040;
  assign new_n17771_ = ys__n30216 & ys__n33521;
  assign new_n17772_ = ~ys__n18128 & ~new_n17771_;
  assign new_n17773_ = ~ys__n33515 & ~new_n17772_;
  assign ys__n18136 = ~new_n17742_ & new_n17773_;
  assign new_n17775_ = ~ys__n17878 & ~ys__n17879;
  assign new_n17776_ = ~ys__n17881 & ~ys__n17882;
  assign new_n17777_ = new_n17775_ & new_n17776_;
  assign new_n17778_ = ~ys__n17872 & ~ys__n17873;
  assign new_n17779_ = ~ys__n17875 & ~ys__n17876;
  assign new_n17780_ = new_n17778_ & new_n17779_;
  assign new_n17781_ = new_n17777_ & new_n17780_;
  assign new_n17782_ = ~ys__n17890 & ~ys__n17891;
  assign new_n17783_ = ~ys__n17893 & ~ys__n17894;
  assign new_n17784_ = new_n17782_ & new_n17783_;
  assign new_n17785_ = ~ys__n17884 & ~ys__n17885;
  assign new_n17786_ = ~ys__n17887 & ~ys__n17888;
  assign new_n17787_ = new_n17785_ & new_n17786_;
  assign new_n17788_ = new_n17784_ & new_n17787_;
  assign new_n17789_ = new_n17781_ & new_n17788_;
  assign new_n17790_ = ~ys__n17827 & ~ys__n17828;
  assign new_n17791_ = ~ys__n17830 & ~ys__n17831;
  assign new_n17792_ = new_n17790_ & new_n17791_;
  assign new_n17793_ = ~ys__n17833 & ~ys__n17834;
  assign new_n17794_ = ~ys__n17836 & ~ys__n17837;
  assign new_n17795_ = new_n17793_ & new_n17794_;
  assign new_n17796_ = new_n17792_ & new_n17795_;
  assign new_n17797_ = ~ys__n17866 & ~ys__n17867;
  assign new_n17798_ = ~ys__n17869 & ~ys__n17870;
  assign new_n17799_ = new_n17797_ & new_n17798_;
  assign new_n17800_ = ~ys__n17845 & ~ys__n17846;
  assign new_n17801_ = ~ys__n17848 & ~ys__n17849;
  assign new_n17802_ = new_n17800_ & new_n17801_;
  assign new_n17803_ = new_n17799_ & new_n17802_;
  assign new_n17804_ = new_n17796_ & new_n17803_;
  assign new_n17805_ = new_n17789_ & new_n17804_;
  assign new_n17806_ = ~ys__n17803 & ~ys__n17804;
  assign new_n17807_ = ~ys__n17806 & ~ys__n17807;
  assign new_n17808_ = new_n17806_ & new_n17807_;
  assign new_n17809_ = ~ys__n17809 & ~ys__n17810;
  assign new_n17810_ = ~ys__n17812 & ~ys__n17813;
  assign new_n17811_ = new_n17809_ & new_n17810_;
  assign new_n17812_ = new_n17808_ & new_n17811_;
  assign new_n17813_ = ~ys__n17815 & ~ys__n17816;
  assign new_n17814_ = ~ys__n17818 & ~ys__n17819;
  assign new_n17815_ = new_n17813_ & new_n17814_;
  assign new_n17816_ = ~ys__n17821 & ~ys__n17822;
  assign new_n17817_ = ~ys__n17824 & ~ys__n17825;
  assign new_n17818_ = new_n17816_ & new_n17817_;
  assign new_n17819_ = new_n17815_ & new_n17818_;
  assign new_n17820_ = new_n17812_ & new_n17819_;
  assign new_n17821_ = ~ys__n17902 & ~ys__n17903;
  assign new_n17822_ = ~ys__n17905 & ~ys__n17906;
  assign new_n17823_ = new_n17821_ & new_n17822_;
  assign new_n17824_ = ~ys__n17896 & ~ys__n17897;
  assign new_n17825_ = ~ys__n17899 & ~ys__n17900;
  assign new_n17826_ = new_n17824_ & new_n17825_;
  assign new_n17827_ = new_n17823_ & new_n17826_;
  assign new_n17828_ = ~ys__n17839 & ~ys__n17840;
  assign new_n17829_ = ~ys__n17842 & ~ys__n17843;
  assign new_n17830_ = new_n17828_ & new_n17829_;
  assign new_n17831_ = ~ys__n17908 & ~ys__n17909;
  assign new_n17832_ = ~ys__n17911 & ~ys__n17912;
  assign new_n17833_ = new_n17831_ & new_n17832_;
  assign new_n17834_ = new_n17830_ & new_n17833_;
  assign new_n17835_ = new_n17827_ & new_n17834_;
  assign new_n17836_ = new_n17820_ & new_n17835_;
  assign new_n17837_ = new_n17805_ & new_n17836_;
  assign ys__n30330 = ys__n17912 & ~ys__n18156;
  assign new_n17839_ = ~ys__n404 & ys__n30330;
  assign new_n17840_ = ys__n404 & ~ys__n30330;
  assign new_n17841_ = ~new_n17839_ & ~new_n17840_;
  assign ys__n18154 = new_n17837_ | ~new_n17841_;
  assign ys__n18165 = ys__n948 & ~new_n17402_;
  assign new_n17844_ = ~ys__n326 & ys__n332;
  assign new_n17845_ = new_n13456_ & new_n17844_;
  assign new_n17846_ = ~ys__n336 & new_n17845_;
  assign new_n17847_ = new_n13454_ & new_n17844_;
  assign new_n17848_ = ~ys__n336 & new_n17847_;
  assign new_n17849_ = ~new_n17846_ & ~new_n17848_;
  assign ys__n18169 = ys__n598 & ~new_n17849_;
  assign new_n17851_ = ys__n26279 & ~ys__n18169;
  assign new_n17852_ = ys__n26437 & ~ys__n30941;
  assign new_n17853_ = ys__n18169 & new_n17852_;
  assign ys__n18170 = new_n17851_ | new_n17853_;
  assign new_n17855_ = new_n13447_ & new_n17844_;
  assign new_n17856_ = ~ys__n336 & new_n17855_;
  assign new_n17857_ = ~new_n17846_ & ~new_n17856_;
  assign new_n17858_ = ys__n598 & ys__n18173;
  assign ys__n18174 = ~new_n17857_ & new_n17858_;
  assign new_n17860_ = new_n13450_ & new_n17844_;
  assign new_n17861_ = ~ys__n336 & new_n17860_;
  assign new_n17862_ = ~new_n17846_ & ~new_n17861_;
  assign ys__n18176 = new_n17858_ & ~new_n17862_;
  assign ys__n18178 = ~ys__n18208 & new_n15156_;
  assign new_n17865_ = ~ys__n1508 & ~ys__n1509;
  assign new_n17866_ = ~ys__n1511 & new_n17865_;
  assign new_n17867_ = ys__n20035 & new_n17866_;
  assign new_n17868_ = ys__n23326 & ys__n28027;
  assign new_n17869_ = ~new_n11876_ & ~new_n11879_;
  assign new_n17870_ = ys__n23320 & ys__n28024;
  assign new_n17871_ = ys__n23318 & ys__n28023;
  assign new_n17872_ = ~new_n11872_ & new_n17871_;
  assign new_n17873_ = ~new_n17870_ & ~new_n17872_;
  assign new_n17874_ = new_n17869_ & ~new_n17873_;
  assign new_n17875_ = ys__n23324 & ys__n28026;
  assign new_n17876_ = ys__n23322 & ys__n28025;
  assign new_n17877_ = ~new_n11879_ & new_n17876_;
  assign new_n17878_ = ~new_n17875_ & ~new_n17877_;
  assign new_n17879_ = ~new_n17874_ & new_n17878_;
  assign new_n17880_ = ~new_n11869_ & ~new_n11872_;
  assign new_n17881_ = new_n17869_ & new_n17880_;
  assign new_n17882_ = ~new_n11830_ & ~new_n11833_;
  assign new_n17883_ = ~new_n11823_ & ~new_n11826_;
  assign new_n17884_ = new_n17882_ & new_n17883_;
  assign new_n17885_ = ~new_n11845_ & ~new_n11848_;
  assign new_n17886_ = ys__n23304 & ys__n28016;
  assign new_n17887_ = ys__n23302 & ys__n28015;
  assign new_n17888_ = ~new_n11841_ & new_n17887_;
  assign new_n17889_ = ~new_n17886_ & ~new_n17888_;
  assign new_n17890_ = new_n17885_ & ~new_n17889_;
  assign new_n17891_ = ys__n23308 & ys__n28018;
  assign new_n17892_ = ys__n23306 & ys__n28017;
  assign new_n17893_ = ~new_n11848_ & new_n17892_;
  assign new_n17894_ = ~new_n17891_ & ~new_n17893_;
  assign new_n17895_ = ~new_n17890_ & new_n17894_;
  assign new_n17896_ = new_n17884_ & ~new_n17895_;
  assign new_n17897_ = ys__n23312 & ys__n28020;
  assign new_n17898_ = ys__n23310 & ys__n28019;
  assign new_n17899_ = ~new_n11826_ & new_n17898_;
  assign new_n17900_ = ~new_n17897_ & ~new_n17899_;
  assign new_n17901_ = new_n17882_ & ~new_n17900_;
  assign new_n17902_ = ys__n23316 & ys__n28022;
  assign new_n17903_ = ys__n23314 & ys__n28021;
  assign new_n17904_ = ~new_n11833_ & new_n17903_;
  assign new_n17905_ = ~new_n17902_ & ~new_n17904_;
  assign new_n17906_ = ~new_n17901_ & new_n17905_;
  assign new_n17907_ = ~new_n17896_ & new_n17906_;
  assign new_n17908_ = ~new_n11838_ & ~new_n11841_;
  assign new_n17909_ = new_n17885_ & new_n17908_;
  assign new_n17910_ = new_n17884_ & new_n17909_;
  assign new_n17911_ = ys__n23272 & ys__n27857;
  assign new_n17912_ = ~new_n11904_ & new_n17743_;
  assign new_n17913_ = ~new_n17911_ & ~new_n17912_;
  assign new_n17914_ = ~new_n11908_ & ~new_n11911_;
  assign new_n17915_ = ~new_n17913_ & new_n17914_;
  assign new_n17916_ = ys__n23276 & ys__n27861;
  assign new_n17917_ = ys__n23274 & ys__n27859;
  assign new_n17918_ = ~new_n11911_ & new_n17917_;
  assign new_n17919_ = ~new_n17916_ & ~new_n17918_;
  assign new_n17920_ = ~new_n17915_ & new_n17919_;
  assign new_n17921_ = ~new_n11893_ & ~new_n11896_;
  assign new_n17922_ = ~new_n11886_ & ~new_n11889_;
  assign new_n17923_ = new_n17921_ & new_n17922_;
  assign new_n17924_ = ~new_n17920_ & new_n17923_;
  assign new_n17925_ = ys__n23280 & ys__n27865;
  assign new_n17926_ = ys__n23278 & ys__n27863;
  assign new_n17927_ = ~new_n11889_ & new_n17926_;
  assign new_n17928_ = ~new_n17925_ & ~new_n17927_;
  assign new_n17929_ = new_n17921_ & ~new_n17928_;
  assign new_n17930_ = ys__n23284 & ys__n27869;
  assign new_n17931_ = ys__n23282 & ys__n27867;
  assign new_n17932_ = ~new_n11896_ & new_n17931_;
  assign new_n17933_ = ~new_n17930_ & ~new_n17932_;
  assign new_n17934_ = ~new_n17929_ & new_n17933_;
  assign new_n17935_ = ~new_n17924_ & new_n17934_;
  assign new_n17936_ = ~new_n11924_ & ~new_n11927_;
  assign new_n17937_ = ~new_n11917_ & ~new_n11920_;
  assign new_n17938_ = new_n17936_ & new_n17937_;
  assign new_n17939_ = ~new_n11939_ & ~new_n11942_;
  assign new_n17940_ = ~new_n11932_ & ~new_n11935_;
  assign new_n17941_ = new_n17939_ & new_n17940_;
  assign new_n17942_ = new_n17938_ & new_n17941_;
  assign new_n17943_ = ~new_n17935_ & new_n17942_;
  assign new_n17944_ = ys__n23288 & ys__n27873;
  assign new_n17945_ = ys__n23286 & ys__n27871;
  assign new_n17946_ = ~new_n11935_ & new_n17945_;
  assign new_n17947_ = ~new_n17944_ & ~new_n17946_;
  assign new_n17948_ = new_n17939_ & ~new_n17947_;
  assign new_n17949_ = ys__n23292 & ys__n27877;
  assign new_n17950_ = ys__n23290 & ys__n27875;
  assign new_n17951_ = ~new_n11942_ & new_n17950_;
  assign new_n17952_ = ~new_n17949_ & ~new_n17951_;
  assign new_n17953_ = ~new_n17948_ & new_n17952_;
  assign new_n17954_ = new_n17938_ & ~new_n17953_;
  assign new_n17955_ = ys__n23296 & ys__n27881;
  assign new_n17956_ = ys__n23294 & ys__n27879;
  assign new_n17957_ = ~new_n11920_ & new_n17956_;
  assign new_n17958_ = ~new_n17955_ & ~new_n17957_;
  assign new_n17959_ = new_n17936_ & ~new_n17958_;
  assign new_n17960_ = ys__n23300 & ys__n27885;
  assign new_n17961_ = ys__n23298 & ys__n27883;
  assign new_n17962_ = ~new_n11927_ & new_n17961_;
  assign new_n17963_ = ~new_n17960_ & ~new_n17962_;
  assign new_n17964_ = ~new_n17959_ & new_n17963_;
  assign new_n17965_ = ~new_n17954_ & new_n17964_;
  assign new_n17966_ = ~new_n17943_ & new_n17965_;
  assign new_n17967_ = new_n17910_ & ~new_n17966_;
  assign new_n17968_ = new_n17907_ & ~new_n17967_;
  assign new_n17969_ = new_n17881_ & ~new_n17968_;
  assign new_n17970_ = new_n17879_ & ~new_n17969_;
  assign new_n17971_ = ~new_n11854_ & ~new_n17970_;
  assign new_n17972_ = ~new_n17868_ & ~new_n17971_;
  assign new_n17973_ = new_n11857_ & ~new_n17972_;
  assign new_n17974_ = ~new_n11857_ & new_n17972_;
  assign new_n17975_ = ~new_n17973_ & ~new_n17974_;
  assign new_n17976_ = ~new_n17866_ & ~new_n17975_;
  assign ys__n18214 = new_n17867_ | new_n17976_;
  assign new_n17978_ = ys__n23328 & ys__n28028;
  assign new_n17979_ = ~new_n11857_ & new_n17868_;
  assign new_n17980_ = ~new_n17978_ & ~new_n17979_;
  assign new_n17981_ = ~new_n11854_ & ~new_n11857_;
  assign new_n17982_ = ~new_n17970_ & new_n17981_;
  assign new_n17983_ = new_n17980_ & ~new_n17982_;
  assign new_n17984_ = new_n11861_ & ~new_n17983_;
  assign new_n17985_ = ~new_n11861_ & new_n17983_;
  assign new_n17986_ = ~new_n17984_ & ~new_n17985_;
  assign new_n17987_ = ~new_n17866_ & ~new_n17986_;
  assign ys__n18216 = new_n17867_ | new_n17987_;
  assign ys__n18217 = ys__n874 & ys__n18216;
  assign new_n17990_ = ys__n23330 & ys__n28029;
  assign new_n17991_ = ~new_n11861_ & ~new_n17983_;
  assign new_n17992_ = ~new_n17990_ & ~new_n17991_;
  assign new_n17993_ = new_n11864_ & ~new_n17992_;
  assign new_n17994_ = ~new_n11864_ & new_n17992_;
  assign new_n17995_ = ~new_n17993_ & ~new_n17994_;
  assign new_n17996_ = ~new_n17866_ & ~new_n17995_;
  assign ys__n18218 = new_n17867_ | new_n17996_;
  assign ys__n18241 = ~ys__n33548 & ys__n4764;
  assign new_n17999_ = ys__n18242 & ~ys__n18241;
  assign new_n18000_ = ys__n98 & ys__n18241;
  assign new_n18001_ = ~new_n17999_ & ~new_n18000_;
  assign ys__n18223 = ys__n874 & ~new_n18001_;
  assign new_n18003_ = ~ys__n18227 & ys__n18214;
  assign new_n18004_ = ys__n18226 & ys__n18227;
  assign new_n18005_ = ~new_n18003_ & ~new_n18004_;
  assign new_n18006_ = ys__n874 & ~new_n18005_;
  assign new_n18007_ = ~ys__n18227 & ys__n18218;
  assign new_n18008_ = ys__n18231 & ys__n18227;
  assign new_n18009_ = ~new_n18007_ & ~new_n18008_;
  assign new_n18010_ = ys__n874 & ~new_n18009_;
  assign new_n18011_ = new_n18006_ & ~new_n18010_;
  assign new_n18012_ = ~ys__n18227 & ys__n18216;
  assign new_n18013_ = ys__n18229 & ys__n18227;
  assign new_n18014_ = ~new_n18012_ & ~new_n18013_;
  assign ys__n18238 = ys__n874 & ~new_n18014_;
  assign new_n18016_ = new_n18006_ & ys__n18238;
  assign new_n18017_ = new_n18010_ & new_n18016_;
  assign ys__n18236 = new_n18011_ | new_n18017_;
  assign new_n18019_ = ~new_n18010_ & ~ys__n18238;
  assign new_n18020_ = new_n18010_ & ys__n18238;
  assign ys__n18239 = new_n18019_ | new_n18020_;
  assign new_n18022_ = ys__n29886 & ~new_n11737_;
  assign new_n18023_ = ~new_n11735_ & new_n18022_;
  assign new_n18024_ = ~ys__n23764 & new_n18023_;
  assign new_n18025_ = ys__n29902 & ~new_n11737_;
  assign new_n18026_ = ~new_n11735_ & new_n18025_;
  assign new_n18027_ = ~ys__n22466 & new_n18026_;
  assign new_n18028_ = ys__n22466 & new_n18023_;
  assign new_n18029_ = ~new_n18027_ & ~new_n18028_;
  assign new_n18030_ = ys__n23764 & ~new_n18029_;
  assign new_n18031_ = ~new_n18024_ & ~new_n18030_;
  assign ys__n25388 = new_n12000_ & ~new_n18031_;
  assign new_n18033_ = ~ys__n19256 & ys__n25388;
  assign new_n18034_ = ys__n530 & ys__n19256;
  assign new_n18035_ = ~new_n18033_ & ~new_n18034_;
  assign ys__n18251 = ys__n874 & ~new_n18035_;
  assign new_n18037_ = ys__n29893 & ~new_n11737_;
  assign new_n18038_ = ~new_n11735_ & new_n18037_;
  assign new_n18039_ = ~ys__n23764 & new_n18038_;
  assign new_n18040_ = ys__n29909 & ~new_n11737_;
  assign new_n18041_ = ~new_n11735_ & new_n18040_;
  assign new_n18042_ = ~ys__n22466 & new_n18041_;
  assign new_n18043_ = ys__n22466 & new_n18038_;
  assign new_n18044_ = ~new_n18042_ & ~new_n18043_;
  assign new_n18045_ = ys__n23764 & ~new_n18044_;
  assign new_n18046_ = ~new_n18039_ & ~new_n18045_;
  assign ys__n25432 = new_n12000_ & ~new_n18046_;
  assign new_n18048_ = ~ys__n19256 & ys__n25432;
  assign new_n18049_ = ys__n640 & ys__n19256;
  assign new_n18050_ = ~new_n18048_ & ~new_n18049_;
  assign ys__n18360 = ~ys__n874 | new_n18050_;
  assign new_n18052_ = ~new_n13277_ & ys__n18360;
  assign ys__n18268 = new_n13261_ & new_n18052_;
  assign ys__n18273 = ys__n18271 | ys__n4414;
  assign new_n18055_ = ~ys__n846 & ~ys__n4185;
  assign new_n18056_ = ~ys__n4625 & new_n18055_;
  assign new_n18057_ = new_n12175_ & new_n18056_;
  assign new_n18058_ = new_n13361_ & new_n18057_;
  assign new_n18059_ = ~ys__n4613 & new_n18058_;
  assign ys__n18303 = ys__n38522 | new_n18059_;
  assign new_n18061_ = ~ys__n18317 & ~ys__n33300;
  assign new_n18062_ = ys__n37692 & new_n18061_;
  assign new_n18063_ = ys__n3214 & ys__n33311;
  assign new_n18064_ = ~new_n13232_ & new_n18063_;
  assign new_n18065_ = ~ys__n37692 & ~new_n18064_;
  assign new_n18066_ = ys__n18317 & ~new_n18065_;
  assign ys__n18321 = new_n18062_ | new_n18066_;
  assign new_n18068_ = ys__n863 & ~new_n13242_;
  assign new_n18069_ = ys__n842 & new_n13242_;
  assign ys__n18329 = new_n18068_ | new_n18069_;
  assign new_n18071_ = ys__n844 & ys__n863;
  assign new_n18072_ = ~new_n13242_ & new_n18071_;
  assign new_n18073_ = ys__n840 & new_n13242_;
  assign ys__n18331 = new_n18072_ | new_n18073_;
  assign new_n18075_ = ys__n842 & ys__n863;
  assign new_n18076_ = ~new_n13242_ & new_n18075_;
  assign new_n18077_ = ys__n838 & new_n13242_;
  assign ys__n18333 = new_n18076_ | new_n18077_;
  assign new_n18079_ = ys__n840 & ys__n863;
  assign new_n18080_ = ~new_n13242_ & new_n18079_;
  assign new_n18081_ = ys__n836 & new_n13242_;
  assign ys__n18335 = new_n18080_ | new_n18081_;
  assign new_n18083_ = ys__n838 & ys__n863;
  assign new_n18084_ = ~new_n13242_ & new_n18083_;
  assign new_n18085_ = ys__n834 & new_n13242_;
  assign ys__n18337 = new_n18084_ | new_n18085_;
  assign new_n18087_ = ys__n836 & ys__n863;
  assign new_n18088_ = ~new_n13242_ & new_n18087_;
  assign new_n18089_ = ys__n832 & new_n13242_;
  assign ys__n18339 = new_n18088_ | new_n18089_;
  assign new_n18091_ = ys__n834 & ys__n863;
  assign new_n18092_ = ~new_n13242_ & new_n18091_;
  assign new_n18093_ = ys__n830 & new_n13242_;
  assign ys__n18341 = new_n18092_ | new_n18093_;
  assign new_n18095_ = ys__n832 & ys__n863;
  assign new_n18096_ = ~new_n13242_ & new_n18095_;
  assign new_n18097_ = ys__n858 & new_n13242_;
  assign ys__n18343 = new_n18096_ | new_n18097_;
  assign new_n18099_ = ys__n830 & ys__n863;
  assign new_n18100_ = ~new_n13242_ & new_n18099_;
  assign new_n18101_ = ys__n856 & new_n13242_;
  assign ys__n18345 = new_n18100_ | new_n18101_;
  assign new_n18103_ = ys__n858 & ys__n863;
  assign new_n18104_ = ~new_n13242_ & new_n18103_;
  assign new_n18105_ = ys__n854 & new_n13242_;
  assign ys__n18347 = new_n18104_ | new_n18105_;
  assign new_n18107_ = ys__n856 & ys__n863;
  assign new_n18108_ = ~new_n13242_ & new_n18107_;
  assign new_n18109_ = ys__n852 & new_n13242_;
  assign ys__n18349 = new_n18108_ | new_n18109_;
  assign new_n18111_ = ys__n854 & ys__n863;
  assign new_n18112_ = ~new_n13242_ & new_n18111_;
  assign new_n18113_ = ys__n850 & new_n13242_;
  assign ys__n18351 = new_n18112_ | new_n18113_;
  assign new_n18115_ = ys__n852 & ys__n863;
  assign new_n18116_ = ~new_n13242_ & new_n18115_;
  assign new_n18117_ = ys__n848 & new_n13242_;
  assign ys__n18353 = new_n18116_ | new_n18117_;
  assign new_n18119_ = ys__n850 & ys__n863;
  assign new_n18120_ = ~new_n13242_ & new_n18119_;
  assign new_n18121_ = ys__n846 & new_n13242_;
  assign ys__n18355 = new_n18120_ | new_n18121_;
  assign new_n18123_ = ys__n848 & ys__n863;
  assign new_n18124_ = ~new_n13242_ & new_n18123_;
  assign new_n18125_ = ys__n116 & new_n13242_;
  assign ys__n18357 = new_n18124_ | new_n18125_;
  assign new_n18127_ = ys__n18378 & ~ys__n18078;
  assign new_n18128_ = ~ys__n18393 & ys__n18544;
  assign new_n18129_ = ys__n19156 & ys__n18287;
  assign new_n18130_ = ~ys__n18284 & new_n18129_;
  assign new_n18131_ = ys__n18749 & ~new_n12256_;
  assign new_n18132_ = ~ys__n33552 & ~new_n12255_;
  assign new_n18133_ = ~ys__n18759 & ~new_n18132_;
  assign new_n18134_ = ~ys__n38894 & ~new_n18133_;
  assign new_n18135_ = ~ys__n38861 & ~new_n18133_;
  assign new_n18136_ = ~new_n18134_ & ~new_n18135_;
  assign new_n18137_ = ~ys__n38893 & ~new_n18133_;
  assign new_n18138_ = ~ys__n38862 & ~new_n18133_;
  assign new_n18139_ = new_n18137_ & new_n18138_;
  assign new_n18140_ = new_n18136_ & new_n18139_;
  assign new_n18141_ = ~new_n18137_ & ~new_n18138_;
  assign new_n18142_ = new_n18136_ & new_n18141_;
  assign new_n18143_ = new_n18134_ & new_n18135_;
  assign new_n18144_ = new_n18141_ & new_n18143_;
  assign new_n18145_ = ~new_n18142_ & ~new_n18144_;
  assign ys__n18750 = new_n18140_ | ~new_n18145_;
  assign new_n18147_ = new_n12256_ & ys__n18750;
  assign ys__n18751 = new_n18131_ | new_n18147_;
  assign new_n18149_ = ys__n18284 & ys__n18751;
  assign new_n18150_ = ~new_n18130_ & ~new_n18149_;
  assign new_n18151_ = ~ys__n18281 & ~new_n18150_;
  assign new_n18152_ = ~ys__n18281 & ~new_n18151_;
  assign new_n18153_ = ~ys__n18278 & ~new_n18152_;
  assign new_n18154_ = ~ys__n35049 & ys__n46214;
  assign new_n18155_ = ys__n30957 & ~new_n18154_;
  assign new_n18156_ = ys__n26557 & ~ys__n26558;
  assign new_n18157_ = ~ys__n26557 & ys__n26558;
  assign new_n18158_ = ~new_n18156_ & ~new_n18157_;
  assign new_n18159_ = new_n18154_ & ~new_n18158_;
  assign ys__n19149 = new_n18155_ | new_n18159_;
  assign new_n18161_ = ys__n18278 & ys__n19149;
  assign ys__n18545 = new_n18153_ | new_n18161_;
  assign new_n18163_ = ys__n18393 & ys__n18545;
  assign new_n18164_ = ~new_n18128_ & ~new_n18163_;
  assign new_n18165_ = ys__n18078 & ~new_n18164_;
  assign ys__n18380 = new_n18127_ | new_n18165_;
  assign new_n18167_ = ys__n18381 & ~ys__n18078;
  assign new_n18168_ = ~ys__n18393 & ys__n18546;
  assign new_n18169_ = ys__n19157 & ys__n18287;
  assign new_n18170_ = ~ys__n18284 & new_n18169_;
  assign new_n18171_ = ys__n18752 & ~new_n12256_;
  assign ys__n18753 = new_n18142_ & ys__n18750;
  assign new_n18173_ = new_n12256_ & ys__n18753;
  assign ys__n18754 = new_n18171_ | new_n18173_;
  assign new_n18175_ = ys__n18284 & ys__n18754;
  assign new_n18176_ = ~new_n18170_ & ~new_n18175_;
  assign new_n18177_ = ~ys__n18281 & ~new_n18176_;
  assign new_n18178_ = ~ys__n18281 & ~new_n18177_;
  assign new_n18179_ = ~ys__n18278 & ~new_n18178_;
  assign new_n18180_ = ys__n30960 & ~new_n18154_;
  assign new_n18181_ = ys__n26558 & new_n18154_;
  assign ys__n19151 = new_n18180_ | new_n18181_;
  assign new_n18183_ = ys__n18278 & ys__n19151;
  assign ys__n18547 = new_n18179_ | new_n18183_;
  assign new_n18185_ = ys__n18393 & ys__n18547;
  assign new_n18186_ = ~new_n18168_ & ~new_n18185_;
  assign new_n18187_ = ys__n18078 & ~new_n18186_;
  assign ys__n18383 = new_n18167_ | new_n18187_;
  assign new_n18189_ = ys__n18384 & ~ys__n18078;
  assign new_n18190_ = ys__n18208 & ~ys__n18393;
  assign new_n18191_ = ys__n18284 & ~ys__n18281;
  assign new_n18192_ = ~ys__n18281 & ~new_n18191_;
  assign new_n18193_ = ~ys__n18278 & ~new_n18192_;
  assign new_n18194_ = ys__n30961 & ~new_n18154_;
  assign new_n18195_ = ys__n26559 & new_n18154_;
  assign ys__n19159 = new_n18194_ | new_n18195_;
  assign new_n18197_ = ys__n18278 & ys__n19159;
  assign ys__n18555 = new_n18193_ | new_n18197_;
  assign new_n18199_ = ys__n18393 & ys__n18555;
  assign new_n18200_ = ~new_n18190_ & ~new_n18199_;
  assign new_n18201_ = ys__n18078 & ~new_n18200_;
  assign ys__n33324 = ~new_n18189_ & ~new_n18201_;
  assign new_n18203_ = ys__n18389 & ~ys__n18078;
  assign new_n18204_ = ~ys__n18393 & ys__n18556;
  assign new_n18205_ = ys__n18755 & ~new_n12256_;
  assign new_n18206_ = ~ys__n38864 & ~new_n12249_;
  assign new_n18207_ = ~ys__n24675 & ~ys__n18759;
  assign new_n18208_ = ~new_n18206_ & new_n18207_;
  assign new_n18209_ = new_n12256_ & new_n18208_;
  assign ys__n18757 = new_n18205_ | new_n18209_;
  assign new_n18211_ = ~ys__n18281 & ys__n18757;
  assign new_n18212_ = ys__n18284 & new_n18211_;
  assign new_n18213_ = ys__n18647 & ~new_n12259_;
  assign new_n18214_ = ys__n96 & ~ys__n98;
  assign new_n18215_ = ys__n100 & new_n18214_;
  assign new_n18216_ = ys__n78 & ys__n96;
  assign new_n18217_ = ys__n98 & ys__n100;
  assign new_n18218_ = new_n18216_ & new_n18217_;
  assign new_n18219_ = ys__n70 & ys__n72;
  assign new_n18220_ = ys__n74 & ys__n76;
  assign new_n18221_ = new_n18219_ & new_n18220_;
  assign new_n18222_ = new_n18218_ & new_n18221_;
  assign new_n18223_ = ~new_n18215_ & ~new_n18222_;
  assign new_n18224_ = new_n12259_ & ~new_n18223_;
  assign ys__n18649 = new_n18213_ | new_n18224_;
  assign new_n18226_ = ys__n18281 & ~ys__n18649;
  assign new_n18227_ = ~new_n18212_ & ~new_n18226_;
  assign ys__n18557 = ~ys__n18278 & ~new_n18227_;
  assign new_n18229_ = ys__n18393 & ys__n18557;
  assign new_n18230_ = ~new_n18204_ & ~new_n18229_;
  assign new_n18231_ = ys__n18078 & ~new_n18230_;
  assign ys__n33317 = ~new_n18203_ & ~new_n18231_;
  assign new_n18233_ = ys__n18956 & ys__n18287;
  assign new_n18234_ = ~ys__n18284 & new_n18233_;
  assign new_n18235_ = ys__n24615 & ~ys__n4764;
  assign new_n18236_ = ys__n24616 & ys__n4764;
  assign ys__n18764 = new_n18235_ | new_n18236_;
  assign new_n18238_ = ~ys__n18071 & ys__n18764;
  assign new_n18239_ = ys__n18071 & ys__n18765;
  assign new_n18240_ = ~new_n18238_ & ~new_n18239_;
  assign new_n18241_ = ~new_n12256_ & ~new_n18240_;
  assign new_n18242_ = ys__n24616 & ~ys__n24675;
  assign new_n18243_ = ys__n24674 & ys__n24675;
  assign new_n18244_ = ~new_n18242_ & ~new_n18243_;
  assign ys__n18654 = ~new_n18133_ & ~new_n18244_;
  assign new_n18246_ = new_n12256_ & ys__n18654;
  assign ys__n18655 = new_n18241_ | new_n18246_;
  assign new_n18248_ = ys__n18284 & ys__n18655;
  assign new_n18249_ = ~new_n18234_ & ~new_n18248_;
  assign new_n18250_ = ~ys__n18281 & ~new_n18249_;
  assign ys__n18559 = ys__n18558 & ~new_n12259_;
  assign new_n18252_ = ys__n18281 & ys__n18559;
  assign new_n18253_ = ~new_n18250_ & ~new_n18252_;
  assign new_n18254_ = ~ys__n18278 & ~new_n18253_;
  assign new_n18255_ = ys__n18829 & ys__n18278;
  assign ys__n18392 = new_n18254_ | new_n18255_;
  assign new_n18257_ = ys__n6112 & ~ys__n18393;
  assign new_n18258_ = ys__n18393 & ys__n18392;
  assign ys__n18394 = new_n18257_ | new_n18258_;
  assign new_n18260_ = ys__n18957 & ys__n18287;
  assign new_n18261_ = ~ys__n18284 & new_n18260_;
  assign new_n18262_ = ys__n24617 & ~ys__n4764;
  assign new_n18263_ = ys__n24618 & ys__n4764;
  assign ys__n18766 = new_n18262_ | new_n18263_;
  assign new_n18265_ = ~ys__n18071 & ys__n18766;
  assign new_n18266_ = ys__n18071 & ys__n18767;
  assign new_n18267_ = ~new_n18265_ & ~new_n18266_;
  assign new_n18268_ = ~new_n12256_ & ~new_n18267_;
  assign new_n18269_ = ys__n24618 & ~ys__n24675;
  assign new_n18270_ = ys__n24675 & ys__n24677;
  assign new_n18271_ = ~new_n18269_ & ~new_n18270_;
  assign ys__n18657 = ~new_n18133_ & ~new_n18271_;
  assign new_n18273_ = new_n12256_ & ys__n18657;
  assign ys__n18658 = new_n18268_ | new_n18273_;
  assign new_n18275_ = ys__n18284 & ys__n18658;
  assign new_n18276_ = ~new_n18261_ & ~new_n18275_;
  assign new_n18277_ = ~ys__n18281 & ~new_n18276_;
  assign ys__n18561 = ys__n18560 & ~new_n12259_;
  assign new_n18279_ = ys__n18281 & ys__n18561;
  assign new_n18280_ = ~new_n18277_ & ~new_n18279_;
  assign new_n18281_ = ~ys__n18278 & ~new_n18280_;
  assign new_n18282_ = ys__n18831 & ys__n18278;
  assign ys__n18395 = new_n18281_ | new_n18282_;
  assign new_n18284_ = ys__n6113 & ~ys__n18393;
  assign new_n18285_ = ys__n18393 & ys__n18395;
  assign ys__n18396 = new_n18284_ | new_n18285_;
  assign new_n18287_ = ys__n18958 & ys__n18287;
  assign new_n18288_ = ~ys__n18284 & new_n18287_;
  assign new_n18289_ = ys__n24619 & ~ys__n4764;
  assign new_n18290_ = ys__n24620 & ys__n4764;
  assign ys__n18768 = new_n18289_ | new_n18290_;
  assign new_n18292_ = ~ys__n18071 & ys__n18768;
  assign new_n18293_ = ys__n18071 & ys__n18769;
  assign new_n18294_ = ~new_n18292_ & ~new_n18293_;
  assign new_n18295_ = ~new_n12256_ & ~new_n18294_;
  assign new_n18296_ = ys__n24620 & ~ys__n24675;
  assign new_n18297_ = ys__n24675 & ys__n24679;
  assign new_n18298_ = ~new_n18296_ & ~new_n18297_;
  assign new_n18299_ = ys__n24107 & new_n18208_;
  assign ys__n18660 = ~new_n18298_ & ~new_n18299_;
  assign new_n18301_ = new_n12256_ & ys__n18660;
  assign ys__n18661 = new_n18295_ | new_n18301_;
  assign new_n18303_ = ys__n18284 & ys__n18661;
  assign new_n18304_ = ~new_n18288_ & ~new_n18303_;
  assign new_n18305_ = ~ys__n18281 & ~new_n18304_;
  assign new_n18306_ = ys__n18562 & ~new_n12259_;
  assign new_n18307_ = ys__n24107 & new_n18223_;
  assign new_n18308_ = ys__n38896 & new_n12259_;
  assign new_n18309_ = ~new_n18307_ & new_n18308_;
  assign ys__n18564 = new_n18306_ | new_n18309_;
  assign new_n18311_ = ys__n18281 & ys__n18564;
  assign new_n18312_ = ~new_n18305_ & ~new_n18311_;
  assign new_n18313_ = ~ys__n18278 & ~new_n18312_;
  assign new_n18314_ = ys__n18833 & ys__n18278;
  assign ys__n18397 = new_n18313_ | new_n18314_;
  assign new_n18316_ = ys__n172 & ~ys__n18393;
  assign new_n18317_ = ys__n18393 & ys__n18397;
  assign ys__n18398 = new_n18316_ | new_n18317_;
  assign new_n18319_ = ys__n18959 & ys__n18287;
  assign new_n18320_ = ~ys__n18284 & new_n18319_;
  assign new_n18321_ = ys__n24621 & ~ys__n4764;
  assign new_n18322_ = ys__n24622 & ys__n4764;
  assign ys__n18770 = new_n18321_ | new_n18322_;
  assign new_n18324_ = ~ys__n18071 & ys__n18770;
  assign new_n18325_ = ys__n18071 & ys__n18771;
  assign new_n18326_ = ~new_n18324_ & ~new_n18325_;
  assign new_n18327_ = ~new_n12256_ & ~new_n18326_;
  assign new_n18328_ = ys__n24622 & ~ys__n24675;
  assign new_n18329_ = ys__n24675 & ys__n24681;
  assign new_n18330_ = ~new_n18328_ & ~new_n18329_;
  assign ys__n18663 = ~new_n18299_ & ~new_n18330_;
  assign new_n18332_ = new_n12256_ & ys__n18663;
  assign ys__n18664 = new_n18327_ | new_n18332_;
  assign new_n18334_ = ys__n18284 & ys__n18664;
  assign new_n18335_ = ~new_n18320_ & ~new_n18334_;
  assign new_n18336_ = ~ys__n18281 & ~new_n18335_;
  assign new_n18337_ = ys__n18565 & ~new_n12259_;
  assign new_n18338_ = ys__n38897 & new_n12259_;
  assign new_n18339_ = ~new_n18307_ & new_n18338_;
  assign ys__n18567 = new_n18337_ | new_n18339_;
  assign new_n18341_ = ys__n18281 & ys__n18567;
  assign new_n18342_ = ~new_n18336_ & ~new_n18341_;
  assign new_n18343_ = ~ys__n18278 & ~new_n18342_;
  assign new_n18344_ = ys__n18835 & ys__n18278;
  assign ys__n18399 = new_n18343_ | new_n18344_;
  assign new_n18346_ = ys__n338 & ~ys__n18393;
  assign new_n18347_ = ys__n18393 & ys__n18399;
  assign ys__n18400 = new_n18346_ | new_n18347_;
  assign new_n18349_ = ys__n18960 & ys__n18287;
  assign new_n18350_ = ~ys__n18284 & new_n18349_;
  assign new_n18351_ = ys__n24623 & ~ys__n4764;
  assign new_n18352_ = ys__n24624 & ys__n4764;
  assign ys__n18772 = new_n18351_ | new_n18352_;
  assign new_n18354_ = ~ys__n18071 & ys__n18772;
  assign new_n18355_ = ys__n18071 & ys__n18773;
  assign new_n18356_ = ~new_n18354_ & ~new_n18355_;
  assign new_n18357_ = ~new_n12256_ & ~new_n18356_;
  assign new_n18358_ = ys__n24624 & ~ys__n24675;
  assign new_n18359_ = ys__n24675 & ys__n24683;
  assign ys__n18666 = new_n18358_ | new_n18359_;
  assign new_n18361_ = new_n12256_ & ys__n18666;
  assign ys__n18667 = new_n18357_ | new_n18361_;
  assign new_n18363_ = ys__n18284 & ys__n18667;
  assign new_n18364_ = ~new_n18350_ & ~new_n18363_;
  assign new_n18365_ = ~ys__n18281 & ~new_n18364_;
  assign new_n18366_ = ys__n18568 & ~new_n12259_;
  assign new_n18367_ = ys__n18569 & new_n12259_;
  assign ys__n18570 = new_n18366_ | new_n18367_;
  assign new_n18369_ = ys__n18281 & ys__n18570;
  assign new_n18370_ = ~new_n18365_ & ~new_n18369_;
  assign new_n18371_ = ~ys__n18278 & ~new_n18370_;
  assign new_n18372_ = ys__n18837 & ys__n18278;
  assign ys__n18401 = new_n18371_ | new_n18372_;
  assign new_n18374_ = ys__n22 & ~ys__n18393;
  assign new_n18375_ = ys__n18393 & ys__n18401;
  assign ys__n18402 = new_n18374_ | new_n18375_;
  assign new_n18377_ = ys__n18961 & ys__n18287;
  assign new_n18378_ = ~ys__n18284 & new_n18377_;
  assign new_n18379_ = ys__n24625 & ~ys__n4764;
  assign new_n18380_ = ys__n24626 & ys__n4764;
  assign ys__n18774 = new_n18379_ | new_n18380_;
  assign new_n18382_ = ~ys__n18071 & ys__n18774;
  assign new_n18383_ = ys__n18071 & ys__n18775;
  assign new_n18384_ = ~new_n18382_ & ~new_n18383_;
  assign new_n18385_ = ~new_n12256_ & ~new_n18384_;
  assign new_n18386_ = ys__n24626 & ~ys__n24675;
  assign new_n18387_ = ys__n24675 & ys__n24684;
  assign ys__n18669 = new_n18386_ | new_n18387_;
  assign new_n18389_ = new_n12256_ & ys__n18669;
  assign ys__n18670 = new_n18385_ | new_n18389_;
  assign new_n18391_ = ys__n18284 & ys__n18670;
  assign new_n18392_ = ~new_n18378_ & ~new_n18391_;
  assign new_n18393_ = ~ys__n18281 & ~new_n18392_;
  assign new_n18394_ = ys__n18571 & ~new_n12259_;
  assign new_n18395_ = ys__n18572 & new_n12259_;
  assign ys__n18573 = new_n18394_ | new_n18395_;
  assign new_n18397_ = ys__n18281 & ys__n18573;
  assign new_n18398_ = ~new_n18393_ & ~new_n18397_;
  assign new_n18399_ = ~ys__n18278 & ~new_n18398_;
  assign new_n18400_ = ys__n18839 & ys__n18278;
  assign ys__n18403 = new_n18399_ | new_n18400_;
  assign new_n18402_ = ys__n316 & ~ys__n18393;
  assign new_n18403_ = ys__n18393 & ys__n18403;
  assign ys__n18404 = new_n18402_ | new_n18403_;
  assign new_n18405_ = ys__n18962 & ys__n18287;
  assign new_n18406_ = ~ys__n18284 & new_n18405_;
  assign new_n18407_ = ys__n24627 & ~ys__n4764;
  assign new_n18408_ = ys__n24628 & ys__n4764;
  assign ys__n18776 = new_n18407_ | new_n18408_;
  assign new_n18410_ = ~ys__n18071 & ys__n18776;
  assign new_n18411_ = ys__n18071 & ys__n18777;
  assign new_n18412_ = ~new_n18410_ & ~new_n18411_;
  assign new_n18413_ = ~new_n12256_ & ~new_n18412_;
  assign new_n18414_ = ys__n24628 & ~ys__n24675;
  assign new_n18415_ = ys__n24675 & ys__n24685;
  assign ys__n18672 = new_n18414_ | new_n18415_;
  assign new_n18417_ = new_n12256_ & ys__n18672;
  assign ys__n18673 = new_n18413_ | new_n18417_;
  assign new_n18419_ = ys__n18284 & ys__n18673;
  assign new_n18420_ = ~new_n18406_ & ~new_n18419_;
  assign new_n18421_ = ~ys__n18281 & ~new_n18420_;
  assign new_n18422_ = ys__n18574 & ~new_n12259_;
  assign new_n18423_ = ys__n18575 & new_n12259_;
  assign ys__n18576 = new_n18422_ | new_n18423_;
  assign new_n18425_ = ys__n18281 & ys__n18576;
  assign new_n18426_ = ~new_n18421_ & ~new_n18425_;
  assign new_n18427_ = ~ys__n18278 & ~new_n18426_;
  assign new_n18428_ = ys__n18841 & ys__n18278;
  assign ys__n18405 = new_n18427_ | new_n18428_;
  assign new_n18430_ = ys__n6115 & ~ys__n18393;
  assign new_n18431_ = ys__n18393 & ys__n18405;
  assign ys__n18406 = new_n18430_ | new_n18431_;
  assign new_n18433_ = ys__n18963 & ys__n18287;
  assign new_n18434_ = ~ys__n18284 & new_n18433_;
  assign new_n18435_ = ys__n24629 & ~ys__n4764;
  assign new_n18436_ = ys__n24630 & ys__n4764;
  assign ys__n18778 = new_n18435_ | new_n18436_;
  assign new_n18438_ = ~ys__n18071 & ys__n18778;
  assign new_n18439_ = ys__n18071 & ys__n18779;
  assign new_n18440_ = ~new_n18438_ & ~new_n18439_;
  assign new_n18441_ = ~new_n12256_ & ~new_n18440_;
  assign new_n18442_ = ys__n24630 & ~ys__n24675;
  assign new_n18443_ = ys__n24675 & ys__n24686;
  assign ys__n18675 = new_n18442_ | new_n18443_;
  assign new_n18445_ = new_n12256_ & ys__n18675;
  assign ys__n18676 = new_n18441_ | new_n18445_;
  assign new_n18447_ = ys__n18284 & ys__n18676;
  assign new_n18448_ = ~new_n18434_ & ~new_n18447_;
  assign new_n18449_ = ~ys__n18281 & ~new_n18448_;
  assign new_n18450_ = ys__n18577 & ~new_n12259_;
  assign new_n18451_ = ys__n18578 & new_n12259_;
  assign ys__n18579 = new_n18450_ | new_n18451_;
  assign new_n18453_ = ys__n18281 & ys__n18579;
  assign new_n18454_ = ~new_n18449_ & ~new_n18453_;
  assign new_n18455_ = ~ys__n18278 & ~new_n18454_;
  assign new_n18456_ = ys__n18843 & ys__n18278;
  assign ys__n18407 = new_n18455_ | new_n18456_;
  assign new_n18458_ = ys__n44 & ~ys__n18393;
  assign new_n18459_ = ys__n18393 & ys__n18407;
  assign ys__n18408 = new_n18458_ | new_n18459_;
  assign new_n18461_ = ys__n18964 & ys__n18287;
  assign new_n18462_ = ~ys__n18284 & new_n18461_;
  assign new_n18463_ = ys__n24631 & ~ys__n4764;
  assign new_n18464_ = ys__n24632 & ys__n4764;
  assign ys__n18780 = new_n18463_ | new_n18464_;
  assign new_n18466_ = ~ys__n18071 & ys__n18780;
  assign new_n18467_ = ys__n18071 & ys__n18781;
  assign new_n18468_ = ~new_n18466_ & ~new_n18467_;
  assign new_n18469_ = ~new_n12256_ & ~new_n18468_;
  assign new_n18470_ = ys__n24632 & ~ys__n24675;
  assign new_n18471_ = ys__n24675 & ys__n24687;
  assign ys__n18678 = new_n18470_ | new_n18471_;
  assign new_n18473_ = new_n12256_ & ys__n18678;
  assign ys__n18679 = new_n18469_ | new_n18473_;
  assign new_n18475_ = ys__n18284 & ys__n18679;
  assign new_n18476_ = ~new_n18462_ & ~new_n18475_;
  assign new_n18477_ = ~ys__n18281 & ~new_n18476_;
  assign new_n18478_ = ys__n18580 & ~new_n12259_;
  assign new_n18479_ = ys__n18581 & new_n12259_;
  assign ys__n18582 = new_n18478_ | new_n18479_;
  assign new_n18481_ = ys__n18281 & ys__n18582;
  assign new_n18482_ = ~new_n18477_ & ~new_n18481_;
  assign new_n18483_ = ~ys__n18278 & ~new_n18482_;
  assign new_n18484_ = ys__n18845 & ys__n18278;
  assign ys__n18409 = new_n18483_ | new_n18484_;
  assign new_n18486_ = ys__n340 & ~ys__n18393;
  assign new_n18487_ = ys__n18393 & ys__n18409;
  assign ys__n18410 = new_n18486_ | new_n18487_;
  assign new_n18489_ = ys__n18965 & ys__n18287;
  assign new_n18490_ = ~ys__n18284 & new_n18489_;
  assign new_n18491_ = ys__n24633 & ~ys__n4764;
  assign new_n18492_ = ys__n24634 & ys__n4764;
  assign ys__n18782 = new_n18491_ | new_n18492_;
  assign new_n18494_ = ~ys__n18071 & ys__n18782;
  assign new_n18495_ = ys__n18071 & ys__n18783;
  assign new_n18496_ = ~new_n18494_ & ~new_n18495_;
  assign new_n18497_ = ~new_n12256_ & ~new_n18496_;
  assign new_n18498_ = ys__n24634 & ~ys__n24675;
  assign new_n18499_ = ys__n24675 & ys__n24688;
  assign ys__n18681 = new_n18498_ | new_n18499_;
  assign new_n18501_ = new_n12256_ & ys__n18681;
  assign ys__n18682 = new_n18497_ | new_n18501_;
  assign new_n18503_ = ys__n18284 & ys__n18682;
  assign new_n18504_ = ~new_n18490_ & ~new_n18503_;
  assign new_n18505_ = ~ys__n18281 & ~new_n18504_;
  assign new_n18506_ = ys__n18583 & ~new_n12259_;
  assign new_n18507_ = ys__n18584 & new_n12259_;
  assign ys__n18585 = new_n18506_ | new_n18507_;
  assign new_n18509_ = ys__n18281 & ys__n18585;
  assign new_n18510_ = ~new_n18505_ & ~new_n18509_;
  assign new_n18511_ = ~ys__n18278 & ~new_n18510_;
  assign new_n18512_ = ys__n18847 & ys__n18278;
  assign ys__n18411 = new_n18511_ | new_n18512_;
  assign new_n18514_ = ys__n46 & ~ys__n18393;
  assign new_n18515_ = ys__n18393 & ys__n18411;
  assign ys__n18412 = new_n18514_ | new_n18515_;
  assign new_n18517_ = ys__n18966 & ys__n18287;
  assign new_n18518_ = ~ys__n18284 & new_n18517_;
  assign new_n18519_ = ys__n24635 & ~ys__n4764;
  assign new_n18520_ = ys__n24636 & ys__n4764;
  assign ys__n18784 = new_n18519_ | new_n18520_;
  assign new_n18522_ = ~ys__n18071 & ys__n18784;
  assign new_n18523_ = ys__n18071 & ys__n18785;
  assign new_n18524_ = ~new_n18522_ & ~new_n18523_;
  assign new_n18525_ = ~new_n12256_ & ~new_n18524_;
  assign new_n18526_ = ys__n24636 & ~ys__n24675;
  assign new_n18527_ = ys__n24675 & ys__n24689;
  assign ys__n18684 = new_n18526_ | new_n18527_;
  assign new_n18529_ = new_n12256_ & ys__n18684;
  assign ys__n18685 = new_n18525_ | new_n18529_;
  assign new_n18531_ = ys__n18284 & ys__n18685;
  assign new_n18532_ = ~new_n18518_ & ~new_n18531_;
  assign new_n18533_ = ~ys__n18281 & ~new_n18532_;
  assign new_n18534_ = ys__n18586 & ~new_n12259_;
  assign new_n18535_ = ys__n18587 & new_n12259_;
  assign ys__n18588 = new_n18534_ | new_n18535_;
  assign new_n18537_ = ys__n18281 & ys__n18588;
  assign new_n18538_ = ~new_n18533_ & ~new_n18537_;
  assign new_n18539_ = ~ys__n18278 & ~new_n18538_;
  assign new_n18540_ = ys__n18849 & ys__n18278;
  assign ys__n18413 = new_n18539_ | new_n18540_;
  assign new_n18542_ = ys__n6118 & ~ys__n18393;
  assign new_n18543_ = ys__n18393 & ys__n18413;
  assign ys__n18414 = new_n18542_ | new_n18543_;
  assign new_n18545_ = ys__n18967 & ys__n18287;
  assign new_n18546_ = ~ys__n18284 & new_n18545_;
  assign new_n18547_ = ys__n24637 & ~ys__n4764;
  assign new_n18548_ = ys__n24638 & ys__n4764;
  assign ys__n18786 = new_n18547_ | new_n18548_;
  assign new_n18550_ = ~ys__n18071 & ys__n18786;
  assign new_n18551_ = ys__n18071 & ys__n18787;
  assign new_n18552_ = ~new_n18550_ & ~new_n18551_;
  assign new_n18553_ = ~new_n12256_ & ~new_n18552_;
  assign new_n18554_ = ys__n24638 & ~ys__n24675;
  assign new_n18555_ = ys__n24675 & ys__n24690;
  assign ys__n18687 = new_n18554_ | new_n18555_;
  assign new_n18557_ = new_n12256_ & ys__n18687;
  assign ys__n18688 = new_n18553_ | new_n18557_;
  assign new_n18559_ = ys__n18284 & ys__n18688;
  assign new_n18560_ = ~new_n18546_ & ~new_n18559_;
  assign new_n18561_ = ~ys__n18281 & ~new_n18560_;
  assign new_n18562_ = ys__n18589 & ~new_n12259_;
  assign new_n18563_ = ys__n18590 & new_n12259_;
  assign ys__n18591 = new_n18562_ | new_n18563_;
  assign new_n18565_ = ys__n18281 & ys__n18591;
  assign new_n18566_ = ~new_n18561_ & ~new_n18565_;
  assign new_n18567_ = ~ys__n18278 & ~new_n18566_;
  assign new_n18568_ = ys__n18851 & ys__n18278;
  assign ys__n18415 = new_n18567_ | new_n18568_;
  assign new_n18570_ = ys__n6119 & ~ys__n18393;
  assign new_n18571_ = ys__n18393 & ys__n18415;
  assign ys__n18416 = new_n18570_ | new_n18571_;
  assign new_n18573_ = ys__n18968 & ys__n18287;
  assign new_n18574_ = ~ys__n18284 & new_n18573_;
  assign new_n18575_ = ys__n24639 & ~ys__n4764;
  assign new_n18576_ = ys__n24640 & ys__n4764;
  assign ys__n18788 = new_n18575_ | new_n18576_;
  assign new_n18578_ = ~ys__n18071 & ys__n18788;
  assign new_n18579_ = ys__n18071 & ys__n18789;
  assign new_n18580_ = ~new_n18578_ & ~new_n18579_;
  assign new_n18581_ = ~new_n12256_ & ~new_n18580_;
  assign new_n18582_ = ys__n24640 & ~ys__n24675;
  assign new_n18583_ = ys__n24675 & ys__n24691;
  assign ys__n18690 = new_n18582_ | new_n18583_;
  assign new_n18585_ = new_n12256_ & ys__n18690;
  assign ys__n18691 = new_n18581_ | new_n18585_;
  assign new_n18587_ = ys__n18284 & ys__n18691;
  assign new_n18588_ = ~new_n18574_ & ~new_n18587_;
  assign new_n18589_ = ~ys__n18281 & ~new_n18588_;
  assign new_n18590_ = ys__n18592 & ~new_n12259_;
  assign new_n18591_ = ys__n18593 & new_n12259_;
  assign ys__n18594 = new_n18590_ | new_n18591_;
  assign new_n18593_ = ys__n18281 & ys__n18594;
  assign new_n18594_ = ~new_n18589_ & ~new_n18593_;
  assign new_n18595_ = ~ys__n18278 & ~new_n18594_;
  assign new_n18596_ = ys__n18853 & ys__n18278;
  assign ys__n18417 = new_n18595_ | new_n18596_;
  assign new_n18598_ = ys__n6120 & ~ys__n18393;
  assign new_n18599_ = ys__n18393 & ys__n18417;
  assign ys__n18418 = new_n18598_ | new_n18599_;
  assign new_n18601_ = ys__n18969 & ys__n18287;
  assign new_n18602_ = ~ys__n18284 & new_n18601_;
  assign new_n18603_ = ys__n24641 & ~ys__n4764;
  assign new_n18604_ = ys__n24642 & ys__n4764;
  assign ys__n18790 = new_n18603_ | new_n18604_;
  assign new_n18606_ = ~ys__n18071 & ys__n18790;
  assign new_n18607_ = ys__n18071 & ys__n18791;
  assign new_n18608_ = ~new_n18606_ & ~new_n18607_;
  assign new_n18609_ = ~new_n12256_ & ~new_n18608_;
  assign new_n18610_ = ys__n24642 & ~ys__n24675;
  assign new_n18611_ = ys__n24675 & ys__n24692;
  assign ys__n18693 = new_n18610_ | new_n18611_;
  assign new_n18613_ = new_n12256_ & ys__n18693;
  assign ys__n18694 = new_n18609_ | new_n18613_;
  assign new_n18615_ = ys__n18284 & ys__n18694;
  assign new_n18616_ = ~new_n18602_ & ~new_n18615_;
  assign new_n18617_ = ~ys__n18281 & ~new_n18616_;
  assign new_n18618_ = ys__n18595 & ~new_n12259_;
  assign new_n18619_ = ys__n18596 & new_n12259_;
  assign ys__n18597 = new_n18618_ | new_n18619_;
  assign new_n18621_ = ys__n18281 & ys__n18597;
  assign new_n18622_ = ~new_n18617_ & ~new_n18621_;
  assign new_n18623_ = ~ys__n18278 & ~new_n18622_;
  assign new_n18624_ = ys__n18855 & ys__n18278;
  assign ys__n18419 = new_n18623_ | new_n18624_;
  assign new_n18626_ = ys__n6121 & ~ys__n18393;
  assign new_n18627_ = ys__n18393 & ys__n18419;
  assign ys__n18420 = new_n18626_ | new_n18627_;
  assign new_n18629_ = ys__n18970 & ys__n18287;
  assign new_n18630_ = ~ys__n18284 & new_n18629_;
  assign new_n18631_ = ys__n24643 & ~ys__n4764;
  assign new_n18632_ = ys__n24644 & ys__n4764;
  assign ys__n18792 = new_n18631_ | new_n18632_;
  assign new_n18634_ = ~ys__n18071 & ys__n18792;
  assign new_n18635_ = ys__n18071 & ys__n18793;
  assign new_n18636_ = ~new_n18634_ & ~new_n18635_;
  assign new_n18637_ = ~new_n12256_ & ~new_n18636_;
  assign new_n18638_ = ys__n24644 & ~ys__n24675;
  assign new_n18639_ = ys__n24675 & ys__n24693;
  assign ys__n18696 = new_n18638_ | new_n18639_;
  assign new_n18641_ = new_n12256_ & ys__n18696;
  assign ys__n18697 = new_n18637_ | new_n18641_;
  assign new_n18643_ = ys__n18284 & ys__n18697;
  assign new_n18644_ = ~new_n18630_ & ~new_n18643_;
  assign new_n18645_ = ~ys__n18281 & ~new_n18644_;
  assign new_n18646_ = ys__n18598 & ~new_n12259_;
  assign new_n18647_ = ys__n18599 & new_n12259_;
  assign ys__n18600 = new_n18646_ | new_n18647_;
  assign new_n18649_ = ys__n18281 & ys__n18600;
  assign new_n18650_ = ~new_n18645_ & ~new_n18649_;
  assign new_n18651_ = ~ys__n18278 & ~new_n18650_;
  assign new_n18652_ = ys__n18857 & ys__n18278;
  assign ys__n18421 = new_n18651_ | new_n18652_;
  assign new_n18654_ = ys__n6123 & ~ys__n18393;
  assign new_n18655_ = ys__n18393 & ys__n18421;
  assign ys__n18422 = new_n18654_ | new_n18655_;
  assign new_n18657_ = ys__n18971 & ys__n18287;
  assign new_n18658_ = ~ys__n18284 & new_n18657_;
  assign new_n18659_ = ys__n24645 & ~ys__n4764;
  assign new_n18660_ = ys__n24646 & ys__n4764;
  assign ys__n18794 = new_n18659_ | new_n18660_;
  assign new_n18662_ = ~ys__n18071 & ys__n18794;
  assign new_n18663_ = ys__n18071 & ys__n18795;
  assign new_n18664_ = ~new_n18662_ & ~new_n18663_;
  assign new_n18665_ = ~new_n12256_ & ~new_n18664_;
  assign new_n18666_ = ys__n24646 & ~ys__n24675;
  assign new_n18667_ = ys__n24675 & ys__n24694;
  assign ys__n18699 = new_n18666_ | new_n18667_;
  assign new_n18669_ = new_n12256_ & ys__n18699;
  assign ys__n18700 = new_n18665_ | new_n18669_;
  assign new_n18671_ = ys__n18284 & ys__n18700;
  assign new_n18672_ = ~new_n18658_ & ~new_n18671_;
  assign new_n18673_ = ~ys__n18281 & ~new_n18672_;
  assign new_n18674_ = ys__n18601 & ~new_n12259_;
  assign new_n18675_ = ys__n18602 & new_n12259_;
  assign ys__n18603 = new_n18674_ | new_n18675_;
  assign new_n18677_ = ys__n18281 & ys__n18603;
  assign new_n18678_ = ~new_n18673_ & ~new_n18677_;
  assign new_n18679_ = ~ys__n18278 & ~new_n18678_;
  assign new_n18680_ = ys__n18859 & ys__n18278;
  assign ys__n18423 = new_n18679_ | new_n18680_;
  assign new_n18682_ = ys__n6124 & ~ys__n18393;
  assign new_n18683_ = ys__n18393 & ys__n18423;
  assign ys__n18424 = new_n18682_ | new_n18683_;
  assign new_n18685_ = ys__n18972 & ys__n18287;
  assign new_n18686_ = ~ys__n18284 & new_n18685_;
  assign new_n18687_ = ys__n24647 & ~ys__n4764;
  assign new_n18688_ = ys__n24648 & ys__n4764;
  assign ys__n18796 = new_n18687_ | new_n18688_;
  assign new_n18690_ = ~ys__n18071 & ys__n18796;
  assign new_n18691_ = ys__n18071 & ys__n18797;
  assign new_n18692_ = ~new_n18690_ & ~new_n18691_;
  assign new_n18693_ = ~new_n12256_ & ~new_n18692_;
  assign new_n18694_ = ys__n24648 & ~ys__n24675;
  assign new_n18695_ = ys__n24675 & ys__n24695;
  assign ys__n18702 = new_n18694_ | new_n18695_;
  assign new_n18697_ = new_n12256_ & ys__n18702;
  assign ys__n18703 = new_n18693_ | new_n18697_;
  assign new_n18699_ = ys__n18284 & ys__n18703;
  assign new_n18700_ = ~new_n18686_ & ~new_n18699_;
  assign new_n18701_ = ~ys__n18281 & ~new_n18700_;
  assign new_n18702_ = ys__n18604 & ~new_n12259_;
  assign new_n18703_ = ys__n18605 & new_n12259_;
  assign ys__n18606 = new_n18702_ | new_n18703_;
  assign new_n18705_ = ys__n18281 & ys__n18606;
  assign new_n18706_ = ~new_n18701_ & ~new_n18705_;
  assign new_n18707_ = ~ys__n18278 & ~new_n18706_;
  assign new_n18708_ = ys__n18861 & ys__n18278;
  assign ys__n18425 = new_n18707_ | new_n18708_;
  assign new_n18710_ = ys__n6126 & ~ys__n18393;
  assign new_n18711_ = ys__n18393 & ys__n18425;
  assign ys__n18426 = new_n18710_ | new_n18711_;
  assign new_n18713_ = ys__n18973 & ys__n18287;
  assign new_n18714_ = ~ys__n18284 & new_n18713_;
  assign new_n18715_ = ys__n24649 & ~ys__n4764;
  assign new_n18716_ = ys__n24650 & ys__n4764;
  assign ys__n18798 = new_n18715_ | new_n18716_;
  assign new_n18718_ = ~ys__n18071 & ys__n18798;
  assign new_n18719_ = ys__n18071 & ys__n18799;
  assign new_n18720_ = ~new_n18718_ & ~new_n18719_;
  assign new_n18721_ = ~new_n12256_ & ~new_n18720_;
  assign new_n18722_ = ys__n24650 & ~ys__n24675;
  assign new_n18723_ = ys__n24675 & ys__n24696;
  assign ys__n18705 = new_n18722_ | new_n18723_;
  assign new_n18725_ = new_n12256_ & ys__n18705;
  assign ys__n18706 = new_n18721_ | new_n18725_;
  assign new_n18727_ = ys__n18284 & ys__n18706;
  assign new_n18728_ = ~new_n18714_ & ~new_n18727_;
  assign new_n18729_ = ~ys__n18281 & ~new_n18728_;
  assign new_n18730_ = ys__n18607 & ~new_n12259_;
  assign new_n18731_ = ys__n18608 & new_n12259_;
  assign ys__n18609 = new_n18730_ | new_n18731_;
  assign new_n18733_ = ys__n18281 & ys__n18609;
  assign new_n18734_ = ~new_n18729_ & ~new_n18733_;
  assign new_n18735_ = ~ys__n18278 & ~new_n18734_;
  assign new_n18736_ = ys__n18863 & ys__n18278;
  assign ys__n18427 = new_n18735_ | new_n18736_;
  assign new_n18738_ = ys__n6127 & ~ys__n18393;
  assign new_n18739_ = ys__n18393 & ys__n18427;
  assign ys__n18428 = new_n18738_ | new_n18739_;
  assign new_n18741_ = ys__n18974 & ys__n18287;
  assign new_n18742_ = ~ys__n18284 & new_n18741_;
  assign new_n18743_ = ys__n24651 & ~ys__n4764;
  assign new_n18744_ = ys__n24652 & ys__n4764;
  assign ys__n18800 = new_n18743_ | new_n18744_;
  assign new_n18746_ = ~ys__n18071 & ys__n18800;
  assign new_n18747_ = ys__n18071 & ys__n18801;
  assign new_n18748_ = ~new_n18746_ & ~new_n18747_;
  assign new_n18749_ = ~new_n12256_ & ~new_n18748_;
  assign new_n18750_ = ys__n24652 & ~ys__n24675;
  assign new_n18751_ = ys__n24675 & ys__n24697;
  assign ys__n18708 = new_n18750_ | new_n18751_;
  assign new_n18753_ = new_n12256_ & ys__n18708;
  assign ys__n18709 = new_n18749_ | new_n18753_;
  assign new_n18755_ = ys__n18284 & ys__n18709;
  assign new_n18756_ = ~new_n18742_ & ~new_n18755_;
  assign new_n18757_ = ~ys__n18281 & ~new_n18756_;
  assign new_n18758_ = ys__n18610 & ~new_n12259_;
  assign new_n18759_ = ys__n18611 & new_n12259_;
  assign ys__n18612 = new_n18758_ | new_n18759_;
  assign new_n18761_ = ys__n18281 & ys__n18612;
  assign new_n18762_ = ~new_n18757_ & ~new_n18761_;
  assign new_n18763_ = ~ys__n18278 & ~new_n18762_;
  assign new_n18764_ = ys__n18865 & ys__n18278;
  assign ys__n18429 = new_n18763_ | new_n18764_;
  assign new_n18766_ = ys__n6129 & ~ys__n18393;
  assign new_n18767_ = ys__n18393 & ys__n18429;
  assign ys__n18430 = new_n18766_ | new_n18767_;
  assign new_n18769_ = ys__n18975 & ys__n18287;
  assign new_n18770_ = ~ys__n18284 & new_n18769_;
  assign new_n18771_ = ys__n24653 & ~ys__n4764;
  assign new_n18772_ = ys__n24654 & ys__n4764;
  assign ys__n18802 = new_n18771_ | new_n18772_;
  assign new_n18774_ = ~ys__n18071 & ys__n18802;
  assign new_n18775_ = ys__n18071 & ys__n18803;
  assign new_n18776_ = ~new_n18774_ & ~new_n18775_;
  assign new_n18777_ = ~new_n12256_ & ~new_n18776_;
  assign new_n18778_ = ys__n24654 & ~ys__n24675;
  assign new_n18779_ = ys__n24675 & ys__n24698;
  assign ys__n18711 = new_n18778_ | new_n18779_;
  assign new_n18781_ = new_n12256_ & ys__n18711;
  assign ys__n18712 = new_n18777_ | new_n18781_;
  assign new_n18783_ = ys__n18284 & ys__n18712;
  assign new_n18784_ = ~new_n18770_ & ~new_n18783_;
  assign new_n18785_ = ~ys__n18281 & ~new_n18784_;
  assign new_n18786_ = ys__n18613 & ~new_n12259_;
  assign new_n18787_ = ys__n18614 & new_n12259_;
  assign ys__n18615 = new_n18786_ | new_n18787_;
  assign new_n18789_ = ys__n18281 & ys__n18615;
  assign new_n18790_ = ~new_n18785_ & ~new_n18789_;
  assign new_n18791_ = ~ys__n18278 & ~new_n18790_;
  assign new_n18792_ = ys__n18867 & ys__n18278;
  assign ys__n18431 = new_n18791_ | new_n18792_;
  assign new_n18794_ = ys__n6130 & ~ys__n18393;
  assign new_n18795_ = ys__n18393 & ys__n18431;
  assign ys__n18432 = new_n18794_ | new_n18795_;
  assign new_n18797_ = ys__n18976 & ys__n18287;
  assign new_n18798_ = ~ys__n18284 & new_n18797_;
  assign new_n18799_ = ys__n24655 & ~ys__n4764;
  assign new_n18800_ = ys__n24656 & ys__n4764;
  assign ys__n18804 = new_n18799_ | new_n18800_;
  assign new_n18802_ = ~ys__n18071 & ys__n18804;
  assign new_n18803_ = ys__n18071 & ys__n18805;
  assign new_n18804_ = ~new_n18802_ & ~new_n18803_;
  assign new_n18805_ = ~new_n12256_ & ~new_n18804_;
  assign new_n18806_ = ys__n24656 & ~ys__n24675;
  assign new_n18807_ = ys__n24675 & ys__n24699;
  assign ys__n18714 = new_n18806_ | new_n18807_;
  assign new_n18809_ = new_n12256_ & ys__n18714;
  assign ys__n18715 = new_n18805_ | new_n18809_;
  assign new_n18811_ = ys__n18284 & ys__n18715;
  assign new_n18812_ = ~new_n18798_ & ~new_n18811_;
  assign new_n18813_ = ~ys__n18281 & ~new_n18812_;
  assign new_n18814_ = ys__n18616 & ~new_n12259_;
  assign new_n18815_ = ys__n18617 & new_n12259_;
  assign ys__n18618 = new_n18814_ | new_n18815_;
  assign new_n18817_ = ys__n18281 & ys__n18618;
  assign new_n18818_ = ~new_n18813_ & ~new_n18817_;
  assign new_n18819_ = ~ys__n18278 & ~new_n18818_;
  assign new_n18820_ = ys__n18869 & ys__n18278;
  assign ys__n18433 = new_n18819_ | new_n18820_;
  assign new_n18822_ = ys__n42 & ~ys__n18393;
  assign new_n18823_ = ys__n18393 & ys__n18433;
  assign ys__n18434 = new_n18822_ | new_n18823_;
  assign new_n18825_ = ys__n40 & ~ys__n18393;
  assign new_n18826_ = ys__n18393 & ys__n806;
  assign ys__n18435 = new_n18825_ | new_n18826_;
  assign new_n18828_ = ys__n6133 & ~ys__n18393;
  assign new_n18829_ = ys__n18393 & ys__n3250;
  assign ys__n18436 = new_n18828_ | new_n18829_;
  assign new_n18831_ = ys__n6134 & ~ys__n18393;
  assign new_n18832_ = ys__n18393 & ys__n3252;
  assign ys__n18437 = new_n18831_ | new_n18832_;
  assign new_n18834_ = ys__n38 & ~ys__n18393;
  assign new_n18835_ = ys__n18393 & ys__n804;
  assign ys__n18438 = new_n18834_ | new_n18835_;
  assign new_n18837_ = ys__n36 & ~ys__n18393;
  assign new_n18838_ = ys__n18393 & ys__n802;
  assign ys__n18439 = new_n18837_ | new_n18838_;
  assign new_n18840_ = ys__n34 & ~ys__n18393;
  assign new_n18841_ = ys__n18393 & ys__n800;
  assign ys__n18440 = new_n18840_ | new_n18841_;
  assign new_n18843_ = ys__n32 & ~ys__n18393;
  assign new_n18844_ = ys__n18393 & ys__n798;
  assign ys__n18441 = new_n18843_ | new_n18844_;
  assign new_n18846_ = ys__n30 & ~ys__n18393;
  assign new_n18847_ = ys__n18393 & ys__n796;
  assign ys__n18442 = new_n18846_ | new_n18847_;
  assign new_n18849_ = ys__n28 & ~ys__n18393;
  assign new_n18850_ = ys__n18393 & ys__n810;
  assign ys__n18443 = new_n18849_ | new_n18850_;
  assign new_n18852_ = ys__n26 & ~ys__n18393;
  assign new_n18853_ = ys__n18393 & ys__n808;
  assign ys__n18444 = new_n18852_ | new_n18853_;
  assign new_n18855_ = ys__n24 & ~ys__n18393;
  assign new_n18856_ = ys__n18393 & ys__n812;
  assign ys__n18445 = new_n18855_ | new_n18856_;
  assign new_n18858_ = ys__n19116 & ~ys__n18281;
  assign new_n18859_ = ~ys__n18278 & new_n18858_;
  assign new_n18860_ = ys__n18287 & new_n18859_;
  assign new_n18861_ = ~ys__n18284 & new_n18860_;
  assign new_n18862_ = ys__n18989 & ys__n18278;
  assign ys__n18449 = new_n18861_ | new_n18862_;
  assign new_n18864_ = ~ys__n18393 & ys__n18448;
  assign new_n18865_ = ys__n18393 & ys__n18449;
  assign ys__n18450 = new_n18864_ | new_n18865_;
  assign new_n18867_ = ys__n19117 & ~ys__n18281;
  assign new_n18868_ = ~ys__n18278 & new_n18867_;
  assign new_n18869_ = ys__n18287 & new_n18868_;
  assign new_n18870_ = ~ys__n18284 & new_n18869_;
  assign new_n18871_ = ys__n18991 & ys__n18278;
  assign ys__n18452 = new_n18870_ | new_n18871_;
  assign new_n18873_ = ~ys__n18393 & ys__n18451;
  assign new_n18874_ = ys__n18393 & ys__n18452;
  assign ys__n18453 = new_n18873_ | new_n18874_;
  assign new_n18876_ = ys__n19118 & ~ys__n18281;
  assign new_n18877_ = ~ys__n18278 & new_n18876_;
  assign new_n18878_ = ys__n18287 & new_n18877_;
  assign new_n18879_ = ~ys__n18284 & new_n18878_;
  assign new_n18880_ = ys__n18993 & ys__n18278;
  assign ys__n18455 = new_n18879_ | new_n18880_;
  assign new_n18882_ = ~ys__n18393 & ys__n18454;
  assign new_n18883_ = ys__n18393 & ys__n18455;
  assign ys__n18456 = new_n18882_ | new_n18883_;
  assign new_n18885_ = ys__n19119 & ~ys__n18281;
  assign new_n18886_ = ~ys__n18278 & new_n18885_;
  assign new_n18887_ = ys__n18287 & new_n18886_;
  assign new_n18888_ = ~ys__n18284 & new_n18887_;
  assign new_n18889_ = ys__n18995 & ys__n18278;
  assign ys__n18458 = new_n18888_ | new_n18889_;
  assign new_n18891_ = ~ys__n18393 & ys__n18457;
  assign new_n18892_ = ys__n18393 & ys__n18458;
  assign ys__n18459 = new_n18891_ | new_n18892_;
  assign new_n18894_ = ys__n19120 & ~ys__n18281;
  assign new_n18895_ = ~ys__n18278 & new_n18894_;
  assign new_n18896_ = ys__n18287 & new_n18895_;
  assign new_n18897_ = ~ys__n18284 & new_n18896_;
  assign new_n18898_ = ys__n18997 & ys__n18278;
  assign ys__n18461 = new_n18897_ | new_n18898_;
  assign new_n18900_ = ~ys__n18393 & ys__n18460;
  assign new_n18901_ = ys__n18393 & ys__n18461;
  assign ys__n18462 = new_n18900_ | new_n18901_;
  assign new_n18903_ = ys__n19121 & ~ys__n18281;
  assign new_n18904_ = ~ys__n18278 & new_n18903_;
  assign new_n18905_ = ys__n18287 & new_n18904_;
  assign new_n18906_ = ~ys__n18284 & new_n18905_;
  assign new_n18907_ = ys__n18999 & ys__n18278;
  assign ys__n18464 = new_n18906_ | new_n18907_;
  assign new_n18909_ = ~ys__n18393 & ys__n18463;
  assign new_n18910_ = ys__n18393 & ys__n18464;
  assign ys__n18465 = new_n18909_ | new_n18910_;
  assign new_n18912_ = ys__n19122 & ~ys__n18281;
  assign new_n18913_ = ~ys__n18278 & new_n18912_;
  assign new_n18914_ = ys__n18287 & new_n18913_;
  assign new_n18915_ = ~ys__n18284 & new_n18914_;
  assign new_n18916_ = ys__n19001 & ys__n18278;
  assign ys__n18467 = new_n18915_ | new_n18916_;
  assign new_n18918_ = ~ys__n18393 & ys__n18466;
  assign new_n18919_ = ys__n18393 & ys__n18467;
  assign ys__n18468 = new_n18918_ | new_n18919_;
  assign new_n18921_ = ys__n19123 & ~ys__n18281;
  assign new_n18922_ = ~ys__n18278 & new_n18921_;
  assign new_n18923_ = ys__n18287 & new_n18922_;
  assign new_n18924_ = ~ys__n18284 & new_n18923_;
  assign new_n18925_ = ys__n19003 & ys__n18278;
  assign ys__n18470 = new_n18924_ | new_n18925_;
  assign new_n18927_ = ~ys__n18393 & ys__n18469;
  assign new_n18928_ = ys__n18393 & ys__n18470;
  assign ys__n18471 = new_n18927_ | new_n18928_;
  assign new_n18930_ = ys__n19124 & ~ys__n18281;
  assign new_n18931_ = ~ys__n18278 & new_n18930_;
  assign new_n18932_ = ys__n18287 & new_n18931_;
  assign new_n18933_ = ~ys__n18284 & new_n18932_;
  assign new_n18934_ = ys__n19005 & ys__n18278;
  assign ys__n18473 = new_n18933_ | new_n18934_;
  assign new_n18936_ = ~ys__n18393 & ys__n18472;
  assign new_n18937_ = ys__n18393 & ys__n18473;
  assign ys__n18474 = new_n18936_ | new_n18937_;
  assign new_n18939_ = ys__n19125 & ~ys__n18281;
  assign new_n18940_ = ~ys__n18278 & new_n18939_;
  assign new_n18941_ = ys__n18287 & new_n18940_;
  assign new_n18942_ = ~ys__n18284 & new_n18941_;
  assign new_n18943_ = ys__n19007 & ys__n18278;
  assign ys__n18476 = new_n18942_ | new_n18943_;
  assign new_n18945_ = ~ys__n18393 & ys__n18475;
  assign new_n18946_ = ys__n18393 & ys__n18476;
  assign ys__n18477 = new_n18945_ | new_n18946_;
  assign new_n18948_ = ys__n19126 & ~ys__n18281;
  assign new_n18949_ = ~ys__n18278 & new_n18948_;
  assign new_n18950_ = ys__n18287 & new_n18949_;
  assign new_n18951_ = ~ys__n18284 & new_n18950_;
  assign new_n18952_ = ys__n19009 & ys__n18278;
  assign ys__n18479 = new_n18951_ | new_n18952_;
  assign new_n18954_ = ~ys__n18393 & ys__n18478;
  assign new_n18955_ = ys__n18393 & ys__n18479;
  assign ys__n18480 = new_n18954_ | new_n18955_;
  assign new_n18957_ = ys__n19127 & ~ys__n18281;
  assign new_n18958_ = ~ys__n18278 & new_n18957_;
  assign new_n18959_ = ys__n18287 & new_n18958_;
  assign new_n18960_ = ~ys__n18284 & new_n18959_;
  assign new_n18961_ = ys__n19011 & ys__n18278;
  assign ys__n18482 = new_n18960_ | new_n18961_;
  assign new_n18963_ = ~ys__n18393 & ys__n18481;
  assign new_n18964_ = ys__n18393 & ys__n18482;
  assign ys__n18483 = new_n18963_ | new_n18964_;
  assign new_n18966_ = ys__n19128 & ~ys__n18281;
  assign new_n18967_ = ~ys__n18278 & new_n18966_;
  assign new_n18968_ = ys__n18287 & new_n18967_;
  assign new_n18969_ = ~ys__n18284 & new_n18968_;
  assign new_n18970_ = ys__n19013 & ys__n18278;
  assign ys__n18485 = new_n18969_ | new_n18970_;
  assign new_n18972_ = ~ys__n18393 & ys__n18484;
  assign new_n18973_ = ys__n18393 & ys__n18485;
  assign ys__n18486 = new_n18972_ | new_n18973_;
  assign new_n18975_ = ys__n19129 & ~ys__n18281;
  assign new_n18976_ = ~ys__n18278 & new_n18975_;
  assign new_n18977_ = ys__n18287 & new_n18976_;
  assign new_n18978_ = ~ys__n18284 & new_n18977_;
  assign new_n18979_ = ys__n19015 & ys__n18278;
  assign ys__n18488 = new_n18978_ | new_n18979_;
  assign new_n18981_ = ~ys__n18393 & ys__n18487;
  assign new_n18982_ = ys__n18393 & ys__n18488;
  assign ys__n18489 = new_n18981_ | new_n18982_;
  assign new_n18984_ = ys__n19130 & ~ys__n18281;
  assign new_n18985_ = ~ys__n18278 & new_n18984_;
  assign new_n18986_ = ys__n18287 & new_n18985_;
  assign new_n18987_ = ~ys__n18284 & new_n18986_;
  assign new_n18988_ = ys__n19017 & ys__n18278;
  assign ys__n18491 = new_n18987_ | new_n18988_;
  assign new_n18990_ = ~ys__n18393 & ys__n18490;
  assign new_n18991_ = ys__n18393 & ys__n18491;
  assign ys__n18492 = new_n18990_ | new_n18991_;
  assign new_n18993_ = ys__n19131 & ~ys__n18281;
  assign new_n18994_ = ~ys__n18278 & new_n18993_;
  assign new_n18995_ = ys__n18287 & new_n18994_;
  assign new_n18996_ = ~ys__n18284 & new_n18995_;
  assign new_n18997_ = ys__n19019 & ys__n18278;
  assign ys__n18494 = new_n18996_ | new_n18997_;
  assign new_n18999_ = ~ys__n18393 & ys__n18493;
  assign new_n19000_ = ys__n18393 & ys__n18494;
  assign ys__n18495 = new_n18999_ | new_n19000_;
  assign new_n19002_ = ys__n19132 & ~ys__n18281;
  assign new_n19003_ = ~ys__n18278 & new_n19002_;
  assign new_n19004_ = ys__n18287 & new_n19003_;
  assign new_n19005_ = ~ys__n18284 & new_n19004_;
  assign new_n19006_ = ys__n19021 & ys__n18278;
  assign ys__n18497 = new_n19005_ | new_n19006_;
  assign new_n19008_ = ~ys__n18393 & ys__n18496;
  assign new_n19009_ = ys__n18393 & ys__n18497;
  assign ys__n18498 = new_n19008_ | new_n19009_;
  assign new_n19011_ = ys__n19133 & ~ys__n18281;
  assign new_n19012_ = ~ys__n18278 & new_n19011_;
  assign new_n19013_ = ys__n18287 & new_n19012_;
  assign new_n19014_ = ~ys__n18284 & new_n19013_;
  assign new_n19015_ = ys__n19023 & ys__n18278;
  assign ys__n18500 = new_n19014_ | new_n19015_;
  assign new_n19017_ = ~ys__n18393 & ys__n18499;
  assign new_n19018_ = ys__n18393 & ys__n18500;
  assign ys__n18501 = new_n19017_ | new_n19018_;
  assign new_n19020_ = ys__n19134 & ~ys__n18281;
  assign new_n19021_ = ~ys__n18278 & new_n19020_;
  assign new_n19022_ = ys__n18287 & new_n19021_;
  assign new_n19023_ = ~ys__n18284 & new_n19022_;
  assign new_n19024_ = ys__n19025 & ys__n18278;
  assign ys__n18503 = new_n19023_ | new_n19024_;
  assign new_n19026_ = ~ys__n18393 & ys__n18502;
  assign new_n19027_ = ys__n18393 & ys__n18503;
  assign ys__n18504 = new_n19026_ | new_n19027_;
  assign new_n19029_ = ys__n19135 & ~ys__n18281;
  assign new_n19030_ = ~ys__n18278 & new_n19029_;
  assign new_n19031_ = ys__n18287 & new_n19030_;
  assign new_n19032_ = ~ys__n18284 & new_n19031_;
  assign new_n19033_ = ys__n19027 & ys__n18278;
  assign ys__n18506 = new_n19032_ | new_n19033_;
  assign new_n19035_ = ~ys__n18393 & ys__n18505;
  assign new_n19036_ = ys__n18393 & ys__n18506;
  assign ys__n18507 = new_n19035_ | new_n19036_;
  assign new_n19038_ = ys__n19136 & ~ys__n18281;
  assign new_n19039_ = ~ys__n18278 & new_n19038_;
  assign new_n19040_ = ys__n18287 & new_n19039_;
  assign new_n19041_ = ~ys__n18284 & new_n19040_;
  assign new_n19042_ = ys__n19029 & ys__n18278;
  assign ys__n18509 = new_n19041_ | new_n19042_;
  assign new_n19044_ = ~ys__n18393 & ys__n18508;
  assign new_n19045_ = ys__n18393 & ys__n18509;
  assign ys__n18510 = new_n19044_ | new_n19045_;
  assign new_n19047_ = ys__n19137 & ~ys__n18281;
  assign new_n19048_ = ~ys__n18278 & new_n19047_;
  assign new_n19049_ = ys__n18287 & new_n19048_;
  assign new_n19050_ = ~ys__n18284 & new_n19049_;
  assign new_n19051_ = ys__n19031 & ys__n18278;
  assign ys__n18512 = new_n19050_ | new_n19051_;
  assign new_n19053_ = ~ys__n18393 & ys__n18511;
  assign new_n19054_ = ys__n18393 & ys__n18512;
  assign ys__n18513 = new_n19053_ | new_n19054_;
  assign new_n19056_ = ys__n19138 & ~ys__n18281;
  assign new_n19057_ = ~ys__n18278 & new_n19056_;
  assign new_n19058_ = ys__n18287 & new_n19057_;
  assign new_n19059_ = ~ys__n18284 & new_n19058_;
  assign new_n19060_ = ys__n19033 & ys__n18278;
  assign ys__n18515 = new_n19059_ | new_n19060_;
  assign new_n19062_ = ~ys__n18393 & ys__n18514;
  assign new_n19063_ = ys__n18393 & ys__n18515;
  assign ys__n18516 = new_n19062_ | new_n19063_;
  assign new_n19065_ = ys__n19139 & ~ys__n18281;
  assign new_n19066_ = ~ys__n18278 & new_n19065_;
  assign new_n19067_ = ys__n18287 & new_n19066_;
  assign new_n19068_ = ~ys__n18284 & new_n19067_;
  assign new_n19069_ = ys__n19035 & ys__n18278;
  assign ys__n18518 = new_n19068_ | new_n19069_;
  assign new_n19071_ = ~ys__n18393 & ys__n18517;
  assign new_n19072_ = ys__n18393 & ys__n18518;
  assign ys__n18519 = new_n19071_ | new_n19072_;
  assign new_n19074_ = ys__n19140 & ~ys__n18281;
  assign new_n19075_ = ~ys__n18278 & new_n19074_;
  assign new_n19076_ = ys__n18287 & new_n19075_;
  assign new_n19077_ = ~ys__n18284 & new_n19076_;
  assign new_n19078_ = ys__n19037 & ys__n18278;
  assign ys__n18521 = new_n19077_ | new_n19078_;
  assign new_n19080_ = ~ys__n18393 & ys__n18520;
  assign new_n19081_ = ys__n18393 & ys__n18521;
  assign ys__n18522 = new_n19080_ | new_n19081_;
  assign new_n19083_ = ys__n19141 & ~ys__n18281;
  assign new_n19084_ = ~ys__n18278 & new_n19083_;
  assign new_n19085_ = ys__n18287 & new_n19084_;
  assign new_n19086_ = ~ys__n18284 & new_n19085_;
  assign new_n19087_ = ys__n19039 & ys__n18278;
  assign ys__n18524 = new_n19086_ | new_n19087_;
  assign new_n19089_ = ~ys__n18393 & ys__n18523;
  assign new_n19090_ = ys__n18393 & ys__n18524;
  assign ys__n18525 = new_n19089_ | new_n19090_;
  assign new_n19092_ = ys__n19142 & ~ys__n18281;
  assign new_n19093_ = ~ys__n18278 & new_n19092_;
  assign new_n19094_ = ys__n18287 & new_n19093_;
  assign new_n19095_ = ~ys__n18284 & new_n19094_;
  assign new_n19096_ = ys__n19041 & ys__n18278;
  assign ys__n18527 = new_n19095_ | new_n19096_;
  assign new_n19098_ = ~ys__n18393 & ys__n18526;
  assign new_n19099_ = ys__n18393 & ys__n18527;
  assign ys__n18528 = new_n19098_ | new_n19099_;
  assign new_n19101_ = ys__n19143 & ~ys__n18281;
  assign new_n19102_ = ~ys__n18278 & new_n19101_;
  assign new_n19103_ = ys__n18287 & new_n19102_;
  assign new_n19104_ = ~ys__n18284 & new_n19103_;
  assign new_n19105_ = ys__n19043 & ys__n18278;
  assign ys__n18530 = new_n19104_ | new_n19105_;
  assign new_n19107_ = ~ys__n18393 & ys__n18529;
  assign new_n19108_ = ys__n18393 & ys__n18530;
  assign ys__n18531 = new_n19107_ | new_n19108_;
  assign new_n19110_ = ys__n19144 & ~ys__n18281;
  assign new_n19111_ = ~ys__n18278 & new_n19110_;
  assign new_n19112_ = ys__n18287 & new_n19111_;
  assign new_n19113_ = ~ys__n18284 & new_n19112_;
  assign new_n19114_ = ys__n19045 & ys__n18278;
  assign ys__n18533 = new_n19113_ | new_n19114_;
  assign new_n19116_ = ~ys__n18393 & ys__n18532;
  assign new_n19117_ = ys__n18393 & ys__n18533;
  assign ys__n18534 = new_n19116_ | new_n19117_;
  assign new_n19119_ = ys__n19145 & ~ys__n18281;
  assign new_n19120_ = ~ys__n18278 & new_n19119_;
  assign new_n19121_ = ys__n18287 & new_n19120_;
  assign new_n19122_ = ~ys__n18284 & new_n19121_;
  assign new_n19123_ = ys__n19047 & ys__n18278;
  assign ys__n18536 = new_n19122_ | new_n19123_;
  assign new_n19125_ = ~ys__n18393 & ys__n18535;
  assign new_n19126_ = ys__n18393 & ys__n18536;
  assign ys__n18537 = new_n19125_ | new_n19126_;
  assign new_n19128_ = ys__n19146 & ~ys__n18281;
  assign new_n19129_ = ~ys__n18278 & new_n19128_;
  assign new_n19130_ = ys__n18287 & new_n19129_;
  assign new_n19131_ = ~ys__n18284 & new_n19130_;
  assign new_n19132_ = ys__n19049 & ys__n18278;
  assign ys__n18539 = new_n19131_ | new_n19132_;
  assign new_n19134_ = ~ys__n18393 & ys__n18538;
  assign new_n19135_ = ys__n18393 & ys__n18539;
  assign ys__n18540 = new_n19134_ | new_n19135_;
  assign new_n19137_ = ys__n19147 & ~ys__n18281;
  assign new_n19138_ = ~ys__n18278 & new_n19137_;
  assign new_n19139_ = ys__n18287 & new_n19138_;
  assign new_n19140_ = ~ys__n18284 & new_n19139_;
  assign new_n19141_ = ys__n19051 & ys__n18278;
  assign ys__n18542 = new_n19140_ | new_n19141_;
  assign new_n19143_ = ~ys__n18393 & ys__n18541;
  assign new_n19144_ = ys__n18393 & ys__n18542;
  assign ys__n18543 = new_n19143_ | new_n19144_;
  assign new_n19146_ = ys__n18281 & ~ys__n18278;
  assign ys__n18548 = ys__n18278 | new_n19146_;
  assign new_n19148_ = ys__n18065 & ~ys__n18393;
  assign new_n19149_ = ys__n18393 & ys__n18548;
  assign ys__n18549 = new_n19148_ | new_n19149_;
  assign new_n19151_ = ys__n19166 & ys__n18287;
  assign new_n19152_ = ~ys__n18284 & new_n19151_;
  assign new_n19153_ = ys__n18758 & ~new_n12256_;
  assign new_n19154_ = ys__n18759 & new_n12256_;
  assign ys__n18760 = new_n19153_ | new_n19154_;
  assign new_n19156_ = ys__n18284 & ys__n18760;
  assign new_n19157_ = ~new_n19152_ & ~new_n19156_;
  assign new_n19158_ = ~ys__n18281 & ~new_n19157_;
  assign new_n19159_ = ys__n18281 & ys__n18649;
  assign new_n19160_ = ~new_n19158_ & ~new_n19159_;
  assign ys__n18550 = ~ys__n18278 & ~new_n19160_;
  assign new_n19162_ = ys__n18059 & ~ys__n18393;
  assign new_n19163_ = ys__n18393 & ys__n18550;
  assign ys__n18551 = new_n19162_ | new_n19163_;
  assign ys__n19183 = ~new_n13277_ & ~ys__n18360;
  assign new_n19166_ = ~new_n13277_ & ~ys__n19183;
  assign new_n19167_ = new_n13204_ & ~new_n13261_;
  assign new_n19168_ = ~new_n19166_ & new_n19167_;
  assign new_n19169_ = new_n13204_ & ~new_n19168_;
  assign new_n19170_ = ~ys__n2 & ~new_n19169_;
  assign new_n19171_ = ~new_n13204_ & new_n13277_;
  assign new_n19172_ = new_n13277_ & ys__n18360;
  assign new_n19173_ = new_n13277_ & ~new_n19172_;
  assign new_n19174_ = new_n13261_ & ~new_n19173_;
  assign new_n19175_ = new_n13261_ & ~new_n19174_;
  assign new_n19176_ = new_n13204_ & ~new_n19175_;
  assign new_n19177_ = ~new_n19171_ & ~new_n19176_;
  assign new_n19178_ = ys__n2 & ~new_n19177_;
  assign ys__n18553 = new_n19170_ | new_n19178_;
  assign new_n19180_ = ys__n18277 & ~ys__n18393;
  assign new_n19181_ = ys__n18393 & ys__n18278;
  assign ys__n18554 = new_n19180_ | new_n19181_;
  assign new_n19183_ = ys__n18650 & ~new_n12259_;
  assign new_n19184_ = ys__n18651 & new_n12259_;
  assign ys__n18652 = new_n19183_ | new_n19184_;
  assign new_n19186_ = ys__n18761 & ~new_n12256_;
  assign new_n19187_ = ys__n18762 & new_n12256_;
  assign ys__n18763 = new_n19186_ | new_n19187_;
  assign new_n19189_ = ys__n124 & ~ys__n18303;
  assign new_n19190_ = ys__n4615 & ys__n18303;
  assign new_n19191_ = ~new_n19189_ & ~new_n19190_;
  assign ys__n19173 = ys__n874 & ~new_n19191_;
  assign new_n19193_ = ys__n126 & ~ys__n18303;
  assign new_n19194_ = ys__n714 & ys__n18303;
  assign new_n19195_ = ~new_n19193_ & ~new_n19194_;
  assign new_n19196_ = ys__n874 & ~new_n19195_;
  assign new_n19197_ = ys__n122 & ~ys__n18303;
  assign new_n19198_ = ys__n716 & ys__n18303;
  assign new_n19199_ = ~new_n19197_ & ~new_n19198_;
  assign new_n19200_ = ys__n874 & ~new_n19199_;
  assign new_n19201_ = new_n19196_ & ~new_n19200_;
  assign new_n19202_ = ys__n19173 & new_n19196_;
  assign new_n19203_ = new_n19200_ & new_n19202_;
  assign ys__n19177 = new_n19201_ | new_n19203_;
  assign new_n19205_ = ~ys__n19173 & ~new_n19200_;
  assign new_n19206_ = ys__n19173 & new_n19200_;
  assign ys__n19178 = new_n19205_ | new_n19206_;
  assign new_n19208_ = ys__n826 & new_n12861_;
  assign new_n19209_ = ~new_n12865_ & new_n19208_;
  assign new_n19210_ = ys__n822 & new_n12865_;
  assign ys__n19227 = new_n19209_ | new_n19210_;
  assign new_n19212_ = ys__n824 & new_n12861_;
  assign new_n19213_ = ~new_n12865_ & new_n19212_;
  assign new_n19214_ = ys__n820 & new_n12865_;
  assign ys__n19229 = new_n19213_ | new_n19214_;
  assign new_n19216_ = ys__n822 & new_n12861_;
  assign new_n19217_ = ~new_n12865_ & new_n19216_;
  assign new_n19218_ = ys__n818 & new_n12865_;
  assign ys__n19231 = new_n19217_ | new_n19218_;
  assign new_n19220_ = ys__n820 & new_n12861_;
  assign new_n19221_ = ~new_n12865_ & new_n19220_;
  assign new_n19222_ = ys__n816 & new_n12865_;
  assign ys__n19233 = new_n19221_ | new_n19222_;
  assign new_n19224_ = ys__n818 & new_n12861_;
  assign new_n19225_ = ~new_n12865_ & new_n19224_;
  assign new_n19226_ = ys__n1301 & new_n12865_;
  assign ys__n19235 = new_n19225_ | new_n19226_;
  assign new_n19228_ = ~ys__n27737 & ys__n732;
  assign new_n19229_ = new_n12860_ & new_n19228_;
  assign new_n19230_ = ~ys__n730 & new_n19229_;
  assign new_n19231_ = ~ys__n27737 & ~new_n12860_;
  assign new_n19232_ = ys__n4603 & new_n19231_;
  assign ys__n19239 = new_n19230_ | new_n19232_;
  assign new_n19234_ = ys__n19245 & ~ys__n19251;
  assign new_n19235_ = ~new_n11994_ & ~new_n19234_;
  assign new_n19236_ = ~ys__n19253 & ~new_n19235_;
  assign ys__n19254 = new_n11992_ | new_n19236_;
  assign new_n19238_ = ys__n19251 & new_n11968_;
  assign ys__n19257 = new_n12006_ | new_n19238_;
  assign new_n19240_ = ys__n140 & ~ys__n19259;
  assign new_n19241_ = ys__n19259 & ~ys__n19261;
  assign new_n19242_ = ~new_n19240_ & ~new_n19241_;
  assign new_n19243_ = ~ys__n19263 & ~new_n19242_;
  assign new_n19244_ = ys__n19263 & ys__n3039;
  assign ys__n19264 = new_n19243_ | new_n19244_;
  assign new_n19246_ = ys__n19259 & ys__n19261;
  assign new_n19247_ = ~ys__n19263 & new_n19246_;
  assign new_n19248_ = ys__n19263 & ~ys__n3039;
  assign ys__n19266 = new_n19247_ | new_n19248_;
  assign new_n19250_ = ~ys__n1505 & ~ys__n1506;
  assign new_n19251_ = ys__n19843 & ys__n19844;
  assign new_n19252_ = new_n19250_ & new_n19251_;
  assign new_n19253_ = ys__n23335 & ys__n27857;
  assign new_n19254_ = ~new_n11899_ & ~new_n19253_;
  assign new_n19255_ = ~ys__n23272 & ~new_n19254_;
  assign new_n19256_ = ~ys__n23335 & ys__n27859;
  assign new_n19257_ = ys__n23335 & ys__n27861;
  assign new_n19258_ = ~new_n19256_ & ~new_n19257_;
  assign new_n19259_ = ys__n23272 & ~new_n19258_;
  assign new_n19260_ = ~new_n19255_ & ~new_n19259_;
  assign new_n19261_ = ~ys__n23274 & ~new_n19260_;
  assign new_n19262_ = ~ys__n23335 & ys__n27863;
  assign new_n19263_ = ys__n23335 & ys__n27865;
  assign new_n19264_ = ~new_n19262_ & ~new_n19263_;
  assign new_n19265_ = ~ys__n23272 & ~new_n19264_;
  assign new_n19266_ = ~ys__n23335 & ys__n27867;
  assign new_n19267_ = ys__n23335 & ys__n27869;
  assign new_n19268_ = ~new_n19266_ & ~new_n19267_;
  assign new_n19269_ = ys__n23272 & ~new_n19268_;
  assign new_n19270_ = ~new_n19265_ & ~new_n19269_;
  assign new_n19271_ = ys__n23274 & ~new_n19270_;
  assign new_n19272_ = ~new_n19261_ & ~new_n19271_;
  assign new_n19273_ = ~ys__n23276 & ~new_n19272_;
  assign new_n19274_ = ~ys__n23335 & ys__n27871;
  assign new_n19275_ = ys__n23335 & ys__n27873;
  assign new_n19276_ = ~new_n19274_ & ~new_n19275_;
  assign new_n19277_ = ~ys__n23272 & ~new_n19276_;
  assign new_n19278_ = ~ys__n23335 & ys__n27875;
  assign new_n19279_ = ys__n23335 & ys__n27877;
  assign new_n19280_ = ~new_n19278_ & ~new_n19279_;
  assign new_n19281_ = ys__n23272 & ~new_n19280_;
  assign new_n19282_ = ~new_n19277_ & ~new_n19281_;
  assign new_n19283_ = ~ys__n23274 & ~new_n19282_;
  assign new_n19284_ = ~ys__n23335 & ys__n27879;
  assign new_n19285_ = ys__n23335 & ys__n27881;
  assign new_n19286_ = ~new_n19284_ & ~new_n19285_;
  assign new_n19287_ = ~ys__n23272 & ~new_n19286_;
  assign new_n19288_ = ~ys__n23335 & ys__n27883;
  assign new_n19289_ = ys__n23335 & ys__n27885;
  assign new_n19290_ = ~new_n19288_ & ~new_n19289_;
  assign new_n19291_ = ys__n23272 & ~new_n19290_;
  assign new_n19292_ = ~new_n19287_ & ~new_n19291_;
  assign new_n19293_ = ys__n23274 & ~new_n19292_;
  assign new_n19294_ = ~new_n19283_ & ~new_n19293_;
  assign new_n19295_ = ys__n23276 & ~new_n19294_;
  assign new_n19296_ = ~new_n19273_ & ~new_n19295_;
  assign new_n19297_ = ~ys__n23278 & ~new_n19296_;
  assign new_n19298_ = ~ys__n23335 & ys__n28015;
  assign new_n19299_ = ys__n23335 & ys__n28016;
  assign new_n19300_ = ~new_n19298_ & ~new_n19299_;
  assign new_n19301_ = ~ys__n23272 & ~new_n19300_;
  assign new_n19302_ = ~ys__n23335 & ys__n28017;
  assign new_n19303_ = ys__n23335 & ys__n28018;
  assign new_n19304_ = ~new_n19302_ & ~new_n19303_;
  assign new_n19305_ = ys__n23272 & ~new_n19304_;
  assign new_n19306_ = ~new_n19301_ & ~new_n19305_;
  assign new_n19307_ = ~ys__n23274 & ~new_n19306_;
  assign new_n19308_ = ~ys__n23335 & ys__n28019;
  assign new_n19309_ = ys__n23335 & ys__n28020;
  assign new_n19310_ = ~new_n19308_ & ~new_n19309_;
  assign new_n19311_ = ~ys__n23272 & ~new_n19310_;
  assign new_n19312_ = ~ys__n23335 & ys__n28021;
  assign new_n19313_ = ys__n23335 & ys__n28022;
  assign new_n19314_ = ~new_n19312_ & ~new_n19313_;
  assign new_n19315_ = ys__n23272 & ~new_n19314_;
  assign new_n19316_ = ~new_n19311_ & ~new_n19315_;
  assign new_n19317_ = ys__n23274 & ~new_n19316_;
  assign new_n19318_ = ~new_n19307_ & ~new_n19317_;
  assign new_n19319_ = ~ys__n23276 & ~new_n19318_;
  assign new_n19320_ = ~ys__n23335 & ys__n28023;
  assign new_n19321_ = ys__n23335 & ys__n28024;
  assign new_n19322_ = ~new_n19320_ & ~new_n19321_;
  assign new_n19323_ = ~ys__n23272 & ~new_n19322_;
  assign new_n19324_ = ~ys__n23335 & ys__n28025;
  assign new_n19325_ = ys__n23335 & ys__n28026;
  assign new_n19326_ = ~new_n19324_ & ~new_n19325_;
  assign new_n19327_ = ys__n23272 & ~new_n19326_;
  assign new_n19328_ = ~new_n19323_ & ~new_n19327_;
  assign new_n19329_ = ~ys__n23274 & ~new_n19328_;
  assign new_n19330_ = ~ys__n23335 & ys__n28027;
  assign new_n19331_ = ys__n23335 & ys__n28028;
  assign new_n19332_ = ~new_n19330_ & ~new_n19331_;
  assign new_n19333_ = ~ys__n23272 & ~new_n19332_;
  assign new_n19334_ = ~ys__n23335 & ys__n28029;
  assign new_n19335_ = ys__n23335 & ys__n28030;
  assign new_n19336_ = ~new_n19334_ & ~new_n19335_;
  assign new_n19337_ = ys__n23272 & ~new_n19336_;
  assign new_n19338_ = ~new_n19333_ & ~new_n19337_;
  assign new_n19339_ = ys__n23274 & ~new_n19338_;
  assign new_n19340_ = ~new_n19329_ & ~new_n19339_;
  assign new_n19341_ = ys__n23276 & ~new_n19340_;
  assign new_n19342_ = ~new_n19319_ & ~new_n19341_;
  assign new_n19343_ = ys__n23278 & ~new_n19342_;
  assign new_n19344_ = ~new_n19297_ & ~new_n19343_;
  assign new_n19345_ = ~new_n19250_ & ~new_n19344_;
  assign new_n19346_ = ~new_n19252_ & ~new_n19345_;
  assign new_n19347_ = ~ys__n1502 & ~ys__n1503;
  assign new_n19348_ = ~new_n19346_ & new_n19347_;
  assign new_n19349_ = ~ys__n23272 & new_n11899_;
  assign new_n19350_ = ~ys__n23274 & new_n19349_;
  assign new_n19351_ = ~ys__n23276 & new_n19350_;
  assign new_n19352_ = ys__n1502 & ~ys__n23278;
  assign new_n19353_ = ~new_n19347_ & new_n19352_;
  assign new_n19354_ = new_n19351_ & new_n19353_;
  assign new_n19355_ = ~new_n19348_ & ~new_n19354_;
  assign new_n19356_ = ~ys__n1495 & ~ys__n1496;
  assign new_n19357_ = ~ys__n1498 & ~ys__n1499;
  assign new_n19358_ = new_n19356_ & new_n19357_;
  assign new_n19359_ = ~new_n19355_ & new_n19358_;
  assign new_n19360_ = ~ys__n1498 & ys__n1499;
  assign new_n19361_ = ~new_n11901_ & new_n19360_;
  assign new_n19362_ = ~ys__n23335 & ~ys__n27855;
  assign new_n19363_ = ys__n1498 & new_n19362_;
  assign new_n19364_ = ~new_n19361_ & ~new_n19363_;
  assign new_n19365_ = ~ys__n1496 & ~new_n19364_;
  assign new_n19366_ = ys__n1496 & ~new_n19362_;
  assign new_n19367_ = ~new_n19365_ & ~new_n19366_;
  assign new_n19368_ = ~ys__n1495 & ~new_n19367_;
  assign new_n19369_ = ys__n1495 & new_n17743_;
  assign new_n19370_ = ~new_n19368_ & ~new_n19369_;
  assign new_n19371_ = ~new_n19358_ & ~new_n19370_;
  assign new_n19372_ = ~new_n19359_ & ~new_n19371_;
  assign new_n19373_ = ~ys__n1492 & ~ys__n1493;
  assign new_n19374_ = ~new_n19372_ & new_n19373_;
  assign new_n19375_ = ~ys__n1492 & ys__n23332;
  assign new_n19376_ = ~ys__n1492 & ys__n28030;
  assign new_n19377_ = ~new_n19375_ & ~new_n19376_;
  assign new_n19378_ = new_n19375_ & new_n19376_;
  assign new_n19379_ = ~new_n19377_ & ~new_n19378_;
  assign new_n19380_ = ~ys__n23272 & ~ys__n27857;
  assign new_n19381_ = ~new_n17911_ & ~new_n19380_;
  assign new_n19382_ = ~new_n17743_ & ~new_n19362_;
  assign new_n19383_ = ~new_n11900_ & new_n19382_;
  assign new_n19384_ = ~new_n19381_ & ~new_n19383_;
  assign new_n19385_ = ~new_n11903_ & ~new_n19384_;
  assign new_n19386_ = ~ys__n23276 & ~ys__n27861;
  assign new_n19387_ = ~new_n17916_ & ~new_n19386_;
  assign new_n19388_ = ~ys__n23274 & ~ys__n27859;
  assign new_n19389_ = ~new_n17917_ & ~new_n19388_;
  assign new_n19390_ = ~new_n19387_ & ~new_n19389_;
  assign new_n19391_ = ~new_n19385_ & new_n19390_;
  assign new_n19392_ = new_n11907_ & ~new_n19387_;
  assign new_n19393_ = ~new_n11910_ & ~new_n19392_;
  assign new_n19394_ = ~new_n19391_ & new_n19393_;
  assign new_n19395_ = ~ys__n23284 & ~ys__n27869;
  assign new_n19396_ = ~new_n17930_ & ~new_n19395_;
  assign new_n19397_ = ~ys__n23282 & ~ys__n27867;
  assign new_n19398_ = ~new_n17931_ & ~new_n19397_;
  assign new_n19399_ = ~new_n19396_ & ~new_n19398_;
  assign new_n19400_ = ~ys__n23280 & ~ys__n27865;
  assign new_n19401_ = ~new_n17925_ & ~new_n19400_;
  assign new_n19402_ = ~ys__n23278 & ~ys__n27863;
  assign new_n19403_ = ~new_n17926_ & ~new_n19402_;
  assign new_n19404_ = ~new_n19401_ & ~new_n19403_;
  assign new_n19405_ = new_n19399_ & new_n19404_;
  assign new_n19406_ = ~new_n19394_ & new_n19405_;
  assign new_n19407_ = new_n11885_ & ~new_n19401_;
  assign new_n19408_ = ~new_n11888_ & ~new_n19407_;
  assign new_n19409_ = new_n19399_ & ~new_n19408_;
  assign new_n19410_ = new_n11892_ & ~new_n19396_;
  assign new_n19411_ = ~new_n11895_ & ~new_n19410_;
  assign new_n19412_ = ~new_n19409_ & new_n19411_;
  assign new_n19413_ = ~new_n19406_ & new_n19412_;
  assign new_n19414_ = ~ys__n23300 & ~ys__n27885;
  assign new_n19415_ = ~new_n17960_ & ~new_n19414_;
  assign new_n19416_ = ~ys__n23298 & ~ys__n27883;
  assign new_n19417_ = ~new_n17961_ & ~new_n19416_;
  assign new_n19418_ = ~new_n19415_ & ~new_n19417_;
  assign new_n19419_ = ~ys__n23296 & ~ys__n27881;
  assign new_n19420_ = ~new_n17955_ & ~new_n19419_;
  assign new_n19421_ = ~ys__n23294 & ~ys__n27879;
  assign new_n19422_ = ~new_n17956_ & ~new_n19421_;
  assign new_n19423_ = ~new_n19420_ & ~new_n19422_;
  assign new_n19424_ = new_n19418_ & new_n19423_;
  assign new_n19425_ = ~ys__n23292 & ~ys__n27877;
  assign new_n19426_ = ~new_n17949_ & ~new_n19425_;
  assign new_n19427_ = ~ys__n23290 & ~ys__n27875;
  assign new_n19428_ = ~new_n17950_ & ~new_n19427_;
  assign new_n19429_ = ~new_n19426_ & ~new_n19428_;
  assign new_n19430_ = ~ys__n23288 & ~ys__n27873;
  assign new_n19431_ = ~new_n17944_ & ~new_n19430_;
  assign new_n19432_ = ~ys__n23286 & ~ys__n27871;
  assign new_n19433_ = ~new_n17945_ & ~new_n19432_;
  assign new_n19434_ = ~new_n19431_ & ~new_n19433_;
  assign new_n19435_ = new_n19429_ & new_n19434_;
  assign new_n19436_ = new_n19424_ & new_n19435_;
  assign new_n19437_ = ~new_n19413_ & new_n19436_;
  assign new_n19438_ = new_n11931_ & ~new_n19431_;
  assign new_n19439_ = ~new_n11934_ & ~new_n19438_;
  assign new_n19440_ = new_n19429_ & ~new_n19439_;
  assign new_n19441_ = new_n11938_ & ~new_n19426_;
  assign new_n19442_ = ~new_n11941_ & ~new_n19441_;
  assign new_n19443_ = ~new_n19440_ & new_n19442_;
  assign new_n19444_ = new_n19424_ & ~new_n19443_;
  assign new_n19445_ = new_n11916_ & ~new_n19420_;
  assign new_n19446_ = ~new_n11919_ & ~new_n19445_;
  assign new_n19447_ = new_n19418_ & ~new_n19446_;
  assign new_n19448_ = new_n11923_ & ~new_n19415_;
  assign new_n19449_ = ~new_n11926_ & ~new_n19448_;
  assign new_n19450_ = ~new_n19447_ & new_n19449_;
  assign new_n19451_ = ~new_n19444_ & new_n19450_;
  assign new_n19452_ = ~new_n19437_ & new_n19451_;
  assign new_n19453_ = ~ys__n23332 & ~ys__n28030;
  assign new_n19454_ = ys__n23332 & ys__n28030;
  assign new_n19455_ = ~new_n19453_ & ~new_n19454_;
  assign new_n19456_ = ~ys__n23330 & ~ys__n28029;
  assign new_n19457_ = ~new_n17990_ & ~new_n19456_;
  assign new_n19458_ = ~new_n19455_ & ~new_n19457_;
  assign new_n19459_ = ~ys__n23328 & ~ys__n28028;
  assign new_n19460_ = ~new_n17978_ & ~new_n19459_;
  assign new_n19461_ = ~ys__n23326 & ~ys__n28027;
  assign new_n19462_ = ~new_n17868_ & ~new_n19461_;
  assign new_n19463_ = ~new_n19460_ & ~new_n19462_;
  assign new_n19464_ = new_n19458_ & new_n19463_;
  assign new_n19465_ = ~ys__n23324 & ~ys__n28026;
  assign new_n19466_ = ~new_n17875_ & ~new_n19465_;
  assign new_n19467_ = ~ys__n23322 & ~ys__n28025;
  assign new_n19468_ = ~new_n17876_ & ~new_n19467_;
  assign new_n19469_ = ~new_n19466_ & ~new_n19468_;
  assign new_n19470_ = ~ys__n23320 & ~ys__n28024;
  assign new_n19471_ = ~new_n17870_ & ~new_n19470_;
  assign new_n19472_ = ~ys__n23318 & ~ys__n28023;
  assign new_n19473_ = ~new_n17871_ & ~new_n19472_;
  assign new_n19474_ = ~new_n19471_ & ~new_n19473_;
  assign new_n19475_ = new_n19469_ & new_n19474_;
  assign new_n19476_ = new_n19464_ & new_n19475_;
  assign new_n19477_ = ~ys__n23316 & ~ys__n28022;
  assign new_n19478_ = ~new_n17902_ & ~new_n19477_;
  assign new_n19479_ = ~ys__n23314 & ~ys__n28021;
  assign new_n19480_ = ~new_n17903_ & ~new_n19479_;
  assign new_n19481_ = ~new_n19478_ & ~new_n19480_;
  assign new_n19482_ = ~ys__n23312 & ~ys__n28020;
  assign new_n19483_ = ~new_n17897_ & ~new_n19482_;
  assign new_n19484_ = ~ys__n23310 & ~ys__n28019;
  assign new_n19485_ = ~new_n17898_ & ~new_n19484_;
  assign new_n19486_ = ~new_n19483_ & ~new_n19485_;
  assign new_n19487_ = new_n19481_ & new_n19486_;
  assign new_n19488_ = ~ys__n23308 & ~ys__n28018;
  assign new_n19489_ = ~new_n17891_ & ~new_n19488_;
  assign new_n19490_ = ~ys__n23306 & ~ys__n28017;
  assign new_n19491_ = ~new_n17892_ & ~new_n19490_;
  assign new_n19492_ = ~new_n19489_ & ~new_n19491_;
  assign new_n19493_ = ~ys__n23304 & ~ys__n28016;
  assign new_n19494_ = ~new_n17886_ & ~new_n19493_;
  assign new_n19495_ = ~ys__n23302 & ~ys__n28015;
  assign new_n19496_ = ~new_n17887_ & ~new_n19495_;
  assign new_n19497_ = ~new_n19494_ & ~new_n19496_;
  assign new_n19498_ = new_n19492_ & new_n19497_;
  assign new_n19499_ = new_n19487_ & new_n19498_;
  assign new_n19500_ = new_n19476_ & new_n19499_;
  assign new_n19501_ = ~new_n19452_ & new_n19500_;
  assign new_n19502_ = new_n11837_ & ~new_n19494_;
  assign new_n19503_ = ~new_n11840_ & ~new_n19502_;
  assign new_n19504_ = new_n19492_ & ~new_n19503_;
  assign new_n19505_ = new_n11844_ & ~new_n19489_;
  assign new_n19506_ = ~new_n11847_ & ~new_n19505_;
  assign new_n19507_ = ~new_n19504_ & new_n19506_;
  assign new_n19508_ = new_n19487_ & ~new_n19507_;
  assign new_n19509_ = new_n11822_ & ~new_n19483_;
  assign new_n19510_ = ~new_n11825_ & ~new_n19509_;
  assign new_n19511_ = new_n19481_ & ~new_n19510_;
  assign new_n19512_ = new_n11829_ & ~new_n19478_;
  assign new_n19513_ = ~new_n11832_ & ~new_n19512_;
  assign new_n19514_ = ~new_n19511_ & new_n19513_;
  assign new_n19515_ = ~new_n19508_ & new_n19514_;
  assign new_n19516_ = new_n19476_ & ~new_n19515_;
  assign new_n19517_ = new_n11868_ & ~new_n19471_;
  assign new_n19518_ = ~new_n11871_ & ~new_n19517_;
  assign new_n19519_ = new_n19469_ & ~new_n19518_;
  assign new_n19520_ = new_n11875_ & ~new_n19466_;
  assign new_n19521_ = ~new_n11878_ & ~new_n19520_;
  assign new_n19522_ = ~new_n19519_ & new_n19521_;
  assign new_n19523_ = new_n19464_ & ~new_n19522_;
  assign new_n19524_ = new_n11853_ & ~new_n19460_;
  assign new_n19525_ = ~new_n11856_ & ~new_n19524_;
  assign new_n19526_ = new_n19458_ & ~new_n19525_;
  assign new_n19527_ = new_n11860_ & ~new_n19455_;
  assign new_n19528_ = ~new_n11863_ & ~new_n19527_;
  assign new_n19529_ = ~new_n19526_ & new_n19528_;
  assign new_n19530_ = ~new_n19523_ & new_n19529_;
  assign new_n19531_ = ~new_n19516_ & new_n19530_;
  assign new_n19532_ = ~new_n19501_ & new_n19531_;
  assign new_n19533_ = new_n19379_ & ~new_n19532_;
  assign new_n19534_ = ~new_n19379_ & new_n19532_;
  assign new_n19535_ = ~new_n19533_ & ~new_n19534_;
  assign new_n19536_ = ~ys__n1489 & ~new_n19535_;
  assign new_n19537_ = ~new_n19375_ & new_n19376_;
  assign new_n19538_ = new_n19375_ & ~new_n19376_;
  assign new_n19539_ = ~new_n19537_ & ~new_n19538_;
  assign new_n19540_ = ~new_n11861_ & ~new_n11864_;
  assign new_n19541_ = new_n17981_ & new_n19540_;
  assign new_n19542_ = new_n17881_ & new_n19541_;
  assign new_n19543_ = new_n17910_ & new_n19542_;
  assign new_n19544_ = ~new_n17966_ & new_n19543_;
  assign new_n19545_ = ~new_n17907_ & new_n19542_;
  assign new_n19546_ = ~new_n17879_ & new_n19541_;
  assign new_n19547_ = ~new_n17980_ & new_n19540_;
  assign new_n19548_ = ~new_n11864_ & new_n17990_;
  assign new_n19549_ = ~new_n19454_ & ~new_n19548_;
  assign new_n19550_ = ~new_n19547_ & new_n19549_;
  assign new_n19551_ = ~new_n19546_ & new_n19550_;
  assign new_n19552_ = ~new_n19545_ & new_n19551_;
  assign new_n19553_ = ~new_n19544_ & new_n19552_;
  assign new_n19554_ = new_n19539_ & ~new_n19553_;
  assign new_n19555_ = ~new_n19539_ & new_n19553_;
  assign new_n19556_ = ~new_n19554_ & ~new_n19555_;
  assign new_n19557_ = ys__n1489 & ~new_n19556_;
  assign new_n19558_ = ~new_n19536_ & ~new_n19557_;
  assign new_n19559_ = ~new_n19373_ & ~new_n19558_;
  assign new_n19560_ = ~new_n19374_ & ~new_n19559_;
  assign new_n19561_ = ~ys__n1489 & ~ys__n1490;
  assign new_n19562_ = ~new_n19560_ & new_n19561_;
  assign new_n19563_ = ~ys__n1489 & new_n19382_;
  assign new_n19564_ = ys__n1489 & ~new_n11901_;
  assign new_n19565_ = ~new_n19563_ & ~new_n19564_;
  assign new_n19566_ = ~new_n19561_ & ~new_n19565_;
  assign new_n19567_ = ~new_n19562_ & ~new_n19566_;
  assign new_n19568_ = ~ys__n19973 & ~new_n19567_;
  assign new_n19569_ = ys__n19972 & ys__n19973;
  assign new_n19570_ = ~new_n19568_ & ~new_n19569_;
  assign new_n19571_ = ~ys__n352 & ~new_n19570_;
  assign new_n19572_ = ~ys__n220 & ys__n47026;
  assign new_n19573_ = ys__n222 & ys__n248;
  assign new_n19574_ = new_n19572_ & new_n19573_;
  assign new_n19575_ = ys__n222 & ~ys__n248;
  assign new_n19576_ = ~ys__n220 & ys__n47074;
  assign new_n19577_ = new_n19575_ & new_n19576_;
  assign new_n19578_ = ~ys__n222 & ys__n248;
  assign new_n19579_ = ~ys__n220 & ys__n47010;
  assign new_n19580_ = new_n19578_ & new_n19579_;
  assign new_n19581_ = ~new_n19577_ & ~new_n19580_;
  assign new_n19582_ = ~new_n19574_ & new_n19581_;
  assign new_n19583_ = ~new_n19575_ & ~new_n19578_;
  assign new_n19584_ = ~ys__n222 & ~ys__n248;
  assign new_n19585_ = ~new_n19573_ & ~new_n19584_;
  assign new_n19586_ = new_n19583_ & new_n19585_;
  assign new_n19587_ = ys__n352 & ~new_n19586_;
  assign new_n19588_ = ~new_n19582_ & new_n19587_;
  assign ys__n19878 = new_n19571_ | new_n19588_;
  assign new_n19590_ = ys__n19844 & ys__n19845;
  assign new_n19591_ = new_n19250_ & new_n19590_;
  assign new_n19592_ = ~ys__n23335 & ys__n27857;
  assign new_n19593_ = ys__n23335 & ys__n27859;
  assign new_n19594_ = ~new_n19592_ & ~new_n19593_;
  assign new_n19595_ = ~ys__n23272 & ~new_n19594_;
  assign new_n19596_ = ~ys__n23335 & ys__n27861;
  assign new_n19597_ = ys__n23335 & ys__n27863;
  assign new_n19598_ = ~new_n19596_ & ~new_n19597_;
  assign new_n19599_ = ys__n23272 & ~new_n19598_;
  assign new_n19600_ = ~new_n19595_ & ~new_n19599_;
  assign new_n19601_ = ~ys__n23274 & ~new_n19600_;
  assign new_n19602_ = ~ys__n23335 & ys__n27865;
  assign new_n19603_ = ys__n23335 & ys__n27867;
  assign new_n19604_ = ~new_n19602_ & ~new_n19603_;
  assign new_n19605_ = ~ys__n23272 & ~new_n19604_;
  assign new_n19606_ = ~ys__n23335 & ys__n27869;
  assign new_n19607_ = ys__n23335 & ys__n27871;
  assign new_n19608_ = ~new_n19606_ & ~new_n19607_;
  assign new_n19609_ = ys__n23272 & ~new_n19608_;
  assign new_n19610_ = ~new_n19605_ & ~new_n19609_;
  assign new_n19611_ = ys__n23274 & ~new_n19610_;
  assign new_n19612_ = ~new_n19601_ & ~new_n19611_;
  assign new_n19613_ = ~ys__n23276 & ~new_n19612_;
  assign new_n19614_ = ~ys__n23335 & ys__n27873;
  assign new_n19615_ = ys__n23335 & ys__n27875;
  assign new_n19616_ = ~new_n19614_ & ~new_n19615_;
  assign new_n19617_ = ~ys__n23272 & ~new_n19616_;
  assign new_n19618_ = ~ys__n23335 & ys__n27877;
  assign new_n19619_ = ys__n23335 & ys__n27879;
  assign new_n19620_ = ~new_n19618_ & ~new_n19619_;
  assign new_n19621_ = ys__n23272 & ~new_n19620_;
  assign new_n19622_ = ~new_n19617_ & ~new_n19621_;
  assign new_n19623_ = ~ys__n23274 & ~new_n19622_;
  assign new_n19624_ = ~ys__n23335 & ys__n27881;
  assign new_n19625_ = ys__n23335 & ys__n27883;
  assign new_n19626_ = ~new_n19624_ & ~new_n19625_;
  assign new_n19627_ = ~ys__n23272 & ~new_n19626_;
  assign new_n19628_ = ~ys__n23335 & ys__n27885;
  assign new_n19629_ = ys__n23335 & ys__n28015;
  assign new_n19630_ = ~new_n19628_ & ~new_n19629_;
  assign new_n19631_ = ys__n23272 & ~new_n19630_;
  assign new_n19632_ = ~new_n19627_ & ~new_n19631_;
  assign new_n19633_ = ys__n23274 & ~new_n19632_;
  assign new_n19634_ = ~new_n19623_ & ~new_n19633_;
  assign new_n19635_ = ys__n23276 & ~new_n19634_;
  assign new_n19636_ = ~new_n19613_ & ~new_n19635_;
  assign new_n19637_ = ~ys__n23278 & ~new_n19636_;
  assign new_n19638_ = ~ys__n23335 & ys__n28016;
  assign new_n19639_ = ys__n23335 & ys__n28017;
  assign new_n19640_ = ~new_n19638_ & ~new_n19639_;
  assign new_n19641_ = ~ys__n23272 & ~new_n19640_;
  assign new_n19642_ = ~ys__n23335 & ys__n28018;
  assign new_n19643_ = ys__n23335 & ys__n28019;
  assign new_n19644_ = ~new_n19642_ & ~new_n19643_;
  assign new_n19645_ = ys__n23272 & ~new_n19644_;
  assign new_n19646_ = ~new_n19641_ & ~new_n19645_;
  assign new_n19647_ = ~ys__n23274 & ~new_n19646_;
  assign new_n19648_ = ~ys__n23335 & ys__n28020;
  assign new_n19649_ = ys__n23335 & ys__n28021;
  assign new_n19650_ = ~new_n19648_ & ~new_n19649_;
  assign new_n19651_ = ~ys__n23272 & ~new_n19650_;
  assign new_n19652_ = ~ys__n23335 & ys__n28022;
  assign new_n19653_ = ys__n23335 & ys__n28023;
  assign new_n19654_ = ~new_n19652_ & ~new_n19653_;
  assign new_n19655_ = ys__n23272 & ~new_n19654_;
  assign new_n19656_ = ~new_n19651_ & ~new_n19655_;
  assign new_n19657_ = ys__n23274 & ~new_n19656_;
  assign new_n19658_ = ~new_n19647_ & ~new_n19657_;
  assign new_n19659_ = ~ys__n23276 & ~new_n19658_;
  assign new_n19660_ = ~ys__n23335 & ys__n28024;
  assign new_n19661_ = ys__n23335 & ys__n28025;
  assign new_n19662_ = ~new_n19660_ & ~new_n19661_;
  assign new_n19663_ = ~ys__n23272 & ~new_n19662_;
  assign new_n19664_ = ~ys__n23335 & ys__n28026;
  assign new_n19665_ = ys__n23335 & ys__n28027;
  assign new_n19666_ = ~new_n19664_ & ~new_n19665_;
  assign new_n19667_ = ys__n23272 & ~new_n19666_;
  assign new_n19668_ = ~new_n19663_ & ~new_n19667_;
  assign new_n19669_ = ~ys__n23274 & ~new_n19668_;
  assign new_n19670_ = ~ys__n23335 & ys__n28028;
  assign new_n19671_ = ys__n23335 & ys__n28029;
  assign new_n19672_ = ~new_n19670_ & ~new_n19671_;
  assign new_n19673_ = ~ys__n23272 & ~new_n19672_;
  assign new_n19674_ = ys__n23272 & ys__n28030;
  assign new_n19675_ = ~new_n19673_ & ~new_n19674_;
  assign new_n19676_ = ys__n23274 & ~new_n19675_;
  assign new_n19677_ = ~new_n19669_ & ~new_n19676_;
  assign new_n19678_ = ys__n23276 & ~new_n19677_;
  assign new_n19679_ = ~new_n19659_ & ~new_n19678_;
  assign new_n19680_ = ys__n23278 & ~new_n19679_;
  assign new_n19681_ = ~new_n19637_ & ~new_n19680_;
  assign new_n19682_ = ~ys__n1505 & ~new_n19681_;
  assign new_n19683_ = ~ys__n23335 & ys__n28030;
  assign new_n19684_ = ys__n23272 & new_n19683_;
  assign new_n19685_ = ~new_n19673_ & ~new_n19684_;
  assign new_n19686_ = ys__n23274 & ~new_n19685_;
  assign new_n19687_ = ~new_n19669_ & ~new_n19686_;
  assign new_n19688_ = ys__n23276 & ~new_n19687_;
  assign new_n19689_ = ~new_n19659_ & ~new_n19688_;
  assign new_n19690_ = ys__n23278 & ~new_n19689_;
  assign new_n19691_ = ~new_n19637_ & ~new_n19690_;
  assign new_n19692_ = ys__n1505 & ~new_n19691_;
  assign new_n19693_ = ~new_n19682_ & ~new_n19692_;
  assign new_n19694_ = ~new_n19250_ & ~new_n19693_;
  assign new_n19695_ = ~new_n19591_ & ~new_n19694_;
  assign new_n19696_ = new_n19347_ & ~new_n19695_;
  assign new_n19697_ = ~new_n17743_ & ~new_n19592_;
  assign new_n19698_ = ~ys__n23272 & ~new_n19697_;
  assign new_n19699_ = ~ys__n23274 & new_n19698_;
  assign new_n19700_ = ~ys__n23276 & new_n19699_;
  assign new_n19701_ = new_n19353_ & new_n19700_;
  assign new_n19702_ = ~new_n19696_ & ~new_n19701_;
  assign new_n19703_ = new_n19358_ & ~new_n19702_;
  assign new_n19704_ = ~new_n11904_ & new_n19360_;
  assign new_n19705_ = ys__n1498 & new_n19380_;
  assign new_n19706_ = ~new_n19704_ & ~new_n19705_;
  assign new_n19707_ = ~ys__n1496 & ~new_n19706_;
  assign new_n19708_ = ys__n1496 & ~new_n19380_;
  assign new_n19709_ = ~new_n19707_ & ~new_n19708_;
  assign new_n19710_ = ~ys__n1495 & ~new_n19709_;
  assign new_n19711_ = ys__n1495 & new_n17911_;
  assign new_n19712_ = ~new_n19710_ & ~new_n19711_;
  assign new_n19713_ = ~new_n19358_ & ~new_n19712_;
  assign new_n19714_ = ~new_n19703_ & ~new_n19713_;
  assign new_n19715_ = new_n19373_ & new_n19561_;
  assign new_n19716_ = ~new_n19714_ & new_n19715_;
  assign new_n19717_ = new_n19381_ & ~new_n19383_;
  assign new_n19718_ = ~new_n19381_ & new_n19383_;
  assign new_n19719_ = ~new_n19717_ & ~new_n19718_;
  assign new_n19720_ = ~ys__n1489 & ~new_n19719_;
  assign new_n19721_ = ys__n1489 & ~new_n17746_;
  assign new_n19722_ = ~new_n19720_ & ~new_n19721_;
  assign new_n19723_ = ~new_n19561_ & ~new_n19722_;
  assign new_n19724_ = ~new_n19716_ & ~new_n19723_;
  assign new_n19725_ = ~ys__n19973 & ~new_n19724_;
  assign new_n19726_ = ys__n19973 & ys__n19974;
  assign new_n19727_ = ~new_n19725_ & ~new_n19726_;
  assign new_n19728_ = ~ys__n352 & ~new_n19727_;
  assign new_n19729_ = ~ys__n220 & ys__n47027;
  assign new_n19730_ = new_n19573_ & new_n19729_;
  assign new_n19731_ = ~ys__n220 & ys__n47075;
  assign new_n19732_ = new_n19575_ & new_n19731_;
  assign new_n19733_ = ~ys__n220 & ys__n47011;
  assign new_n19734_ = new_n19578_ & new_n19733_;
  assign new_n19735_ = ~new_n19732_ & ~new_n19734_;
  assign new_n19736_ = ~new_n19730_ & new_n19735_;
  assign new_n19737_ = new_n19587_ & ~new_n19736_;
  assign ys__n19881 = new_n19728_ | new_n19737_;
  assign new_n19739_ = ys__n19844 & ys__n19846;
  assign new_n19740_ = new_n19250_ & new_n19739_;
  assign new_n19741_ = ~ys__n23272 & ~new_n19258_;
  assign new_n19742_ = ys__n23272 & ~new_n19264_;
  assign new_n19743_ = ~new_n19741_ & ~new_n19742_;
  assign new_n19744_ = ~ys__n23274 & ~new_n19743_;
  assign new_n19745_ = ~ys__n23272 & ~new_n19268_;
  assign new_n19746_ = ys__n23272 & ~new_n19276_;
  assign new_n19747_ = ~new_n19745_ & ~new_n19746_;
  assign new_n19748_ = ys__n23274 & ~new_n19747_;
  assign new_n19749_ = ~new_n19744_ & ~new_n19748_;
  assign new_n19750_ = ~ys__n23276 & ~new_n19749_;
  assign new_n19751_ = ~ys__n23272 & ~new_n19280_;
  assign new_n19752_ = ys__n23272 & ~new_n19286_;
  assign new_n19753_ = ~new_n19751_ & ~new_n19752_;
  assign new_n19754_ = ~ys__n23274 & ~new_n19753_;
  assign new_n19755_ = ~ys__n23272 & ~new_n19290_;
  assign new_n19756_ = ys__n23272 & ~new_n19300_;
  assign new_n19757_ = ~new_n19755_ & ~new_n19756_;
  assign new_n19758_ = ys__n23274 & ~new_n19757_;
  assign new_n19759_ = ~new_n19754_ & ~new_n19758_;
  assign new_n19760_ = ys__n23276 & ~new_n19759_;
  assign new_n19761_ = ~new_n19750_ & ~new_n19760_;
  assign new_n19762_ = ~ys__n23278 & ~new_n19761_;
  assign new_n19763_ = ~ys__n23272 & ~new_n19304_;
  assign new_n19764_ = ys__n23272 & ~new_n19310_;
  assign new_n19765_ = ~new_n19763_ & ~new_n19764_;
  assign new_n19766_ = ~ys__n23274 & ~new_n19765_;
  assign new_n19767_ = ~ys__n23272 & ~new_n19314_;
  assign new_n19768_ = ys__n23272 & ~new_n19322_;
  assign new_n19769_ = ~new_n19767_ & ~new_n19768_;
  assign new_n19770_ = ys__n23274 & ~new_n19769_;
  assign new_n19771_ = ~new_n19766_ & ~new_n19770_;
  assign new_n19772_ = ~ys__n23276 & ~new_n19771_;
  assign new_n19773_ = ~ys__n23272 & ~new_n19326_;
  assign new_n19774_ = ys__n23272 & ~new_n19332_;
  assign new_n19775_ = ~new_n19773_ & ~new_n19774_;
  assign new_n19776_ = ~ys__n23274 & ~new_n19775_;
  assign new_n19777_ = ~ys__n23272 & ~new_n19336_;
  assign new_n19778_ = ~new_n19674_ & ~new_n19777_;
  assign new_n19779_ = ys__n23274 & ~new_n19778_;
  assign new_n19780_ = ~new_n19776_ & ~new_n19779_;
  assign new_n19781_ = ys__n23276 & ~new_n19780_;
  assign new_n19782_ = ~new_n19772_ & ~new_n19781_;
  assign new_n19783_ = ys__n23278 & ~new_n19782_;
  assign new_n19784_ = ~new_n19762_ & ~new_n19783_;
  assign new_n19785_ = ~ys__n1505 & ~new_n19784_;
  assign new_n19786_ = ys__n23274 & new_n19777_;
  assign new_n19787_ = ~new_n19776_ & ~new_n19786_;
  assign new_n19788_ = ys__n23276 & ~new_n19787_;
  assign new_n19789_ = ~new_n19772_ & ~new_n19788_;
  assign new_n19790_ = ys__n23278 & ~new_n19789_;
  assign new_n19791_ = ~new_n19762_ & ~new_n19790_;
  assign new_n19792_ = ys__n1505 & ~new_n19791_;
  assign new_n19793_ = ~new_n19785_ & ~new_n19792_;
  assign new_n19794_ = ~new_n19250_ & ~new_n19793_;
  assign new_n19795_ = ~new_n19740_ & ~new_n19794_;
  assign new_n19796_ = new_n19347_ & ~new_n19795_;
  assign new_n19797_ = ~new_n19253_ & ~new_n19256_;
  assign new_n19798_ = ~ys__n23272 & ~new_n19797_;
  assign new_n19799_ = ys__n23272 & new_n11899_;
  assign new_n19800_ = ~new_n19798_ & ~new_n19799_;
  assign new_n19801_ = ~ys__n23274 & ~new_n19800_;
  assign new_n19802_ = ~ys__n23276 & new_n19801_;
  assign new_n19803_ = new_n19353_ & new_n19802_;
  assign new_n19804_ = ~new_n19796_ & ~new_n19803_;
  assign new_n19805_ = new_n19358_ & ~new_n19804_;
  assign new_n19806_ = ~new_n11908_ & new_n19360_;
  assign new_n19807_ = ys__n1498 & new_n19388_;
  assign new_n19808_ = ~new_n19806_ & ~new_n19807_;
  assign new_n19809_ = ~ys__n1496 & ~new_n19808_;
  assign new_n19810_ = ys__n1496 & ~new_n19388_;
  assign new_n19811_ = ~new_n19809_ & ~new_n19810_;
  assign new_n19812_ = ~ys__n1495 & ~new_n19811_;
  assign new_n19813_ = ys__n1495 & new_n17917_;
  assign new_n19814_ = ~new_n19812_ & ~new_n19813_;
  assign new_n19815_ = ~new_n19358_ & ~new_n19814_;
  assign new_n19816_ = ~new_n19805_ & ~new_n19815_;
  assign new_n19817_ = new_n19715_ & ~new_n19816_;
  assign new_n19818_ = ~new_n19385_ & new_n19389_;
  assign new_n19819_ = new_n19385_ & ~new_n19389_;
  assign new_n19820_ = ~new_n19818_ & ~new_n19819_;
  assign new_n19821_ = ~ys__n1489 & ~new_n19820_;
  assign new_n19822_ = new_n11908_ & ~new_n17913_;
  assign new_n19823_ = ~new_n11908_ & new_n17913_;
  assign new_n19824_ = ~new_n19822_ & ~new_n19823_;
  assign new_n19825_ = ys__n1489 & ~new_n19824_;
  assign new_n19826_ = ~new_n19821_ & ~new_n19825_;
  assign new_n19827_ = ~new_n19561_ & ~new_n19826_;
  assign new_n19828_ = ~new_n19817_ & ~new_n19827_;
  assign new_n19829_ = ~ys__n19973 & ~new_n19828_;
  assign new_n19830_ = ys__n19973 & ys__n19975;
  assign new_n19831_ = ~new_n19829_ & ~new_n19830_;
  assign new_n19832_ = ~ys__n352 & ~new_n19831_;
  assign new_n19833_ = ~ys__n220 & ys__n47028;
  assign new_n19834_ = new_n19573_ & new_n19833_;
  assign new_n19835_ = ~ys__n220 & ys__n47076;
  assign new_n19836_ = new_n19575_ & new_n19835_;
  assign new_n19837_ = ~ys__n220 & ys__n47012;
  assign new_n19838_ = new_n19578_ & new_n19837_;
  assign new_n19839_ = ~new_n19836_ & ~new_n19838_;
  assign new_n19840_ = ~new_n19834_ & new_n19839_;
  assign new_n19841_ = new_n19587_ & ~new_n19840_;
  assign ys__n19884 = new_n19832_ | new_n19841_;
  assign new_n19843_ = ys__n19844 & ys__n19847;
  assign new_n19844_ = new_n19250_ & new_n19843_;
  assign new_n19845_ = ~ys__n23272 & ~new_n19598_;
  assign new_n19846_ = ys__n23272 & ~new_n19604_;
  assign new_n19847_ = ~new_n19845_ & ~new_n19846_;
  assign new_n19848_ = ~ys__n23274 & ~new_n19847_;
  assign new_n19849_ = ~ys__n23272 & ~new_n19608_;
  assign new_n19850_ = ys__n23272 & ~new_n19616_;
  assign new_n19851_ = ~new_n19849_ & ~new_n19850_;
  assign new_n19852_ = ys__n23274 & ~new_n19851_;
  assign new_n19853_ = ~new_n19848_ & ~new_n19852_;
  assign new_n19854_ = ~ys__n23276 & ~new_n19853_;
  assign new_n19855_ = ~ys__n23272 & ~new_n19620_;
  assign new_n19856_ = ys__n23272 & ~new_n19626_;
  assign new_n19857_ = ~new_n19855_ & ~new_n19856_;
  assign new_n19858_ = ~ys__n23274 & ~new_n19857_;
  assign new_n19859_ = ~ys__n23272 & ~new_n19630_;
  assign new_n19860_ = ys__n23272 & ~new_n19640_;
  assign new_n19861_ = ~new_n19859_ & ~new_n19860_;
  assign new_n19862_ = ys__n23274 & ~new_n19861_;
  assign new_n19863_ = ~new_n19858_ & ~new_n19862_;
  assign new_n19864_ = ys__n23276 & ~new_n19863_;
  assign new_n19865_ = ~new_n19854_ & ~new_n19864_;
  assign new_n19866_ = ~ys__n23278 & ~new_n19865_;
  assign new_n19867_ = ~ys__n23272 & ~new_n19644_;
  assign new_n19868_ = ys__n23272 & ~new_n19650_;
  assign new_n19869_ = ~new_n19867_ & ~new_n19868_;
  assign new_n19870_ = ~ys__n23274 & ~new_n19869_;
  assign new_n19871_ = ~ys__n23272 & ~new_n19654_;
  assign new_n19872_ = ys__n23272 & ~new_n19662_;
  assign new_n19873_ = ~new_n19871_ & ~new_n19872_;
  assign new_n19874_ = ys__n23274 & ~new_n19873_;
  assign new_n19875_ = ~new_n19870_ & ~new_n19874_;
  assign new_n19876_ = ~ys__n23276 & ~new_n19875_;
  assign new_n19877_ = ~ys__n23272 & ~new_n19666_;
  assign new_n19878_ = ys__n23272 & ~new_n19672_;
  assign new_n19879_ = ~new_n19877_ & ~new_n19878_;
  assign new_n19880_ = ~ys__n23274 & ~new_n19879_;
  assign new_n19881_ = ys__n23274 & ys__n28030;
  assign new_n19882_ = ~new_n19880_ & ~new_n19881_;
  assign new_n19883_ = ys__n23276 & ~new_n19882_;
  assign new_n19884_ = ~new_n19876_ & ~new_n19883_;
  assign new_n19885_ = ys__n23278 & ~new_n19884_;
  assign new_n19886_ = ~new_n19866_ & ~new_n19885_;
  assign new_n19887_ = ~ys__n1505 & ~new_n19886_;
  assign new_n19888_ = ~ys__n23272 & new_n19683_;
  assign new_n19889_ = ys__n23274 & new_n19888_;
  assign new_n19890_ = ~new_n19880_ & ~new_n19889_;
  assign new_n19891_ = ys__n23276 & ~new_n19890_;
  assign new_n19892_ = ~new_n19876_ & ~new_n19891_;
  assign new_n19893_ = ys__n23278 & ~new_n19892_;
  assign new_n19894_ = ~new_n19866_ & ~new_n19893_;
  assign new_n19895_ = ys__n1505 & ~new_n19894_;
  assign new_n19896_ = ~new_n19887_ & ~new_n19895_;
  assign new_n19897_ = ~new_n19250_ & ~new_n19896_;
  assign new_n19898_ = ~new_n19844_ & ~new_n19897_;
  assign new_n19899_ = new_n19347_ & ~new_n19898_;
  assign new_n19900_ = ~new_n19593_ & ~new_n19596_;
  assign new_n19901_ = ~ys__n23272 & ~new_n19900_;
  assign new_n19902_ = ys__n23272 & ~new_n19697_;
  assign new_n19903_ = ~new_n19901_ & ~new_n19902_;
  assign new_n19904_ = ~ys__n23274 & ~new_n19903_;
  assign new_n19905_ = ~ys__n23276 & new_n19904_;
  assign new_n19906_ = new_n19353_ & new_n19905_;
  assign new_n19907_ = ~new_n19899_ & ~new_n19906_;
  assign new_n19908_ = new_n19358_ & ~new_n19907_;
  assign new_n19909_ = ~new_n11911_ & new_n19360_;
  assign new_n19910_ = ys__n1498 & new_n19386_;
  assign new_n19911_ = ~new_n19909_ & ~new_n19910_;
  assign new_n19912_ = ~ys__n1496 & ~new_n19911_;
  assign new_n19913_ = ys__n1496 & ~new_n19386_;
  assign new_n19914_ = ~new_n19912_ & ~new_n19913_;
  assign new_n19915_ = ~ys__n1495 & ~new_n19914_;
  assign new_n19916_ = ys__n1495 & new_n17916_;
  assign new_n19917_ = ~new_n19915_ & ~new_n19916_;
  assign new_n19918_ = ~new_n19358_ & ~new_n19917_;
  assign new_n19919_ = ~new_n19908_ & ~new_n19918_;
  assign new_n19920_ = new_n19715_ & ~new_n19919_;
  assign new_n19921_ = ~new_n19385_ & ~new_n19389_;
  assign new_n19922_ = ~new_n11907_ & ~new_n19921_;
  assign new_n19923_ = new_n19387_ & ~new_n19922_;
  assign new_n19924_ = ~new_n19387_ & new_n19922_;
  assign new_n19925_ = ~new_n19923_ & ~new_n19924_;
  assign new_n19926_ = ~ys__n1489 & ~new_n19925_;
  assign new_n19927_ = ~new_n11908_ & ~new_n17913_;
  assign new_n19928_ = ~new_n17917_ & ~new_n19927_;
  assign new_n19929_ = new_n11911_ & ~new_n19928_;
  assign new_n19930_ = ~new_n11911_ & new_n19928_;
  assign new_n19931_ = ~new_n19929_ & ~new_n19930_;
  assign new_n19932_ = ys__n1489 & ~new_n19931_;
  assign new_n19933_ = ~new_n19926_ & ~new_n19932_;
  assign new_n19934_ = ~new_n19561_ & ~new_n19933_;
  assign new_n19935_ = ~new_n19920_ & ~new_n19934_;
  assign new_n19936_ = ~ys__n19973 & ~new_n19935_;
  assign new_n19937_ = ys__n19973 & ys__n19976;
  assign new_n19938_ = ~new_n19936_ & ~new_n19937_;
  assign new_n19939_ = ~ys__n352 & ~new_n19938_;
  assign new_n19940_ = ~ys__n220 & ys__n47029;
  assign new_n19941_ = new_n19573_ & new_n19940_;
  assign new_n19942_ = ~ys__n220 & ys__n47077;
  assign new_n19943_ = new_n19575_ & new_n19942_;
  assign new_n19944_ = ~ys__n220 & ys__n47013;
  assign new_n19945_ = new_n19578_ & new_n19944_;
  assign new_n19946_ = ~new_n19943_ & ~new_n19945_;
  assign new_n19947_ = ~new_n19941_ & new_n19946_;
  assign new_n19948_ = new_n19587_ & ~new_n19947_;
  assign ys__n19887 = new_n19939_ | new_n19948_;
  assign new_n19950_ = ys__n19844 & ys__n19848;
  assign new_n19951_ = new_n19250_ & new_n19950_;
  assign new_n19952_ = ~ys__n23274 & ~new_n19270_;
  assign new_n19953_ = ys__n23274 & ~new_n19282_;
  assign new_n19954_ = ~new_n19952_ & ~new_n19953_;
  assign new_n19955_ = ~ys__n23276 & ~new_n19954_;
  assign new_n19956_ = ~ys__n23274 & ~new_n19292_;
  assign new_n19957_ = ys__n23274 & ~new_n19306_;
  assign new_n19958_ = ~new_n19956_ & ~new_n19957_;
  assign new_n19959_ = ys__n23276 & ~new_n19958_;
  assign new_n19960_ = ~new_n19955_ & ~new_n19959_;
  assign new_n19961_ = ~ys__n23278 & ~new_n19960_;
  assign new_n19962_ = ~ys__n23274 & ~new_n19316_;
  assign new_n19963_ = ys__n23274 & ~new_n19328_;
  assign new_n19964_ = ~new_n19962_ & ~new_n19963_;
  assign new_n19965_ = ~ys__n23276 & ~new_n19964_;
  assign new_n19966_ = ~ys__n23274 & ~new_n19338_;
  assign new_n19967_ = ~new_n19881_ & ~new_n19966_;
  assign new_n19968_ = ys__n23276 & ~new_n19967_;
  assign new_n19969_ = ~new_n19965_ & ~new_n19968_;
  assign new_n19970_ = ys__n23278 & ~new_n19969_;
  assign new_n19971_ = ~new_n19961_ & ~new_n19970_;
  assign new_n19972_ = ~ys__n1505 & ~new_n19971_;
  assign new_n19973_ = ys__n23276 & new_n19966_;
  assign new_n19974_ = ~new_n19965_ & ~new_n19973_;
  assign new_n19975_ = ys__n23278 & ~new_n19974_;
  assign new_n19976_ = ~new_n19961_ & ~new_n19975_;
  assign new_n19977_ = ys__n1505 & ~new_n19976_;
  assign new_n19978_ = ~new_n19972_ & ~new_n19977_;
  assign new_n19979_ = ~new_n19250_ & ~new_n19978_;
  assign new_n19980_ = ~new_n19951_ & ~new_n19979_;
  assign new_n19981_ = new_n19347_ & ~new_n19980_;
  assign new_n19982_ = ~new_n19257_ & ~new_n19262_;
  assign new_n19983_ = ~ys__n23272 & ~new_n19982_;
  assign new_n19984_ = ys__n23272 & ~new_n19797_;
  assign new_n19985_ = ~new_n19983_ & ~new_n19984_;
  assign new_n19986_ = ~ys__n23274 & ~new_n19985_;
  assign new_n19987_ = ys__n23274 & new_n19349_;
  assign new_n19988_ = ~new_n19986_ & ~new_n19987_;
  assign new_n19989_ = ~ys__n23276 & ~new_n19988_;
  assign new_n19990_ = new_n19353_ & new_n19989_;
  assign new_n19991_ = ~new_n19981_ & ~new_n19990_;
  assign new_n19992_ = new_n19358_ & ~new_n19991_;
  assign new_n19993_ = ~new_n11886_ & new_n19360_;
  assign new_n19994_ = ys__n1498 & new_n19402_;
  assign new_n19995_ = ~new_n19993_ & ~new_n19994_;
  assign new_n19996_ = ~ys__n1496 & ~new_n19995_;
  assign new_n19997_ = ys__n1496 & ~new_n19402_;
  assign new_n19998_ = ~new_n19996_ & ~new_n19997_;
  assign new_n19999_ = ~ys__n1495 & ~new_n19998_;
  assign new_n20000_ = ys__n1495 & new_n17926_;
  assign new_n20001_ = ~new_n19999_ & ~new_n20000_;
  assign new_n20002_ = ~new_n19358_ & ~new_n20001_;
  assign new_n20003_ = ~new_n19992_ & ~new_n20002_;
  assign new_n20004_ = new_n19715_ & ~new_n20003_;
  assign new_n20005_ = ~new_n19394_ & new_n19403_;
  assign new_n20006_ = new_n19394_ & ~new_n19403_;
  assign new_n20007_ = ~new_n20005_ & ~new_n20006_;
  assign new_n20008_ = ~ys__n1489 & ~new_n20007_;
  assign new_n20009_ = new_n11886_ & ~new_n17920_;
  assign new_n20010_ = ~new_n11886_ & new_n17920_;
  assign new_n20011_ = ~new_n20009_ & ~new_n20010_;
  assign new_n20012_ = ys__n1489 & ~new_n20011_;
  assign new_n20013_ = ~new_n20008_ & ~new_n20012_;
  assign new_n20014_ = ~new_n19561_ & ~new_n20013_;
  assign new_n20015_ = ~new_n20004_ & ~new_n20014_;
  assign new_n20016_ = ~ys__n19973 & ~new_n20015_;
  assign new_n20017_ = ys__n19973 & ys__n19977;
  assign new_n20018_ = ~new_n20016_ & ~new_n20017_;
  assign new_n20019_ = ~ys__n352 & ~new_n20018_;
  assign new_n20020_ = ~ys__n220 & ys__n47030;
  assign new_n20021_ = new_n19573_ & new_n20020_;
  assign new_n20022_ = ~ys__n220 & ys__n47078;
  assign new_n20023_ = new_n19575_ & new_n20022_;
  assign new_n20024_ = ~ys__n220 & ys__n47014;
  assign new_n20025_ = new_n19578_ & new_n20024_;
  assign new_n20026_ = ~new_n20023_ & ~new_n20025_;
  assign new_n20027_ = ~new_n20021_ & new_n20026_;
  assign new_n20028_ = new_n19587_ & ~new_n20027_;
  assign ys__n19890 = new_n20019_ | new_n20028_;
  assign new_n20030_ = ys__n19844 & ys__n19849;
  assign new_n20031_ = new_n19250_ & new_n20030_;
  assign new_n20032_ = ~ys__n23274 & ~new_n19610_;
  assign new_n20033_ = ys__n23274 & ~new_n19622_;
  assign new_n20034_ = ~new_n20032_ & ~new_n20033_;
  assign new_n20035_ = ~ys__n23276 & ~new_n20034_;
  assign new_n20036_ = ~ys__n23274 & ~new_n19632_;
  assign new_n20037_ = ys__n23274 & ~new_n19646_;
  assign new_n20038_ = ~new_n20036_ & ~new_n20037_;
  assign new_n20039_ = ys__n23276 & ~new_n20038_;
  assign new_n20040_ = ~new_n20035_ & ~new_n20039_;
  assign new_n20041_ = ~ys__n23278 & ~new_n20040_;
  assign new_n20042_ = ~ys__n23274 & ~new_n19656_;
  assign new_n20043_ = ys__n23274 & ~new_n19668_;
  assign new_n20044_ = ~new_n20042_ & ~new_n20043_;
  assign new_n20045_ = ~ys__n23276 & ~new_n20044_;
  assign new_n20046_ = ~ys__n23274 & ~new_n19675_;
  assign new_n20047_ = ~new_n19881_ & ~new_n20046_;
  assign new_n20048_ = ys__n23276 & ~new_n20047_;
  assign new_n20049_ = ~new_n20045_ & ~new_n20048_;
  assign new_n20050_ = ys__n23278 & ~new_n20049_;
  assign new_n20051_ = ~new_n20041_ & ~new_n20050_;
  assign new_n20052_ = ~ys__n1505 & ~new_n20051_;
  assign new_n20053_ = ~ys__n23274 & ~new_n19685_;
  assign new_n20054_ = ys__n23276 & new_n20053_;
  assign new_n20055_ = ~new_n20045_ & ~new_n20054_;
  assign new_n20056_ = ys__n23278 & ~new_n20055_;
  assign new_n20057_ = ~new_n20041_ & ~new_n20056_;
  assign new_n20058_ = ys__n1505 & ~new_n20057_;
  assign new_n20059_ = ~new_n20052_ & ~new_n20058_;
  assign new_n20060_ = ~new_n19250_ & ~new_n20059_;
  assign new_n20061_ = ~new_n20031_ & ~new_n20060_;
  assign new_n20062_ = new_n19347_ & ~new_n20061_;
  assign new_n20063_ = ~new_n19597_ & ~new_n19602_;
  assign new_n20064_ = ~ys__n23272 & ~new_n20063_;
  assign new_n20065_ = ys__n23272 & ~new_n19900_;
  assign new_n20066_ = ~new_n20064_ & ~new_n20065_;
  assign new_n20067_ = ~ys__n23274 & ~new_n20066_;
  assign new_n20068_ = ys__n23274 & new_n19698_;
  assign new_n20069_ = ~new_n20067_ & ~new_n20068_;
  assign new_n20070_ = ~ys__n23276 & ~new_n20069_;
  assign new_n20071_ = new_n19353_ & new_n20070_;
  assign new_n20072_ = ~new_n20062_ & ~new_n20071_;
  assign new_n20073_ = new_n19358_ & ~new_n20072_;
  assign new_n20074_ = ~new_n11889_ & new_n19360_;
  assign new_n20075_ = ys__n1498 & new_n19400_;
  assign new_n20076_ = ~new_n20074_ & ~new_n20075_;
  assign new_n20077_ = ~ys__n1496 & ~new_n20076_;
  assign new_n20078_ = ys__n1496 & ~new_n19400_;
  assign new_n20079_ = ~new_n20077_ & ~new_n20078_;
  assign new_n20080_ = ~ys__n1495 & ~new_n20079_;
  assign new_n20081_ = ys__n1495 & new_n17925_;
  assign new_n20082_ = ~new_n20080_ & ~new_n20081_;
  assign new_n20083_ = ~new_n19358_ & ~new_n20082_;
  assign new_n20084_ = ~new_n20073_ & ~new_n20083_;
  assign new_n20085_ = new_n19715_ & ~new_n20084_;
  assign new_n20086_ = ~new_n19394_ & ~new_n19403_;
  assign new_n20087_ = ~new_n11885_ & ~new_n20086_;
  assign new_n20088_ = new_n19401_ & ~new_n20087_;
  assign new_n20089_ = ~new_n19401_ & new_n20087_;
  assign new_n20090_ = ~new_n20088_ & ~new_n20089_;
  assign new_n20091_ = ~ys__n1489 & ~new_n20090_;
  assign new_n20092_ = ~new_n11886_ & ~new_n17920_;
  assign new_n20093_ = ~new_n17926_ & ~new_n20092_;
  assign new_n20094_ = new_n11889_ & ~new_n20093_;
  assign new_n20095_ = ~new_n11889_ & new_n20093_;
  assign new_n20096_ = ~new_n20094_ & ~new_n20095_;
  assign new_n20097_ = ys__n1489 & ~new_n20096_;
  assign new_n20098_ = ~new_n20091_ & ~new_n20097_;
  assign new_n20099_ = ~new_n19561_ & ~new_n20098_;
  assign new_n20100_ = ~new_n20085_ & ~new_n20099_;
  assign new_n20101_ = ~ys__n19973 & ~new_n20100_;
  assign new_n20102_ = ys__n19973 & ys__n19978;
  assign new_n20103_ = ~new_n20101_ & ~new_n20102_;
  assign new_n20104_ = ~ys__n352 & ~new_n20103_;
  assign new_n20105_ = ~ys__n220 & ys__n47031;
  assign new_n20106_ = new_n19573_ & new_n20105_;
  assign new_n20107_ = ~ys__n220 & ys__n47079;
  assign new_n20108_ = new_n19575_ & new_n20107_;
  assign new_n20109_ = ~ys__n220 & ys__n47015;
  assign new_n20110_ = new_n19578_ & new_n20109_;
  assign new_n20111_ = ~new_n20108_ & ~new_n20110_;
  assign new_n20112_ = ~new_n20106_ & new_n20111_;
  assign new_n20113_ = new_n19587_ & ~new_n20112_;
  assign ys__n19893 = new_n20104_ | new_n20113_;
  assign new_n20115_ = ys__n19844 & ys__n19850;
  assign new_n20116_ = new_n19250_ & new_n20115_;
  assign new_n20117_ = ~ys__n23274 & ~new_n19747_;
  assign new_n20118_ = ys__n23274 & ~new_n19753_;
  assign new_n20119_ = ~new_n20117_ & ~new_n20118_;
  assign new_n20120_ = ~ys__n23276 & ~new_n20119_;
  assign new_n20121_ = ~ys__n23274 & ~new_n19757_;
  assign new_n20122_ = ys__n23274 & ~new_n19765_;
  assign new_n20123_ = ~new_n20121_ & ~new_n20122_;
  assign new_n20124_ = ys__n23276 & ~new_n20123_;
  assign new_n20125_ = ~new_n20120_ & ~new_n20124_;
  assign new_n20126_ = ~ys__n23278 & ~new_n20125_;
  assign new_n20127_ = ~ys__n23274 & ~new_n19769_;
  assign new_n20128_ = ys__n23274 & ~new_n19775_;
  assign new_n20129_ = ~new_n20127_ & ~new_n20128_;
  assign new_n20130_ = ~ys__n23276 & ~new_n20129_;
  assign new_n20131_ = ~ys__n23274 & ~new_n19778_;
  assign new_n20132_ = ~new_n19881_ & ~new_n20131_;
  assign new_n20133_ = ys__n23276 & ~new_n20132_;
  assign new_n20134_ = ~new_n20130_ & ~new_n20133_;
  assign new_n20135_ = ys__n23278 & ~new_n20134_;
  assign new_n20136_ = ~new_n20126_ & ~new_n20135_;
  assign new_n20137_ = ~ys__n1505 & ~new_n20136_;
  assign new_n20138_ = ~ys__n23274 & new_n19777_;
  assign new_n20139_ = ys__n23276 & new_n20138_;
  assign new_n20140_ = ~new_n20130_ & ~new_n20139_;
  assign new_n20141_ = ys__n23278 & ~new_n20140_;
  assign new_n20142_ = ~new_n20126_ & ~new_n20141_;
  assign new_n20143_ = ys__n1505 & ~new_n20142_;
  assign new_n20144_ = ~new_n20137_ & ~new_n20143_;
  assign new_n20145_ = ~new_n19250_ & ~new_n20144_;
  assign new_n20146_ = ~new_n20116_ & ~new_n20145_;
  assign new_n20147_ = new_n19347_ & ~new_n20146_;
  assign new_n20148_ = ~new_n19263_ & ~new_n19266_;
  assign new_n20149_ = ~ys__n23272 & ~new_n20148_;
  assign new_n20150_ = ys__n23272 & ~new_n19982_;
  assign new_n20151_ = ~new_n20149_ & ~new_n20150_;
  assign new_n20152_ = ~ys__n23274 & ~new_n20151_;
  assign new_n20153_ = ys__n23274 & ~new_n19800_;
  assign new_n20154_ = ~new_n20152_ & ~new_n20153_;
  assign new_n20155_ = ~ys__n23276 & ~new_n20154_;
  assign new_n20156_ = new_n19353_ & new_n20155_;
  assign new_n20157_ = ~new_n20147_ & ~new_n20156_;
  assign new_n20158_ = new_n19358_ & ~new_n20157_;
  assign new_n20159_ = ~new_n11893_ & new_n19360_;
  assign new_n20160_ = ys__n1498 & new_n19397_;
  assign new_n20161_ = ~new_n20159_ & ~new_n20160_;
  assign new_n20162_ = ~ys__n1496 & ~new_n20161_;
  assign new_n20163_ = ys__n1496 & ~new_n19397_;
  assign new_n20164_ = ~new_n20162_ & ~new_n20163_;
  assign new_n20165_ = ~ys__n1495 & ~new_n20164_;
  assign new_n20166_ = ys__n1495 & new_n17931_;
  assign new_n20167_ = ~new_n20165_ & ~new_n20166_;
  assign new_n20168_ = ~new_n19358_ & ~new_n20167_;
  assign new_n20169_ = ~new_n20158_ & ~new_n20168_;
  assign new_n20170_ = new_n19715_ & ~new_n20169_;
  assign new_n20171_ = ~new_n19394_ & new_n19404_;
  assign new_n20172_ = new_n19408_ & ~new_n20171_;
  assign new_n20173_ = new_n19398_ & ~new_n20172_;
  assign new_n20174_ = ~new_n19398_ & new_n20172_;
  assign new_n20175_ = ~new_n20173_ & ~new_n20174_;
  assign new_n20176_ = ~ys__n1489 & ~new_n20175_;
  assign new_n20177_ = ~new_n17920_ & new_n17922_;
  assign new_n20178_ = new_n17928_ & ~new_n20177_;
  assign new_n20179_ = new_n11893_ & ~new_n20178_;
  assign new_n20180_ = ~new_n11893_ & new_n20178_;
  assign new_n20181_ = ~new_n20179_ & ~new_n20180_;
  assign new_n20182_ = ys__n1489 & ~new_n20181_;
  assign new_n20183_ = ~new_n20176_ & ~new_n20182_;
  assign new_n20184_ = ~new_n19561_ & ~new_n20183_;
  assign new_n20185_ = ~new_n20170_ & ~new_n20184_;
  assign new_n20186_ = ~ys__n19973 & ~new_n20185_;
  assign new_n20187_ = ys__n19973 & ys__n19979;
  assign new_n20188_ = ~new_n20186_ & ~new_n20187_;
  assign new_n20189_ = ~ys__n352 & ~new_n20188_;
  assign new_n20190_ = ~ys__n220 & ys__n47032;
  assign new_n20191_ = new_n19573_ & new_n20190_;
  assign new_n20192_ = ~ys__n220 & ys__n47080;
  assign new_n20193_ = new_n19575_ & new_n20192_;
  assign new_n20194_ = ~ys__n220 & ys__n47016;
  assign new_n20195_ = new_n19578_ & new_n20194_;
  assign new_n20196_ = ~new_n20193_ & ~new_n20195_;
  assign new_n20197_ = ~new_n20191_ & new_n20196_;
  assign new_n20198_ = new_n19587_ & ~new_n20197_;
  assign ys__n19896 = new_n20189_ | new_n20198_;
  assign new_n20200_ = ys__n19844 & ys__n19851;
  assign new_n20201_ = new_n19250_ & new_n20200_;
  assign new_n20202_ = ~ys__n23274 & ~new_n19851_;
  assign new_n20203_ = ys__n23274 & ~new_n19857_;
  assign new_n20204_ = ~new_n20202_ & ~new_n20203_;
  assign new_n20205_ = ~ys__n23276 & ~new_n20204_;
  assign new_n20206_ = ~ys__n23274 & ~new_n19861_;
  assign new_n20207_ = ys__n23274 & ~new_n19869_;
  assign new_n20208_ = ~new_n20206_ & ~new_n20207_;
  assign new_n20209_ = ys__n23276 & ~new_n20208_;
  assign new_n20210_ = ~new_n20205_ & ~new_n20209_;
  assign new_n20211_ = ~ys__n23278 & ~new_n20210_;
  assign new_n20212_ = ~ys__n23274 & ~new_n19873_;
  assign new_n20213_ = ys__n23274 & ~new_n19879_;
  assign new_n20214_ = ~new_n20212_ & ~new_n20213_;
  assign new_n20215_ = ~ys__n23276 & ~new_n20214_;
  assign new_n20216_ = ys__n23276 & ys__n28030;
  assign new_n20217_ = ~new_n20215_ & ~new_n20216_;
  assign new_n20218_ = ys__n23278 & ~new_n20217_;
  assign new_n20219_ = ~new_n20211_ & ~new_n20218_;
  assign new_n20220_ = ~ys__n1505 & ~new_n20219_;
  assign new_n20221_ = ~ys__n23274 & new_n19888_;
  assign new_n20222_ = ys__n23276 & new_n20221_;
  assign new_n20223_ = ~new_n20215_ & ~new_n20222_;
  assign new_n20224_ = ys__n23278 & ~new_n20223_;
  assign new_n20225_ = ~new_n20211_ & ~new_n20224_;
  assign new_n20226_ = ys__n1505 & ~new_n20225_;
  assign new_n20227_ = ~new_n20220_ & ~new_n20226_;
  assign new_n20228_ = ~new_n19250_ & ~new_n20227_;
  assign new_n20229_ = ~new_n20201_ & ~new_n20228_;
  assign new_n20230_ = new_n19347_ & ~new_n20229_;
  assign new_n20231_ = ~new_n19603_ & ~new_n19606_;
  assign new_n20232_ = ~ys__n23272 & ~new_n20231_;
  assign new_n20233_ = ys__n23272 & ~new_n20063_;
  assign new_n20234_ = ~new_n20232_ & ~new_n20233_;
  assign new_n20235_ = ~ys__n23274 & ~new_n20234_;
  assign new_n20236_ = ys__n23274 & ~new_n19903_;
  assign new_n20237_ = ~new_n20235_ & ~new_n20236_;
  assign new_n20238_ = ~ys__n23276 & ~new_n20237_;
  assign new_n20239_ = new_n19353_ & new_n20238_;
  assign new_n20240_ = ~new_n20230_ & ~new_n20239_;
  assign new_n20241_ = new_n19358_ & ~new_n20240_;
  assign new_n20242_ = ~new_n11896_ & new_n19360_;
  assign new_n20243_ = ys__n1498 & new_n19395_;
  assign new_n20244_ = ~new_n20242_ & ~new_n20243_;
  assign new_n20245_ = ~ys__n1496 & ~new_n20244_;
  assign new_n20246_ = ys__n1496 & ~new_n19395_;
  assign new_n20247_ = ~new_n20245_ & ~new_n20246_;
  assign new_n20248_ = ~ys__n1495 & ~new_n20247_;
  assign new_n20249_ = ys__n1495 & new_n17930_;
  assign new_n20250_ = ~new_n20248_ & ~new_n20249_;
  assign new_n20251_ = ~new_n19358_ & ~new_n20250_;
  assign new_n20252_ = ~new_n20241_ & ~new_n20251_;
  assign new_n20253_ = new_n19715_ & ~new_n20252_;
  assign new_n20254_ = ~new_n19398_ & ~new_n20172_;
  assign new_n20255_ = ~new_n11892_ & ~new_n20254_;
  assign new_n20256_ = new_n19396_ & ~new_n20255_;
  assign new_n20257_ = ~new_n19396_ & new_n20255_;
  assign new_n20258_ = ~new_n20256_ & ~new_n20257_;
  assign new_n20259_ = ~ys__n1489 & ~new_n20258_;
  assign new_n20260_ = ~new_n11893_ & ~new_n20178_;
  assign new_n20261_ = ~new_n17931_ & ~new_n20260_;
  assign new_n20262_ = new_n11896_ & ~new_n20261_;
  assign new_n20263_ = ~new_n11896_ & new_n20261_;
  assign new_n20264_ = ~new_n20262_ & ~new_n20263_;
  assign new_n20265_ = ys__n1489 & ~new_n20264_;
  assign new_n20266_ = ~new_n20259_ & ~new_n20265_;
  assign new_n20267_ = ~new_n19561_ & ~new_n20266_;
  assign new_n20268_ = ~new_n20253_ & ~new_n20267_;
  assign new_n20269_ = ~ys__n19973 & ~new_n20268_;
  assign new_n20270_ = ys__n19973 & ys__n19980;
  assign new_n20271_ = ~new_n20269_ & ~new_n20270_;
  assign new_n20272_ = ~ys__n352 & ~new_n20271_;
  assign new_n20273_ = ~ys__n220 & ys__n47033;
  assign new_n20274_ = new_n19573_ & new_n20273_;
  assign new_n20275_ = ~ys__n220 & ys__n47081;
  assign new_n20276_ = new_n19575_ & new_n20275_;
  assign new_n20277_ = ~ys__n220 & ys__n47017;
  assign new_n20278_ = new_n19578_ & new_n20277_;
  assign new_n20279_ = ~new_n20276_ & ~new_n20278_;
  assign new_n20280_ = ~new_n20274_ & new_n20279_;
  assign new_n20281_ = new_n19587_ & ~new_n20280_;
  assign ys__n19899 = new_n20272_ | new_n20281_;
  assign new_n20283_ = ys__n19844 & ys__n19852;
  assign new_n20284_ = new_n19250_ & new_n20283_;
  assign new_n20285_ = ~ys__n23276 & ~new_n19294_;
  assign new_n20286_ = ys__n23276 & ~new_n19318_;
  assign new_n20287_ = ~new_n20285_ & ~new_n20286_;
  assign new_n20288_ = ~ys__n23278 & ~new_n20287_;
  assign new_n20289_ = ~ys__n23276 & ~new_n19340_;
  assign new_n20290_ = ~new_n20216_ & ~new_n20289_;
  assign new_n20291_ = ys__n23278 & ~new_n20290_;
  assign new_n20292_ = ~new_n20288_ & ~new_n20291_;
  assign new_n20293_ = ~ys__n1505 & ~new_n20292_;
  assign new_n20294_ = ys__n23278 & new_n20289_;
  assign new_n20295_ = ~new_n20288_ & ~new_n20294_;
  assign new_n20296_ = ys__n1505 & ~new_n20295_;
  assign new_n20297_ = ~new_n20293_ & ~new_n20296_;
  assign new_n20298_ = ~new_n19250_ & ~new_n20297_;
  assign new_n20299_ = ~new_n20284_ & ~new_n20298_;
  assign new_n20300_ = new_n19347_ & ~new_n20299_;
  assign new_n20301_ = ~new_n19267_ & ~new_n19274_;
  assign new_n20302_ = ~ys__n23272 & ~new_n20301_;
  assign new_n20303_ = ys__n23272 & ~new_n20148_;
  assign new_n20304_ = ~new_n20302_ & ~new_n20303_;
  assign new_n20305_ = ~ys__n23274 & ~new_n20304_;
  assign new_n20306_ = ys__n23274 & ~new_n19985_;
  assign new_n20307_ = ~new_n20305_ & ~new_n20306_;
  assign new_n20308_ = ~ys__n23276 & ~new_n20307_;
  assign new_n20309_ = ys__n23276 & new_n19350_;
  assign new_n20310_ = ~new_n20308_ & ~new_n20309_;
  assign new_n20311_ = new_n19353_ & ~new_n20310_;
  assign new_n20312_ = ~new_n20300_ & ~new_n20311_;
  assign new_n20313_ = new_n19358_ & ~new_n20312_;
  assign new_n20314_ = ~new_n11932_ & new_n19360_;
  assign new_n20315_ = ys__n1498 & new_n19432_;
  assign new_n20316_ = ~new_n20314_ & ~new_n20315_;
  assign new_n20317_ = ~ys__n1496 & ~new_n20316_;
  assign new_n20318_ = ys__n1496 & ~new_n19432_;
  assign new_n20319_ = ~new_n20317_ & ~new_n20318_;
  assign new_n20320_ = ~ys__n1495 & ~new_n20319_;
  assign new_n20321_ = ys__n1495 & new_n17945_;
  assign new_n20322_ = ~new_n20320_ & ~new_n20321_;
  assign new_n20323_ = ~new_n19358_ & ~new_n20322_;
  assign new_n20324_ = ~new_n20313_ & ~new_n20323_;
  assign new_n20325_ = new_n19715_ & ~new_n20324_;
  assign new_n20326_ = ~new_n19413_ & new_n19433_;
  assign new_n20327_ = new_n19413_ & ~new_n19433_;
  assign new_n20328_ = ~new_n20326_ & ~new_n20327_;
  assign new_n20329_ = ~ys__n1489 & ~new_n20328_;
  assign new_n20330_ = new_n11932_ & ~new_n17935_;
  assign new_n20331_ = ~new_n11932_ & new_n17935_;
  assign new_n20332_ = ~new_n20330_ & ~new_n20331_;
  assign new_n20333_ = ys__n1489 & ~new_n20332_;
  assign new_n20334_ = ~new_n20329_ & ~new_n20333_;
  assign new_n20335_ = ~new_n19561_ & ~new_n20334_;
  assign new_n20336_ = ~new_n20325_ & ~new_n20335_;
  assign new_n20337_ = ~ys__n19973 & ~new_n20336_;
  assign new_n20338_ = ys__n19973 & ys__n19981;
  assign new_n20339_ = ~new_n20337_ & ~new_n20338_;
  assign new_n20340_ = ~ys__n352 & ~new_n20339_;
  assign new_n20341_ = ~ys__n220 & ys__n47034;
  assign new_n20342_ = new_n19573_ & new_n20341_;
  assign new_n20343_ = ~ys__n220 & ys__n47082;
  assign new_n20344_ = new_n19575_ & new_n20343_;
  assign new_n20345_ = ~ys__n220 & ys__n47018;
  assign new_n20346_ = new_n19578_ & new_n20345_;
  assign new_n20347_ = ~new_n20344_ & ~new_n20346_;
  assign new_n20348_ = ~new_n20342_ & new_n20347_;
  assign new_n20349_ = new_n19587_ & ~new_n20348_;
  assign ys__n19902 = new_n20340_ | new_n20349_;
  assign new_n20351_ = ys__n19844 & ys__n19853;
  assign new_n20352_ = new_n19250_ & new_n20351_;
  assign new_n20353_ = ~ys__n23276 & ~new_n19634_;
  assign new_n20354_ = ys__n23276 & ~new_n19658_;
  assign new_n20355_ = ~new_n20353_ & ~new_n20354_;
  assign new_n20356_ = ~ys__n23278 & ~new_n20355_;
  assign new_n20357_ = ~ys__n23276 & ~new_n19677_;
  assign new_n20358_ = ~new_n20216_ & ~new_n20357_;
  assign new_n20359_ = ys__n23278 & ~new_n20358_;
  assign new_n20360_ = ~new_n20356_ & ~new_n20359_;
  assign new_n20361_ = ~ys__n1505 & ~new_n20360_;
  assign new_n20362_ = ~ys__n23276 & ~new_n19687_;
  assign new_n20363_ = ys__n23278 & new_n20362_;
  assign new_n20364_ = ~new_n20356_ & ~new_n20363_;
  assign new_n20365_ = ys__n1505 & ~new_n20364_;
  assign new_n20366_ = ~new_n20361_ & ~new_n20365_;
  assign new_n20367_ = ~new_n19250_ & ~new_n20366_;
  assign new_n20368_ = ~new_n20352_ & ~new_n20367_;
  assign new_n20369_ = new_n19347_ & ~new_n20368_;
  assign new_n20370_ = ~new_n19607_ & ~new_n19614_;
  assign new_n20371_ = ~ys__n23272 & ~new_n20370_;
  assign new_n20372_ = ys__n23272 & ~new_n20231_;
  assign new_n20373_ = ~new_n20371_ & ~new_n20372_;
  assign new_n20374_ = ~ys__n23274 & ~new_n20373_;
  assign new_n20375_ = ys__n23274 & ~new_n20066_;
  assign new_n20376_ = ~new_n20374_ & ~new_n20375_;
  assign new_n20377_ = ~ys__n23276 & ~new_n20376_;
  assign new_n20378_ = ys__n23276 & new_n19699_;
  assign new_n20379_ = ~new_n20377_ & ~new_n20378_;
  assign new_n20380_ = new_n19353_ & ~new_n20379_;
  assign new_n20381_ = ~new_n20369_ & ~new_n20380_;
  assign new_n20382_ = new_n19358_ & ~new_n20381_;
  assign new_n20383_ = ~new_n11935_ & new_n19360_;
  assign new_n20384_ = ys__n1498 & new_n19430_;
  assign new_n20385_ = ~new_n20383_ & ~new_n20384_;
  assign new_n20386_ = ~ys__n1496 & ~new_n20385_;
  assign new_n20387_ = ys__n1496 & ~new_n19430_;
  assign new_n20388_ = ~new_n20386_ & ~new_n20387_;
  assign new_n20389_ = ~ys__n1495 & ~new_n20388_;
  assign new_n20390_ = ys__n1495 & new_n17944_;
  assign new_n20391_ = ~new_n20389_ & ~new_n20390_;
  assign new_n20392_ = ~new_n19358_ & ~new_n20391_;
  assign new_n20393_ = ~new_n20382_ & ~new_n20392_;
  assign new_n20394_ = new_n19715_ & ~new_n20393_;
  assign new_n20395_ = ~new_n19413_ & ~new_n19433_;
  assign new_n20396_ = ~new_n11931_ & ~new_n20395_;
  assign new_n20397_ = new_n19431_ & ~new_n20396_;
  assign new_n20398_ = ~new_n19431_ & new_n20396_;
  assign new_n20399_ = ~new_n20397_ & ~new_n20398_;
  assign new_n20400_ = ~ys__n1489 & ~new_n20399_;
  assign new_n20401_ = ~new_n11932_ & ~new_n17935_;
  assign new_n20402_ = ~new_n17945_ & ~new_n20401_;
  assign new_n20403_ = new_n11935_ & ~new_n20402_;
  assign new_n20404_ = ~new_n11935_ & new_n20402_;
  assign new_n20405_ = ~new_n20403_ & ~new_n20404_;
  assign new_n20406_ = ys__n1489 & ~new_n20405_;
  assign new_n20407_ = ~new_n20400_ & ~new_n20406_;
  assign new_n20408_ = ~new_n19561_ & ~new_n20407_;
  assign new_n20409_ = ~new_n20394_ & ~new_n20408_;
  assign new_n20410_ = ~ys__n19973 & ~new_n20409_;
  assign new_n20411_ = ys__n19973 & ys__n19982;
  assign new_n20412_ = ~new_n20410_ & ~new_n20411_;
  assign new_n20413_ = ~ys__n352 & ~new_n20412_;
  assign new_n20414_ = ~ys__n220 & ys__n47035;
  assign new_n20415_ = new_n19573_ & new_n20414_;
  assign new_n20416_ = ~ys__n220 & ys__n47083;
  assign new_n20417_ = new_n19575_ & new_n20416_;
  assign new_n20418_ = ~ys__n220 & ys__n47019;
  assign new_n20419_ = new_n19578_ & new_n20418_;
  assign new_n20420_ = ~new_n20417_ & ~new_n20419_;
  assign new_n20421_ = ~new_n20415_ & new_n20420_;
  assign new_n20422_ = new_n19587_ & ~new_n20421_;
  assign ys__n19905 = new_n20413_ | new_n20422_;
  assign new_n20424_ = ys__n19844 & ys__n19854;
  assign new_n20425_ = new_n19250_ & new_n20424_;
  assign new_n20426_ = ~ys__n23276 & ~new_n19759_;
  assign new_n20427_ = ys__n23276 & ~new_n19771_;
  assign new_n20428_ = ~new_n20426_ & ~new_n20427_;
  assign new_n20429_ = ~ys__n23278 & ~new_n20428_;
  assign new_n20430_ = ~ys__n23276 & ~new_n19780_;
  assign new_n20431_ = ~new_n20216_ & ~new_n20430_;
  assign new_n20432_ = ys__n23278 & ~new_n20431_;
  assign new_n20433_ = ~new_n20429_ & ~new_n20432_;
  assign new_n20434_ = ~ys__n1505 & ~new_n20433_;
  assign new_n20435_ = ~ys__n23276 & ~new_n19787_;
  assign new_n20436_ = ys__n23278 & new_n20435_;
  assign new_n20437_ = ~new_n20429_ & ~new_n20436_;
  assign new_n20438_ = ys__n1505 & ~new_n20437_;
  assign new_n20439_ = ~new_n20434_ & ~new_n20438_;
  assign new_n20440_ = ~new_n19250_ & ~new_n20439_;
  assign new_n20441_ = ~new_n20425_ & ~new_n20440_;
  assign new_n20442_ = new_n19347_ & ~new_n20441_;
  assign new_n20443_ = ~new_n19275_ & ~new_n19278_;
  assign new_n20444_ = ~ys__n23272 & ~new_n20443_;
  assign new_n20445_ = ys__n23272 & ~new_n20301_;
  assign new_n20446_ = ~new_n20444_ & ~new_n20445_;
  assign new_n20447_ = ~ys__n23274 & ~new_n20446_;
  assign new_n20448_ = ys__n23274 & ~new_n20151_;
  assign new_n20449_ = ~new_n20447_ & ~new_n20448_;
  assign new_n20450_ = ~ys__n23276 & ~new_n20449_;
  assign new_n20451_ = ys__n23276 & new_n19801_;
  assign new_n20452_ = ~new_n20450_ & ~new_n20451_;
  assign new_n20453_ = new_n19353_ & ~new_n20452_;
  assign new_n20454_ = ~new_n20442_ & ~new_n20453_;
  assign new_n20455_ = new_n19358_ & ~new_n20454_;
  assign new_n20456_ = ~new_n11939_ & new_n19360_;
  assign new_n20457_ = ys__n1498 & new_n19427_;
  assign new_n20458_ = ~new_n20456_ & ~new_n20457_;
  assign new_n20459_ = ~ys__n1496 & ~new_n20458_;
  assign new_n20460_ = ys__n1496 & ~new_n19427_;
  assign new_n20461_ = ~new_n20459_ & ~new_n20460_;
  assign new_n20462_ = ~ys__n1495 & ~new_n20461_;
  assign new_n20463_ = ys__n1495 & new_n17950_;
  assign new_n20464_ = ~new_n20462_ & ~new_n20463_;
  assign new_n20465_ = ~new_n19358_ & ~new_n20464_;
  assign new_n20466_ = ~new_n20455_ & ~new_n20465_;
  assign new_n20467_ = new_n19715_ & ~new_n20466_;
  assign new_n20468_ = ~new_n19413_ & new_n19434_;
  assign new_n20469_ = new_n19439_ & ~new_n20468_;
  assign new_n20470_ = new_n19428_ & ~new_n20469_;
  assign new_n20471_ = ~new_n19428_ & new_n20469_;
  assign new_n20472_ = ~new_n20470_ & ~new_n20471_;
  assign new_n20473_ = ~ys__n1489 & ~new_n20472_;
  assign new_n20474_ = ~new_n17935_ & new_n17940_;
  assign new_n20475_ = new_n17947_ & ~new_n20474_;
  assign new_n20476_ = new_n11939_ & ~new_n20475_;
  assign new_n20477_ = ~new_n11939_ & new_n20475_;
  assign new_n20478_ = ~new_n20476_ & ~new_n20477_;
  assign new_n20479_ = ys__n1489 & ~new_n20478_;
  assign new_n20480_ = ~new_n20473_ & ~new_n20479_;
  assign new_n20481_ = ~new_n19561_ & ~new_n20480_;
  assign new_n20482_ = ~new_n20467_ & ~new_n20481_;
  assign new_n20483_ = ~ys__n19973 & ~new_n20482_;
  assign new_n20484_ = ys__n19973 & ys__n19983;
  assign new_n20485_ = ~new_n20483_ & ~new_n20484_;
  assign new_n20486_ = ~ys__n352 & ~new_n20485_;
  assign new_n20487_ = ~ys__n220 & ys__n47036;
  assign new_n20488_ = new_n19573_ & new_n20487_;
  assign new_n20489_ = ~ys__n220 & ys__n47084;
  assign new_n20490_ = new_n19575_ & new_n20489_;
  assign new_n20491_ = ~ys__n220 & ys__n47020;
  assign new_n20492_ = new_n19578_ & new_n20491_;
  assign new_n20493_ = ~new_n20490_ & ~new_n20492_;
  assign new_n20494_ = ~new_n20488_ & new_n20493_;
  assign new_n20495_ = new_n19587_ & ~new_n20494_;
  assign ys__n19908 = new_n20486_ | new_n20495_;
  assign new_n20497_ = ys__n19844 & ys__n19855;
  assign new_n20498_ = new_n19250_ & new_n20497_;
  assign new_n20499_ = ~ys__n23276 & ~new_n19863_;
  assign new_n20500_ = ys__n23276 & ~new_n19875_;
  assign new_n20501_ = ~new_n20499_ & ~new_n20500_;
  assign new_n20502_ = ~ys__n23278 & ~new_n20501_;
  assign new_n20503_ = ~ys__n23276 & ~new_n19882_;
  assign new_n20504_ = ~new_n20216_ & ~new_n20503_;
  assign new_n20505_ = ys__n23278 & ~new_n20504_;
  assign new_n20506_ = ~new_n20502_ & ~new_n20505_;
  assign new_n20507_ = ~ys__n1505 & ~new_n20506_;
  assign new_n20508_ = ~ys__n23276 & ~new_n19890_;
  assign new_n20509_ = ys__n23278 & new_n20508_;
  assign new_n20510_ = ~new_n20502_ & ~new_n20509_;
  assign new_n20511_ = ys__n1505 & ~new_n20510_;
  assign new_n20512_ = ~new_n20507_ & ~new_n20511_;
  assign new_n20513_ = ~new_n19250_ & ~new_n20512_;
  assign new_n20514_ = ~new_n20498_ & ~new_n20513_;
  assign new_n20515_ = new_n19347_ & ~new_n20514_;
  assign new_n20516_ = ~new_n19615_ & ~new_n19618_;
  assign new_n20517_ = ~ys__n23272 & ~new_n20516_;
  assign new_n20518_ = ys__n23272 & ~new_n20370_;
  assign new_n20519_ = ~new_n20517_ & ~new_n20518_;
  assign new_n20520_ = ~ys__n23274 & ~new_n20519_;
  assign new_n20521_ = ys__n23274 & ~new_n20234_;
  assign new_n20522_ = ~new_n20520_ & ~new_n20521_;
  assign new_n20523_ = ~ys__n23276 & ~new_n20522_;
  assign new_n20524_ = ys__n23276 & new_n19904_;
  assign new_n20525_ = ~new_n20523_ & ~new_n20524_;
  assign new_n20526_ = new_n19353_ & ~new_n20525_;
  assign new_n20527_ = ~new_n20515_ & ~new_n20526_;
  assign new_n20528_ = new_n19358_ & ~new_n20527_;
  assign new_n20529_ = ~new_n11942_ & new_n19360_;
  assign new_n20530_ = ys__n1498 & new_n19425_;
  assign new_n20531_ = ~new_n20529_ & ~new_n20530_;
  assign new_n20532_ = ~ys__n1496 & ~new_n20531_;
  assign new_n20533_ = ys__n1496 & ~new_n19425_;
  assign new_n20534_ = ~new_n20532_ & ~new_n20533_;
  assign new_n20535_ = ~ys__n1495 & ~new_n20534_;
  assign new_n20536_ = ys__n1495 & new_n17949_;
  assign new_n20537_ = ~new_n20535_ & ~new_n20536_;
  assign new_n20538_ = ~new_n19358_ & ~new_n20537_;
  assign new_n20539_ = ~new_n20528_ & ~new_n20538_;
  assign new_n20540_ = new_n19715_ & ~new_n20539_;
  assign new_n20541_ = ~new_n19428_ & ~new_n20469_;
  assign new_n20542_ = ~new_n11938_ & ~new_n20541_;
  assign new_n20543_ = new_n19426_ & ~new_n20542_;
  assign new_n20544_ = ~new_n19426_ & new_n20542_;
  assign new_n20545_ = ~new_n20543_ & ~new_n20544_;
  assign new_n20546_ = ~ys__n1489 & ~new_n20545_;
  assign new_n20547_ = ~new_n11939_ & ~new_n20475_;
  assign new_n20548_ = ~new_n17950_ & ~new_n20547_;
  assign new_n20549_ = new_n11942_ & ~new_n20548_;
  assign new_n20550_ = ~new_n11942_ & new_n20548_;
  assign new_n20551_ = ~new_n20549_ & ~new_n20550_;
  assign new_n20552_ = ys__n1489 & ~new_n20551_;
  assign new_n20553_ = ~new_n20546_ & ~new_n20552_;
  assign new_n20554_ = ~new_n19561_ & ~new_n20553_;
  assign new_n20555_ = ~new_n20540_ & ~new_n20554_;
  assign new_n20556_ = ~ys__n19973 & ~new_n20555_;
  assign new_n20557_ = ys__n19973 & ys__n19984;
  assign new_n20558_ = ~new_n20556_ & ~new_n20557_;
  assign new_n20559_ = ~ys__n352 & ~new_n20558_;
  assign new_n20560_ = ~ys__n220 & ys__n47037;
  assign new_n20561_ = new_n19573_ & new_n20560_;
  assign new_n20562_ = ~ys__n220 & ys__n47085;
  assign new_n20563_ = new_n19575_ & new_n20562_;
  assign new_n20564_ = ~ys__n220 & ys__n47021;
  assign new_n20565_ = new_n19578_ & new_n20564_;
  assign new_n20566_ = ~new_n20563_ & ~new_n20565_;
  assign new_n20567_ = ~new_n20561_ & new_n20566_;
  assign new_n20568_ = new_n19587_ & ~new_n20567_;
  assign ys__n19911 = new_n20559_ | new_n20568_;
  assign new_n20570_ = ys__n19844 & ys__n19856;
  assign new_n20571_ = new_n19250_ & new_n20570_;
  assign new_n20572_ = ~ys__n23276 & ~new_n19958_;
  assign new_n20573_ = ys__n23276 & ~new_n19964_;
  assign new_n20574_ = ~new_n20572_ & ~new_n20573_;
  assign new_n20575_ = ~ys__n23278 & ~new_n20574_;
  assign new_n20576_ = ~ys__n23276 & ~new_n19967_;
  assign new_n20577_ = ~new_n20216_ & ~new_n20576_;
  assign new_n20578_ = ys__n23278 & ~new_n20577_;
  assign new_n20579_ = ~new_n20575_ & ~new_n20578_;
  assign new_n20580_ = ~ys__n1505 & ~new_n20579_;
  assign new_n20581_ = ~ys__n23276 & new_n19966_;
  assign new_n20582_ = ys__n23278 & new_n20581_;
  assign new_n20583_ = ~new_n20575_ & ~new_n20582_;
  assign new_n20584_ = ys__n1505 & ~new_n20583_;
  assign new_n20585_ = ~new_n20580_ & ~new_n20584_;
  assign new_n20586_ = ~new_n19250_ & ~new_n20585_;
  assign new_n20587_ = ~new_n20571_ & ~new_n20586_;
  assign new_n20588_ = new_n19347_ & ~new_n20587_;
  assign new_n20589_ = ~new_n19279_ & ~new_n19284_;
  assign new_n20590_ = ~ys__n23272 & ~new_n20589_;
  assign new_n20591_ = ys__n23272 & ~new_n20443_;
  assign new_n20592_ = ~new_n20590_ & ~new_n20591_;
  assign new_n20593_ = ~ys__n23274 & ~new_n20592_;
  assign new_n20594_ = ys__n23274 & ~new_n20304_;
  assign new_n20595_ = ~new_n20593_ & ~new_n20594_;
  assign new_n20596_ = ~ys__n23276 & ~new_n20595_;
  assign new_n20597_ = ys__n23276 & ~new_n19988_;
  assign new_n20598_ = ~new_n20596_ & ~new_n20597_;
  assign new_n20599_ = new_n19353_ & ~new_n20598_;
  assign new_n20600_ = ~new_n20588_ & ~new_n20599_;
  assign new_n20601_ = new_n19358_ & ~new_n20600_;
  assign new_n20602_ = ~new_n11917_ & new_n19360_;
  assign new_n20603_ = ys__n1498 & new_n19421_;
  assign new_n20604_ = ~new_n20602_ & ~new_n20603_;
  assign new_n20605_ = ~ys__n1496 & ~new_n20604_;
  assign new_n20606_ = ys__n1496 & ~new_n19421_;
  assign new_n20607_ = ~new_n20605_ & ~new_n20606_;
  assign new_n20608_ = ~ys__n1495 & ~new_n20607_;
  assign new_n20609_ = ys__n1495 & new_n17956_;
  assign new_n20610_ = ~new_n20608_ & ~new_n20609_;
  assign new_n20611_ = ~new_n19358_ & ~new_n20610_;
  assign new_n20612_ = ~new_n20601_ & ~new_n20611_;
  assign new_n20613_ = new_n19715_ & ~new_n20612_;
  assign new_n20614_ = ~new_n19413_ & new_n19435_;
  assign new_n20615_ = new_n19443_ & ~new_n20614_;
  assign new_n20616_ = new_n19422_ & ~new_n20615_;
  assign new_n20617_ = ~new_n19422_ & new_n20615_;
  assign new_n20618_ = ~new_n20616_ & ~new_n20617_;
  assign new_n20619_ = ~ys__n1489 & ~new_n20618_;
  assign new_n20620_ = ~new_n17935_ & new_n17941_;
  assign new_n20621_ = new_n17953_ & ~new_n20620_;
  assign new_n20622_ = new_n11917_ & ~new_n20621_;
  assign new_n20623_ = ~new_n11917_ & new_n20621_;
  assign new_n20624_ = ~new_n20622_ & ~new_n20623_;
  assign new_n20625_ = ys__n1489 & ~new_n20624_;
  assign new_n20626_ = ~new_n20619_ & ~new_n20625_;
  assign new_n20627_ = ~new_n19561_ & ~new_n20626_;
  assign new_n20628_ = ~new_n20613_ & ~new_n20627_;
  assign new_n20629_ = ~ys__n19973 & ~new_n20628_;
  assign new_n20630_ = ys__n19973 & ys__n19985;
  assign new_n20631_ = ~new_n20629_ & ~new_n20630_;
  assign new_n20632_ = ~ys__n352 & ~new_n20631_;
  assign new_n20633_ = ~ys__n220 & ys__n47038;
  assign new_n20634_ = new_n19573_ & new_n20633_;
  assign new_n20635_ = ~ys__n220 & ys__n47086;
  assign new_n20636_ = new_n19575_ & new_n20635_;
  assign new_n20637_ = ~ys__n220 & ys__n47022;
  assign new_n20638_ = new_n19578_ & new_n20637_;
  assign new_n20639_ = ~new_n20636_ & ~new_n20638_;
  assign new_n20640_ = ~new_n20634_ & new_n20639_;
  assign new_n20641_ = new_n19587_ & ~new_n20640_;
  assign ys__n19914 = new_n20632_ | new_n20641_;
  assign new_n20643_ = ys__n19844 & ys__n19857;
  assign new_n20644_ = new_n19250_ & new_n20643_;
  assign new_n20645_ = ~ys__n23276 & ~new_n20038_;
  assign new_n20646_ = ys__n23276 & ~new_n20044_;
  assign new_n20647_ = ~new_n20645_ & ~new_n20646_;
  assign new_n20648_ = ~ys__n23278 & ~new_n20647_;
  assign new_n20649_ = ~ys__n23276 & ~new_n20047_;
  assign new_n20650_ = ~new_n20216_ & ~new_n20649_;
  assign new_n20651_ = ys__n23278 & ~new_n20650_;
  assign new_n20652_ = ~new_n20648_ & ~new_n20651_;
  assign new_n20653_ = ~ys__n1505 & ~new_n20652_;
  assign new_n20654_ = ~ys__n23276 & new_n20053_;
  assign new_n20655_ = ys__n23278 & new_n20654_;
  assign new_n20656_ = ~new_n20648_ & ~new_n20655_;
  assign new_n20657_ = ys__n1505 & ~new_n20656_;
  assign new_n20658_ = ~new_n20653_ & ~new_n20657_;
  assign new_n20659_ = ~new_n19250_ & ~new_n20658_;
  assign new_n20660_ = ~new_n20644_ & ~new_n20659_;
  assign new_n20661_ = new_n19347_ & ~new_n20660_;
  assign new_n20662_ = ~new_n19619_ & ~new_n19624_;
  assign new_n20663_ = ~ys__n23272 & ~new_n20662_;
  assign new_n20664_ = ys__n23272 & ~new_n20516_;
  assign new_n20665_ = ~new_n20663_ & ~new_n20664_;
  assign new_n20666_ = ~ys__n23274 & ~new_n20665_;
  assign new_n20667_ = ys__n23274 & ~new_n20373_;
  assign new_n20668_ = ~new_n20666_ & ~new_n20667_;
  assign new_n20669_ = ~ys__n23276 & ~new_n20668_;
  assign new_n20670_ = ys__n23276 & ~new_n20069_;
  assign new_n20671_ = ~new_n20669_ & ~new_n20670_;
  assign new_n20672_ = new_n19353_ & ~new_n20671_;
  assign new_n20673_ = ~new_n20661_ & ~new_n20672_;
  assign new_n20674_ = new_n19358_ & ~new_n20673_;
  assign new_n20675_ = ~new_n11920_ & new_n19360_;
  assign new_n20676_ = ys__n1498 & new_n19419_;
  assign new_n20677_ = ~new_n20675_ & ~new_n20676_;
  assign new_n20678_ = ~ys__n1496 & ~new_n20677_;
  assign new_n20679_ = ys__n1496 & ~new_n19419_;
  assign new_n20680_ = ~new_n20678_ & ~new_n20679_;
  assign new_n20681_ = ~ys__n1495 & ~new_n20680_;
  assign new_n20682_ = ys__n1495 & new_n17955_;
  assign new_n20683_ = ~new_n20681_ & ~new_n20682_;
  assign new_n20684_ = ~new_n19358_ & ~new_n20683_;
  assign new_n20685_ = ~new_n20674_ & ~new_n20684_;
  assign new_n20686_ = new_n19715_ & ~new_n20685_;
  assign new_n20687_ = ~new_n19422_ & ~new_n20615_;
  assign new_n20688_ = ~new_n11916_ & ~new_n20687_;
  assign new_n20689_ = new_n19420_ & ~new_n20688_;
  assign new_n20690_ = ~new_n19420_ & new_n20688_;
  assign new_n20691_ = ~new_n20689_ & ~new_n20690_;
  assign new_n20692_ = ~ys__n1489 & ~new_n20691_;
  assign new_n20693_ = ~new_n11917_ & ~new_n20621_;
  assign new_n20694_ = ~new_n17956_ & ~new_n20693_;
  assign new_n20695_ = new_n11920_ & ~new_n20694_;
  assign new_n20696_ = ~new_n11920_ & new_n20694_;
  assign new_n20697_ = ~new_n20695_ & ~new_n20696_;
  assign new_n20698_ = ys__n1489 & ~new_n20697_;
  assign new_n20699_ = ~new_n20692_ & ~new_n20698_;
  assign new_n20700_ = ~new_n19561_ & ~new_n20699_;
  assign new_n20701_ = ~new_n20686_ & ~new_n20700_;
  assign new_n20702_ = ~ys__n19973 & ~new_n20701_;
  assign new_n20703_ = ys__n19973 & ys__n19986;
  assign new_n20704_ = ~new_n20702_ & ~new_n20703_;
  assign new_n20705_ = ~ys__n352 & ~new_n20704_;
  assign new_n20706_ = ~ys__n220 & ys__n47039;
  assign new_n20707_ = new_n19573_ & new_n20706_;
  assign new_n20708_ = ~ys__n220 & ys__n47087;
  assign new_n20709_ = new_n19575_ & new_n20708_;
  assign new_n20710_ = ~ys__n220 & ys__n47023;
  assign new_n20711_ = new_n19578_ & new_n20710_;
  assign new_n20712_ = ~new_n20709_ & ~new_n20711_;
  assign new_n20713_ = ~new_n20707_ & new_n20712_;
  assign new_n20714_ = new_n19587_ & ~new_n20713_;
  assign ys__n19917 = new_n20705_ | new_n20714_;
  assign new_n20716_ = ys__n19844 & ys__n19858;
  assign new_n20717_ = new_n19250_ & new_n20716_;
  assign new_n20718_ = ~ys__n23276 & ~new_n20123_;
  assign new_n20719_ = ys__n23276 & ~new_n20129_;
  assign new_n20720_ = ~new_n20718_ & ~new_n20719_;
  assign new_n20721_ = ~ys__n23278 & ~new_n20720_;
  assign new_n20722_ = ~ys__n23276 & ~new_n20132_;
  assign new_n20723_ = ~new_n20216_ & ~new_n20722_;
  assign new_n20724_ = ys__n23278 & ~new_n20723_;
  assign new_n20725_ = ~new_n20721_ & ~new_n20724_;
  assign new_n20726_ = ~ys__n1505 & ~new_n20725_;
  assign new_n20727_ = ~ys__n23276 & new_n20138_;
  assign new_n20728_ = ys__n23278 & new_n20727_;
  assign new_n20729_ = ~new_n20721_ & ~new_n20728_;
  assign new_n20730_ = ys__n1505 & ~new_n20729_;
  assign new_n20731_ = ~new_n20726_ & ~new_n20730_;
  assign new_n20732_ = ~new_n19250_ & ~new_n20731_;
  assign new_n20733_ = ~new_n20717_ & ~new_n20732_;
  assign new_n20734_ = new_n19347_ & ~new_n20733_;
  assign new_n20735_ = ~new_n19285_ & ~new_n19288_;
  assign new_n20736_ = ~ys__n23272 & ~new_n20735_;
  assign new_n20737_ = ys__n23272 & ~new_n20589_;
  assign new_n20738_ = ~new_n20736_ & ~new_n20737_;
  assign new_n20739_ = ~ys__n23274 & ~new_n20738_;
  assign new_n20740_ = ys__n23274 & ~new_n20446_;
  assign new_n20741_ = ~new_n20739_ & ~new_n20740_;
  assign new_n20742_ = ~ys__n23276 & ~new_n20741_;
  assign new_n20743_ = ys__n23276 & ~new_n20154_;
  assign new_n20744_ = ~new_n20742_ & ~new_n20743_;
  assign new_n20745_ = new_n19353_ & ~new_n20744_;
  assign new_n20746_ = ~new_n20734_ & ~new_n20745_;
  assign new_n20747_ = new_n19358_ & ~new_n20746_;
  assign new_n20748_ = ~new_n11924_ & new_n19360_;
  assign new_n20749_ = ys__n1498 & new_n19416_;
  assign new_n20750_ = ~new_n20748_ & ~new_n20749_;
  assign new_n20751_ = ~ys__n1496 & ~new_n20750_;
  assign new_n20752_ = ys__n1496 & ~new_n19416_;
  assign new_n20753_ = ~new_n20751_ & ~new_n20752_;
  assign new_n20754_ = ~ys__n1495 & ~new_n20753_;
  assign new_n20755_ = ys__n1495 & new_n17961_;
  assign new_n20756_ = ~new_n20754_ & ~new_n20755_;
  assign new_n20757_ = ~new_n19358_ & ~new_n20756_;
  assign new_n20758_ = ~new_n20747_ & ~new_n20757_;
  assign new_n20759_ = new_n19715_ & ~new_n20758_;
  assign new_n20760_ = new_n19423_ & ~new_n20615_;
  assign new_n20761_ = new_n19446_ & ~new_n20760_;
  assign new_n20762_ = new_n19417_ & ~new_n20761_;
  assign new_n20763_ = ~new_n19417_ & new_n20761_;
  assign new_n20764_ = ~new_n20762_ & ~new_n20763_;
  assign new_n20765_ = ~ys__n1489 & ~new_n20764_;
  assign new_n20766_ = new_n17937_ & ~new_n20621_;
  assign new_n20767_ = new_n17958_ & ~new_n20766_;
  assign new_n20768_ = new_n11924_ & ~new_n20767_;
  assign new_n20769_ = ~new_n11924_ & new_n20767_;
  assign new_n20770_ = ~new_n20768_ & ~new_n20769_;
  assign new_n20771_ = ys__n1489 & ~new_n20770_;
  assign new_n20772_ = ~new_n20765_ & ~new_n20771_;
  assign new_n20773_ = ~new_n19561_ & ~new_n20772_;
  assign new_n20774_ = ~new_n20759_ & ~new_n20773_;
  assign new_n20775_ = ~ys__n19973 & ~new_n20774_;
  assign new_n20776_ = ys__n19973 & ys__n19987;
  assign new_n20777_ = ~new_n20775_ & ~new_n20776_;
  assign new_n20778_ = ~ys__n352 & ~new_n20777_;
  assign new_n20779_ = ~ys__n220 & ys__n47040;
  assign new_n20780_ = new_n19573_ & new_n20779_;
  assign new_n20781_ = ~ys__n220 & ys__n47088;
  assign new_n20782_ = new_n19575_ & new_n20781_;
  assign new_n20783_ = ~ys__n220 & ys__n47024;
  assign new_n20784_ = new_n19578_ & new_n20783_;
  assign new_n20785_ = ~new_n20782_ & ~new_n20784_;
  assign new_n20786_ = ~new_n20780_ & new_n20785_;
  assign new_n20787_ = new_n19587_ & ~new_n20786_;
  assign ys__n19920 = new_n20778_ | new_n20787_;
  assign new_n20789_ = ys__n19844 & ys__n19859;
  assign new_n20790_ = new_n19250_ & new_n20789_;
  assign new_n20791_ = ~ys__n23276 & ~new_n20208_;
  assign new_n20792_ = ys__n23276 & ~new_n20214_;
  assign new_n20793_ = ~new_n20791_ & ~new_n20792_;
  assign new_n20794_ = ~ys__n23278 & ~new_n20793_;
  assign new_n20795_ = ys__n23278 & ys__n28030;
  assign new_n20796_ = ~new_n20794_ & ~new_n20795_;
  assign new_n20797_ = ~ys__n1505 & ~new_n20796_;
  assign new_n20798_ = ~ys__n23276 & new_n20221_;
  assign new_n20799_ = ys__n23278 & new_n20798_;
  assign new_n20800_ = ~new_n20794_ & ~new_n20799_;
  assign new_n20801_ = ys__n1505 & ~new_n20800_;
  assign new_n20802_ = ~new_n20797_ & ~new_n20801_;
  assign new_n20803_ = ~new_n19250_ & ~new_n20802_;
  assign new_n20804_ = ~new_n20790_ & ~new_n20803_;
  assign new_n20805_ = new_n19347_ & ~new_n20804_;
  assign new_n20806_ = ~new_n19625_ & ~new_n19628_;
  assign new_n20807_ = ~ys__n23272 & ~new_n20806_;
  assign new_n20808_ = ys__n23272 & ~new_n20662_;
  assign new_n20809_ = ~new_n20807_ & ~new_n20808_;
  assign new_n20810_ = ~ys__n23274 & ~new_n20809_;
  assign new_n20811_ = ys__n23274 & ~new_n20519_;
  assign new_n20812_ = ~new_n20810_ & ~new_n20811_;
  assign new_n20813_ = ~ys__n23276 & ~new_n20812_;
  assign new_n20814_ = ys__n23276 & ~new_n20237_;
  assign new_n20815_ = ~new_n20813_ & ~new_n20814_;
  assign new_n20816_ = new_n19353_ & ~new_n20815_;
  assign new_n20817_ = ~new_n20805_ & ~new_n20816_;
  assign new_n20818_ = new_n19358_ & ~new_n20817_;
  assign new_n20819_ = ~new_n11927_ & new_n19360_;
  assign new_n20820_ = ys__n1498 & new_n19414_;
  assign new_n20821_ = ~new_n20819_ & ~new_n20820_;
  assign new_n20822_ = ~ys__n1496 & ~new_n20821_;
  assign new_n20823_ = ys__n1496 & ~new_n19414_;
  assign new_n20824_ = ~new_n20822_ & ~new_n20823_;
  assign new_n20825_ = ~ys__n1495 & ~new_n20824_;
  assign new_n20826_ = ys__n1495 & new_n17960_;
  assign new_n20827_ = ~new_n20825_ & ~new_n20826_;
  assign new_n20828_ = ~new_n19358_ & ~new_n20827_;
  assign new_n20829_ = ~new_n20818_ & ~new_n20828_;
  assign new_n20830_ = new_n19715_ & ~new_n20829_;
  assign new_n20831_ = ~new_n19417_ & ~new_n20761_;
  assign new_n20832_ = ~new_n11923_ & ~new_n20831_;
  assign new_n20833_ = new_n19415_ & ~new_n20832_;
  assign new_n20834_ = ~new_n19415_ & new_n20832_;
  assign new_n20835_ = ~new_n20833_ & ~new_n20834_;
  assign new_n20836_ = ~ys__n1489 & ~new_n20835_;
  assign new_n20837_ = ~new_n11924_ & ~new_n20767_;
  assign new_n20838_ = ~new_n17961_ & ~new_n20837_;
  assign new_n20839_ = new_n11927_ & ~new_n20838_;
  assign new_n20840_ = ~new_n11927_ & new_n20838_;
  assign new_n20841_ = ~new_n20839_ & ~new_n20840_;
  assign new_n20842_ = ys__n1489 & ~new_n20841_;
  assign new_n20843_ = ~new_n20836_ & ~new_n20842_;
  assign new_n20844_ = ~new_n19561_ & ~new_n20843_;
  assign new_n20845_ = ~new_n20830_ & ~new_n20844_;
  assign new_n20846_ = ~ys__n19973 & ~new_n20845_;
  assign new_n20847_ = ys__n19973 & ys__n19988;
  assign new_n20848_ = ~new_n20846_ & ~new_n20847_;
  assign new_n20849_ = ~ys__n352 & ~new_n20848_;
  assign new_n20850_ = ~ys__n220 & ys__n47041;
  assign new_n20851_ = new_n19573_ & new_n20850_;
  assign new_n20852_ = ~ys__n220 & ys__n47089;
  assign new_n20853_ = new_n19575_ & new_n20852_;
  assign new_n20854_ = ~ys__n220 & ys__n47025;
  assign new_n20855_ = new_n19578_ & new_n20854_;
  assign new_n20856_ = ~new_n20853_ & ~new_n20855_;
  assign new_n20857_ = ~new_n20851_ & new_n20856_;
  assign new_n20858_ = new_n19587_ & ~new_n20857_;
  assign ys__n19923 = new_n20849_ | new_n20858_;
  assign new_n20860_ = ys__n19844 & ys__n19860;
  assign new_n20861_ = new_n19250_ & new_n20860_;
  assign new_n20862_ = ~ys__n23278 & ~new_n19342_;
  assign new_n20863_ = ~new_n20795_ & ~new_n20862_;
  assign new_n20864_ = ~ys__n1505 & ~new_n20863_;
  assign new_n20865_ = ys__n1505 & new_n20862_;
  assign new_n20866_ = ~new_n20864_ & ~new_n20865_;
  assign new_n20867_ = ~new_n19250_ & ~new_n20866_;
  assign new_n20868_ = ~new_n20861_ & ~new_n20867_;
  assign new_n20869_ = new_n19347_ & ~new_n20868_;
  assign new_n20870_ = ~ys__n1502 & ys__n27855;
  assign new_n20871_ = ~new_n19289_ & ~new_n19298_;
  assign new_n20872_ = ~ys__n23272 & ~new_n20871_;
  assign new_n20873_ = ys__n23272 & ~new_n20735_;
  assign new_n20874_ = ~new_n20872_ & ~new_n20873_;
  assign new_n20875_ = ~ys__n23274 & ~new_n20874_;
  assign new_n20876_ = ys__n23274 & ~new_n20592_;
  assign new_n20877_ = ~new_n20875_ & ~new_n20876_;
  assign new_n20878_ = ~ys__n23276 & ~new_n20877_;
  assign new_n20879_ = ys__n23276 & ~new_n20307_;
  assign new_n20880_ = ~new_n20878_ & ~new_n20879_;
  assign new_n20881_ = ~ys__n23278 & ~new_n20880_;
  assign new_n20882_ = ys__n23278 & new_n19351_;
  assign new_n20883_ = ~new_n20881_ & ~new_n20882_;
  assign new_n20884_ = ys__n1502 & ~new_n20883_;
  assign new_n20885_ = ~new_n20870_ & ~new_n20884_;
  assign new_n20886_ = ~new_n19347_ & ~new_n20885_;
  assign new_n20887_ = ~new_n20869_ & ~new_n20886_;
  assign new_n20888_ = new_n19358_ & ~new_n20887_;
  assign new_n20889_ = ~new_n11838_ & new_n19360_;
  assign new_n20890_ = ys__n1498 & new_n19495_;
  assign new_n20891_ = ~new_n20889_ & ~new_n20890_;
  assign new_n20892_ = ~ys__n1496 & ~new_n20891_;
  assign new_n20893_ = ys__n1496 & ~new_n19495_;
  assign new_n20894_ = ~new_n20892_ & ~new_n20893_;
  assign new_n20895_ = ~ys__n1495 & ~new_n20894_;
  assign new_n20896_ = ys__n1495 & new_n17887_;
  assign new_n20897_ = ~new_n20895_ & ~new_n20896_;
  assign new_n20898_ = ~new_n19358_ & ~new_n20897_;
  assign new_n20899_ = ~new_n20888_ & ~new_n20898_;
  assign new_n20900_ = new_n19715_ & ~new_n20899_;
  assign new_n20901_ = ~new_n19452_ & new_n19496_;
  assign new_n20902_ = new_n19452_ & ~new_n19496_;
  assign new_n20903_ = ~new_n20901_ & ~new_n20902_;
  assign new_n20904_ = ~ys__n1489 & ~new_n20903_;
  assign new_n20905_ = new_n11838_ & ~new_n17966_;
  assign new_n20906_ = ~new_n11838_ & new_n17966_;
  assign new_n20907_ = ~new_n20905_ & ~new_n20906_;
  assign new_n20908_ = ys__n1489 & ~new_n20907_;
  assign new_n20909_ = ~new_n20904_ & ~new_n20908_;
  assign new_n20910_ = ~new_n19561_ & ~new_n20909_;
  assign new_n20911_ = ~new_n20900_ & ~new_n20910_;
  assign new_n20912_ = ~ys__n19973 & ~new_n20911_;
  assign new_n20913_ = ys__n19973 & ys__n19989;
  assign new_n20914_ = ~new_n20912_ & ~new_n20913_;
  assign new_n20915_ = ~ys__n352 & ~new_n20914_;
  assign new_n20916_ = ~ys__n220 & ys__n47090;
  assign new_n20917_ = new_n19573_ & new_n20916_;
  assign new_n20918_ = new_n19575_ & new_n20916_;
  assign new_n20919_ = new_n19572_ & new_n19578_;
  assign new_n20920_ = ~new_n20918_ & ~new_n20919_;
  assign new_n20921_ = ~new_n20917_ & new_n20920_;
  assign new_n20922_ = new_n19587_ & ~new_n20921_;
  assign ys__n19926 = new_n20915_ | new_n20922_;
  assign new_n20924_ = ys__n19844 & ys__n19861;
  assign new_n20925_ = new_n19250_ & new_n20924_;
  assign new_n20926_ = ~ys__n23278 & ~new_n19679_;
  assign new_n20927_ = ~new_n20795_ & ~new_n20926_;
  assign new_n20928_ = ~ys__n1505 & ~new_n20927_;
  assign new_n20929_ = ys__n1505 & ~ys__n23278;
  assign new_n20930_ = ~new_n19689_ & new_n20929_;
  assign new_n20931_ = ~new_n20928_ & ~new_n20930_;
  assign new_n20932_ = ~new_n19250_ & ~new_n20931_;
  assign new_n20933_ = ~new_n20925_ & ~new_n20932_;
  assign new_n20934_ = new_n19347_ & ~new_n20933_;
  assign new_n20935_ = ~ys__n1502 & ys__n27857;
  assign new_n20936_ = ~new_n19629_ & ~new_n19638_;
  assign new_n20937_ = ~ys__n23272 & ~new_n20936_;
  assign new_n20938_ = ys__n23272 & ~new_n20806_;
  assign new_n20939_ = ~new_n20937_ & ~new_n20938_;
  assign new_n20940_ = ~ys__n23274 & ~new_n20939_;
  assign new_n20941_ = ys__n23274 & ~new_n20665_;
  assign new_n20942_ = ~new_n20940_ & ~new_n20941_;
  assign new_n20943_ = ~ys__n23276 & ~new_n20942_;
  assign new_n20944_ = ys__n23276 & ~new_n20376_;
  assign new_n20945_ = ~new_n20943_ & ~new_n20944_;
  assign new_n20946_ = ~ys__n23278 & ~new_n20945_;
  assign new_n20947_ = ys__n23278 & new_n19700_;
  assign new_n20948_ = ~new_n20946_ & ~new_n20947_;
  assign new_n20949_ = ys__n1502 & ~new_n20948_;
  assign new_n20950_ = ~new_n20935_ & ~new_n20949_;
  assign new_n20951_ = ~new_n19347_ & ~new_n20950_;
  assign new_n20952_ = ~new_n20934_ & ~new_n20951_;
  assign new_n20953_ = new_n19358_ & ~new_n20952_;
  assign new_n20954_ = ~new_n11841_ & new_n19360_;
  assign new_n20955_ = ys__n1498 & new_n19493_;
  assign new_n20956_ = ~new_n20954_ & ~new_n20955_;
  assign new_n20957_ = ~ys__n1496 & ~new_n20956_;
  assign new_n20958_ = ys__n1496 & ~new_n19493_;
  assign new_n20959_ = ~new_n20957_ & ~new_n20958_;
  assign new_n20960_ = ~ys__n1495 & ~new_n20959_;
  assign new_n20961_ = ys__n1495 & new_n17886_;
  assign new_n20962_ = ~new_n20960_ & ~new_n20961_;
  assign new_n20963_ = ~new_n19358_ & ~new_n20962_;
  assign new_n20964_ = ~new_n20953_ & ~new_n20963_;
  assign new_n20965_ = new_n19715_ & ~new_n20964_;
  assign new_n20966_ = ~new_n19452_ & ~new_n19496_;
  assign new_n20967_ = ~new_n11837_ & ~new_n20966_;
  assign new_n20968_ = new_n19494_ & ~new_n20967_;
  assign new_n20969_ = ~new_n19494_ & new_n20967_;
  assign new_n20970_ = ~new_n20968_ & ~new_n20969_;
  assign new_n20971_ = ~ys__n1489 & ~new_n20970_;
  assign new_n20972_ = ~new_n11838_ & ~new_n17966_;
  assign new_n20973_ = ~new_n17887_ & ~new_n20972_;
  assign new_n20974_ = new_n11841_ & ~new_n20973_;
  assign new_n20975_ = ~new_n11841_ & new_n20973_;
  assign new_n20976_ = ~new_n20974_ & ~new_n20975_;
  assign new_n20977_ = ys__n1489 & ~new_n20976_;
  assign new_n20978_ = ~new_n20971_ & ~new_n20977_;
  assign new_n20979_ = ~new_n19561_ & ~new_n20978_;
  assign new_n20980_ = ~new_n20965_ & ~new_n20979_;
  assign new_n20981_ = ~ys__n19973 & ~new_n20980_;
  assign new_n20982_ = ys__n19973 & ys__n19990;
  assign new_n20983_ = ~new_n20981_ & ~new_n20982_;
  assign new_n20984_ = ~ys__n352 & ~new_n20983_;
  assign new_n20985_ = ~ys__n220 & ys__n47091;
  assign new_n20986_ = new_n19573_ & new_n20985_;
  assign new_n20987_ = new_n19575_ & new_n20985_;
  assign new_n20988_ = new_n19578_ & new_n19729_;
  assign new_n20989_ = ~new_n20987_ & ~new_n20988_;
  assign new_n20990_ = ~new_n20986_ & new_n20989_;
  assign new_n20991_ = new_n19587_ & ~new_n20990_;
  assign ys__n19929 = new_n20984_ | new_n20991_;
  assign new_n20993_ = ys__n19844 & ys__n19862;
  assign new_n20994_ = new_n19250_ & new_n20993_;
  assign new_n20995_ = ~ys__n23278 & ~new_n19782_;
  assign new_n20996_ = ~new_n20795_ & ~new_n20995_;
  assign new_n20997_ = ~ys__n1505 & ~new_n20996_;
  assign new_n20998_ = ~new_n19789_ & new_n20929_;
  assign new_n20999_ = ~new_n20997_ & ~new_n20998_;
  assign new_n21000_ = ~new_n19250_ & ~new_n20999_;
  assign new_n21001_ = ~new_n20994_ & ~new_n21000_;
  assign new_n21002_ = new_n19347_ & ~new_n21001_;
  assign new_n21003_ = ~ys__n1502 & ys__n27859;
  assign new_n21004_ = ~new_n19299_ & ~new_n19302_;
  assign new_n21005_ = ~ys__n23272 & ~new_n21004_;
  assign new_n21006_ = ys__n23272 & ~new_n20871_;
  assign new_n21007_ = ~new_n21005_ & ~new_n21006_;
  assign new_n21008_ = ~ys__n23274 & ~new_n21007_;
  assign new_n21009_ = ys__n23274 & ~new_n20738_;
  assign new_n21010_ = ~new_n21008_ & ~new_n21009_;
  assign new_n21011_ = ~ys__n23276 & ~new_n21010_;
  assign new_n21012_ = ys__n23276 & ~new_n20449_;
  assign new_n21013_ = ~new_n21011_ & ~new_n21012_;
  assign new_n21014_ = ~ys__n23278 & ~new_n21013_;
  assign new_n21015_ = ys__n23278 & new_n19802_;
  assign new_n21016_ = ~new_n21014_ & ~new_n21015_;
  assign new_n21017_ = ys__n1502 & ~new_n21016_;
  assign new_n21018_ = ~new_n21003_ & ~new_n21017_;
  assign new_n21019_ = ~new_n19347_ & ~new_n21018_;
  assign new_n21020_ = ~new_n21002_ & ~new_n21019_;
  assign new_n21021_ = new_n19358_ & ~new_n21020_;
  assign new_n21022_ = ~new_n11845_ & new_n19360_;
  assign new_n21023_ = ys__n1498 & new_n19490_;
  assign new_n21024_ = ~new_n21022_ & ~new_n21023_;
  assign new_n21025_ = ~ys__n1496 & ~new_n21024_;
  assign new_n21026_ = ys__n1496 & ~new_n19490_;
  assign new_n21027_ = ~new_n21025_ & ~new_n21026_;
  assign new_n21028_ = ~ys__n1495 & ~new_n21027_;
  assign new_n21029_ = ys__n1495 & new_n17892_;
  assign new_n21030_ = ~new_n21028_ & ~new_n21029_;
  assign new_n21031_ = ~new_n19358_ & ~new_n21030_;
  assign new_n21032_ = ~new_n21021_ & ~new_n21031_;
  assign new_n21033_ = new_n19715_ & ~new_n21032_;
  assign new_n21034_ = ~new_n19452_ & new_n19497_;
  assign new_n21035_ = new_n19503_ & ~new_n21034_;
  assign new_n21036_ = new_n19491_ & ~new_n21035_;
  assign new_n21037_ = ~new_n19491_ & new_n21035_;
  assign new_n21038_ = ~new_n21036_ & ~new_n21037_;
  assign new_n21039_ = ~ys__n1489 & ~new_n21038_;
  assign new_n21040_ = new_n17908_ & ~new_n17966_;
  assign new_n21041_ = new_n17889_ & ~new_n21040_;
  assign new_n21042_ = new_n11845_ & ~new_n21041_;
  assign new_n21043_ = ~new_n11845_ & new_n21041_;
  assign new_n21044_ = ~new_n21042_ & ~new_n21043_;
  assign new_n21045_ = ys__n1489 & ~new_n21044_;
  assign new_n21046_ = ~new_n21039_ & ~new_n21045_;
  assign new_n21047_ = ~new_n19561_ & ~new_n21046_;
  assign new_n21048_ = ~new_n21033_ & ~new_n21047_;
  assign new_n21049_ = ~ys__n19973 & ~new_n21048_;
  assign new_n21050_ = ys__n19973 & ys__n19991;
  assign new_n21051_ = ~new_n21049_ & ~new_n21050_;
  assign new_n21052_ = ~ys__n352 & ~new_n21051_;
  assign new_n21053_ = ~ys__n220 & ys__n47092;
  assign new_n21054_ = new_n19573_ & new_n21053_;
  assign new_n21055_ = new_n19575_ & new_n21053_;
  assign new_n21056_ = new_n19578_ & new_n19833_;
  assign new_n21057_ = ~new_n21055_ & ~new_n21056_;
  assign new_n21058_ = ~new_n21054_ & new_n21057_;
  assign new_n21059_ = new_n19587_ & ~new_n21058_;
  assign ys__n19932 = new_n21052_ | new_n21059_;
  assign new_n21061_ = ys__n19844 & ys__n19863;
  assign new_n21062_ = new_n19250_ & new_n21061_;
  assign new_n21063_ = ~ys__n23278 & ~new_n19884_;
  assign new_n21064_ = ~new_n20795_ & ~new_n21063_;
  assign new_n21065_ = ~ys__n1505 & ~new_n21064_;
  assign new_n21066_ = ~new_n19892_ & new_n20929_;
  assign new_n21067_ = ~new_n21065_ & ~new_n21066_;
  assign new_n21068_ = ~new_n19250_ & ~new_n21067_;
  assign new_n21069_ = ~new_n21062_ & ~new_n21068_;
  assign new_n21070_ = new_n19347_ & ~new_n21069_;
  assign new_n21071_ = ~ys__n1502 & ys__n27861;
  assign new_n21072_ = ~new_n19639_ & ~new_n19642_;
  assign new_n21073_ = ~ys__n23272 & ~new_n21072_;
  assign new_n21074_ = ys__n23272 & ~new_n20936_;
  assign new_n21075_ = ~new_n21073_ & ~new_n21074_;
  assign new_n21076_ = ~ys__n23274 & ~new_n21075_;
  assign new_n21077_ = ys__n23274 & ~new_n20809_;
  assign new_n21078_ = ~new_n21076_ & ~new_n21077_;
  assign new_n21079_ = ~ys__n23276 & ~new_n21078_;
  assign new_n21080_ = ys__n23276 & ~new_n20522_;
  assign new_n21081_ = ~new_n21079_ & ~new_n21080_;
  assign new_n21082_ = ~ys__n23278 & ~new_n21081_;
  assign new_n21083_ = ys__n23278 & new_n19905_;
  assign new_n21084_ = ~new_n21082_ & ~new_n21083_;
  assign new_n21085_ = ys__n1502 & ~new_n21084_;
  assign new_n21086_ = ~new_n21071_ & ~new_n21085_;
  assign new_n21087_ = ~new_n19347_ & ~new_n21086_;
  assign new_n21088_ = ~new_n21070_ & ~new_n21087_;
  assign new_n21089_ = new_n19358_ & ~new_n21088_;
  assign new_n21090_ = ~new_n11848_ & new_n19360_;
  assign new_n21091_ = ys__n1498 & new_n19488_;
  assign new_n21092_ = ~new_n21090_ & ~new_n21091_;
  assign new_n21093_ = ~ys__n1496 & ~new_n21092_;
  assign new_n21094_ = ys__n1496 & ~new_n19488_;
  assign new_n21095_ = ~new_n21093_ & ~new_n21094_;
  assign new_n21096_ = ~ys__n1495 & ~new_n21095_;
  assign new_n21097_ = ys__n1495 & new_n17891_;
  assign new_n21098_ = ~new_n21096_ & ~new_n21097_;
  assign new_n21099_ = ~new_n19358_ & ~new_n21098_;
  assign new_n21100_ = ~new_n21089_ & ~new_n21099_;
  assign new_n21101_ = new_n19715_ & ~new_n21100_;
  assign new_n21102_ = ~new_n19491_ & ~new_n21035_;
  assign new_n21103_ = ~new_n11844_ & ~new_n21102_;
  assign new_n21104_ = new_n19489_ & ~new_n21103_;
  assign new_n21105_ = ~new_n19489_ & new_n21103_;
  assign new_n21106_ = ~new_n21104_ & ~new_n21105_;
  assign new_n21107_ = ~ys__n1489 & ~new_n21106_;
  assign new_n21108_ = ~new_n11845_ & ~new_n21041_;
  assign new_n21109_ = ~new_n17892_ & ~new_n21108_;
  assign new_n21110_ = new_n11848_ & ~new_n21109_;
  assign new_n21111_ = ~new_n11848_ & new_n21109_;
  assign new_n21112_ = ~new_n21110_ & ~new_n21111_;
  assign new_n21113_ = ys__n1489 & ~new_n21112_;
  assign new_n21114_ = ~new_n21107_ & ~new_n21113_;
  assign new_n21115_ = ~new_n19561_ & ~new_n21114_;
  assign new_n21116_ = ~new_n21101_ & ~new_n21115_;
  assign new_n21117_ = ~ys__n19973 & ~new_n21116_;
  assign new_n21118_ = ys__n19973 & ys__n19992;
  assign new_n21119_ = ~new_n21117_ & ~new_n21118_;
  assign new_n21120_ = ~ys__n352 & ~new_n21119_;
  assign new_n21121_ = ~ys__n220 & ys__n47093;
  assign new_n21122_ = new_n19573_ & new_n21121_;
  assign new_n21123_ = new_n19575_ & new_n21121_;
  assign new_n21124_ = new_n19578_ & new_n19940_;
  assign new_n21125_ = ~new_n21123_ & ~new_n21124_;
  assign new_n21126_ = ~new_n21122_ & new_n21125_;
  assign new_n21127_ = new_n19587_ & ~new_n21126_;
  assign ys__n19935 = new_n21120_ | new_n21127_;
  assign new_n21129_ = ys__n19844 & ys__n19864;
  assign new_n21130_ = new_n19250_ & new_n21129_;
  assign new_n21131_ = ~ys__n23278 & ~new_n19969_;
  assign new_n21132_ = ~new_n20795_ & ~new_n21131_;
  assign new_n21133_ = ~ys__n1505 & ~new_n21132_;
  assign new_n21134_ = ~new_n19974_ & new_n20929_;
  assign new_n21135_ = ~new_n21133_ & ~new_n21134_;
  assign new_n21136_ = ~new_n19250_ & ~new_n21135_;
  assign new_n21137_ = ~new_n21130_ & ~new_n21136_;
  assign new_n21138_ = new_n19347_ & ~new_n21137_;
  assign new_n21139_ = ~ys__n1502 & ys__n27863;
  assign new_n21140_ = ~new_n19303_ & ~new_n19308_;
  assign new_n21141_ = ~ys__n23272 & ~new_n21140_;
  assign new_n21142_ = ys__n23272 & ~new_n21004_;
  assign new_n21143_ = ~new_n21141_ & ~new_n21142_;
  assign new_n21144_ = ~ys__n23274 & ~new_n21143_;
  assign new_n21145_ = ys__n23274 & ~new_n20874_;
  assign new_n21146_ = ~new_n21144_ & ~new_n21145_;
  assign new_n21147_ = ~ys__n23276 & ~new_n21146_;
  assign new_n21148_ = ys__n23276 & ~new_n20595_;
  assign new_n21149_ = ~new_n21147_ & ~new_n21148_;
  assign new_n21150_ = ~ys__n23278 & ~new_n21149_;
  assign new_n21151_ = ys__n23278 & new_n19989_;
  assign new_n21152_ = ~new_n21150_ & ~new_n21151_;
  assign new_n21153_ = ys__n1502 & ~new_n21152_;
  assign new_n21154_ = ~new_n21139_ & ~new_n21153_;
  assign new_n21155_ = ~new_n19347_ & ~new_n21154_;
  assign new_n21156_ = ~new_n21138_ & ~new_n21155_;
  assign new_n21157_ = new_n19358_ & ~new_n21156_;
  assign new_n21158_ = ~new_n11823_ & new_n19360_;
  assign new_n21159_ = ys__n1498 & new_n19484_;
  assign new_n21160_ = ~new_n21158_ & ~new_n21159_;
  assign new_n21161_ = ~ys__n1496 & ~new_n21160_;
  assign new_n21162_ = ys__n1496 & ~new_n19484_;
  assign new_n21163_ = ~new_n21161_ & ~new_n21162_;
  assign new_n21164_ = ~ys__n1495 & ~new_n21163_;
  assign new_n21165_ = ys__n1495 & new_n17898_;
  assign new_n21166_ = ~new_n21164_ & ~new_n21165_;
  assign new_n21167_ = ~new_n19358_ & ~new_n21166_;
  assign new_n21168_ = ~new_n21157_ & ~new_n21167_;
  assign new_n21169_ = new_n19715_ & ~new_n21168_;
  assign new_n21170_ = ~new_n19452_ & new_n19498_;
  assign new_n21171_ = new_n19507_ & ~new_n21170_;
  assign new_n21172_ = new_n19485_ & ~new_n21171_;
  assign new_n21173_ = ~new_n19485_ & new_n21171_;
  assign new_n21174_ = ~new_n21172_ & ~new_n21173_;
  assign new_n21175_ = ~ys__n1489 & ~new_n21174_;
  assign new_n21176_ = new_n17909_ & ~new_n17966_;
  assign new_n21177_ = new_n17895_ & ~new_n21176_;
  assign new_n21178_ = new_n11823_ & ~new_n21177_;
  assign new_n21179_ = ~new_n11823_ & new_n21177_;
  assign new_n21180_ = ~new_n21178_ & ~new_n21179_;
  assign new_n21181_ = ys__n1489 & ~new_n21180_;
  assign new_n21182_ = ~new_n21175_ & ~new_n21181_;
  assign new_n21183_ = ~new_n19561_ & ~new_n21182_;
  assign new_n21184_ = ~new_n21169_ & ~new_n21183_;
  assign new_n21185_ = ~ys__n19973 & ~new_n21184_;
  assign new_n21186_ = ys__n19973 & ys__n19993;
  assign new_n21187_ = ~new_n21185_ & ~new_n21186_;
  assign new_n21188_ = ~ys__n352 & ~new_n21187_;
  assign new_n21189_ = ~ys__n220 & ys__n47094;
  assign new_n21190_ = new_n19573_ & new_n21189_;
  assign new_n21191_ = new_n19575_ & new_n21189_;
  assign new_n21192_ = new_n19578_ & new_n20020_;
  assign new_n21193_ = ~new_n21191_ & ~new_n21192_;
  assign new_n21194_ = ~new_n21190_ & new_n21193_;
  assign new_n21195_ = new_n19587_ & ~new_n21194_;
  assign ys__n19938 = new_n21188_ | new_n21195_;
  assign new_n21197_ = ys__n19844 & ys__n19865;
  assign new_n21198_ = new_n19250_ & new_n21197_;
  assign new_n21199_ = ~ys__n23278 & ~new_n20049_;
  assign new_n21200_ = ~new_n20795_ & ~new_n21199_;
  assign new_n21201_ = ~ys__n1505 & ~new_n21200_;
  assign new_n21202_ = ~new_n20055_ & new_n20929_;
  assign new_n21203_ = ~new_n21201_ & ~new_n21202_;
  assign new_n21204_ = ~new_n19250_ & ~new_n21203_;
  assign new_n21205_ = ~new_n21198_ & ~new_n21204_;
  assign new_n21206_ = new_n19347_ & ~new_n21205_;
  assign new_n21207_ = ~ys__n1502 & ys__n27865;
  assign new_n21208_ = ~new_n19643_ & ~new_n19648_;
  assign new_n21209_ = ~ys__n23272 & ~new_n21208_;
  assign new_n21210_ = ys__n23272 & ~new_n21072_;
  assign new_n21211_ = ~new_n21209_ & ~new_n21210_;
  assign new_n21212_ = ~ys__n23274 & ~new_n21211_;
  assign new_n21213_ = ys__n23274 & ~new_n20939_;
  assign new_n21214_ = ~new_n21212_ & ~new_n21213_;
  assign new_n21215_ = ~ys__n23276 & ~new_n21214_;
  assign new_n21216_ = ys__n23276 & ~new_n20668_;
  assign new_n21217_ = ~new_n21215_ & ~new_n21216_;
  assign new_n21218_ = ~ys__n23278 & ~new_n21217_;
  assign new_n21219_ = ys__n23278 & new_n20070_;
  assign new_n21220_ = ~new_n21218_ & ~new_n21219_;
  assign new_n21221_ = ys__n1502 & ~new_n21220_;
  assign new_n21222_ = ~new_n21207_ & ~new_n21221_;
  assign new_n21223_ = ~new_n19347_ & ~new_n21222_;
  assign new_n21224_ = ~new_n21206_ & ~new_n21223_;
  assign new_n21225_ = new_n19358_ & ~new_n21224_;
  assign new_n21226_ = ~new_n11826_ & new_n19360_;
  assign new_n21227_ = ys__n1498 & new_n19482_;
  assign new_n21228_ = ~new_n21226_ & ~new_n21227_;
  assign new_n21229_ = ~ys__n1496 & ~new_n21228_;
  assign new_n21230_ = ys__n1496 & ~new_n19482_;
  assign new_n21231_ = ~new_n21229_ & ~new_n21230_;
  assign new_n21232_ = ~ys__n1495 & ~new_n21231_;
  assign new_n21233_ = ys__n1495 & new_n17897_;
  assign new_n21234_ = ~new_n21232_ & ~new_n21233_;
  assign new_n21235_ = ~new_n19358_ & ~new_n21234_;
  assign new_n21236_ = ~new_n21225_ & ~new_n21235_;
  assign new_n21237_ = new_n19715_ & ~new_n21236_;
  assign new_n21238_ = ~new_n19485_ & ~new_n21171_;
  assign new_n21239_ = ~new_n11822_ & ~new_n21238_;
  assign new_n21240_ = new_n19483_ & ~new_n21239_;
  assign new_n21241_ = ~new_n19483_ & new_n21239_;
  assign new_n21242_ = ~new_n21240_ & ~new_n21241_;
  assign new_n21243_ = ~ys__n1489 & ~new_n21242_;
  assign new_n21244_ = ~new_n11823_ & ~new_n21177_;
  assign new_n21245_ = ~new_n17898_ & ~new_n21244_;
  assign new_n21246_ = new_n11826_ & ~new_n21245_;
  assign new_n21247_ = ~new_n11826_ & new_n21245_;
  assign new_n21248_ = ~new_n21246_ & ~new_n21247_;
  assign new_n21249_ = ys__n1489 & ~new_n21248_;
  assign new_n21250_ = ~new_n21243_ & ~new_n21249_;
  assign new_n21251_ = ~new_n19561_ & ~new_n21250_;
  assign new_n21252_ = ~new_n21237_ & ~new_n21251_;
  assign new_n21253_ = ~ys__n19973 & ~new_n21252_;
  assign new_n21254_ = ys__n19973 & ys__n19994;
  assign new_n21255_ = ~new_n21253_ & ~new_n21254_;
  assign new_n21256_ = ~ys__n352 & ~new_n21255_;
  assign new_n21257_ = ~ys__n220 & ys__n47095;
  assign new_n21258_ = new_n19573_ & new_n21257_;
  assign new_n21259_ = new_n19575_ & new_n21257_;
  assign new_n21260_ = new_n19578_ & new_n20105_;
  assign new_n21261_ = ~new_n21259_ & ~new_n21260_;
  assign new_n21262_ = ~new_n21258_ & new_n21261_;
  assign new_n21263_ = new_n19587_ & ~new_n21262_;
  assign ys__n19941 = new_n21256_ | new_n21263_;
  assign new_n21265_ = ys__n19844 & ys__n19866;
  assign new_n21266_ = new_n19250_ & new_n21265_;
  assign new_n21267_ = ~ys__n23278 & ~new_n20134_;
  assign new_n21268_ = ~new_n20795_ & ~new_n21267_;
  assign new_n21269_ = ~ys__n1505 & ~new_n21268_;
  assign new_n21270_ = ~new_n20140_ & new_n20929_;
  assign new_n21271_ = ~new_n21269_ & ~new_n21270_;
  assign new_n21272_ = ~new_n19250_ & ~new_n21271_;
  assign new_n21273_ = ~new_n21266_ & ~new_n21272_;
  assign new_n21274_ = new_n19347_ & ~new_n21273_;
  assign new_n21275_ = ~ys__n1502 & ys__n27867;
  assign new_n21276_ = ~new_n19309_ & ~new_n19312_;
  assign new_n21277_ = ~ys__n23272 & ~new_n21276_;
  assign new_n21278_ = ys__n23272 & ~new_n21140_;
  assign new_n21279_ = ~new_n21277_ & ~new_n21278_;
  assign new_n21280_ = ~ys__n23274 & ~new_n21279_;
  assign new_n21281_ = ys__n23274 & ~new_n21007_;
  assign new_n21282_ = ~new_n21280_ & ~new_n21281_;
  assign new_n21283_ = ~ys__n23276 & ~new_n21282_;
  assign new_n21284_ = ys__n23276 & ~new_n20741_;
  assign new_n21285_ = ~new_n21283_ & ~new_n21284_;
  assign new_n21286_ = ~ys__n23278 & ~new_n21285_;
  assign new_n21287_ = ys__n23278 & new_n20155_;
  assign new_n21288_ = ~new_n21286_ & ~new_n21287_;
  assign new_n21289_ = ys__n1502 & ~new_n21288_;
  assign new_n21290_ = ~new_n21275_ & ~new_n21289_;
  assign new_n21291_ = ~new_n19347_ & ~new_n21290_;
  assign new_n21292_ = ~new_n21274_ & ~new_n21291_;
  assign new_n21293_ = new_n19358_ & ~new_n21292_;
  assign new_n21294_ = ~new_n11830_ & new_n19360_;
  assign new_n21295_ = ys__n1498 & new_n19479_;
  assign new_n21296_ = ~new_n21294_ & ~new_n21295_;
  assign new_n21297_ = ~ys__n1496 & ~new_n21296_;
  assign new_n21298_ = ys__n1496 & ~new_n19479_;
  assign new_n21299_ = ~new_n21297_ & ~new_n21298_;
  assign new_n21300_ = ~ys__n1495 & ~new_n21299_;
  assign new_n21301_ = ys__n1495 & new_n17903_;
  assign new_n21302_ = ~new_n21300_ & ~new_n21301_;
  assign new_n21303_ = ~new_n19358_ & ~new_n21302_;
  assign new_n21304_ = ~new_n21293_ & ~new_n21303_;
  assign new_n21305_ = new_n19715_ & ~new_n21304_;
  assign new_n21306_ = new_n19486_ & ~new_n21171_;
  assign new_n21307_ = new_n19510_ & ~new_n21306_;
  assign new_n21308_ = new_n19480_ & ~new_n21307_;
  assign new_n21309_ = ~new_n19480_ & new_n21307_;
  assign new_n21310_ = ~new_n21308_ & ~new_n21309_;
  assign new_n21311_ = ~ys__n1489 & ~new_n21310_;
  assign new_n21312_ = new_n17883_ & ~new_n21177_;
  assign new_n21313_ = new_n17900_ & ~new_n21312_;
  assign new_n21314_ = new_n11830_ & ~new_n21313_;
  assign new_n21315_ = ~new_n11830_ & new_n21313_;
  assign new_n21316_ = ~new_n21314_ & ~new_n21315_;
  assign new_n21317_ = ys__n1489 & ~new_n21316_;
  assign new_n21318_ = ~new_n21311_ & ~new_n21317_;
  assign new_n21319_ = ~new_n19561_ & ~new_n21318_;
  assign new_n21320_ = ~new_n21305_ & ~new_n21319_;
  assign new_n21321_ = ~ys__n19973 & ~new_n21320_;
  assign new_n21322_ = ys__n19973 & ys__n19995;
  assign new_n21323_ = ~new_n21321_ & ~new_n21322_;
  assign new_n21324_ = ~ys__n352 & ~new_n21323_;
  assign new_n21325_ = ~ys__n220 & ys__n47096;
  assign new_n21326_ = new_n19573_ & new_n21325_;
  assign new_n21327_ = new_n19575_ & new_n21325_;
  assign new_n21328_ = new_n19578_ & new_n20190_;
  assign new_n21329_ = ~new_n21327_ & ~new_n21328_;
  assign new_n21330_ = ~new_n21326_ & new_n21329_;
  assign new_n21331_ = new_n19587_ & ~new_n21330_;
  assign ys__n19944 = new_n21324_ | new_n21331_;
  assign new_n21333_ = ys__n19844 & ys__n19867;
  assign new_n21334_ = new_n19250_ & new_n21333_;
  assign new_n21335_ = ~ys__n23278 & ~new_n20217_;
  assign new_n21336_ = ~new_n20795_ & ~new_n21335_;
  assign new_n21337_ = ~ys__n1505 & ~new_n21336_;
  assign new_n21338_ = ~new_n20223_ & new_n20929_;
  assign new_n21339_ = ~new_n21337_ & ~new_n21338_;
  assign new_n21340_ = ~new_n19250_ & ~new_n21339_;
  assign new_n21341_ = ~new_n21334_ & ~new_n21340_;
  assign new_n21342_ = new_n19347_ & ~new_n21341_;
  assign new_n21343_ = ~ys__n1502 & ys__n27869;
  assign new_n21344_ = ~new_n19649_ & ~new_n19652_;
  assign new_n21345_ = ~ys__n23272 & ~new_n21344_;
  assign new_n21346_ = ys__n23272 & ~new_n21208_;
  assign new_n21347_ = ~new_n21345_ & ~new_n21346_;
  assign new_n21348_ = ~ys__n23274 & ~new_n21347_;
  assign new_n21349_ = ys__n23274 & ~new_n21075_;
  assign new_n21350_ = ~new_n21348_ & ~new_n21349_;
  assign new_n21351_ = ~ys__n23276 & ~new_n21350_;
  assign new_n21352_ = ys__n23276 & ~new_n20812_;
  assign new_n21353_ = ~new_n21351_ & ~new_n21352_;
  assign new_n21354_ = ~ys__n23278 & ~new_n21353_;
  assign new_n21355_ = ys__n23278 & new_n20238_;
  assign new_n21356_ = ~new_n21354_ & ~new_n21355_;
  assign new_n21357_ = ys__n1502 & ~new_n21356_;
  assign new_n21358_ = ~new_n21343_ & ~new_n21357_;
  assign new_n21359_ = ~new_n19347_ & ~new_n21358_;
  assign new_n21360_ = ~new_n21342_ & ~new_n21359_;
  assign new_n21361_ = new_n19358_ & ~new_n21360_;
  assign new_n21362_ = ~new_n11833_ & new_n19360_;
  assign new_n21363_ = ys__n1498 & new_n19477_;
  assign new_n21364_ = ~new_n21362_ & ~new_n21363_;
  assign new_n21365_ = ~ys__n1496 & ~new_n21364_;
  assign new_n21366_ = ys__n1496 & ~new_n19477_;
  assign new_n21367_ = ~new_n21365_ & ~new_n21366_;
  assign new_n21368_ = ~ys__n1495 & ~new_n21367_;
  assign new_n21369_ = ys__n1495 & new_n17902_;
  assign new_n21370_ = ~new_n21368_ & ~new_n21369_;
  assign new_n21371_ = ~new_n19358_ & ~new_n21370_;
  assign new_n21372_ = ~new_n21361_ & ~new_n21371_;
  assign new_n21373_ = new_n19715_ & ~new_n21372_;
  assign new_n21374_ = ~new_n19480_ & ~new_n21307_;
  assign new_n21375_ = ~new_n11829_ & ~new_n21374_;
  assign new_n21376_ = new_n19478_ & ~new_n21375_;
  assign new_n21377_ = ~new_n19478_ & new_n21375_;
  assign new_n21378_ = ~new_n21376_ & ~new_n21377_;
  assign new_n21379_ = ~ys__n1489 & ~new_n21378_;
  assign new_n21380_ = ~new_n11830_ & ~new_n21313_;
  assign new_n21381_ = ~new_n17903_ & ~new_n21380_;
  assign new_n21382_ = new_n11833_ & ~new_n21381_;
  assign new_n21383_ = ~new_n11833_ & new_n21381_;
  assign new_n21384_ = ~new_n21382_ & ~new_n21383_;
  assign new_n21385_ = ys__n1489 & ~new_n21384_;
  assign new_n21386_ = ~new_n21379_ & ~new_n21385_;
  assign new_n21387_ = ~new_n19561_ & ~new_n21386_;
  assign new_n21388_ = ~new_n21373_ & ~new_n21387_;
  assign new_n21389_ = ~ys__n19973 & ~new_n21388_;
  assign new_n21390_ = ys__n19973 & ys__n19996;
  assign new_n21391_ = ~new_n21389_ & ~new_n21390_;
  assign new_n21392_ = ~ys__n352 & ~new_n21391_;
  assign new_n21393_ = ~ys__n220 & ys__n47097;
  assign new_n21394_ = new_n19573_ & new_n21393_;
  assign new_n21395_ = new_n19575_ & new_n21393_;
  assign new_n21396_ = new_n19578_ & new_n20273_;
  assign new_n21397_ = ~new_n21395_ & ~new_n21396_;
  assign new_n21398_ = ~new_n21394_ & new_n21397_;
  assign new_n21399_ = new_n19587_ & ~new_n21398_;
  assign ys__n19947 = new_n21392_ | new_n21399_;
  assign new_n21401_ = ys__n19844 & ys__n19868;
  assign new_n21402_ = new_n19250_ & new_n21401_;
  assign new_n21403_ = ~ys__n23278 & ~new_n20290_;
  assign new_n21404_ = ~new_n20795_ & ~new_n21403_;
  assign new_n21405_ = ~ys__n1505 & ~new_n21404_;
  assign new_n21406_ = new_n20289_ & new_n20929_;
  assign new_n21407_ = ~new_n21405_ & ~new_n21406_;
  assign new_n21408_ = ~new_n19250_ & ~new_n21407_;
  assign new_n21409_ = ~new_n21402_ & ~new_n21408_;
  assign new_n21410_ = new_n19347_ & ~new_n21409_;
  assign new_n21411_ = ~ys__n1502 & ys__n27871;
  assign new_n21412_ = ~new_n19313_ & ~new_n19320_;
  assign new_n21413_ = ~ys__n23272 & ~new_n21412_;
  assign new_n21414_ = ys__n23272 & ~new_n21276_;
  assign new_n21415_ = ~new_n21413_ & ~new_n21414_;
  assign new_n21416_ = ~ys__n23274 & ~new_n21415_;
  assign new_n21417_ = ys__n23274 & ~new_n21143_;
  assign new_n21418_ = ~new_n21416_ & ~new_n21417_;
  assign new_n21419_ = ~ys__n23276 & ~new_n21418_;
  assign new_n21420_ = ys__n23276 & ~new_n20877_;
  assign new_n21421_ = ~new_n21419_ & ~new_n21420_;
  assign new_n21422_ = ~ys__n23278 & ~new_n21421_;
  assign new_n21423_ = ys__n23278 & ~new_n20310_;
  assign new_n21424_ = ~new_n21422_ & ~new_n21423_;
  assign new_n21425_ = ys__n1502 & ~new_n21424_;
  assign new_n21426_ = ~new_n21411_ & ~new_n21425_;
  assign new_n21427_ = ~new_n19347_ & ~new_n21426_;
  assign new_n21428_ = ~new_n21410_ & ~new_n21427_;
  assign new_n21429_ = new_n19358_ & ~new_n21428_;
  assign new_n21430_ = ~new_n11869_ & new_n19360_;
  assign new_n21431_ = ys__n1498 & new_n19472_;
  assign new_n21432_ = ~new_n21430_ & ~new_n21431_;
  assign new_n21433_ = ~ys__n1496 & ~new_n21432_;
  assign new_n21434_ = ys__n1496 & ~new_n19472_;
  assign new_n21435_ = ~new_n21433_ & ~new_n21434_;
  assign new_n21436_ = ~ys__n1495 & ~new_n21435_;
  assign new_n21437_ = ys__n1495 & new_n17871_;
  assign new_n21438_ = ~new_n21436_ & ~new_n21437_;
  assign new_n21439_ = ~new_n19358_ & ~new_n21438_;
  assign new_n21440_ = ~new_n21429_ & ~new_n21439_;
  assign new_n21441_ = new_n19715_ & ~new_n21440_;
  assign new_n21442_ = ~new_n19452_ & new_n19499_;
  assign new_n21443_ = new_n19515_ & ~new_n21442_;
  assign new_n21444_ = new_n19473_ & ~new_n21443_;
  assign new_n21445_ = ~new_n19473_ & new_n21443_;
  assign new_n21446_ = ~new_n21444_ & ~new_n21445_;
  assign new_n21447_ = ~ys__n1489 & ~new_n21446_;
  assign new_n21448_ = new_n11869_ & ~new_n17968_;
  assign new_n21449_ = ~new_n11869_ & new_n17968_;
  assign new_n21450_ = ~new_n21448_ & ~new_n21449_;
  assign new_n21451_ = ys__n1489 & ~new_n21450_;
  assign new_n21452_ = ~new_n21447_ & ~new_n21451_;
  assign new_n21453_ = ~new_n19561_ & ~new_n21452_;
  assign new_n21454_ = ~new_n21441_ & ~new_n21453_;
  assign new_n21455_ = ~ys__n19973 & ~new_n21454_;
  assign new_n21456_ = ys__n19973 & ys__n19997;
  assign new_n21457_ = ~new_n21455_ & ~new_n21456_;
  assign new_n21458_ = ~ys__n352 & ~new_n21457_;
  assign new_n21459_ = ~ys__n220 & ys__n47098;
  assign new_n21460_ = new_n19573_ & new_n21459_;
  assign new_n21461_ = new_n19575_ & new_n21459_;
  assign new_n21462_ = new_n19578_ & new_n20341_;
  assign new_n21463_ = ~new_n21461_ & ~new_n21462_;
  assign new_n21464_ = ~new_n21460_ & new_n21463_;
  assign new_n21465_ = new_n19587_ & ~new_n21464_;
  assign ys__n19950 = new_n21458_ | new_n21465_;
  assign new_n21467_ = ys__n19844 & ys__n19869;
  assign new_n21468_ = new_n19250_ & new_n21467_;
  assign new_n21469_ = ~ys__n23278 & ~new_n20358_;
  assign new_n21470_ = ~new_n20795_ & ~new_n21469_;
  assign new_n21471_ = ~ys__n1505 & ~new_n21470_;
  assign new_n21472_ = new_n20362_ & new_n20929_;
  assign new_n21473_ = ~new_n21471_ & ~new_n21472_;
  assign new_n21474_ = ~new_n19250_ & ~new_n21473_;
  assign new_n21475_ = ~new_n21468_ & ~new_n21474_;
  assign new_n21476_ = new_n19347_ & ~new_n21475_;
  assign new_n21477_ = ~ys__n1502 & ys__n27873;
  assign new_n21478_ = ~new_n19653_ & ~new_n19660_;
  assign new_n21479_ = ~ys__n23272 & ~new_n21478_;
  assign new_n21480_ = ys__n23272 & ~new_n21344_;
  assign new_n21481_ = ~new_n21479_ & ~new_n21480_;
  assign new_n21482_ = ~ys__n23274 & ~new_n21481_;
  assign new_n21483_ = ys__n23274 & ~new_n21211_;
  assign new_n21484_ = ~new_n21482_ & ~new_n21483_;
  assign new_n21485_ = ~ys__n23276 & ~new_n21484_;
  assign new_n21486_ = ys__n23276 & ~new_n20942_;
  assign new_n21487_ = ~new_n21485_ & ~new_n21486_;
  assign new_n21488_ = ~ys__n23278 & ~new_n21487_;
  assign new_n21489_ = ys__n23278 & ~new_n20379_;
  assign new_n21490_ = ~new_n21488_ & ~new_n21489_;
  assign new_n21491_ = ys__n1502 & ~new_n21490_;
  assign new_n21492_ = ~new_n21477_ & ~new_n21491_;
  assign new_n21493_ = ~new_n19347_ & ~new_n21492_;
  assign new_n21494_ = ~new_n21476_ & ~new_n21493_;
  assign new_n21495_ = new_n19358_ & ~new_n21494_;
  assign new_n21496_ = ~new_n11872_ & new_n19360_;
  assign new_n21497_ = ys__n1498 & new_n19470_;
  assign new_n21498_ = ~new_n21496_ & ~new_n21497_;
  assign new_n21499_ = ~ys__n1496 & ~new_n21498_;
  assign new_n21500_ = ys__n1496 & ~new_n19470_;
  assign new_n21501_ = ~new_n21499_ & ~new_n21500_;
  assign new_n21502_ = ~ys__n1495 & ~new_n21501_;
  assign new_n21503_ = ys__n1495 & new_n17870_;
  assign new_n21504_ = ~new_n21502_ & ~new_n21503_;
  assign new_n21505_ = ~new_n19358_ & ~new_n21504_;
  assign new_n21506_ = ~new_n21495_ & ~new_n21505_;
  assign new_n21507_ = new_n19715_ & ~new_n21506_;
  assign new_n21508_ = ~new_n19473_ & ~new_n21443_;
  assign new_n21509_ = ~new_n11868_ & ~new_n21508_;
  assign new_n21510_ = new_n19471_ & ~new_n21509_;
  assign new_n21511_ = ~new_n19471_ & new_n21509_;
  assign new_n21512_ = ~new_n21510_ & ~new_n21511_;
  assign new_n21513_ = ~ys__n1489 & ~new_n21512_;
  assign new_n21514_ = ~new_n11869_ & ~new_n17968_;
  assign new_n21515_ = ~new_n17871_ & ~new_n21514_;
  assign new_n21516_ = new_n11872_ & ~new_n21515_;
  assign new_n21517_ = ~new_n11872_ & new_n21515_;
  assign new_n21518_ = ~new_n21516_ & ~new_n21517_;
  assign new_n21519_ = ys__n1489 & ~new_n21518_;
  assign new_n21520_ = ~new_n21513_ & ~new_n21519_;
  assign new_n21521_ = ~new_n19561_ & ~new_n21520_;
  assign new_n21522_ = ~new_n21507_ & ~new_n21521_;
  assign new_n21523_ = ~ys__n19973 & ~new_n21522_;
  assign new_n21524_ = ys__n19973 & ys__n19998;
  assign new_n21525_ = ~new_n21523_ & ~new_n21524_;
  assign new_n21526_ = ~ys__n352 & ~new_n21525_;
  assign new_n21527_ = ~ys__n220 & ys__n47099;
  assign new_n21528_ = new_n19573_ & new_n21527_;
  assign new_n21529_ = new_n19575_ & new_n21527_;
  assign new_n21530_ = new_n19578_ & new_n20414_;
  assign new_n21531_ = ~new_n21529_ & ~new_n21530_;
  assign new_n21532_ = ~new_n21528_ & new_n21531_;
  assign new_n21533_ = new_n19587_ & ~new_n21532_;
  assign ys__n19953 = new_n21526_ | new_n21533_;
  assign new_n21535_ = ys__n19844 & ys__n19870;
  assign new_n21536_ = new_n19250_ & new_n21535_;
  assign new_n21537_ = ~ys__n23278 & ~new_n20431_;
  assign new_n21538_ = ~new_n20795_ & ~new_n21537_;
  assign new_n21539_ = ~ys__n1505 & ~new_n21538_;
  assign new_n21540_ = new_n20435_ & new_n20929_;
  assign new_n21541_ = ~new_n21539_ & ~new_n21540_;
  assign new_n21542_ = ~new_n19250_ & ~new_n21541_;
  assign new_n21543_ = ~new_n21536_ & ~new_n21542_;
  assign new_n21544_ = new_n19347_ & ~new_n21543_;
  assign new_n21545_ = ~ys__n1502 & ys__n27875;
  assign new_n21546_ = ~new_n19321_ & ~new_n19324_;
  assign new_n21547_ = ~ys__n23272 & ~new_n21546_;
  assign new_n21548_ = ys__n23272 & ~new_n21412_;
  assign new_n21549_ = ~new_n21547_ & ~new_n21548_;
  assign new_n21550_ = ~ys__n23274 & ~new_n21549_;
  assign new_n21551_ = ys__n23274 & ~new_n21279_;
  assign new_n21552_ = ~new_n21550_ & ~new_n21551_;
  assign new_n21553_ = ~ys__n23276 & ~new_n21552_;
  assign new_n21554_ = ys__n23276 & ~new_n21010_;
  assign new_n21555_ = ~new_n21553_ & ~new_n21554_;
  assign new_n21556_ = ~ys__n23278 & ~new_n21555_;
  assign new_n21557_ = ys__n23278 & ~new_n20452_;
  assign new_n21558_ = ~new_n21556_ & ~new_n21557_;
  assign new_n21559_ = ys__n1502 & ~new_n21558_;
  assign new_n21560_ = ~new_n21545_ & ~new_n21559_;
  assign new_n21561_ = ~new_n19347_ & ~new_n21560_;
  assign new_n21562_ = ~new_n21544_ & ~new_n21561_;
  assign new_n21563_ = new_n19358_ & ~new_n21562_;
  assign new_n21564_ = ~new_n11876_ & new_n19360_;
  assign new_n21565_ = ys__n1498 & new_n19467_;
  assign new_n21566_ = ~new_n21564_ & ~new_n21565_;
  assign new_n21567_ = ~ys__n1496 & ~new_n21566_;
  assign new_n21568_ = ys__n1496 & ~new_n19467_;
  assign new_n21569_ = ~new_n21567_ & ~new_n21568_;
  assign new_n21570_ = ~ys__n1495 & ~new_n21569_;
  assign new_n21571_ = ys__n1495 & new_n17876_;
  assign new_n21572_ = ~new_n21570_ & ~new_n21571_;
  assign new_n21573_ = ~new_n19358_ & ~new_n21572_;
  assign new_n21574_ = ~new_n21563_ & ~new_n21573_;
  assign new_n21575_ = new_n19715_ & ~new_n21574_;
  assign new_n21576_ = new_n19474_ & ~new_n21443_;
  assign new_n21577_ = new_n19518_ & ~new_n21576_;
  assign new_n21578_ = new_n19468_ & ~new_n21577_;
  assign new_n21579_ = ~new_n19468_ & new_n21577_;
  assign new_n21580_ = ~new_n21578_ & ~new_n21579_;
  assign new_n21581_ = ~ys__n1489 & ~new_n21580_;
  assign new_n21582_ = new_n17880_ & ~new_n17968_;
  assign new_n21583_ = new_n17873_ & ~new_n21582_;
  assign new_n21584_ = new_n11876_ & ~new_n21583_;
  assign new_n21585_ = ~new_n11876_ & new_n21583_;
  assign new_n21586_ = ~new_n21584_ & ~new_n21585_;
  assign new_n21587_ = ys__n1489 & ~new_n21586_;
  assign new_n21588_ = ~new_n21581_ & ~new_n21587_;
  assign new_n21589_ = ~new_n19561_ & ~new_n21588_;
  assign new_n21590_ = ~new_n21575_ & ~new_n21589_;
  assign new_n21591_ = ~ys__n19973 & ~new_n21590_;
  assign new_n21592_ = ys__n19973 & ys__n19999;
  assign new_n21593_ = ~new_n21591_ & ~new_n21592_;
  assign new_n21594_ = ~ys__n352 & ~new_n21593_;
  assign new_n21595_ = ~ys__n220 & ys__n47100;
  assign new_n21596_ = new_n19573_ & new_n21595_;
  assign new_n21597_ = new_n19575_ & new_n21595_;
  assign new_n21598_ = new_n19578_ & new_n20487_;
  assign new_n21599_ = ~new_n21597_ & ~new_n21598_;
  assign new_n21600_ = ~new_n21596_ & new_n21599_;
  assign new_n21601_ = new_n19587_ & ~new_n21600_;
  assign ys__n19956 = new_n21594_ | new_n21601_;
  assign new_n21603_ = ys__n19844 & ys__n19871;
  assign new_n21604_ = new_n19250_ & new_n21603_;
  assign new_n21605_ = ~ys__n23278 & ~new_n20504_;
  assign new_n21606_ = ~new_n20795_ & ~new_n21605_;
  assign new_n21607_ = ~ys__n1505 & ~new_n21606_;
  assign new_n21608_ = new_n20508_ & new_n20929_;
  assign new_n21609_ = ~new_n21607_ & ~new_n21608_;
  assign new_n21610_ = ~new_n19250_ & ~new_n21609_;
  assign new_n21611_ = ~new_n21604_ & ~new_n21610_;
  assign new_n21612_ = new_n19347_ & ~new_n21611_;
  assign new_n21613_ = ~ys__n1502 & ys__n27877;
  assign new_n21614_ = ~new_n19661_ & ~new_n19664_;
  assign new_n21615_ = ~ys__n23272 & ~new_n21614_;
  assign new_n21616_ = ys__n23272 & ~new_n21478_;
  assign new_n21617_ = ~new_n21615_ & ~new_n21616_;
  assign new_n21618_ = ~ys__n23274 & ~new_n21617_;
  assign new_n21619_ = ys__n23274 & ~new_n21347_;
  assign new_n21620_ = ~new_n21618_ & ~new_n21619_;
  assign new_n21621_ = ~ys__n23276 & ~new_n21620_;
  assign new_n21622_ = ys__n23276 & ~new_n21078_;
  assign new_n21623_ = ~new_n21621_ & ~new_n21622_;
  assign new_n21624_ = ~ys__n23278 & ~new_n21623_;
  assign new_n21625_ = ys__n23278 & ~new_n20525_;
  assign new_n21626_ = ~new_n21624_ & ~new_n21625_;
  assign new_n21627_ = ys__n1502 & ~new_n21626_;
  assign new_n21628_ = ~new_n21613_ & ~new_n21627_;
  assign new_n21629_ = ~new_n19347_ & ~new_n21628_;
  assign new_n21630_ = ~new_n21612_ & ~new_n21629_;
  assign new_n21631_ = new_n19358_ & ~new_n21630_;
  assign new_n21632_ = ~new_n11879_ & new_n19360_;
  assign new_n21633_ = ys__n1498 & new_n19465_;
  assign new_n21634_ = ~new_n21632_ & ~new_n21633_;
  assign new_n21635_ = ~ys__n1496 & ~new_n21634_;
  assign new_n21636_ = ys__n1496 & ~new_n19465_;
  assign new_n21637_ = ~new_n21635_ & ~new_n21636_;
  assign new_n21638_ = ~ys__n1495 & ~new_n21637_;
  assign new_n21639_ = ys__n1495 & new_n17875_;
  assign new_n21640_ = ~new_n21638_ & ~new_n21639_;
  assign new_n21641_ = ~new_n19358_ & ~new_n21640_;
  assign new_n21642_ = ~new_n21631_ & ~new_n21641_;
  assign new_n21643_ = new_n19715_ & ~new_n21642_;
  assign new_n21644_ = ~new_n19468_ & ~new_n21577_;
  assign new_n21645_ = ~new_n11875_ & ~new_n21644_;
  assign new_n21646_ = new_n19466_ & ~new_n21645_;
  assign new_n21647_ = ~new_n19466_ & new_n21645_;
  assign new_n21648_ = ~new_n21646_ & ~new_n21647_;
  assign new_n21649_ = ~ys__n1489 & ~new_n21648_;
  assign new_n21650_ = ~new_n11876_ & ~new_n21583_;
  assign new_n21651_ = ~new_n17876_ & ~new_n21650_;
  assign new_n21652_ = new_n11879_ & ~new_n21651_;
  assign new_n21653_ = ~new_n11879_ & new_n21651_;
  assign new_n21654_ = ~new_n21652_ & ~new_n21653_;
  assign new_n21655_ = ys__n1489 & ~new_n21654_;
  assign new_n21656_ = ~new_n21649_ & ~new_n21655_;
  assign new_n21657_ = ~new_n19561_ & ~new_n21656_;
  assign new_n21658_ = ~new_n21643_ & ~new_n21657_;
  assign new_n21659_ = ~ys__n19973 & ~new_n21658_;
  assign new_n21660_ = ys__n19973 & ys__n20000;
  assign new_n21661_ = ~new_n21659_ & ~new_n21660_;
  assign new_n21662_ = ~ys__n352 & ~new_n21661_;
  assign new_n21663_ = ~ys__n220 & ys__n47101;
  assign new_n21664_ = new_n19573_ & new_n21663_;
  assign new_n21665_ = new_n19575_ & new_n21663_;
  assign new_n21666_ = new_n19578_ & new_n20560_;
  assign new_n21667_ = ~new_n21665_ & ~new_n21666_;
  assign new_n21668_ = ~new_n21664_ & new_n21667_;
  assign new_n21669_ = new_n19587_ & ~new_n21668_;
  assign ys__n19959 = new_n21662_ | new_n21669_;
  assign new_n21671_ = ys__n19844 & ys__n19872;
  assign new_n21672_ = new_n19250_ & new_n21671_;
  assign new_n21673_ = ~ys__n23278 & ~new_n20577_;
  assign new_n21674_ = ~new_n20795_ & ~new_n21673_;
  assign new_n21675_ = ~ys__n1505 & ~new_n21674_;
  assign new_n21676_ = new_n20581_ & new_n20929_;
  assign new_n21677_ = ~new_n21675_ & ~new_n21676_;
  assign new_n21678_ = ~new_n19250_ & ~new_n21677_;
  assign new_n21679_ = ~new_n21672_ & ~new_n21678_;
  assign new_n21680_ = new_n19347_ & ~new_n21679_;
  assign new_n21681_ = ~ys__n1502 & ys__n27879;
  assign new_n21682_ = ~new_n19325_ & ~new_n19330_;
  assign new_n21683_ = ~ys__n23272 & ~new_n21682_;
  assign new_n21684_ = ys__n23272 & ~new_n21546_;
  assign new_n21685_ = ~new_n21683_ & ~new_n21684_;
  assign new_n21686_ = ~ys__n23274 & ~new_n21685_;
  assign new_n21687_ = ys__n23274 & ~new_n21415_;
  assign new_n21688_ = ~new_n21686_ & ~new_n21687_;
  assign new_n21689_ = ~ys__n23276 & ~new_n21688_;
  assign new_n21690_ = ys__n23276 & ~new_n21146_;
  assign new_n21691_ = ~new_n21689_ & ~new_n21690_;
  assign new_n21692_ = ~ys__n23278 & ~new_n21691_;
  assign new_n21693_ = ys__n23278 & ~new_n20598_;
  assign new_n21694_ = ~new_n21692_ & ~new_n21693_;
  assign new_n21695_ = ys__n1502 & ~new_n21694_;
  assign new_n21696_ = ~new_n21681_ & ~new_n21695_;
  assign new_n21697_ = ~new_n19347_ & ~new_n21696_;
  assign new_n21698_ = ~new_n21680_ & ~new_n21697_;
  assign new_n21699_ = new_n19358_ & ~new_n21698_;
  assign new_n21700_ = ~new_n11854_ & new_n19360_;
  assign new_n21701_ = ys__n1498 & new_n19461_;
  assign new_n21702_ = ~new_n21700_ & ~new_n21701_;
  assign new_n21703_ = ~ys__n1496 & ~new_n21702_;
  assign new_n21704_ = ys__n1496 & ~new_n19461_;
  assign new_n21705_ = ~new_n21703_ & ~new_n21704_;
  assign new_n21706_ = ~ys__n1495 & ~new_n21705_;
  assign new_n21707_ = ys__n1495 & new_n17868_;
  assign new_n21708_ = ~new_n21706_ & ~new_n21707_;
  assign new_n21709_ = ~new_n19358_ & ~new_n21708_;
  assign new_n21710_ = ~new_n21699_ & ~new_n21709_;
  assign new_n21711_ = new_n19715_ & ~new_n21710_;
  assign new_n21712_ = new_n19475_ & ~new_n21443_;
  assign new_n21713_ = new_n19522_ & ~new_n21712_;
  assign new_n21714_ = new_n19462_ & ~new_n21713_;
  assign new_n21715_ = ~new_n19462_ & new_n21713_;
  assign new_n21716_ = ~new_n21714_ & ~new_n21715_;
  assign new_n21717_ = ~ys__n1489 & ~new_n21716_;
  assign new_n21718_ = new_n11854_ & ~new_n17970_;
  assign new_n21719_ = ~new_n11854_ & new_n17970_;
  assign new_n21720_ = ~new_n21718_ & ~new_n21719_;
  assign new_n21721_ = ys__n1489 & ~new_n21720_;
  assign new_n21722_ = ~new_n21717_ & ~new_n21721_;
  assign new_n21723_ = ~new_n19561_ & ~new_n21722_;
  assign new_n21724_ = ~new_n21711_ & ~new_n21723_;
  assign new_n21725_ = ~ys__n19973 & ~new_n21724_;
  assign new_n21726_ = ys__n19973 & ys__n20001;
  assign new_n21727_ = ~new_n21725_ & ~new_n21726_;
  assign new_n21728_ = ~ys__n352 & ~new_n21727_;
  assign new_n21729_ = ~ys__n220 & ys__n47102;
  assign new_n21730_ = new_n19573_ & new_n21729_;
  assign new_n21731_ = new_n19575_ & new_n21729_;
  assign new_n21732_ = new_n19578_ & new_n20633_;
  assign new_n21733_ = ~new_n21731_ & ~new_n21732_;
  assign new_n21734_ = ~new_n21730_ & new_n21733_;
  assign new_n21735_ = new_n19587_ & ~new_n21734_;
  assign ys__n19962 = new_n21728_ | new_n21735_;
  assign new_n21737_ = ys__n19844 & ys__n19873;
  assign new_n21738_ = new_n19250_ & new_n21737_;
  assign new_n21739_ = ~ys__n23278 & ~new_n20650_;
  assign new_n21740_ = ~new_n20795_ & ~new_n21739_;
  assign new_n21741_ = ~ys__n1505 & ~new_n21740_;
  assign new_n21742_ = new_n20654_ & new_n20929_;
  assign new_n21743_ = ~new_n21741_ & ~new_n21742_;
  assign new_n21744_ = ~new_n19250_ & ~new_n21743_;
  assign new_n21745_ = ~new_n21738_ & ~new_n21744_;
  assign new_n21746_ = new_n19347_ & ~new_n21745_;
  assign new_n21747_ = ~ys__n1502 & ys__n27881;
  assign new_n21748_ = ~new_n19665_ & ~new_n19670_;
  assign new_n21749_ = ~ys__n23272 & ~new_n21748_;
  assign new_n21750_ = ys__n23272 & ~new_n21614_;
  assign new_n21751_ = ~new_n21749_ & ~new_n21750_;
  assign new_n21752_ = ~ys__n23274 & ~new_n21751_;
  assign new_n21753_ = ys__n23274 & ~new_n21481_;
  assign new_n21754_ = ~new_n21752_ & ~new_n21753_;
  assign new_n21755_ = ~ys__n23276 & ~new_n21754_;
  assign new_n21756_ = ys__n23276 & ~new_n21214_;
  assign new_n21757_ = ~new_n21755_ & ~new_n21756_;
  assign new_n21758_ = ~ys__n23278 & ~new_n21757_;
  assign new_n21759_ = ys__n23278 & ~new_n20671_;
  assign new_n21760_ = ~new_n21758_ & ~new_n21759_;
  assign new_n21761_ = ys__n1502 & ~new_n21760_;
  assign new_n21762_ = ~new_n21747_ & ~new_n21761_;
  assign new_n21763_ = ~new_n19347_ & ~new_n21762_;
  assign new_n21764_ = ~new_n21746_ & ~new_n21763_;
  assign new_n21765_ = new_n19358_ & ~new_n21764_;
  assign new_n21766_ = ~new_n11857_ & new_n19360_;
  assign new_n21767_ = ys__n1498 & new_n19459_;
  assign new_n21768_ = ~new_n21766_ & ~new_n21767_;
  assign new_n21769_ = ~ys__n1496 & ~new_n21768_;
  assign new_n21770_ = ys__n1496 & ~new_n19459_;
  assign new_n21771_ = ~new_n21769_ & ~new_n21770_;
  assign new_n21772_ = ~ys__n1495 & ~new_n21771_;
  assign new_n21773_ = ys__n1495 & new_n17978_;
  assign new_n21774_ = ~new_n21772_ & ~new_n21773_;
  assign new_n21775_ = ~new_n19358_ & ~new_n21774_;
  assign new_n21776_ = ~new_n21765_ & ~new_n21775_;
  assign new_n21777_ = new_n19715_ & ~new_n21776_;
  assign new_n21778_ = ~new_n19462_ & ~new_n21713_;
  assign new_n21779_ = ~new_n11853_ & ~new_n21778_;
  assign new_n21780_ = new_n19460_ & ~new_n21779_;
  assign new_n21781_ = ~new_n19460_ & new_n21779_;
  assign new_n21782_ = ~new_n21780_ & ~new_n21781_;
  assign new_n21783_ = ~ys__n1489 & ~new_n21782_;
  assign new_n21784_ = ys__n1489 & ~new_n17975_;
  assign new_n21785_ = ~new_n21783_ & ~new_n21784_;
  assign new_n21786_ = ~new_n19561_ & ~new_n21785_;
  assign new_n21787_ = ~new_n21777_ & ~new_n21786_;
  assign new_n21788_ = ~ys__n19973 & ~new_n21787_;
  assign new_n21789_ = ys__n19973 & ys__n20002;
  assign new_n21790_ = ~new_n21788_ & ~new_n21789_;
  assign new_n21791_ = ~ys__n352 & ~new_n21790_;
  assign new_n21792_ = ~ys__n220 & ys__n47103;
  assign new_n21793_ = new_n19573_ & new_n21792_;
  assign new_n21794_ = new_n19575_ & new_n21792_;
  assign new_n21795_ = new_n19578_ & new_n20706_;
  assign new_n21796_ = ~new_n21794_ & ~new_n21795_;
  assign new_n21797_ = ~new_n21793_ & new_n21796_;
  assign new_n21798_ = new_n19587_ & ~new_n21797_;
  assign ys__n19965 = new_n21791_ | new_n21798_;
  assign new_n21800_ = ys__n19844 & ys__n19874;
  assign new_n21801_ = new_n19250_ & new_n21800_;
  assign new_n21802_ = ~ys__n23278 & ~new_n20723_;
  assign new_n21803_ = ~new_n20795_ & ~new_n21802_;
  assign new_n21804_ = ~ys__n1505 & ~new_n21803_;
  assign new_n21805_ = new_n20727_ & new_n20929_;
  assign new_n21806_ = ~new_n21804_ & ~new_n21805_;
  assign new_n21807_ = ~new_n19250_ & ~new_n21806_;
  assign new_n21808_ = ~new_n21801_ & ~new_n21807_;
  assign new_n21809_ = new_n19347_ & ~new_n21808_;
  assign new_n21810_ = ~ys__n1502 & ys__n27883;
  assign new_n21811_ = ~new_n19331_ & ~new_n19334_;
  assign new_n21812_ = ~ys__n23272 & ~new_n21811_;
  assign new_n21813_ = ys__n23272 & ~new_n21682_;
  assign new_n21814_ = ~new_n21812_ & ~new_n21813_;
  assign new_n21815_ = ~ys__n23274 & ~new_n21814_;
  assign new_n21816_ = ys__n23274 & ~new_n21549_;
  assign new_n21817_ = ~new_n21815_ & ~new_n21816_;
  assign new_n21818_ = ~ys__n23276 & ~new_n21817_;
  assign new_n21819_ = ys__n23276 & ~new_n21282_;
  assign new_n21820_ = ~new_n21818_ & ~new_n21819_;
  assign new_n21821_ = ~ys__n23278 & ~new_n21820_;
  assign new_n21822_ = ys__n23278 & ~new_n20744_;
  assign new_n21823_ = ~new_n21821_ & ~new_n21822_;
  assign new_n21824_ = ys__n1502 & ~new_n21823_;
  assign new_n21825_ = ~new_n21810_ & ~new_n21824_;
  assign new_n21826_ = ~new_n19347_ & ~new_n21825_;
  assign new_n21827_ = ~new_n21809_ & ~new_n21826_;
  assign new_n21828_ = new_n19358_ & ~new_n21827_;
  assign new_n21829_ = ~new_n11861_ & new_n19360_;
  assign new_n21830_ = ys__n1498 & new_n19456_;
  assign new_n21831_ = ~new_n21829_ & ~new_n21830_;
  assign new_n21832_ = ~ys__n1496 & ~new_n21831_;
  assign new_n21833_ = ys__n1496 & ~new_n19456_;
  assign new_n21834_ = ~new_n21832_ & ~new_n21833_;
  assign new_n21835_ = ~ys__n1495 & ~new_n21834_;
  assign new_n21836_ = ys__n1495 & new_n17990_;
  assign new_n21837_ = ~new_n21835_ & ~new_n21836_;
  assign new_n21838_ = ~new_n19358_ & ~new_n21837_;
  assign new_n21839_ = ~new_n21828_ & ~new_n21838_;
  assign new_n21840_ = new_n19715_ & ~new_n21839_;
  assign new_n21841_ = new_n19463_ & ~new_n21713_;
  assign new_n21842_ = new_n19525_ & ~new_n21841_;
  assign new_n21843_ = new_n19457_ & ~new_n21842_;
  assign new_n21844_ = ~new_n19457_ & new_n21842_;
  assign new_n21845_ = ~new_n21843_ & ~new_n21844_;
  assign new_n21846_ = ~ys__n1489 & ~new_n21845_;
  assign new_n21847_ = ys__n1489 & ~new_n17986_;
  assign new_n21848_ = ~new_n21846_ & ~new_n21847_;
  assign new_n21849_ = ~new_n19561_ & ~new_n21848_;
  assign new_n21850_ = ~new_n21840_ & ~new_n21849_;
  assign new_n21851_ = ~ys__n19973 & ~new_n21850_;
  assign new_n21852_ = ys__n19973 & ys__n20003;
  assign new_n21853_ = ~new_n21851_ & ~new_n21852_;
  assign new_n21854_ = ~ys__n352 & ~new_n21853_;
  assign new_n21855_ = ~ys__n220 & ys__n47104;
  assign new_n21856_ = new_n19573_ & new_n21855_;
  assign new_n21857_ = new_n19575_ & new_n21855_;
  assign new_n21858_ = new_n19578_ & new_n20779_;
  assign new_n21859_ = ~new_n21857_ & ~new_n21858_;
  assign new_n21860_ = ~new_n21856_ & new_n21859_;
  assign new_n21861_ = new_n19587_ & ~new_n21860_;
  assign ys__n19968 = new_n21854_ | new_n21861_;
  assign new_n21863_ = ys__n19844 & ys__n19875;
  assign new_n21864_ = new_n19250_ & new_n21863_;
  assign new_n21865_ = ~ys__n1505 & ys__n28030;
  assign new_n21866_ = new_n20798_ & new_n20929_;
  assign new_n21867_ = ~new_n21865_ & ~new_n21866_;
  assign new_n21868_ = ~new_n19250_ & ~new_n21867_;
  assign new_n21869_ = ~new_n21864_ & ~new_n21868_;
  assign new_n21870_ = new_n19347_ & ~new_n21869_;
  assign new_n21871_ = ~ys__n1502 & ys__n27885;
  assign new_n21872_ = ~new_n19671_ & ~new_n19683_;
  assign new_n21873_ = ~ys__n23272 & ~new_n21872_;
  assign new_n21874_ = ys__n23272 & ~new_n21748_;
  assign new_n21875_ = ~new_n21873_ & ~new_n21874_;
  assign new_n21876_ = ~ys__n23274 & ~new_n21875_;
  assign new_n21877_ = ys__n23274 & ~new_n21617_;
  assign new_n21878_ = ~new_n21876_ & ~new_n21877_;
  assign new_n21879_ = ~ys__n23276 & ~new_n21878_;
  assign new_n21880_ = ys__n23276 & ~new_n21350_;
  assign new_n21881_ = ~new_n21879_ & ~new_n21880_;
  assign new_n21882_ = ~ys__n23278 & ~new_n21881_;
  assign new_n21883_ = ys__n23278 & ~new_n20815_;
  assign new_n21884_ = ~new_n21882_ & ~new_n21883_;
  assign new_n21885_ = ys__n1502 & ~new_n21884_;
  assign new_n21886_ = ~new_n21871_ & ~new_n21885_;
  assign new_n21887_ = ~new_n19347_ & ~new_n21886_;
  assign new_n21888_ = ~new_n21870_ & ~new_n21887_;
  assign new_n21889_ = new_n19358_ & ~new_n21888_;
  assign new_n21890_ = ~new_n11864_ & new_n19360_;
  assign new_n21891_ = ys__n1498 & new_n19453_;
  assign new_n21892_ = ~new_n21890_ & ~new_n21891_;
  assign new_n21893_ = ~ys__n1496 & ~new_n21892_;
  assign new_n21894_ = ys__n1496 & ~new_n19453_;
  assign new_n21895_ = ~new_n21893_ & ~new_n21894_;
  assign new_n21896_ = ~ys__n1495 & ~new_n21895_;
  assign new_n21897_ = ys__n1495 & new_n19454_;
  assign new_n21898_ = ~new_n21896_ & ~new_n21897_;
  assign new_n21899_ = ~new_n19358_ & ~new_n21898_;
  assign new_n21900_ = ~new_n21889_ & ~new_n21899_;
  assign new_n21901_ = new_n19715_ & ~new_n21900_;
  assign new_n21902_ = ~new_n19457_ & ~new_n21842_;
  assign new_n21903_ = ~new_n11860_ & ~new_n21902_;
  assign new_n21904_ = new_n19455_ & ~new_n21903_;
  assign new_n21905_ = ~new_n19455_ & new_n21903_;
  assign new_n21906_ = ~new_n21904_ & ~new_n21905_;
  assign new_n21907_ = ~ys__n1489 & ~new_n21906_;
  assign new_n21908_ = ys__n1489 & ~new_n17995_;
  assign new_n21909_ = ~new_n21907_ & ~new_n21908_;
  assign new_n21910_ = ~new_n19561_ & ~new_n21909_;
  assign new_n21911_ = ~new_n21901_ & ~new_n21910_;
  assign new_n21912_ = ~ys__n19973 & ~new_n21911_;
  assign new_n21913_ = ys__n19973 & ys__n20004;
  assign new_n21914_ = ~new_n21912_ & ~new_n21913_;
  assign new_n21915_ = ~ys__n352 & ~new_n21914_;
  assign new_n21916_ = ~ys__n220 & ys__n47105;
  assign new_n21917_ = new_n19573_ & new_n21916_;
  assign new_n21918_ = new_n19575_ & new_n21916_;
  assign new_n21919_ = new_n19578_ & new_n20850_;
  assign new_n21920_ = ~new_n21918_ & ~new_n21919_;
  assign new_n21921_ = ~new_n21917_ & new_n21920_;
  assign new_n21922_ = new_n19587_ & ~new_n21921_;
  assign ys__n19971 = new_n21915_ | new_n21922_;
  assign new_n21924_ = ~new_n11901_ & ~new_n17866_;
  assign ys__n20006 = new_n17867_ | new_n21924_;
  assign new_n21926_ = ~new_n17746_ & ~new_n17866_;
  assign ys__n20007 = new_n17867_ | new_n21926_;
  assign new_n21928_ = ~new_n17866_ & ~new_n19824_;
  assign ys__n20008 = new_n17867_ | new_n21928_;
  assign new_n21930_ = ~new_n17866_ & ~new_n19931_;
  assign ys__n20009 = new_n17867_ | new_n21930_;
  assign new_n21932_ = ~new_n17866_ & ~new_n20011_;
  assign ys__n20010 = new_n17867_ | new_n21932_;
  assign new_n21934_ = ~new_n17866_ & ~new_n20096_;
  assign ys__n20011 = new_n17867_ | new_n21934_;
  assign new_n21936_ = ~new_n17866_ & ~new_n20181_;
  assign ys__n20012 = new_n17867_ | new_n21936_;
  assign new_n21938_ = ~new_n17866_ & ~new_n20264_;
  assign ys__n20013 = new_n17867_ | new_n21938_;
  assign new_n21940_ = ~new_n17866_ & ~new_n20332_;
  assign ys__n20014 = new_n17867_ | new_n21940_;
  assign new_n21942_ = ~new_n17866_ & ~new_n20405_;
  assign ys__n20015 = new_n17867_ | new_n21942_;
  assign new_n21944_ = ~new_n17866_ & ~new_n20478_;
  assign ys__n20016 = new_n17867_ | new_n21944_;
  assign new_n21946_ = ~new_n17866_ & ~new_n20551_;
  assign ys__n20017 = new_n17867_ | new_n21946_;
  assign new_n21948_ = ~new_n17866_ & ~new_n20624_;
  assign ys__n20018 = new_n17867_ | new_n21948_;
  assign new_n21950_ = ~new_n17866_ & ~new_n20697_;
  assign ys__n20019 = new_n17867_ | new_n21950_;
  assign new_n21952_ = ~new_n17866_ & ~new_n20770_;
  assign ys__n20020 = new_n17867_ | new_n21952_;
  assign new_n21954_ = ~new_n17866_ & ~new_n20841_;
  assign ys__n20021 = new_n17867_ | new_n21954_;
  assign new_n21956_ = ~new_n17866_ & ~new_n20907_;
  assign ys__n20022 = new_n17867_ | new_n21956_;
  assign new_n21958_ = ~new_n17866_ & ~new_n20976_;
  assign ys__n20023 = new_n17867_ | new_n21958_;
  assign new_n21960_ = ~new_n17866_ & ~new_n21044_;
  assign ys__n20024 = new_n17867_ | new_n21960_;
  assign new_n21962_ = ~new_n17866_ & ~new_n21112_;
  assign ys__n20025 = new_n17867_ | new_n21962_;
  assign new_n21964_ = ~new_n17866_ & ~new_n21180_;
  assign ys__n20026 = new_n17867_ | new_n21964_;
  assign new_n21966_ = ~new_n17866_ & ~new_n21248_;
  assign ys__n20027 = new_n17867_ | new_n21966_;
  assign new_n21968_ = ~new_n17866_ & ~new_n21316_;
  assign ys__n20028 = new_n17867_ | new_n21968_;
  assign new_n21970_ = ~new_n17866_ & ~new_n21384_;
  assign ys__n20029 = new_n17867_ | new_n21970_;
  assign new_n21972_ = ~new_n17866_ & ~new_n21450_;
  assign ys__n20030 = new_n17867_ | new_n21972_;
  assign new_n21974_ = ~new_n17866_ & ~new_n21518_;
  assign ys__n20031 = new_n17867_ | new_n21974_;
  assign new_n21976_ = ~new_n17866_ & ~new_n21586_;
  assign ys__n20032 = new_n17867_ | new_n21976_;
  assign new_n21978_ = ~new_n17866_ & ~new_n21654_;
  assign ys__n20033 = new_n17867_ | new_n21978_;
  assign new_n21980_ = ~new_n17866_ & ~new_n21720_;
  assign ys__n20034 = new_n17867_ | new_n21980_;
  assign new_n21982_ = ys__n1508 & new_n17750_;
  assign new_n21983_ = ~new_n17753_ & new_n21982_;
  assign ys__n20038 = new_n17766_ | new_n21983_;
  assign new_n21985_ = ys__n1508 & new_n17747_;
  assign new_n21986_ = ~new_n17753_ & new_n21985_;
  assign ys__n20043 = new_n17759_ | new_n21986_;
  assign new_n21988_ = ~new_n17747_ & ~new_n17750_;
  assign new_n21989_ = ~new_n17751_ & new_n21988_;
  assign new_n21990_ = ~new_n17748_ & new_n21989_;
  assign new_n21991_ = new_n17754_ & ~new_n21989_;
  assign new_n21992_ = ~new_n21990_ & new_n21991_;
  assign new_n21993_ = ~new_n17748_ & ~new_n17751_;
  assign new_n21994_ = new_n21988_ & new_n21993_;
  assign new_n21995_ = ys__n1509 & ~new_n21988_;
  assign new_n21996_ = ~new_n21994_ & new_n21995_;
  assign new_n21997_ = ~new_n21992_ & ~new_n21996_;
  assign ys__n20053 = ~ys__n1508 & ~new_n21997_;
  assign new_n21999_ = ~ys__n1511 & ys__n20035;
  assign new_n22000_ = ys__n20058 & new_n21999_;
  assign new_n22001_ = ys__n1511 & ys__n20058;
  assign new_n22002_ = ~new_n22000_ & ~new_n22001_;
  assign new_n22003_ = ~ys__n1509 & ~new_n22002_;
  assign new_n22004_ = ys__n1509 & ys__n20058;
  assign new_n22005_ = ~new_n22003_ & ~new_n22004_;
  assign new_n22006_ = ~ys__n1508 & ~new_n22005_;
  assign new_n22007_ = ys__n1508 & ys__n20058;
  assign ys__n20059 = new_n22006_ | new_n22007_;
  assign new_n22009_ = ys__n20061 & new_n21999_;
  assign new_n22010_ = ys__n1511 & ys__n20061;
  assign new_n22011_ = ~new_n22009_ & ~new_n22010_;
  assign new_n22012_ = ~ys__n1509 & ~new_n22011_;
  assign new_n22013_ = ys__n1509 & ys__n20061;
  assign new_n22014_ = ~new_n22012_ & ~new_n22013_;
  assign new_n22015_ = ~ys__n1508 & ~new_n22014_;
  assign new_n22016_ = ys__n1508 & ys__n20061;
  assign ys__n20062 = new_n22015_ | new_n22016_;
  assign new_n22018_ = ys__n20064 & new_n21999_;
  assign new_n22019_ = ys__n1511 & ys__n20064;
  assign new_n22020_ = ~new_n22018_ & ~new_n22019_;
  assign new_n22021_ = ~ys__n1509 & ~new_n22020_;
  assign new_n22022_ = ys__n1509 & ys__n20064;
  assign new_n22023_ = ~new_n22021_ & ~new_n22022_;
  assign new_n22024_ = ~ys__n1508 & ~new_n22023_;
  assign new_n22025_ = ys__n1508 & ys__n20064;
  assign ys__n20065 = new_n22024_ | new_n22025_;
  assign new_n22027_ = ys__n20067 & new_n21999_;
  assign new_n22028_ = ys__n1511 & ys__n20067;
  assign new_n22029_ = ~new_n22027_ & ~new_n22028_;
  assign new_n22030_ = ~ys__n1509 & ~new_n22029_;
  assign new_n22031_ = ys__n1509 & ys__n20067;
  assign new_n22032_ = ~new_n22030_ & ~new_n22031_;
  assign new_n22033_ = ~ys__n1508 & ~new_n22032_;
  assign new_n22034_ = ys__n1508 & ys__n20067;
  assign ys__n20068 = new_n22033_ | new_n22034_;
  assign new_n22036_ = ys__n20070 & new_n21999_;
  assign new_n22037_ = ys__n1511 & ys__n20070;
  assign new_n22038_ = ~new_n22036_ & ~new_n22037_;
  assign new_n22039_ = ~ys__n1509 & ~new_n22038_;
  assign new_n22040_ = ys__n1509 & ys__n20070;
  assign new_n22041_ = ~new_n22039_ & ~new_n22040_;
  assign new_n22042_ = ~ys__n1508 & ~new_n22041_;
  assign new_n22043_ = ys__n1508 & ys__n20070;
  assign ys__n20071 = new_n22042_ | new_n22043_;
  assign new_n22045_ = ys__n20073 & new_n21999_;
  assign new_n22046_ = ys__n1511 & ys__n20073;
  assign new_n22047_ = ~new_n22045_ & ~new_n22046_;
  assign new_n22048_ = ~ys__n1509 & ~new_n22047_;
  assign new_n22049_ = ys__n1509 & ys__n20073;
  assign new_n22050_ = ~new_n22048_ & ~new_n22049_;
  assign new_n22051_ = ~ys__n1508 & ~new_n22050_;
  assign new_n22052_ = ys__n1508 & ys__n20073;
  assign ys__n20074 = new_n22051_ | new_n22052_;
  assign new_n22054_ = ys__n20076 & new_n21999_;
  assign new_n22055_ = ys__n1511 & ys__n20076;
  assign new_n22056_ = ~new_n22054_ & ~new_n22055_;
  assign new_n22057_ = ~ys__n1509 & ~new_n22056_;
  assign new_n22058_ = ys__n1509 & ys__n20076;
  assign new_n22059_ = ~new_n22057_ & ~new_n22058_;
  assign new_n22060_ = ~ys__n1508 & ~new_n22059_;
  assign new_n22061_ = ys__n1508 & ys__n20076;
  assign ys__n20077 = new_n22060_ | new_n22061_;
  assign new_n22063_ = ys__n20079 & new_n21999_;
  assign new_n22064_ = ys__n1511 & ys__n20079;
  assign new_n22065_ = ~new_n22063_ & ~new_n22064_;
  assign new_n22066_ = ~ys__n1509 & ~new_n22065_;
  assign new_n22067_ = ys__n1509 & ys__n20079;
  assign new_n22068_ = ~new_n22066_ & ~new_n22067_;
  assign new_n22069_ = ~ys__n1508 & ~new_n22068_;
  assign new_n22070_ = ys__n1508 & ys__n20079;
  assign ys__n20080 = new_n22069_ | new_n22070_;
  assign new_n22072_ = ys__n20138 & new_n21999_;
  assign new_n22073_ = ys__n1511 & ys__n20138;
  assign new_n22074_ = ~new_n22072_ & ~new_n22073_;
  assign new_n22075_ = ~ys__n1509 & ~new_n22074_;
  assign new_n22076_ = ys__n1509 & ys__n20138;
  assign new_n22077_ = ~new_n22075_ & ~new_n22076_;
  assign new_n22078_ = ~ys__n1508 & ~new_n22077_;
  assign ys__n20082 = new_n22007_ | new_n22078_;
  assign new_n22080_ = ys__n20140 & new_n21999_;
  assign new_n22081_ = ys__n1511 & ys__n20140;
  assign new_n22082_ = ~new_n22080_ & ~new_n22081_;
  assign new_n22083_ = ~ys__n1509 & ~new_n22082_;
  assign new_n22084_ = ys__n1509 & ys__n20140;
  assign new_n22085_ = ~new_n22083_ & ~new_n22084_;
  assign new_n22086_ = ~ys__n1508 & ~new_n22085_;
  assign ys__n20084 = new_n22016_ | new_n22086_;
  assign new_n22088_ = ys__n20142 & new_n21999_;
  assign new_n22089_ = ys__n1511 & ys__n20142;
  assign new_n22090_ = ~new_n22088_ & ~new_n22089_;
  assign new_n22091_ = ~ys__n1509 & ~new_n22090_;
  assign new_n22092_ = ys__n1509 & ys__n20142;
  assign new_n22093_ = ~new_n22091_ & ~new_n22092_;
  assign new_n22094_ = ~ys__n1508 & ~new_n22093_;
  assign ys__n20086 = new_n22025_ | new_n22094_;
  assign new_n22096_ = ys__n20144 & new_n21999_;
  assign new_n22097_ = ys__n1511 & ys__n20144;
  assign new_n22098_ = ~new_n22096_ & ~new_n22097_;
  assign new_n22099_ = ~ys__n1509 & ~new_n22098_;
  assign new_n22100_ = ys__n1509 & ys__n20144;
  assign new_n22101_ = ~new_n22099_ & ~new_n22100_;
  assign new_n22102_ = ~ys__n1508 & ~new_n22101_;
  assign ys__n20088 = new_n22034_ | new_n22102_;
  assign new_n22104_ = ys__n20146 & new_n21999_;
  assign new_n22105_ = ys__n1511 & ys__n20146;
  assign new_n22106_ = ~new_n22104_ & ~new_n22105_;
  assign new_n22107_ = ~ys__n1509 & ~new_n22106_;
  assign new_n22108_ = ys__n1509 & ys__n20146;
  assign new_n22109_ = ~new_n22107_ & ~new_n22108_;
  assign new_n22110_ = ~ys__n1508 & ~new_n22109_;
  assign ys__n20090 = new_n22043_ | new_n22110_;
  assign new_n22112_ = ys__n20148 & new_n21999_;
  assign new_n22113_ = ys__n1511 & ys__n20148;
  assign new_n22114_ = ~new_n22112_ & ~new_n22113_;
  assign new_n22115_ = ~ys__n1509 & ~new_n22114_;
  assign new_n22116_ = ys__n1509 & ys__n20148;
  assign new_n22117_ = ~new_n22115_ & ~new_n22116_;
  assign new_n22118_ = ~ys__n1508 & ~new_n22117_;
  assign ys__n20092 = new_n22052_ | new_n22118_;
  assign new_n22120_ = ys__n20150 & new_n21999_;
  assign new_n22121_ = ys__n1511 & ys__n20150;
  assign new_n22122_ = ~new_n22120_ & ~new_n22121_;
  assign new_n22123_ = ~ys__n1509 & ~new_n22122_;
  assign new_n22124_ = ys__n1509 & ys__n20150;
  assign new_n22125_ = ~new_n22123_ & ~new_n22124_;
  assign new_n22126_ = ~ys__n1508 & ~new_n22125_;
  assign ys__n20094 = new_n22061_ | new_n22126_;
  assign new_n22128_ = ys__n20152 & new_n21999_;
  assign new_n22129_ = ys__n1511 & ys__n20152;
  assign new_n22130_ = ~new_n22128_ & ~new_n22129_;
  assign new_n22131_ = ~ys__n1509 & ~new_n22130_;
  assign new_n22132_ = ys__n1509 & ys__n20152;
  assign new_n22133_ = ~new_n22131_ & ~new_n22132_;
  assign new_n22134_ = ~ys__n1508 & ~new_n22133_;
  assign ys__n20096 = new_n22070_ | new_n22134_;
  assign new_n22136_ = ys__n20186 & new_n21999_;
  assign new_n22137_ = ys__n1511 & ys__n20186;
  assign new_n22138_ = ~new_n22136_ & ~new_n22137_;
  assign new_n22139_ = ~ys__n1509 & ~new_n22138_;
  assign new_n22140_ = ~new_n22004_ & ~new_n22139_;
  assign new_n22141_ = ~ys__n1508 & ~new_n22140_;
  assign ys__n20098 = new_n22007_ | new_n22141_;
  assign new_n22143_ = ys__n20188 & new_n21999_;
  assign new_n22144_ = ys__n1511 & ys__n20188;
  assign new_n22145_ = ~new_n22143_ & ~new_n22144_;
  assign new_n22146_ = ~ys__n1509 & ~new_n22145_;
  assign new_n22147_ = ~new_n22013_ & ~new_n22146_;
  assign new_n22148_ = ~ys__n1508 & ~new_n22147_;
  assign ys__n20100 = new_n22016_ | new_n22148_;
  assign new_n22150_ = ys__n20190 & new_n21999_;
  assign new_n22151_ = ys__n1511 & ys__n20190;
  assign new_n22152_ = ~new_n22150_ & ~new_n22151_;
  assign new_n22153_ = ~ys__n1509 & ~new_n22152_;
  assign new_n22154_ = ~new_n22022_ & ~new_n22153_;
  assign new_n22155_ = ~ys__n1508 & ~new_n22154_;
  assign ys__n20102 = new_n22025_ | new_n22155_;
  assign new_n22157_ = ys__n20192 & new_n21999_;
  assign new_n22158_ = ys__n1511 & ys__n20192;
  assign new_n22159_ = ~new_n22157_ & ~new_n22158_;
  assign new_n22160_ = ~ys__n1509 & ~new_n22159_;
  assign new_n22161_ = ~new_n22031_ & ~new_n22160_;
  assign new_n22162_ = ~ys__n1508 & ~new_n22161_;
  assign ys__n20104 = new_n22034_ | new_n22162_;
  assign new_n22164_ = ys__n20194 & new_n21999_;
  assign new_n22165_ = ys__n1511 & ys__n20194;
  assign new_n22166_ = ~new_n22164_ & ~new_n22165_;
  assign new_n22167_ = ~ys__n1509 & ~new_n22166_;
  assign new_n22168_ = ~new_n22040_ & ~new_n22167_;
  assign new_n22169_ = ~ys__n1508 & ~new_n22168_;
  assign ys__n20106 = new_n22043_ | new_n22169_;
  assign new_n22171_ = ys__n20196 & new_n21999_;
  assign new_n22172_ = ys__n1511 & ys__n20196;
  assign new_n22173_ = ~new_n22171_ & ~new_n22172_;
  assign new_n22174_ = ~ys__n1509 & ~new_n22173_;
  assign new_n22175_ = ~new_n22049_ & ~new_n22174_;
  assign new_n22176_ = ~ys__n1508 & ~new_n22175_;
  assign ys__n20108 = new_n22052_ | new_n22176_;
  assign new_n22178_ = ys__n20198 & new_n21999_;
  assign new_n22179_ = ys__n1511 & ys__n20198;
  assign new_n22180_ = ~new_n22178_ & ~new_n22179_;
  assign new_n22181_ = ~ys__n1509 & ~new_n22180_;
  assign new_n22182_ = ~new_n22058_ & ~new_n22181_;
  assign new_n22183_ = ~ys__n1508 & ~new_n22182_;
  assign ys__n20110 = new_n22061_ | new_n22183_;
  assign new_n22185_ = ys__n20200 & new_n21999_;
  assign new_n22186_ = ys__n1511 & ys__n20200;
  assign new_n22187_ = ~new_n22185_ & ~new_n22186_;
  assign new_n22188_ = ~ys__n1509 & ~new_n22187_;
  assign new_n22189_ = ~new_n22067_ & ~new_n22188_;
  assign new_n22190_ = ~ys__n1508 & ~new_n22189_;
  assign ys__n20112 = new_n22070_ | new_n22190_;
  assign new_n22192_ = ys__n20202 & new_n21999_;
  assign new_n22193_ = ys__n1511 & ys__n20202;
  assign new_n22194_ = ~new_n22192_ & ~new_n22193_;
  assign new_n22195_ = ~ys__n1509 & ~new_n22194_;
  assign new_n22196_ = ~new_n22076_ & ~new_n22195_;
  assign new_n22197_ = ~ys__n1508 & ~new_n22196_;
  assign ys__n20114 = new_n22007_ | new_n22197_;
  assign new_n22199_ = ys__n20204 & new_n21999_;
  assign new_n22200_ = ys__n1511 & ys__n20204;
  assign new_n22201_ = ~new_n22199_ & ~new_n22200_;
  assign new_n22202_ = ~ys__n1509 & ~new_n22201_;
  assign new_n22203_ = ~new_n22084_ & ~new_n22202_;
  assign new_n22204_ = ~ys__n1508 & ~new_n22203_;
  assign ys__n20116 = new_n22016_ | new_n22204_;
  assign new_n22206_ = ys__n20206 & new_n21999_;
  assign new_n22207_ = ys__n1511 & ys__n20206;
  assign new_n22208_ = ~new_n22206_ & ~new_n22207_;
  assign new_n22209_ = ~ys__n1509 & ~new_n22208_;
  assign new_n22210_ = ~new_n22092_ & ~new_n22209_;
  assign new_n22211_ = ~ys__n1508 & ~new_n22210_;
  assign ys__n20118 = new_n22025_ | new_n22211_;
  assign new_n22213_ = ys__n20208 & new_n21999_;
  assign new_n22214_ = ys__n1511 & ys__n20208;
  assign new_n22215_ = ~new_n22213_ & ~new_n22214_;
  assign new_n22216_ = ~ys__n1509 & ~new_n22215_;
  assign new_n22217_ = ~new_n22100_ & ~new_n22216_;
  assign new_n22218_ = ~ys__n1508 & ~new_n22217_;
  assign ys__n20120 = new_n22034_ | new_n22218_;
  assign new_n22220_ = ys__n20210 & new_n21999_;
  assign new_n22221_ = ys__n1511 & ys__n20210;
  assign new_n22222_ = ~new_n22220_ & ~new_n22221_;
  assign new_n22223_ = ~ys__n1509 & ~new_n22222_;
  assign new_n22224_ = ~new_n22108_ & ~new_n22223_;
  assign new_n22225_ = ~ys__n1508 & ~new_n22224_;
  assign ys__n20122 = new_n22043_ | new_n22225_;
  assign new_n22227_ = ys__n20212 & new_n21999_;
  assign new_n22228_ = ys__n1511 & ys__n20212;
  assign new_n22229_ = ~new_n22227_ & ~new_n22228_;
  assign new_n22230_ = ~ys__n1509 & ~new_n22229_;
  assign new_n22231_ = ~new_n22116_ & ~new_n22230_;
  assign new_n22232_ = ~ys__n1508 & ~new_n22231_;
  assign ys__n20124 = new_n22052_ | new_n22232_;
  assign new_n22234_ = ys__n20214 & new_n21999_;
  assign new_n22235_ = ys__n1511 & ys__n20214;
  assign new_n22236_ = ~new_n22234_ & ~new_n22235_;
  assign new_n22237_ = ~ys__n1509 & ~new_n22236_;
  assign new_n22238_ = ~new_n22124_ & ~new_n22237_;
  assign new_n22239_ = ~ys__n1508 & ~new_n22238_;
  assign ys__n20126 = new_n22061_ | new_n22239_;
  assign new_n22241_ = ys__n20216 & new_n21999_;
  assign new_n22242_ = ys__n1511 & ys__n20216;
  assign new_n22243_ = ~new_n22241_ & ~new_n22242_;
  assign new_n22244_ = ~ys__n1509 & ~new_n22243_;
  assign new_n22245_ = ~new_n22132_ & ~new_n22244_;
  assign new_n22246_ = ~ys__n1508 & ~new_n22245_;
  assign ys__n20128 = new_n22070_ | new_n22246_;
  assign new_n22248_ = ys__n23077 & ~new_n13442_;
  assign new_n22249_ = new_n13439_ & new_n22248_;
  assign new_n22250_ = ys__n23014 & new_n13442_;
  assign new_n22251_ = ~new_n22249_ & ~new_n22250_;
  assign new_n22252_ = ~new_n13440_ & ~new_n22251_;
  assign new_n22253_ = ys__n22918 & new_n13440_;
  assign ys__n22919 = new_n22252_ | new_n22253_;
  assign new_n22255_ = ys__n23078 & ~new_n13442_;
  assign new_n22256_ = new_n13439_ & new_n22255_;
  assign new_n22257_ = ys__n23016 & new_n13442_;
  assign new_n22258_ = ~new_n22256_ & ~new_n22257_;
  assign new_n22259_ = ~new_n13440_ & ~new_n22258_;
  assign new_n22260_ = ys__n22921 & new_n13440_;
  assign ys__n22922 = new_n22259_ | new_n22260_;
  assign new_n22262_ = ys__n23079 & ~new_n13442_;
  assign new_n22263_ = new_n13439_ & new_n22262_;
  assign new_n22264_ = ys__n23018 & new_n13442_;
  assign new_n22265_ = ~new_n22263_ & ~new_n22264_;
  assign new_n22266_ = ~new_n13440_ & ~new_n22265_;
  assign new_n22267_ = ys__n22924 & new_n13440_;
  assign ys__n22925 = new_n22266_ | new_n22267_;
  assign new_n22269_ = ys__n23080 & ~new_n13442_;
  assign new_n22270_ = new_n13439_ & new_n22269_;
  assign new_n22271_ = ys__n23020 & new_n13442_;
  assign new_n22272_ = ~new_n22270_ & ~new_n22271_;
  assign new_n22273_ = ~new_n13440_ & ~new_n22272_;
  assign new_n22274_ = ys__n22927 & new_n13440_;
  assign ys__n22928 = new_n22273_ | new_n22274_;
  assign new_n22276_ = ys__n23081 & ~new_n13442_;
  assign new_n22277_ = new_n13439_ & new_n22276_;
  assign new_n22278_ = ys__n23022 & new_n13442_;
  assign new_n22279_ = ~new_n22277_ & ~new_n22278_;
  assign new_n22280_ = ~new_n13440_ & ~new_n22279_;
  assign new_n22281_ = ys__n22930 & new_n13440_;
  assign ys__n22931 = new_n22280_ | new_n22281_;
  assign new_n22283_ = ys__n23082 & ~new_n13442_;
  assign new_n22284_ = new_n13439_ & new_n22283_;
  assign new_n22285_ = ys__n23024 & new_n13442_;
  assign new_n22286_ = ~new_n22284_ & ~new_n22285_;
  assign new_n22287_ = ~new_n13440_ & ~new_n22286_;
  assign new_n22288_ = ys__n22933 & new_n13440_;
  assign ys__n22934 = new_n22287_ | new_n22288_;
  assign new_n22290_ = ys__n23083 & ~new_n13442_;
  assign new_n22291_ = new_n13439_ & new_n22290_;
  assign new_n22292_ = ys__n23026 & new_n13442_;
  assign new_n22293_ = ~new_n22291_ & ~new_n22292_;
  assign new_n22294_ = ~new_n13440_ & ~new_n22293_;
  assign new_n22295_ = ys__n22936 & new_n13440_;
  assign ys__n22937 = new_n22294_ | new_n22295_;
  assign new_n22297_ = ys__n23084 & ~new_n13442_;
  assign new_n22298_ = new_n13439_ & new_n22297_;
  assign new_n22299_ = ys__n23028 & new_n13442_;
  assign new_n22300_ = ~new_n22298_ & ~new_n22299_;
  assign new_n22301_ = ~new_n13440_ & ~new_n22300_;
  assign new_n22302_ = ys__n22939 & new_n13440_;
  assign ys__n22940 = new_n22301_ | new_n22302_;
  assign new_n22304_ = ys__n23085 & ~new_n13442_;
  assign new_n22305_ = new_n13439_ & new_n22304_;
  assign new_n22306_ = ys__n23030 & new_n13442_;
  assign new_n22307_ = ~new_n22305_ & ~new_n22306_;
  assign new_n22308_ = ~new_n13440_ & ~new_n22307_;
  assign new_n22309_ = ys__n22942 & new_n13440_;
  assign ys__n22943 = new_n22308_ | new_n22309_;
  assign new_n22311_ = ys__n23086 & ~new_n13442_;
  assign new_n22312_ = new_n13439_ & new_n22311_;
  assign new_n22313_ = ys__n23032 & new_n13442_;
  assign new_n22314_ = ~new_n22312_ & ~new_n22313_;
  assign new_n22315_ = ~new_n13440_ & ~new_n22314_;
  assign new_n22316_ = ys__n22945 & new_n13440_;
  assign ys__n22946 = new_n22315_ | new_n22316_;
  assign new_n22318_ = ys__n23087 & ~new_n13442_;
  assign new_n22319_ = new_n13439_ & new_n22318_;
  assign new_n22320_ = ys__n23034 & new_n13442_;
  assign new_n22321_ = ~new_n22319_ & ~new_n22320_;
  assign new_n22322_ = ~new_n13440_ & ~new_n22321_;
  assign new_n22323_ = ys__n22948 & new_n13440_;
  assign ys__n22949 = new_n22322_ | new_n22323_;
  assign new_n22325_ = ys__n23088 & ~new_n13442_;
  assign new_n22326_ = new_n13439_ & new_n22325_;
  assign new_n22327_ = ys__n23036 & new_n13442_;
  assign new_n22328_ = ~new_n22326_ & ~new_n22327_;
  assign new_n22329_ = ~new_n13440_ & ~new_n22328_;
  assign new_n22330_ = ys__n22951 & new_n13440_;
  assign ys__n22952 = new_n22329_ | new_n22330_;
  assign new_n22332_ = ys__n23089 & ~new_n13442_;
  assign new_n22333_ = new_n13439_ & new_n22332_;
  assign new_n22334_ = ys__n23038 & new_n13442_;
  assign new_n22335_ = ~new_n22333_ & ~new_n22334_;
  assign new_n22336_ = ~new_n13440_ & ~new_n22335_;
  assign new_n22337_ = ys__n22954 & new_n13440_;
  assign ys__n22955 = new_n22336_ | new_n22337_;
  assign new_n22339_ = ys__n23090 & ~new_n13442_;
  assign new_n22340_ = new_n13439_ & new_n22339_;
  assign new_n22341_ = ys__n23040 & new_n13442_;
  assign new_n22342_ = ~new_n22340_ & ~new_n22341_;
  assign new_n22343_ = ~new_n13440_ & ~new_n22342_;
  assign new_n22344_ = ys__n22957 & new_n13440_;
  assign ys__n22958 = new_n22343_ | new_n22344_;
  assign new_n22346_ = ys__n23091 & ~new_n13442_;
  assign new_n22347_ = new_n13439_ & new_n22346_;
  assign new_n22348_ = ys__n23042 & new_n13442_;
  assign new_n22349_ = ~new_n22347_ & ~new_n22348_;
  assign new_n22350_ = ~new_n13440_ & ~new_n22349_;
  assign new_n22351_ = ys__n22960 & new_n13440_;
  assign ys__n22961 = new_n22350_ | new_n22351_;
  assign new_n22353_ = ys__n23092 & ~new_n13442_;
  assign new_n22354_ = new_n13439_ & new_n22353_;
  assign new_n22355_ = ys__n23044 & new_n13442_;
  assign new_n22356_ = ~new_n22354_ & ~new_n22355_;
  assign new_n22357_ = ~new_n13440_ & ~new_n22356_;
  assign new_n22358_ = ys__n22963 & new_n13440_;
  assign ys__n22964 = new_n22357_ | new_n22358_;
  assign new_n22360_ = ys__n23093 & ~new_n13442_;
  assign new_n22361_ = new_n13439_ & new_n22360_;
  assign new_n22362_ = ys__n23046 & new_n13442_;
  assign new_n22363_ = ~new_n22361_ & ~new_n22362_;
  assign new_n22364_ = ~new_n13440_ & ~new_n22363_;
  assign new_n22365_ = ys__n22966 & new_n13440_;
  assign ys__n22967 = new_n22364_ | new_n22365_;
  assign new_n22367_ = ys__n23094 & ~new_n13442_;
  assign new_n22368_ = new_n13439_ & new_n22367_;
  assign new_n22369_ = ys__n23048 & new_n13442_;
  assign new_n22370_ = ~new_n22368_ & ~new_n22369_;
  assign new_n22371_ = ~new_n13440_ & ~new_n22370_;
  assign new_n22372_ = ys__n22969 & new_n13440_;
  assign ys__n22970 = new_n22371_ | new_n22372_;
  assign new_n22374_ = ys__n23095 & ~new_n13442_;
  assign new_n22375_ = new_n13439_ & new_n22374_;
  assign new_n22376_ = ys__n23050 & new_n13442_;
  assign new_n22377_ = ~new_n22375_ & ~new_n22376_;
  assign new_n22378_ = ~new_n13440_ & ~new_n22377_;
  assign new_n22379_ = ys__n22972 & new_n13440_;
  assign ys__n22973 = new_n22378_ | new_n22379_;
  assign new_n22381_ = ys__n23096 & ~new_n13442_;
  assign new_n22382_ = new_n13439_ & new_n22381_;
  assign new_n22383_ = ys__n23052 & new_n13442_;
  assign new_n22384_ = ~new_n22382_ & ~new_n22383_;
  assign new_n22385_ = ~new_n13440_ & ~new_n22384_;
  assign new_n22386_ = ys__n22975 & new_n13440_;
  assign ys__n22976 = new_n22385_ | new_n22386_;
  assign new_n22388_ = ys__n23097 & ~new_n13442_;
  assign new_n22389_ = new_n13439_ & new_n22388_;
  assign new_n22390_ = ys__n23054 & new_n13442_;
  assign new_n22391_ = ~new_n22389_ & ~new_n22390_;
  assign new_n22392_ = ~new_n13440_ & ~new_n22391_;
  assign new_n22393_ = ys__n22978 & new_n13440_;
  assign ys__n22979 = new_n22392_ | new_n22393_;
  assign new_n22395_ = ys__n23098 & ~new_n13442_;
  assign new_n22396_ = new_n13439_ & new_n22395_;
  assign new_n22397_ = ys__n23056 & new_n13442_;
  assign new_n22398_ = ~new_n22396_ & ~new_n22397_;
  assign new_n22399_ = ~new_n13440_ & ~new_n22398_;
  assign new_n22400_ = ys__n22981 & new_n13440_;
  assign ys__n22982 = new_n22399_ | new_n22400_;
  assign new_n22402_ = ys__n23099 & ~new_n13442_;
  assign new_n22403_ = new_n13439_ & new_n22402_;
  assign new_n22404_ = ys__n23058 & new_n13442_;
  assign new_n22405_ = ~new_n22403_ & ~new_n22404_;
  assign new_n22406_ = ~new_n13440_ & ~new_n22405_;
  assign new_n22407_ = ys__n22984 & new_n13440_;
  assign ys__n22985 = new_n22406_ | new_n22407_;
  assign new_n22409_ = ys__n23100 & ~new_n13442_;
  assign new_n22410_ = new_n13439_ & new_n22409_;
  assign new_n22411_ = ys__n23060 & new_n13442_;
  assign new_n22412_ = ~new_n22410_ & ~new_n22411_;
  assign new_n22413_ = ~new_n13440_ & ~new_n22412_;
  assign new_n22414_ = ys__n22987 & new_n13440_;
  assign ys__n22988 = new_n22413_ | new_n22414_;
  assign new_n22416_ = ys__n23101 & ~new_n13442_;
  assign new_n22417_ = new_n13439_ & new_n22416_;
  assign new_n22418_ = ys__n23062 & new_n13442_;
  assign new_n22419_ = ~new_n22417_ & ~new_n22418_;
  assign new_n22420_ = ~new_n13440_ & ~new_n22419_;
  assign new_n22421_ = ys__n22990 & new_n13440_;
  assign ys__n22991 = new_n22420_ | new_n22421_;
  assign new_n22423_ = ys__n23102 & ~new_n13442_;
  assign new_n22424_ = new_n13439_ & new_n22423_;
  assign new_n22425_ = ys__n23064 & new_n13442_;
  assign new_n22426_ = ~new_n22424_ & ~new_n22425_;
  assign new_n22427_ = ~new_n13440_ & ~new_n22426_;
  assign new_n22428_ = ys__n22993 & new_n13440_;
  assign ys__n22994 = new_n22427_ | new_n22428_;
  assign new_n22430_ = ys__n23103 & ~new_n13442_;
  assign new_n22431_ = new_n13439_ & new_n22430_;
  assign new_n22432_ = ys__n23066 & new_n13442_;
  assign new_n22433_ = ~new_n22431_ & ~new_n22432_;
  assign new_n22434_ = ~new_n13440_ & ~new_n22433_;
  assign new_n22435_ = ys__n22996 & new_n13440_;
  assign ys__n22997 = new_n22434_ | new_n22435_;
  assign new_n22437_ = ys__n23104 & ~new_n13442_;
  assign new_n22438_ = new_n13439_ & new_n22437_;
  assign new_n22439_ = ys__n23068 & new_n13442_;
  assign new_n22440_ = ~new_n22438_ & ~new_n22439_;
  assign new_n22441_ = ~new_n13440_ & ~new_n22440_;
  assign new_n22442_ = ys__n22999 & new_n13440_;
  assign ys__n23000 = new_n22441_ | new_n22442_;
  assign new_n22444_ = ys__n23105 & ~new_n13442_;
  assign new_n22445_ = new_n13439_ & new_n22444_;
  assign new_n22446_ = ys__n23070 & new_n13442_;
  assign new_n22447_ = ~new_n22445_ & ~new_n22446_;
  assign new_n22448_ = ~new_n13440_ & ~new_n22447_;
  assign new_n22449_ = ys__n23002 & new_n13440_;
  assign ys__n23003 = new_n22448_ | new_n22449_;
  assign new_n22451_ = ys__n23106 & ~new_n13442_;
  assign new_n22452_ = new_n13439_ & new_n22451_;
  assign new_n22453_ = ys__n23072 & new_n13442_;
  assign new_n22454_ = ~new_n22452_ & ~new_n22453_;
  assign new_n22455_ = ~new_n13440_ & ~new_n22454_;
  assign new_n22456_ = ys__n23005 & new_n13440_;
  assign ys__n23006 = new_n22455_ | new_n22456_;
  assign new_n22458_ = ys__n23107 & ~new_n13442_;
  assign new_n22459_ = new_n13439_ & new_n22458_;
  assign new_n22460_ = ys__n23074 & new_n13442_;
  assign new_n22461_ = ~new_n22459_ & ~new_n22460_;
  assign new_n22462_ = ~new_n13440_ & ~new_n22461_;
  assign new_n22463_ = ys__n23008 & new_n13440_;
  assign ys__n23009 = new_n22462_ | new_n22463_;
  assign new_n22465_ = ys__n23108 & ~new_n13442_;
  assign new_n22466_ = new_n13439_ & new_n22465_;
  assign new_n22467_ = ys__n23076 & new_n13442_;
  assign new_n22468_ = ~new_n22466_ & ~new_n22467_;
  assign new_n22469_ = ~new_n13440_ & ~new_n22468_;
  assign new_n22470_ = ys__n23011 & new_n13440_;
  assign ys__n23012 = new_n22469_ | new_n22470_;
  assign new_n22472_ = ys__n18240 & ~ys__n18241;
  assign new_n22473_ = ys__n100 & ys__n18241;
  assign new_n22474_ = ~new_n22472_ & ~new_n22473_;
  assign new_n22475_ = ys__n874 & ~new_n22474_;
  assign new_n22476_ = ys__n18243 & ~ys__n18241;
  assign new_n22477_ = ys__n96 & ys__n18241;
  assign new_n22478_ = ~new_n22476_ & ~new_n22477_;
  assign new_n22479_ = ys__n874 & ~new_n22478_;
  assign new_n22480_ = new_n22475_ & ~new_n22479_;
  assign new_n22481_ = ys__n18223 & new_n22475_;
  assign new_n22482_ = new_n22479_ & new_n22481_;
  assign ys__n23263 = new_n22480_ | new_n22482_;
  assign new_n22484_ = ~ys__n18223 & ~new_n22479_;
  assign new_n22485_ = ys__n18223 & new_n22479_;
  assign ys__n23264 = new_n22484_ | new_n22485_;
  assign new_n22487_ = ~ys__n22464 & ys__n23339;
  assign new_n22488_ = ys__n22464 & ~ys__n23339;
  assign ys__n23483 = new_n22487_ | new_n22488_;
  assign new_n22490_ = new_n12410_ & new_n12411_;
  assign new_n22491_ = ~new_n12410_ & ~new_n12411_;
  assign ys__n23485 = new_n22490_ | new_n22491_;
  assign new_n22493_ = ~new_n12410_ & new_n12411_;
  assign new_n22494_ = ~new_n12406_ & ~new_n22493_;
  assign new_n22495_ = ~ys__n23550 & ~new_n22494_;
  assign new_n22496_ = ys__n23550 & new_n22494_;
  assign ys__n23487 = new_n22495_ | new_n22496_;
  assign new_n22498_ = ~ys__n23552 & ~new_n12414_;
  assign new_n22499_ = ys__n23552 & new_n12414_;
  assign ys__n23489 = new_n22498_ | new_n22499_;
  assign new_n22501_ = ys__n23552 & ~new_n12414_;
  assign new_n22502_ = ~ys__n23554 & new_n22501_;
  assign new_n22503_ = ys__n23554 & ~new_n22501_;
  assign ys__n23491 = new_n22502_ | new_n22503_;
  assign new_n22505_ = ~new_n12414_ & new_n12415_;
  assign new_n22506_ = ~ys__n23556 & new_n22505_;
  assign new_n22507_ = ys__n23556 & ~new_n22505_;
  assign ys__n23493 = new_n22506_ | new_n22507_;
  assign new_n22509_ = ys__n23556 & new_n22505_;
  assign new_n22510_ = ~ys__n23558 & new_n22509_;
  assign new_n22511_ = ys__n23558 & ~new_n22509_;
  assign ys__n23495 = new_n22510_ | new_n22511_;
  assign new_n22513_ = ~ys__n23560 & new_n12418_;
  assign new_n22514_ = ys__n23560 & ~new_n12418_;
  assign ys__n23497 = new_n22513_ | new_n22514_;
  assign new_n22516_ = ys__n23560 & new_n12418_;
  assign new_n22517_ = ~ys__n23562 & new_n22516_;
  assign new_n22518_ = ys__n23562 & ~new_n22516_;
  assign ys__n23499 = new_n22517_ | new_n22518_;
  assign new_n22520_ = new_n12418_ & new_n12419_;
  assign new_n22521_ = ~ys__n23564 & new_n22520_;
  assign new_n22522_ = ys__n23564 & ~new_n22520_;
  assign ys__n23501 = new_n22521_ | new_n22522_;
  assign new_n22524_ = ys__n23564 & new_n22520_;
  assign new_n22525_ = ~ys__n23566 & new_n22524_;
  assign new_n22526_ = ys__n23566 & ~new_n22524_;
  assign ys__n23503 = new_n22525_ | new_n22526_;
  assign new_n22528_ = new_n12418_ & new_n12421_;
  assign new_n22529_ = ~ys__n23568 & new_n22528_;
  assign new_n22530_ = ys__n23568 & ~new_n22528_;
  assign ys__n23505 = new_n22529_ | new_n22530_;
  assign new_n22532_ = ys__n23568 & new_n22528_;
  assign new_n22533_ = ~ys__n23570 & new_n22532_;
  assign new_n22534_ = ys__n23570 & ~new_n22532_;
  assign ys__n23507 = new_n22533_ | new_n22534_;
  assign new_n22536_ = new_n12422_ & new_n22528_;
  assign new_n22537_ = ~ys__n23572 & new_n22536_;
  assign new_n22538_ = ys__n23572 & ~new_n22536_;
  assign ys__n23509 = new_n22537_ | new_n22538_;
  assign new_n22540_ = ys__n23572 & new_n22536_;
  assign new_n22541_ = ~ys__n23574 & new_n22540_;
  assign new_n22542_ = ys__n23574 & ~new_n22540_;
  assign ys__n23511 = new_n22541_ | new_n22542_;
  assign new_n22544_ = ys__n420 & ~new_n12426_;
  assign new_n22545_ = ~ys__n420 & new_n12426_;
  assign ys__n23513 = new_n22544_ | new_n22545_;
  assign new_n22547_ = ys__n442 & ~new_n12426_;
  assign new_n22548_ = ys__n420 & ~ys__n442;
  assign new_n22549_ = ~ys__n420 & ys__n442;
  assign new_n22550_ = ~new_n22548_ & ~new_n22549_;
  assign new_n22551_ = new_n12426_ & ~new_n22550_;
  assign ys__n23515 = new_n22547_ | new_n22551_;
  assign new_n22553_ = ys__n440 & ~new_n12426_;
  assign new_n22554_ = ~ys__n440 & new_n12428_;
  assign new_n22555_ = ys__n440 & ~new_n12428_;
  assign new_n22556_ = ~new_n22554_ & ~new_n22555_;
  assign new_n22557_ = new_n12426_ & ~new_n22556_;
  assign ys__n23517 = new_n22553_ | new_n22557_;
  assign new_n22559_ = ys__n444 & ~new_n12426_;
  assign new_n22560_ = ys__n440 & new_n12428_;
  assign new_n22561_ = ~ys__n444 & new_n22560_;
  assign new_n22562_ = ys__n444 & ~new_n22560_;
  assign new_n22563_ = ~new_n22561_ & ~new_n22562_;
  assign new_n22564_ = new_n12426_ & ~new_n22563_;
  assign ys__n23519 = new_n22559_ | new_n22564_;
  assign new_n22566_ = ys__n438 & ~new_n12426_;
  assign new_n22567_ = ~ys__n438 & new_n12430_;
  assign new_n22568_ = ys__n438 & ~new_n12430_;
  assign new_n22569_ = ~new_n22567_ & ~new_n22568_;
  assign new_n22570_ = new_n12426_ & ~new_n22569_;
  assign ys__n23521 = new_n22566_ | new_n22570_;
  assign new_n22572_ = ys__n446 & ~new_n12426_;
  assign new_n22573_ = ys__n438 & new_n12430_;
  assign new_n22574_ = ~ys__n446 & new_n22573_;
  assign new_n22575_ = ys__n446 & ~new_n22573_;
  assign new_n22576_ = ~new_n22574_ & ~new_n22575_;
  assign new_n22577_ = new_n12426_ & ~new_n22576_;
  assign ys__n23523 = new_n22572_ | new_n22577_;
  assign new_n22579_ = ys__n434 & ~new_n12426_;
  assign new_n22580_ = new_n12430_ & new_n12431_;
  assign new_n22581_ = ~ys__n434 & new_n22580_;
  assign new_n22582_ = ys__n434 & ~new_n22580_;
  assign new_n22583_ = ~new_n22581_ & ~new_n22582_;
  assign new_n22584_ = new_n12426_ & ~new_n22583_;
  assign ys__n23525 = new_n22579_ | new_n22584_;
  assign new_n22586_ = ys__n436 & ~new_n12426_;
  assign new_n22587_ = ys__n434 & new_n22580_;
  assign new_n22588_ = ~ys__n436 & new_n22587_;
  assign new_n22589_ = ys__n436 & ~new_n22587_;
  assign new_n22590_ = ~new_n22588_ & ~new_n22589_;
  assign new_n22591_ = new_n12426_ & ~new_n22590_;
  assign ys__n23527 = new_n22586_ | new_n22591_;
  assign new_n22593_ = ys__n432 & ~new_n12426_;
  assign new_n22594_ = ~ys__n432 & new_n12434_;
  assign new_n22595_ = ys__n432 & ~new_n12434_;
  assign new_n22596_ = ~new_n22594_ & ~new_n22595_;
  assign new_n22597_ = new_n12426_ & ~new_n22596_;
  assign ys__n23529 = new_n22593_ | new_n22597_;
  assign new_n22599_ = ys__n448 & ~new_n12426_;
  assign new_n22600_ = ys__n432 & new_n12434_;
  assign new_n22601_ = ~ys__n448 & new_n22600_;
  assign new_n22602_ = ys__n448 & ~new_n22600_;
  assign new_n22603_ = ~new_n22601_ & ~new_n22602_;
  assign new_n22604_ = new_n12426_ & ~new_n22603_;
  assign ys__n23531 = new_n22599_ | new_n22604_;
  assign new_n22606_ = ys__n428 & ~new_n12426_;
  assign new_n22607_ = new_n12434_ & new_n12435_;
  assign new_n22608_ = ~ys__n428 & new_n22607_;
  assign new_n22609_ = ys__n428 & ~new_n22607_;
  assign new_n22610_ = ~new_n22608_ & ~new_n22609_;
  assign new_n22611_ = new_n12426_ & ~new_n22610_;
  assign ys__n23533 = new_n22606_ | new_n22611_;
  assign new_n22613_ = ys__n430 & ~new_n12426_;
  assign new_n22614_ = ys__n428 & new_n22607_;
  assign new_n22615_ = ~ys__n430 & new_n22614_;
  assign new_n22616_ = ys__n430 & ~new_n22614_;
  assign new_n22617_ = ~new_n22615_ & ~new_n22616_;
  assign new_n22618_ = new_n12426_ & ~new_n22617_;
  assign ys__n23535 = new_n22613_ | new_n22618_;
  assign new_n22620_ = ys__n426 & ~new_n12426_;
  assign new_n22621_ = ~ys__n426 & new_n12438_;
  assign new_n22622_ = ys__n426 & ~new_n12438_;
  assign new_n22623_ = ~new_n22621_ & ~new_n22622_;
  assign new_n22624_ = new_n12426_ & ~new_n22623_;
  assign ys__n23537 = new_n22620_ | new_n22624_;
  assign new_n22626_ = ~ys__n256 & ~ys__n18101;
  assign new_n22627_ = ~ys__n18105 & ~ys__n18106;
  assign new_n22628_ = new_n22626_ & new_n22627_;
  assign new_n22629_ = ~ys__n4566 & new_n22628_;
  assign new_n22630_ = ~new_n11954_ & ~new_n12762_;
  assign new_n22631_ = new_n11954_ & ~new_n12762_;
  assign new_n22632_ = ~new_n12762_ & ~new_n22630_;
  assign new_n22633_ = ~new_n22631_ & new_n22632_;
  assign new_n22634_ = new_n22630_ & ~new_n22633_;
  assign new_n22635_ = ys__n38398 & ~new_n22634_;
  assign new_n22636_ = ~ys__n18111 & ~ys__n18112;
  assign new_n22637_ = ys__n18109 & ~new_n22636_;
  assign new_n22638_ = ~ys__n262 & ~new_n22637_;
  assign new_n22639_ = ~new_n22635_ & ~new_n22638_;
  assign new_n22640_ = ~new_n22635_ & ~new_n22639_;
  assign new_n22641_ = new_n22629_ & ~new_n22640_;
  assign ys__n23635 = ~new_n22629_ | new_n22641_;
  assign new_n22643_ = new_n12314_ & new_n22638_;
  assign new_n22644_ = new_n22629_ & new_n22643_;
  assign new_n22645_ = new_n22631_ & new_n22644_;
  assign new_n22646_ = ~new_n22633_ & new_n22645_;
  assign new_n22647_ = ~new_n22635_ & new_n22646_;
  assign ys__n23636 = ~new_n22629_ | new_n22647_;
  assign new_n22649_ = ~ys__n23840 & ys__n38490;
  assign new_n22650_ = ys__n23840 & ~ys__n38490;
  assign new_n22651_ = ~new_n22649_ & ~new_n22650_;
  assign new_n22652_ = ~ys__n23842 & ys__n38491;
  assign new_n22653_ = ys__n23842 & ~ys__n38491;
  assign new_n22654_ = ~new_n22652_ & ~new_n22653_;
  assign new_n22655_ = new_n22651_ & new_n22654_;
  assign new_n22656_ = ~ys__n23834 & ys__n38487;
  assign new_n22657_ = ys__n23834 & ~ys__n38487;
  assign new_n22658_ = ~new_n22656_ & ~new_n22657_;
  assign new_n22659_ = ~ys__n23836 & ys__n38488;
  assign new_n22660_ = ys__n23836 & ~ys__n38488;
  assign new_n22661_ = ~new_n22659_ & ~new_n22660_;
  assign new_n22662_ = ~ys__n23838 & ys__n38489;
  assign new_n22663_ = ys__n23838 & ~ys__n38489;
  assign new_n22664_ = ~new_n22662_ & ~new_n22663_;
  assign new_n22665_ = new_n22661_ & new_n22664_;
  assign new_n22666_ = new_n22658_ & new_n22665_;
  assign new_n22667_ = new_n22655_ & new_n22666_;
  assign new_n22668_ = ys__n18114 & new_n22667_;
  assign new_n22669_ = ~ys__n296 & ~ys__n2251;
  assign new_n22670_ = ~ys__n2245 & new_n22669_;
  assign new_n22671_ = ~ys__n294 & ~ys__n2247;
  assign new_n22672_ = new_n22670_ & new_n22671_;
  assign new_n22673_ = ys__n23834 & new_n22672_;
  assign new_n22674_ = ~new_n22668_ & new_n22673_;
  assign new_n22675_ = ys__n294 & ~ys__n2247;
  assign new_n22676_ = new_n22670_ & new_n22675_;
  assign new_n22677_ = ys__n296 & ~ys__n2251;
  assign new_n22678_ = ~ys__n2245 & new_n22675_;
  assign new_n22679_ = new_n22677_ & new_n22678_;
  assign new_n22680_ = ~new_n22676_ & ~new_n22679_;
  assign new_n22681_ = ys__n23834 & ~new_n22680_;
  assign new_n22682_ = ys__n29220 & new_n22667_;
  assign new_n22683_ = ~ys__n2245 & new_n22677_;
  assign new_n22684_ = new_n22671_ & new_n22683_;
  assign new_n22685_ = ys__n23834 & new_n22684_;
  assign new_n22686_ = ~new_n22682_ & new_n22685_;
  assign new_n22687_ = ~new_n22681_ & ~new_n22686_;
  assign new_n22688_ = ~new_n22674_ & new_n22687_;
  assign new_n22689_ = ~new_n22672_ & ~new_n22684_;
  assign new_n22690_ = new_n22680_ & new_n22689_;
  assign new_n22691_ = ys__n648 & ~ys__n2239;
  assign new_n22692_ = ~ys__n650 & ~ys__n2233;
  assign new_n22693_ = new_n22691_ & new_n22692_;
  assign new_n22694_ = ys__n644 & ~ys__n646;
  assign new_n22695_ = new_n22693_ & new_n22694_;
  assign new_n22696_ = ~new_n22690_ & new_n22695_;
  assign new_n22697_ = ~new_n22688_ & new_n22696_;
  assign new_n22698_ = ys__n23822 & ~ys__n38491;
  assign new_n22699_ = ys__n23821 & ~ys__n38490;
  assign new_n22700_ = ~ys__n23822 & ys__n38491;
  assign new_n22701_ = ~new_n22699_ & ~new_n22700_;
  assign new_n22702_ = ~new_n22698_ & new_n22701_;
  assign new_n22703_ = ys__n23819 & ~ys__n38488;
  assign new_n22704_ = ~ys__n23820 & ys__n38489;
  assign new_n22705_ = ~new_n22703_ & ~new_n22704_;
  assign new_n22706_ = ys__n23820 & ~ys__n38489;
  assign new_n22707_ = ~ys__n23821 & ys__n38490;
  assign new_n22708_ = ~new_n22706_ & ~new_n22707_;
  assign new_n22709_ = new_n22705_ & new_n22708_;
  assign new_n22710_ = ~ys__n23818 & ys__n38487;
  assign new_n22711_ = ys__n18114 & ~new_n22710_;
  assign new_n22712_ = ys__n23818 & ~ys__n38487;
  assign new_n22713_ = ~ys__n23819 & ys__n38488;
  assign new_n22714_ = ~new_n22712_ & ~new_n22713_;
  assign new_n22715_ = new_n22711_ & new_n22714_;
  assign new_n22716_ = new_n22709_ & new_n22715_;
  assign new_n22717_ = new_n22702_ & new_n22716_;
  assign new_n22718_ = ys__n644 & ys__n646;
  assign new_n22719_ = ys__n650 & ~ys__n2233;
  assign new_n22720_ = new_n22691_ & new_n22719_;
  assign new_n22721_ = new_n22718_ & new_n22720_;
  assign new_n22722_ = ys__n23818 & new_n22721_;
  assign new_n22723_ = ~new_n22717_ & new_n22722_;
  assign new_n22724_ = new_n22693_ & new_n22718_;
  assign new_n22725_ = ys__n23818 & ~new_n22721_;
  assign new_n22726_ = new_n22724_ & new_n22725_;
  assign new_n22727_ = ~new_n22723_ & ~new_n22726_;
  assign new_n22728_ = ~new_n22695_ & ~new_n22727_;
  assign ys__n23795 = new_n22697_ | new_n22728_;
  assign new_n22730_ = ys__n23836 & new_n22672_;
  assign new_n22731_ = ~new_n22668_ & new_n22730_;
  assign new_n22732_ = ys__n23836 & ~new_n22680_;
  assign new_n22733_ = ys__n23836 & new_n22684_;
  assign new_n22734_ = ~new_n22682_ & new_n22733_;
  assign new_n22735_ = ~new_n22732_ & ~new_n22734_;
  assign new_n22736_ = ~new_n22731_ & new_n22735_;
  assign new_n22737_ = new_n22696_ & ~new_n22736_;
  assign new_n22738_ = ys__n23819 & new_n22721_;
  assign new_n22739_ = ~new_n22717_ & new_n22738_;
  assign new_n22740_ = ys__n23819 & ~new_n22721_;
  assign new_n22741_ = new_n22724_ & new_n22740_;
  assign new_n22742_ = ~new_n22739_ & ~new_n22741_;
  assign new_n22743_ = ~new_n22695_ & ~new_n22742_;
  assign ys__n23798 = new_n22737_ | new_n22743_;
  assign new_n22745_ = ys__n23838 & new_n22672_;
  assign new_n22746_ = ~new_n22668_ & new_n22745_;
  assign new_n22747_ = ys__n23838 & ~new_n22680_;
  assign new_n22748_ = ys__n23838 & new_n22684_;
  assign new_n22749_ = ~new_n22682_ & new_n22748_;
  assign new_n22750_ = ~new_n22747_ & ~new_n22749_;
  assign new_n22751_ = ~new_n22746_ & new_n22750_;
  assign new_n22752_ = new_n22696_ & ~new_n22751_;
  assign new_n22753_ = ys__n23820 & new_n22721_;
  assign new_n22754_ = ~new_n22717_ & new_n22753_;
  assign new_n22755_ = ys__n23820 & ~new_n22721_;
  assign new_n22756_ = new_n22724_ & new_n22755_;
  assign new_n22757_ = ~new_n22754_ & ~new_n22756_;
  assign new_n22758_ = ~new_n22695_ & ~new_n22757_;
  assign ys__n23801 = new_n22752_ | new_n22758_;
  assign new_n22760_ = ys__n23840 & new_n22672_;
  assign new_n22761_ = ~new_n22668_ & new_n22760_;
  assign new_n22762_ = ys__n23840 & ~new_n22680_;
  assign new_n22763_ = ys__n23840 & new_n22684_;
  assign new_n22764_ = ~new_n22682_ & new_n22763_;
  assign new_n22765_ = ~new_n22762_ & ~new_n22764_;
  assign new_n22766_ = ~new_n22761_ & new_n22765_;
  assign new_n22767_ = new_n22696_ & ~new_n22766_;
  assign new_n22768_ = ys__n23821 & new_n22721_;
  assign new_n22769_ = ~new_n22717_ & new_n22768_;
  assign new_n22770_ = ys__n23821 & ~new_n22721_;
  assign new_n22771_ = new_n22724_ & new_n22770_;
  assign new_n22772_ = ~new_n22769_ & ~new_n22771_;
  assign new_n22773_ = ~new_n22695_ & ~new_n22772_;
  assign ys__n23804 = new_n22767_ | new_n22773_;
  assign new_n22775_ = ys__n23842 & new_n22672_;
  assign new_n22776_ = ~new_n22668_ & new_n22775_;
  assign new_n22777_ = ys__n23842 & ~new_n22680_;
  assign new_n22778_ = ys__n23842 & new_n22684_;
  assign new_n22779_ = ~new_n22682_ & new_n22778_;
  assign new_n22780_ = ~new_n22777_ & ~new_n22779_;
  assign new_n22781_ = ~new_n22776_ & new_n22780_;
  assign new_n22782_ = new_n22696_ & ~new_n22781_;
  assign new_n22783_ = ys__n23822 & new_n22721_;
  assign new_n22784_ = ~new_n22717_ & new_n22783_;
  assign new_n22785_ = ys__n23822 & ~new_n22721_;
  assign new_n22786_ = new_n22724_ & new_n22785_;
  assign new_n22787_ = ~new_n22784_ & ~new_n22786_;
  assign new_n22788_ = ~new_n22695_ & ~new_n22787_;
  assign ys__n23807 = new_n22782_ | new_n22788_;
  assign new_n22790_ = ~ys__n740 & new_n13284_;
  assign new_n22791_ = ~new_n13564_ & ~new_n22790_;
  assign new_n22792_ = ~new_n13291_ & ~new_n22791_;
  assign new_n22793_ = ~new_n13291_ & ~new_n22792_;
  assign new_n22794_ = ~new_n13280_ & ~new_n22793_;
  assign ys__n23853 = new_n13280_ | new_n22794_;
  assign new_n22796_ = ~ys__n23910 & ys__n38498;
  assign new_n22797_ = ys__n23910 & ~ys__n38498;
  assign new_n22798_ = ~new_n22796_ & ~new_n22797_;
  assign new_n22799_ = ~ys__n23912 & ys__n38499;
  assign new_n22800_ = ys__n23912 & ~ys__n38499;
  assign new_n22801_ = ~new_n22799_ & ~new_n22800_;
  assign new_n22802_ = new_n22798_ & new_n22801_;
  assign new_n22803_ = ~ys__n23904 & ys__n38495;
  assign new_n22804_ = ys__n23904 & ~ys__n38495;
  assign new_n22805_ = ~new_n22803_ & ~new_n22804_;
  assign new_n22806_ = ~ys__n23906 & ys__n38496;
  assign new_n22807_ = ys__n23906 & ~ys__n38496;
  assign new_n22808_ = ~new_n22806_ & ~new_n22807_;
  assign new_n22809_ = ~ys__n23908 & ys__n38497;
  assign new_n22810_ = ys__n23908 & ~ys__n38497;
  assign new_n22811_ = ~new_n22809_ & ~new_n22810_;
  assign new_n22812_ = new_n22808_ & new_n22811_;
  assign new_n22813_ = new_n22805_ & new_n22812_;
  assign new_n22814_ = new_n22802_ & new_n22813_;
  assign new_n22815_ = ys__n18116 & new_n22814_;
  assign new_n22816_ = ~ys__n586 & ~ys__n2312;
  assign new_n22817_ = ~ys__n2306 & new_n22816_;
  assign new_n22818_ = ~ys__n588 & ~ys__n2308;
  assign new_n22819_ = new_n22817_ & new_n22818_;
  assign new_n22820_ = ys__n23904 & new_n22819_;
  assign new_n22821_ = ~new_n22815_ & new_n22820_;
  assign new_n22822_ = ys__n588 & ~ys__n2308;
  assign new_n22823_ = new_n22817_ & new_n22822_;
  assign new_n22824_ = ys__n586 & ~ys__n2312;
  assign new_n22825_ = ~ys__n2306 & new_n22822_;
  assign new_n22826_ = new_n22824_ & new_n22825_;
  assign new_n22827_ = ~new_n22823_ & ~new_n22826_;
  assign new_n22828_ = ys__n23904 & ~new_n22827_;
  assign new_n22829_ = ys__n29533 & new_n22814_;
  assign new_n22830_ = ~ys__n2306 & new_n22824_;
  assign new_n22831_ = new_n22818_ & new_n22830_;
  assign new_n22832_ = ys__n23904 & new_n22831_;
  assign new_n22833_ = ~new_n22829_ & new_n22832_;
  assign new_n22834_ = ~new_n22828_ & ~new_n22833_;
  assign new_n22835_ = ~new_n22821_ & new_n22834_;
  assign new_n22836_ = ~new_n22819_ & ~new_n22831_;
  assign new_n22837_ = new_n22827_ & new_n22836_;
  assign new_n22838_ = ys__n656 & ~ys__n2282;
  assign new_n22839_ = ~ys__n658 & ~ys__n2276;
  assign new_n22840_ = new_n22838_ & new_n22839_;
  assign new_n22841_ = ys__n652 & ~ys__n654;
  assign new_n22842_ = new_n22840_ & new_n22841_;
  assign new_n22843_ = ~new_n22837_ & new_n22842_;
  assign new_n22844_ = ~new_n22835_ & new_n22843_;
  assign new_n22845_ = ys__n23892 & ~ys__n38499;
  assign new_n22846_ = ys__n23891 & ~ys__n38498;
  assign new_n22847_ = ~ys__n23892 & ys__n38499;
  assign new_n22848_ = ~new_n22846_ & ~new_n22847_;
  assign new_n22849_ = ~new_n22845_ & new_n22848_;
  assign new_n22850_ = ys__n23889 & ~ys__n38496;
  assign new_n22851_ = ~ys__n23890 & ys__n38497;
  assign new_n22852_ = ~new_n22850_ & ~new_n22851_;
  assign new_n22853_ = ys__n23890 & ~ys__n38497;
  assign new_n22854_ = ~ys__n23891 & ys__n38498;
  assign new_n22855_ = ~new_n22853_ & ~new_n22854_;
  assign new_n22856_ = new_n22852_ & new_n22855_;
  assign new_n22857_ = ~ys__n23888 & ys__n38495;
  assign new_n22858_ = ys__n18116 & ~new_n22857_;
  assign new_n22859_ = ys__n23888 & ~ys__n38495;
  assign new_n22860_ = ~ys__n23889 & ys__n38496;
  assign new_n22861_ = ~new_n22859_ & ~new_n22860_;
  assign new_n22862_ = new_n22858_ & new_n22861_;
  assign new_n22863_ = new_n22856_ & new_n22862_;
  assign new_n22864_ = new_n22849_ & new_n22863_;
  assign new_n22865_ = ys__n652 & ys__n654;
  assign new_n22866_ = ys__n658 & ~ys__n2276;
  assign new_n22867_ = new_n22838_ & new_n22866_;
  assign new_n22868_ = new_n22865_ & new_n22867_;
  assign new_n22869_ = ys__n23888 & new_n22868_;
  assign new_n22870_ = ~new_n22864_ & new_n22869_;
  assign new_n22871_ = new_n22840_ & new_n22865_;
  assign new_n22872_ = ys__n23888 & ~new_n22868_;
  assign new_n22873_ = new_n22871_ & new_n22872_;
  assign new_n22874_ = ~new_n22870_ & ~new_n22873_;
  assign new_n22875_ = ~new_n22842_ & ~new_n22874_;
  assign ys__n23865 = new_n22844_ | new_n22875_;
  assign new_n22877_ = ys__n23906 & new_n22819_;
  assign new_n22878_ = ~new_n22815_ & new_n22877_;
  assign new_n22879_ = ys__n23906 & ~new_n22827_;
  assign new_n22880_ = ys__n23906 & new_n22831_;
  assign new_n22881_ = ~new_n22829_ & new_n22880_;
  assign new_n22882_ = ~new_n22879_ & ~new_n22881_;
  assign new_n22883_ = ~new_n22878_ & new_n22882_;
  assign new_n22884_ = new_n22843_ & ~new_n22883_;
  assign new_n22885_ = ys__n23889 & new_n22868_;
  assign new_n22886_ = ~new_n22864_ & new_n22885_;
  assign new_n22887_ = ys__n23889 & ~new_n22868_;
  assign new_n22888_ = new_n22871_ & new_n22887_;
  assign new_n22889_ = ~new_n22886_ & ~new_n22888_;
  assign new_n22890_ = ~new_n22842_ & ~new_n22889_;
  assign ys__n23868 = new_n22884_ | new_n22890_;
  assign new_n22892_ = ys__n23908 & new_n22819_;
  assign new_n22893_ = ~new_n22815_ & new_n22892_;
  assign new_n22894_ = ys__n23908 & ~new_n22827_;
  assign new_n22895_ = ys__n23908 & new_n22831_;
  assign new_n22896_ = ~new_n22829_ & new_n22895_;
  assign new_n22897_ = ~new_n22894_ & ~new_n22896_;
  assign new_n22898_ = ~new_n22893_ & new_n22897_;
  assign new_n22899_ = new_n22843_ & ~new_n22898_;
  assign new_n22900_ = ys__n23890 & new_n22868_;
  assign new_n22901_ = ~new_n22864_ & new_n22900_;
  assign new_n22902_ = ys__n23890 & ~new_n22868_;
  assign new_n22903_ = new_n22871_ & new_n22902_;
  assign new_n22904_ = ~new_n22901_ & ~new_n22903_;
  assign new_n22905_ = ~new_n22842_ & ~new_n22904_;
  assign ys__n23871 = new_n22899_ | new_n22905_;
  assign new_n22907_ = ys__n23910 & new_n22819_;
  assign new_n22908_ = ~new_n22815_ & new_n22907_;
  assign new_n22909_ = ys__n23910 & ~new_n22827_;
  assign new_n22910_ = ys__n23910 & new_n22831_;
  assign new_n22911_ = ~new_n22829_ & new_n22910_;
  assign new_n22912_ = ~new_n22909_ & ~new_n22911_;
  assign new_n22913_ = ~new_n22908_ & new_n22912_;
  assign new_n22914_ = new_n22843_ & ~new_n22913_;
  assign new_n22915_ = ys__n23891 & new_n22868_;
  assign new_n22916_ = ~new_n22864_ & new_n22915_;
  assign new_n22917_ = ys__n23891 & ~new_n22868_;
  assign new_n22918_ = new_n22871_ & new_n22917_;
  assign new_n22919_ = ~new_n22916_ & ~new_n22918_;
  assign new_n22920_ = ~new_n22842_ & ~new_n22919_;
  assign ys__n23874 = new_n22914_ | new_n22920_;
  assign new_n22922_ = ys__n23912 & new_n22819_;
  assign new_n22923_ = ~new_n22815_ & new_n22922_;
  assign new_n22924_ = ys__n23912 & ~new_n22827_;
  assign new_n22925_ = ys__n23912 & new_n22831_;
  assign new_n22926_ = ~new_n22829_ & new_n22925_;
  assign new_n22927_ = ~new_n22924_ & ~new_n22926_;
  assign new_n22928_ = ~new_n22923_ & new_n22927_;
  assign new_n22929_ = new_n22843_ & ~new_n22928_;
  assign new_n22930_ = ys__n23892 & new_n22868_;
  assign new_n22931_ = ~new_n22864_ & new_n22930_;
  assign new_n22932_ = ys__n23892 & ~new_n22868_;
  assign new_n22933_ = new_n22871_ & new_n22932_;
  assign new_n22934_ = ~new_n22931_ & ~new_n22933_;
  assign new_n22935_ = ~new_n22842_ & ~new_n22934_;
  assign ys__n23877 = new_n22929_ | new_n22935_;
  assign new_n22937_ = ~ys__n740 & new_n13295_;
  assign new_n22938_ = ~new_n13585_ & ~new_n22937_;
  assign new_n22939_ = ~new_n13302_ & ~new_n22938_;
  assign new_n22940_ = ~new_n13302_ & ~new_n22939_;
  assign new_n22941_ = ~new_n13280_ & ~new_n22940_;
  assign ys__n23921 = new_n13280_ | new_n22941_;
  assign new_n22943_ = ~ys__n23983 & ys__n38506;
  assign new_n22944_ = ys__n23983 & ~ys__n38506;
  assign new_n22945_ = ~new_n22943_ & ~new_n22944_;
  assign new_n22946_ = ~ys__n23985 & ys__n38507;
  assign new_n22947_ = ys__n23985 & ~ys__n38507;
  assign new_n22948_ = ~new_n22946_ & ~new_n22947_;
  assign new_n22949_ = new_n22945_ & new_n22948_;
  assign new_n22950_ = ~ys__n23977 & ys__n38503;
  assign new_n22951_ = ys__n23977 & ~ys__n38503;
  assign new_n22952_ = ~new_n22950_ & ~new_n22951_;
  assign new_n22953_ = ~ys__n23979 & ys__n38504;
  assign new_n22954_ = ys__n23979 & ~ys__n38504;
  assign new_n22955_ = ~new_n22953_ & ~new_n22954_;
  assign new_n22956_ = ~ys__n23981 & ys__n38505;
  assign new_n22957_ = ys__n23981 & ~ys__n38505;
  assign new_n22958_ = ~new_n22956_ & ~new_n22957_;
  assign new_n22959_ = new_n22955_ & new_n22958_;
  assign new_n22960_ = new_n22952_ & new_n22959_;
  assign new_n22961_ = new_n22949_ & new_n22960_;
  assign new_n22962_ = ys__n18118 & new_n22961_;
  assign new_n22963_ = ~ys__n194 & ~ys__n2433;
  assign new_n22964_ = ~ys__n2427 & new_n22963_;
  assign new_n22965_ = ~ys__n304 & ~ys__n2429;
  assign new_n22966_ = new_n22964_ & new_n22965_;
  assign new_n22967_ = ys__n23977 & new_n22966_;
  assign new_n22968_ = ~new_n22962_ & new_n22967_;
  assign new_n22969_ = ys__n304 & ~ys__n2429;
  assign new_n22970_ = new_n22964_ & new_n22969_;
  assign new_n22971_ = ys__n194 & ~ys__n2433;
  assign new_n22972_ = ~ys__n2427 & new_n22969_;
  assign new_n22973_ = new_n22971_ & new_n22972_;
  assign new_n22974_ = ~new_n22970_ & ~new_n22973_;
  assign new_n22975_ = ys__n23977 & ~new_n22974_;
  assign new_n22976_ = ys__n29808 & new_n22961_;
  assign new_n22977_ = ~ys__n2427 & new_n22971_;
  assign new_n22978_ = new_n22965_ & new_n22977_;
  assign new_n22979_ = ys__n23977 & new_n22978_;
  assign new_n22980_ = ~new_n22976_ & new_n22979_;
  assign new_n22981_ = ~new_n22975_ & ~new_n22980_;
  assign new_n22982_ = ~new_n22968_ & new_n22981_;
  assign new_n22983_ = ~new_n22966_ & ~new_n22978_;
  assign new_n22984_ = new_n22974_ & new_n22983_;
  assign new_n22985_ = ys__n662 & ys__n668;
  assign new_n22986_ = ~ys__n660 & ~ys__n666;
  assign new_n22987_ = new_n22985_ & new_n22986_;
  assign new_n22988_ = ys__n626 & ~ys__n664;
  assign new_n22989_ = new_n22987_ & new_n22988_;
  assign new_n22990_ = ~new_n22984_ & new_n22989_;
  assign new_n22991_ = ~new_n22982_ & new_n22990_;
  assign new_n22992_ = ys__n23960 & ~ys__n38507;
  assign new_n22993_ = ys__n23959 & ~ys__n38506;
  assign new_n22994_ = ~ys__n23960 & ys__n38507;
  assign new_n22995_ = ~new_n22993_ & ~new_n22994_;
  assign new_n22996_ = ~new_n22992_ & new_n22995_;
  assign new_n22997_ = ys__n23957 & ~ys__n38504;
  assign new_n22998_ = ~ys__n23958 & ys__n38505;
  assign new_n22999_ = ~new_n22997_ & ~new_n22998_;
  assign new_n23000_ = ys__n23958 & ~ys__n38505;
  assign new_n23001_ = ~ys__n23959 & ys__n38506;
  assign new_n23002_ = ~new_n23000_ & ~new_n23001_;
  assign new_n23003_ = new_n22999_ & new_n23002_;
  assign new_n23004_ = ~ys__n23956 & ys__n38503;
  assign new_n23005_ = ys__n18118 & ~new_n23004_;
  assign new_n23006_ = ys__n23956 & ~ys__n38503;
  assign new_n23007_ = ~ys__n23957 & ys__n38504;
  assign new_n23008_ = ~new_n23006_ & ~new_n23007_;
  assign new_n23009_ = new_n23005_ & new_n23008_;
  assign new_n23010_ = new_n23003_ & new_n23009_;
  assign new_n23011_ = new_n22996_ & new_n23010_;
  assign new_n23012_ = ys__n626 & ys__n664;
  assign new_n23013_ = ~ys__n660 & ys__n666;
  assign new_n23014_ = new_n22985_ & new_n23013_;
  assign new_n23015_ = new_n23012_ & new_n23014_;
  assign new_n23016_ = ys__n23956 & new_n23015_;
  assign new_n23017_ = ~new_n23011_ & new_n23016_;
  assign new_n23018_ = new_n22987_ & new_n23012_;
  assign new_n23019_ = ys__n23956 & ~new_n23015_;
  assign new_n23020_ = new_n23018_ & new_n23019_;
  assign new_n23021_ = ~new_n23017_ & ~new_n23020_;
  assign new_n23022_ = ~new_n22989_ & ~new_n23021_;
  assign ys__n23933 = new_n22991_ | new_n23022_;
  assign new_n23024_ = ys__n23979 & new_n22966_;
  assign new_n23025_ = ~new_n22962_ & new_n23024_;
  assign new_n23026_ = ys__n23979 & ~new_n22974_;
  assign new_n23027_ = ys__n23979 & new_n22978_;
  assign new_n23028_ = ~new_n22976_ & new_n23027_;
  assign new_n23029_ = ~new_n23026_ & ~new_n23028_;
  assign new_n23030_ = ~new_n23025_ & new_n23029_;
  assign new_n23031_ = new_n22990_ & ~new_n23030_;
  assign new_n23032_ = ys__n23957 & new_n23015_;
  assign new_n23033_ = ~new_n23011_ & new_n23032_;
  assign new_n23034_ = ys__n23957 & ~new_n23015_;
  assign new_n23035_ = new_n23018_ & new_n23034_;
  assign new_n23036_ = ~new_n23033_ & ~new_n23035_;
  assign new_n23037_ = ~new_n22989_ & ~new_n23036_;
  assign ys__n23936 = new_n23031_ | new_n23037_;
  assign new_n23039_ = ys__n23981 & new_n22966_;
  assign new_n23040_ = ~new_n22962_ & new_n23039_;
  assign new_n23041_ = ys__n23981 & ~new_n22974_;
  assign new_n23042_ = ys__n23981 & new_n22978_;
  assign new_n23043_ = ~new_n22976_ & new_n23042_;
  assign new_n23044_ = ~new_n23041_ & ~new_n23043_;
  assign new_n23045_ = ~new_n23040_ & new_n23044_;
  assign new_n23046_ = new_n22990_ & ~new_n23045_;
  assign new_n23047_ = ys__n23958 & new_n23015_;
  assign new_n23048_ = ~new_n23011_ & new_n23047_;
  assign new_n23049_ = ys__n23958 & ~new_n23015_;
  assign new_n23050_ = new_n23018_ & new_n23049_;
  assign new_n23051_ = ~new_n23048_ & ~new_n23050_;
  assign new_n23052_ = ~new_n22989_ & ~new_n23051_;
  assign ys__n23939 = new_n23046_ | new_n23052_;
  assign new_n23054_ = ys__n23983 & new_n22966_;
  assign new_n23055_ = ~new_n22962_ & new_n23054_;
  assign new_n23056_ = ys__n23983 & ~new_n22974_;
  assign new_n23057_ = ys__n23983 & new_n22978_;
  assign new_n23058_ = ~new_n22976_ & new_n23057_;
  assign new_n23059_ = ~new_n23056_ & ~new_n23058_;
  assign new_n23060_ = ~new_n23055_ & new_n23059_;
  assign new_n23061_ = new_n22990_ & ~new_n23060_;
  assign new_n23062_ = ys__n23959 & new_n23015_;
  assign new_n23063_ = ~new_n23011_ & new_n23062_;
  assign new_n23064_ = ys__n23959 & ~new_n23015_;
  assign new_n23065_ = new_n23018_ & new_n23064_;
  assign new_n23066_ = ~new_n23063_ & ~new_n23065_;
  assign new_n23067_ = ~new_n22989_ & ~new_n23066_;
  assign ys__n23942 = new_n23061_ | new_n23067_;
  assign new_n23069_ = ys__n23985 & new_n22966_;
  assign new_n23070_ = ~new_n22962_ & new_n23069_;
  assign new_n23071_ = ys__n23985 & ~new_n22974_;
  assign new_n23072_ = ys__n23985 & new_n22978_;
  assign new_n23073_ = ~new_n22976_ & new_n23072_;
  assign new_n23074_ = ~new_n23071_ & ~new_n23073_;
  assign new_n23075_ = ~new_n23070_ & new_n23074_;
  assign new_n23076_ = new_n22990_ & ~new_n23075_;
  assign new_n23077_ = ys__n23960 & new_n23015_;
  assign new_n23078_ = ~new_n23011_ & new_n23077_;
  assign new_n23079_ = ys__n23960 & ~new_n23015_;
  assign new_n23080_ = new_n23018_ & new_n23079_;
  assign new_n23081_ = ~new_n23078_ & ~new_n23080_;
  assign new_n23082_ = ~new_n22989_ & ~new_n23081_;
  assign ys__n23945 = new_n23076_ | new_n23082_;
  assign new_n23084_ = ~ys__n740 & new_n13328_;
  assign new_n23085_ = ~new_n13593_ & ~new_n23084_;
  assign new_n23086_ = ~new_n13335_ & ~new_n23085_;
  assign new_n23087_ = ~new_n13335_ & ~new_n23086_;
  assign new_n23088_ = ~new_n13280_ & ~new_n23087_;
  assign ys__n24099 = new_n13280_ | new_n23088_;
  assign ys__n24101 = ys__n24106 & ~ys__n24107;
  assign new_n23091_ = ~ys__n416 & ~ys__n38526;
  assign new_n23092_ = ys__n416 & ys__n38526;
  assign new_n23093_ = ~new_n23091_ & ~new_n23092_;
  assign new_n23094_ = ~ys__n24112 & ~new_n23093_;
  assign new_n23095_ = ~ys__n418 & ys__n24112;
  assign new_n23096_ = ~new_n23094_ & ~new_n23095_;
  assign new_n23097_ = ~ys__n1029 & ys__n1030;
  assign new_n23098_ = ~new_n23096_ & new_n23097_;
  assign new_n23099_ = ys__n1029 & ys__n24101;
  assign ys__n24102 = new_n23098_ | new_n23099_;
  assign ys__n24104 = ~ys__n24107 & ys__n24108;
  assign new_n23102_ = ys__n416 & ~ys__n686;
  assign new_n23103_ = ~ys__n416 & ys__n686;
  assign ys__n35705 = new_n23102_ | new_n23103_;
  assign new_n23105_ = ~ys__n38527 & ys__n35705;
  assign new_n23106_ = ys__n38527 & ~ys__n35705;
  assign new_n23107_ = ~new_n23105_ & ~new_n23106_;
  assign new_n23108_ = ~ys__n24112 & ~new_n23107_;
  assign new_n23109_ = ys__n418 & ~ys__n35704;
  assign new_n23110_ = ~ys__n418 & ys__n35704;
  assign new_n23111_ = ~new_n23109_ & ~new_n23110_;
  assign new_n23112_ = ys__n24112 & ~new_n23111_;
  assign new_n23113_ = ~new_n23108_ & ~new_n23112_;
  assign new_n23114_ = new_n23097_ & ~new_n23113_;
  assign new_n23115_ = ys__n1029 & ys__n24104;
  assign ys__n24105 = new_n23114_ | new_n23115_;
  assign new_n23117_ = ys__n47663 & new_n12768_;
  assign new_n23118_ = ys__n22826 & ~new_n12314_;
  assign new_n23119_ = new_n12309_ & new_n23118_;
  assign new_n23120_ = ~new_n17417_ & ~new_n23119_;
  assign new_n23121_ = ~new_n12320_ & ~new_n23120_;
  assign new_n23122_ = ys__n23548 & new_n12320_;
  assign new_n23123_ = ~new_n23121_ & ~new_n23122_;
  assign new_n23124_ = ~new_n12404_ & ~new_n23123_;
  assign new_n23125_ = new_n12404_ & ys__n23485;
  assign new_n23126_ = ~new_n23124_ & ~new_n23125_;
  assign new_n23127_ = new_n12458_ & ~new_n23126_;
  assign new_n23128_ = ys__n528 & ~new_n12458_;
  assign new_n23129_ = ~new_n23127_ & ~new_n23128_;
  assign new_n23130_ = ~new_n12477_ & ~new_n23129_;
  assign new_n23131_ = new_n12506_ & new_n12524_;
  assign new_n23132_ = ~new_n12506_ & ~new_n12524_;
  assign new_n23133_ = ~new_n23131_ & ~new_n23132_;
  assign new_n23134_ = new_n12477_ & ~new_n23133_;
  assign new_n23135_ = ~new_n23130_ & ~new_n23134_;
  assign new_n23136_ = new_n12763_ & ~new_n23135_;
  assign new_n23137_ = ~new_n23117_ & ~new_n23136_;
  assign new_n23138_ = new_n12774_ & ~new_n23137_;
  assign new_n23139_ = ys__n47663 & new_n12778_;
  assign new_n23140_ = new_n12776_ & ~new_n23135_;
  assign new_n23141_ = ~new_n23139_ & ~new_n23140_;
  assign new_n23142_ = new_n12784_ & ~new_n23141_;
  assign ys__n24116 = new_n23138_ | new_n23142_;
  assign new_n23144_ = ~ys__n18121 & ys__n24106;
  assign new_n23145_ = ys__n418 & ys__n18121;
  assign new_n23146_ = ~new_n23144_ & ~new_n23145_;
  assign new_n23147_ = new_n12175_ & new_n17031_;
  assign new_n23148_ = new_n13361_ & new_n23147_;
  assign new_n23149_ = ys__n1029 & new_n23148_;
  assign new_n23150_ = ~new_n23146_ & ~new_n23149_;
  assign new_n23151_ = ys__n24116 & new_n23149_;
  assign ys__n24118 = new_n23150_ | new_n23151_;
  assign new_n23153_ = ys__n1036 & ~ys__n1048;
  assign new_n23154_ = ~ys__n24123 & ys__n24124;
  assign new_n23155_ = new_n23153_ & new_n23154_;
  assign new_n23156_ = ys__n1048 & ~ys__n18007;
  assign new_n23157_ = ~new_n23155_ & ~new_n23156_;
  assign new_n23158_ = ~ys__n140 & ~new_n23157_;
  assign ys__n24120 = ys__n140 | new_n23158_;
  assign new_n23160_ = ~ys__n1036 & ~ys__n24123;
  assign new_n23161_ = ys__n24124 & new_n23160_;
  assign ys__n24126 = ys__n24123 | new_n23161_;
  assign new_n23163_ = ys__n1029 & ~ys__n1036;
  assign new_n23164_ = ys__n24131 & new_n23163_;
  assign new_n23165_ = ys__n1036 & ~ys__n24123;
  assign ys__n24130 = new_n23164_ | new_n23165_;
  assign new_n23167_ = ~ys__n18121 & ys__n18122;
  assign new_n23168_ = ~ys__n18124 & new_n23167_;
  assign new_n23169_ = new_n13573_ & new_n23168_;
  assign new_n23170_ = ys__n678 & ys__n680;
  assign new_n23171_ = ys__n682 & ys__n684;
  assign new_n23172_ = new_n23170_ & new_n23171_;
  assign new_n23173_ = ys__n670 & ys__n672;
  assign new_n23174_ = ys__n674 & ys__n676;
  assign new_n23175_ = new_n23173_ & new_n23174_;
  assign new_n23176_ = new_n23172_ & new_n23175_;
  assign new_n23177_ = ~ys__n38524 & ~new_n23176_;
  assign new_n23178_ = ~ys__n33423 & new_n11734_;
  assign new_n23179_ = new_n23148_ & new_n23178_;
  assign new_n23180_ = ~new_n23177_ & new_n23179_;
  assign new_n23181_ = ~ys__n18120 & new_n23180_;
  assign new_n23182_ = ~new_n11731_ & new_n23181_;
  assign ys__n24134 = new_n23169_ | new_n23182_;
  assign new_n23184_ = ~ys__n18122 & ys__n24143;
  assign new_n23185_ = ~ys__n24158 & new_n23184_;
  assign new_n23186_ = ~new_n11989_ & ~new_n23185_;
  assign new_n23187_ = ~ys__n18121 & ~new_n23186_;
  assign new_n23188_ = ys__n416 & ys__n686;
  assign new_n23189_ = ys__n18124 & new_n23188_;
  assign new_n23190_ = ys__n18121 & new_n23189_;
  assign ys__n24140 = new_n23187_ | new_n23190_;
  assign new_n23192_ = ~ys__n1029 & ys__n1038;
  assign new_n23193_ = ~ys__n18120 & new_n23149_;
  assign new_n23194_ = ~new_n11731_ & new_n23193_;
  assign new_n23195_ = ~ys__n33423 & new_n23194_;
  assign new_n23196_ = ~ys__n18120 & ~new_n23195_;
  assign new_n23197_ = ~ys__n18120 & new_n23148_;
  assign new_n23198_ = ~new_n11731_ & new_n23197_;
  assign new_n23199_ = ~new_n23196_ & new_n23198_;
  assign new_n23200_ = ~ys__n24158 & new_n11734_;
  assign new_n23201_ = ~new_n23199_ & new_n23200_;
  assign new_n23202_ = ~new_n23192_ & ~new_n23201_;
  assign new_n23203_ = ~ys__n1036 & ~new_n23202_;
  assign new_n23204_ = ys__n1036 & ys__n24123;
  assign ys__n24145 = new_n23203_ | new_n23204_;
  assign new_n23206_ = ys__n18121 & new_n13573_;
  assign new_n23207_ = ~new_n23189_ & new_n23206_;
  assign new_n23208_ = new_n23177_ & new_n23179_;
  assign new_n23209_ = ~ys__n18120 & new_n23208_;
  assign new_n23210_ = ~new_n11731_ & new_n23209_;
  assign new_n23211_ = new_n23194_ & new_n23210_;
  assign ys__n24149 = new_n23207_ | new_n23211_;
  assign ys__n38521 = ys__n24143 & ys__n24158;
  assign new_n23214_ = new_n13568_ & new_n13573_;
  assign new_n23215_ = ys__n38521 & new_n23214_;
  assign new_n23216_ = ys__n24158 & new_n11734_;
  assign new_n23217_ = ~new_n23194_ & new_n23216_;
  assign ys__n24154 = new_n23215_ | new_n23217_;
  assign new_n23219_ = ~ys__n30974 & ~ys__n33272;
  assign new_n23220_ = ~ys__n33274 & ~ys__n33276;
  assign new_n23221_ = new_n23219_ & new_n23220_;
  assign new_n23222_ = ~ys__n33278 & ~new_n23221_;
  assign new_n23223_ = ~ys__n33274 & new_n23219_;
  assign new_n23224_ = ~ys__n33276 & ~new_n23223_;
  assign new_n23225_ = ys__n33278 & new_n23221_;
  assign new_n23226_ = ~new_n23224_ & ~new_n23225_;
  assign new_n23227_ = ~new_n23222_ & new_n23226_;
  assign new_n23228_ = ys__n30974 & ~ys__n33272;
  assign new_n23229_ = ~ys__n30974 & ys__n33272;
  assign new_n23230_ = ~ys__n30974 & ~new_n23229_;
  assign new_n23231_ = ~new_n23228_ & new_n23230_;
  assign new_n23232_ = ys__n33274 & new_n23219_;
  assign new_n23233_ = ~ys__n33274 & ~new_n23219_;
  assign new_n23234_ = ~new_n23232_ & ~new_n23233_;
  assign new_n23235_ = new_n23231_ & new_n23234_;
  assign new_n23236_ = ~ys__n33278 & new_n23221_;
  assign new_n23237_ = ys__n33276 & new_n23223_;
  assign new_n23238_ = new_n23236_ & ~new_n23237_;
  assign new_n23239_ = new_n23235_ & new_n23238_;
  assign new_n23240_ = new_n23227_ & new_n23239_;
  assign new_n23241_ = ~ys__n38561 & ~new_n23240_;
  assign ys__n24160 = ~ys__n1084 & ~new_n23241_;
  assign ys__n24162 = ~ys__n24107 & ys__n24167;
  assign new_n23244_ = ~ys__n318 & ~ys__n38564;
  assign new_n23245_ = ys__n318 & ys__n38564;
  assign new_n23246_ = ~new_n23244_ & ~new_n23245_;
  assign new_n23247_ = ~ys__n24112 & ~new_n23246_;
  assign new_n23248_ = ~ys__n306 & ys__n24112;
  assign new_n23249_ = ~new_n23247_ & ~new_n23248_;
  assign new_n23250_ = ~ys__n1072 & ys__n1073;
  assign new_n23251_ = ~new_n23249_ & new_n23250_;
  assign new_n23252_ = ys__n1072 & ys__n24162;
  assign ys__n24163 = new_n23251_ | new_n23252_;
  assign ys__n24165 = ~ys__n24107 & ys__n24168;
  assign new_n23255_ = ys__n318 & ~ys__n624;
  assign new_n23256_ = ~ys__n318 & ys__n624;
  assign ys__n38566 = new_n23255_ | new_n23256_;
  assign new_n23258_ = ~ys__n38565 & ys__n38566;
  assign new_n23259_ = ys__n38565 & ~ys__n38566;
  assign new_n23260_ = ~new_n23258_ & ~new_n23259_;
  assign new_n23261_ = ~ys__n24112 & ~new_n23260_;
  assign new_n23262_ = ys__n306 & ~ys__n38568;
  assign new_n23263_ = ~ys__n306 & ys__n38568;
  assign new_n23264_ = ~new_n23262_ & ~new_n23263_;
  assign new_n23265_ = ys__n24112 & ~new_n23264_;
  assign new_n23266_ = ~new_n23261_ & ~new_n23265_;
  assign new_n23267_ = new_n23250_ & ~new_n23266_;
  assign new_n23268_ = ys__n1072 & ys__n24165;
  assign ys__n24166 = new_n23267_ | new_n23268_;
  assign new_n23270_ = ys__n24167 & ~ys__n24177;
  assign new_n23271_ = ys__n306 & ys__n24177;
  assign new_n23272_ = ~new_n23270_ & ~new_n23271_;
  assign new_n23273_ = ys__n1072 & new_n18058_;
  assign new_n23274_ = ~new_n23272_ & ~new_n23273_;
  assign new_n23275_ = ys__n24116 & new_n23273_;
  assign ys__n24176 = new_n23274_ | new_n23275_;
  assign new_n23277_ = ys__n47665 & new_n12768_;
  assign new_n23278_ = ys__n22830 & ~new_n12314_;
  assign new_n23279_ = new_n12309_ & new_n23278_;
  assign new_n23280_ = ~new_n17429_ & ~new_n23279_;
  assign new_n23281_ = ~new_n12320_ & ~new_n23280_;
  assign new_n23282_ = ys__n23552 & new_n12320_;
  assign new_n23283_ = ~new_n23281_ & ~new_n23282_;
  assign new_n23284_ = ~new_n12404_ & ~new_n23283_;
  assign new_n23285_ = new_n12404_ & ys__n23489;
  assign new_n23286_ = ~new_n23284_ & ~new_n23285_;
  assign new_n23287_ = new_n12458_ & ~new_n23286_;
  assign new_n23288_ = ys__n524 & ~new_n12458_;
  assign new_n23289_ = ~new_n23287_ & ~new_n23288_;
  assign new_n23290_ = ~new_n12477_ & ~new_n23289_;
  assign new_n23291_ = ~new_n12531_ & new_n12576_;
  assign new_n23292_ = new_n12531_ & ~new_n12576_;
  assign new_n23293_ = ~new_n23291_ & ~new_n23292_;
  assign new_n23294_ = new_n12477_ & ~new_n23293_;
  assign new_n23295_ = ~new_n23290_ & ~new_n23294_;
  assign new_n23296_ = new_n12763_ & ~new_n23295_;
  assign new_n23297_ = ~new_n23277_ & ~new_n23296_;
  assign new_n23298_ = new_n12774_ & ~new_n23297_;
  assign new_n23299_ = ys__n47665 & new_n12778_;
  assign new_n23300_ = new_n12776_ & ~new_n23295_;
  assign new_n23301_ = ~new_n23299_ & ~new_n23300_;
  assign new_n23302_ = new_n12784_ & ~new_n23301_;
  assign ys__n24179 = new_n23298_ | new_n23302_;
  assign new_n23304_ = ~ys__n1084 & ~ys__n24177;
  assign new_n23305_ = ys__n24197 & new_n23304_;
  assign new_n23306_ = ys__n24177 & ys__n24209;
  assign new_n23307_ = ~new_n23305_ & ~new_n23306_;
  assign new_n23308_ = ~ys__n1078 & ~new_n23307_;
  assign new_n23309_ = ys__n1078 & ys__n24197;
  assign new_n23310_ = ~new_n23308_ & ~new_n23309_;
  assign new_n23311_ = ~new_n23273_ & ~new_n23310_;
  assign new_n23312_ = new_n23273_ & ys__n24179;
  assign ys__n24180 = new_n23311_ | new_n23312_;
  assign new_n23314_ = ys__n47666 & new_n12768_;
  assign new_n23315_ = ys__n22832 & ~new_n12314_;
  assign new_n23316_ = new_n12309_ & new_n23315_;
  assign new_n23317_ = ~new_n17435_ & ~new_n23316_;
  assign new_n23318_ = ~new_n12320_ & ~new_n23317_;
  assign new_n23319_ = ys__n23554 & new_n12320_;
  assign new_n23320_ = ~new_n23318_ & ~new_n23319_;
  assign new_n23321_ = ~new_n12404_ & ~new_n23320_;
  assign new_n23322_ = new_n12404_ & ys__n23491;
  assign new_n23323_ = ~new_n23321_ & ~new_n23322_;
  assign new_n23324_ = new_n12458_ & ~new_n23323_;
  assign new_n23325_ = ys__n522 & ~new_n12458_;
  assign new_n23326_ = ~new_n23324_ & ~new_n23325_;
  assign new_n23327_ = ~new_n12477_ & ~new_n23326_;
  assign new_n23328_ = ~new_n12531_ & ~new_n12576_;
  assign new_n23329_ = ~new_n12581_ & ~new_n23328_;
  assign new_n23330_ = new_n12565_ & ~new_n23329_;
  assign new_n23331_ = ~new_n12565_ & new_n23329_;
  assign new_n23332_ = ~new_n23330_ & ~new_n23331_;
  assign new_n23333_ = new_n12477_ & ~new_n23332_;
  assign new_n23334_ = ~new_n23327_ & ~new_n23333_;
  assign new_n23335_ = new_n12763_ & ~new_n23334_;
  assign new_n23336_ = ~new_n23314_ & ~new_n23335_;
  assign new_n23337_ = new_n12774_ & ~new_n23336_;
  assign new_n23338_ = ys__n47666 & new_n12778_;
  assign new_n23339_ = new_n12776_ & ~new_n23334_;
  assign new_n23340_ = ~new_n23338_ & ~new_n23339_;
  assign new_n23341_ = new_n12784_ & ~new_n23340_;
  assign ys__n24182 = new_n23337_ | new_n23341_;
  assign new_n23343_ = ys__n24199 & new_n23304_;
  assign new_n23344_ = ys__n24177 & ys__n24211;
  assign new_n23345_ = ~new_n23343_ & ~new_n23344_;
  assign new_n23346_ = ~ys__n1078 & ~new_n23345_;
  assign new_n23347_ = ys__n1078 & ys__n24199;
  assign new_n23348_ = ~new_n23346_ & ~new_n23347_;
  assign new_n23349_ = ~new_n23273_ & ~new_n23348_;
  assign new_n23350_ = new_n23273_ & ys__n24182;
  assign ys__n24183 = new_n23349_ | new_n23350_;
  assign new_n23352_ = ys__n47667 & new_n12768_;
  assign new_n23353_ = ys__n22834 & ~new_n12314_;
  assign new_n23354_ = new_n12309_ & new_n23353_;
  assign new_n23355_ = ~new_n17441_ & ~new_n23354_;
  assign new_n23356_ = ~new_n12320_ & ~new_n23355_;
  assign new_n23357_ = ys__n23556 & new_n12320_;
  assign new_n23358_ = ~new_n23356_ & ~new_n23357_;
  assign new_n23359_ = ~new_n12404_ & ~new_n23358_;
  assign new_n23360_ = new_n12404_ & ys__n23493;
  assign new_n23361_ = ~new_n23359_ & ~new_n23360_;
  assign new_n23362_ = new_n12458_ & ~new_n23361_;
  assign new_n23363_ = ys__n530 & ~new_n12458_;
  assign new_n23364_ = ~new_n23362_ & ~new_n23363_;
  assign new_n23365_ = ~new_n12477_ & ~new_n23364_;
  assign new_n23366_ = ~new_n12531_ & new_n12577_;
  assign new_n23367_ = new_n12583_ & ~new_n23366_;
  assign new_n23368_ = new_n12553_ & ~new_n23367_;
  assign new_n23369_ = ~new_n12553_ & new_n23367_;
  assign new_n23370_ = ~new_n23368_ & ~new_n23369_;
  assign new_n23371_ = new_n12477_ & ~new_n23370_;
  assign new_n23372_ = ~new_n23365_ & ~new_n23371_;
  assign new_n23373_ = new_n12763_ & ~new_n23372_;
  assign new_n23374_ = ~new_n23352_ & ~new_n23373_;
  assign new_n23375_ = new_n12774_ & ~new_n23374_;
  assign new_n23376_ = ys__n47667 & new_n12778_;
  assign new_n23377_ = new_n12776_ & ~new_n23372_;
  assign new_n23378_ = ~new_n23376_ & ~new_n23377_;
  assign new_n23379_ = new_n12784_ & ~new_n23378_;
  assign ys__n24185 = new_n23375_ | new_n23379_;
  assign new_n23381_ = ys__n24201 & new_n23304_;
  assign new_n23382_ = ys__n24177 & ys__n24213;
  assign new_n23383_ = ~new_n23381_ & ~new_n23382_;
  assign new_n23384_ = ~ys__n1078 & ~new_n23383_;
  assign new_n23385_ = ys__n1078 & ys__n24201;
  assign new_n23386_ = ~new_n23384_ & ~new_n23385_;
  assign new_n23387_ = ~new_n23273_ & ~new_n23386_;
  assign new_n23388_ = new_n23273_ & ys__n24185;
  assign ys__n24186 = new_n23387_ | new_n23388_;
  assign new_n23390_ = ys__n22836 & ~new_n12314_;
  assign new_n23391_ = new_n12309_ & new_n23390_;
  assign new_n23392_ = ~new_n17447_ & ~new_n23391_;
  assign new_n23393_ = ~new_n12320_ & ~new_n23392_;
  assign new_n23394_ = ys__n23558 & new_n12320_;
  assign new_n23395_ = ~new_n23393_ & ~new_n23394_;
  assign new_n23396_ = ~new_n12404_ & ~new_n23395_;
  assign new_n23397_ = new_n12404_ & ys__n23495;
  assign new_n23398_ = ~new_n23396_ & ~new_n23397_;
  assign new_n23399_ = new_n12458_ & ~new_n23398_;
  assign new_n23400_ = ys__n752 & ~new_n12458_;
  assign new_n23401_ = ~new_n23399_ & ~new_n23400_;
  assign new_n23402_ = ~new_n12477_ & ~new_n23401_;
  assign new_n23403_ = ~new_n12553_ & ~new_n23367_;
  assign new_n23404_ = ~new_n12586_ & ~new_n23403_;
  assign new_n23405_ = new_n12542_ & ~new_n23404_;
  assign new_n23406_ = ~new_n12542_ & new_n23404_;
  assign new_n23407_ = ~new_n23405_ & ~new_n23406_;
  assign new_n23408_ = new_n12477_ & ~new_n23407_;
  assign new_n23409_ = ~new_n23402_ & ~new_n23408_;
  assign new_n23410_ = new_n12763_ & ~new_n23409_;
  assign new_n23411_ = ~ys__n935 & new_n12762_;
  assign new_n23412_ = ys__n47668 & new_n12768_;
  assign new_n23413_ = ~new_n23411_ & ~new_n23412_;
  assign new_n23414_ = ~new_n23410_ & new_n23413_;
  assign new_n23415_ = new_n12774_ & ~new_n23414_;
  assign new_n23416_ = new_n12776_ & ~new_n23409_;
  assign new_n23417_ = ys__n47668 & new_n12778_;
  assign new_n23418_ = ~new_n23411_ & ~new_n23417_;
  assign new_n23419_ = ~new_n23416_ & new_n23418_;
  assign new_n23420_ = new_n12784_ & ~new_n23419_;
  assign ys__n24188 = new_n23415_ | new_n23420_;
  assign new_n23422_ = ys__n24203 & new_n23304_;
  assign new_n23423_ = ys__n24177 & ys__n24215;
  assign new_n23424_ = ~new_n23422_ & ~new_n23423_;
  assign new_n23425_ = ~ys__n1078 & ~new_n23424_;
  assign new_n23426_ = ys__n1078 & ys__n24203;
  assign new_n23427_ = ~new_n23425_ & ~new_n23426_;
  assign new_n23428_ = ~new_n23273_ & ~new_n23427_;
  assign new_n23429_ = new_n23273_ & ys__n24188;
  assign ys__n24189 = new_n23428_ | new_n23429_;
  assign new_n23431_ = ys__n22838 & ~new_n12314_;
  assign new_n23432_ = new_n12309_ & new_n23431_;
  assign new_n23433_ = ~new_n17453_ & ~new_n23432_;
  assign new_n23434_ = ~new_n12320_ & ~new_n23433_;
  assign new_n23435_ = ys__n23560 & new_n12320_;
  assign new_n23436_ = ~new_n23434_ & ~new_n23435_;
  assign new_n23437_ = ~new_n12404_ & ~new_n23436_;
  assign new_n23438_ = new_n12404_ & ys__n23497;
  assign new_n23439_ = ~new_n23437_ & ~new_n23438_;
  assign new_n23440_ = new_n12458_ & ~new_n23439_;
  assign new_n23441_ = ys__n736 & ~new_n12458_;
  assign new_n23442_ = ~new_n23440_ & ~new_n23441_;
  assign new_n23443_ = ~new_n12477_ & ~new_n23442_;
  assign new_n23444_ = ~new_n12590_ & new_n12669_;
  assign new_n23445_ = new_n12590_ & ~new_n12669_;
  assign new_n23446_ = ~new_n23444_ & ~new_n23445_;
  assign new_n23447_ = new_n12477_ & ~new_n23446_;
  assign new_n23448_ = ~new_n23443_ & ~new_n23447_;
  assign new_n23449_ = new_n12763_ & ~new_n23448_;
  assign new_n23450_ = new_n12762_ & new_n12765_;
  assign new_n23451_ = ys__n47669 & new_n12768_;
  assign new_n23452_ = ~new_n23450_ & ~new_n23451_;
  assign new_n23453_ = ~new_n23449_ & new_n23452_;
  assign new_n23454_ = new_n12774_ & ~new_n23453_;
  assign new_n23455_ = new_n12776_ & ~new_n23448_;
  assign new_n23456_ = ys__n47669 & new_n12778_;
  assign new_n23457_ = ~new_n23450_ & ~new_n23456_;
  assign new_n23458_ = ~new_n23455_ & new_n23457_;
  assign new_n23459_ = new_n12784_ & ~new_n23458_;
  assign ys__n24191 = new_n23454_ | new_n23459_;
  assign new_n23461_ = ys__n24205 & new_n23304_;
  assign new_n23462_ = ys__n24177 & ys__n24217;
  assign new_n23463_ = ~new_n23461_ & ~new_n23462_;
  assign new_n23464_ = ~ys__n1078 & ~new_n23463_;
  assign new_n23465_ = ys__n1078 & ys__n24205;
  assign new_n23466_ = ~new_n23464_ & ~new_n23465_;
  assign new_n23467_ = ~new_n23273_ & ~new_n23466_;
  assign new_n23468_ = new_n23273_ & ys__n24191;
  assign ys__n24192 = new_n23467_ | new_n23468_;
  assign new_n23470_ = ys__n22840 & ~new_n12314_;
  assign new_n23471_ = new_n12309_ & new_n23470_;
  assign new_n23472_ = ~new_n17459_ & ~new_n23471_;
  assign new_n23473_ = ~new_n12320_ & ~new_n23472_;
  assign new_n23474_ = ys__n23562 & new_n12320_;
  assign new_n23475_ = ~new_n23473_ & ~new_n23474_;
  assign new_n23476_ = ~new_n12404_ & ~new_n23475_;
  assign new_n23477_ = new_n12404_ & ys__n23499;
  assign new_n23478_ = ~new_n23476_ & ~new_n23477_;
  assign new_n23479_ = new_n12458_ & ~new_n23478_;
  assign new_n23480_ = ys__n4488 & ~new_n12458_;
  assign new_n23481_ = ~new_n23479_ & ~new_n23480_;
  assign new_n23482_ = ~new_n12477_ & ~new_n23481_;
  assign new_n23483_ = ~new_n12590_ & ~new_n12669_;
  assign new_n23484_ = ~new_n12675_ & ~new_n23483_;
  assign new_n23485_ = new_n12659_ & ~new_n23484_;
  assign new_n23486_ = ~new_n12659_ & new_n23484_;
  assign new_n23487_ = ~new_n23485_ & ~new_n23486_;
  assign new_n23488_ = new_n12477_ & ~new_n23487_;
  assign new_n23489_ = ~new_n23482_ & ~new_n23488_;
  assign new_n23490_ = new_n12763_ & ~new_n23489_;
  assign new_n23491_ = ys__n935 & new_n12762_;
  assign new_n23492_ = ys__n47670 & new_n12768_;
  assign new_n23493_ = ~new_n23491_ & ~new_n23492_;
  assign new_n23494_ = ~new_n23490_ & new_n23493_;
  assign new_n23495_ = new_n12774_ & ~new_n23494_;
  assign new_n23496_ = new_n12776_ & ~new_n23489_;
  assign new_n23497_ = ys__n47670 & new_n12778_;
  assign new_n23498_ = ~new_n23491_ & ~new_n23497_;
  assign new_n23499_ = ~new_n23496_ & new_n23498_;
  assign new_n23500_ = new_n12784_ & ~new_n23499_;
  assign ys__n24194 = new_n23495_ | new_n23500_;
  assign new_n23502_ = ~ys__n1084 & ys__n24207;
  assign new_n23503_ = ys__n312 & ys__n1084;
  assign new_n23504_ = ~new_n23502_ & ~new_n23503_;
  assign new_n23505_ = ~ys__n24177 & ~new_n23504_;
  assign new_n23506_ = ys__n24177 & ys__n24219;
  assign new_n23507_ = ~new_n23505_ & ~new_n23506_;
  assign new_n23508_ = ~ys__n1078 & ~new_n23507_;
  assign new_n23509_ = ys__n1078 & ys__n24207;
  assign new_n23510_ = ~new_n23508_ & ~new_n23509_;
  assign new_n23511_ = ~new_n23273_ & ~new_n23510_;
  assign new_n23512_ = new_n23273_ & ys__n24194;
  assign ys__n24195 = new_n23511_ | new_n23512_;
  assign new_n23514_ = ys__n318 & ys__n624;
  assign new_n23515_ = ys__n18124 & new_n23514_;
  assign new_n23516_ = ys__n24177 & ~ys__n1079;
  assign new_n23517_ = ~new_n23515_ & new_n23516_;
  assign new_n23518_ = ys__n38561 & new_n23240_;
  assign new_n23519_ = new_n23273_ & ~new_n23518_;
  assign new_n23520_ = ~ys__n18120 & new_n23519_;
  assign new_n23521_ = new_n11730_ & new_n23520_;
  assign new_n23522_ = ys__n1072 & ~ys__n24228;
  assign new_n23523_ = ~ys__n33442 & new_n23522_;
  assign new_n23524_ = new_n18058_ & new_n23523_;
  assign new_n23525_ = ~ys__n18120 & new_n23524_;
  assign new_n23526_ = new_n23521_ & new_n23525_;
  assign ys__n24222 = new_n23517_ | new_n23526_;
  assign new_n23528_ = ys__n1072 & ~ys__n1076;
  assign new_n23529_ = ys__n24228 & new_n23528_;
  assign new_n23530_ = ys__n1076 & ~ys__n24235;
  assign ys__n24227 = new_n23529_ | new_n23530_;
  assign new_n23532_ = ~ys__n24177 & ys__n24233;
  assign new_n23533_ = ~ys__n24243 & new_n23532_;
  assign new_n23534_ = ys__n24177 & new_n23515_;
  assign ys__n24231 = new_n23533_ | new_n23534_;
  assign new_n23536_ = ~ys__n1072 & ys__n1078;
  assign new_n23537_ = ~ys__n33442 & new_n23521_;
  assign new_n23538_ = ~ys__n18120 & ~new_n23537_;
  assign new_n23539_ = ~ys__n18120 & new_n18058_;
  assign new_n23540_ = ~new_n23538_ & new_n23539_;
  assign new_n23541_ = ~ys__n24243 & new_n23522_;
  assign new_n23542_ = ~new_n23540_ & new_n23541_;
  assign new_n23543_ = ~new_n23536_ & ~new_n23542_;
  assign new_n23544_ = ~ys__n1076 & ~new_n23543_;
  assign new_n23545_ = ys__n1076 & ys__n24235;
  assign ys__n24236 = new_n23544_ | new_n23545_;
  assign ys__n38556 = ys__n24233 & ys__n24243;
  assign new_n23548_ = ~ys__n24177 & ~ys__n1079;
  assign new_n23549_ = ys__n38556 & new_n23548_;
  assign new_n23550_ = ys__n24243 & new_n23522_;
  assign new_n23551_ = ~new_n23521_ & new_n23550_;
  assign ys__n24240 = new_n23549_ | new_n23551_;
  assign new_n23553_ = ~ys__n1084 & ys__n24248;
  assign new_n23554_ = new_n23530_ & new_n23553_;
  assign new_n23555_ = ys__n1084 & ~ys__n18015;
  assign new_n23556_ = ~new_n23554_ & ~new_n23555_;
  assign new_n23557_ = ~ys__n140 & ~new_n23556_;
  assign ys__n24245 = ys__n140 | new_n23557_;
  assign new_n23559_ = ~ys__n1076 & ~ys__n24235;
  assign new_n23560_ = ys__n24248 & new_n23559_;
  assign ys__n24250 = ys__n24235 | new_n23560_;
  assign new_n23562_ = ~ys__n24464 & ys__n24483;
  assign new_n23563_ = ys__n24464 & new_n17716_;
  assign new_n23564_ = ~new_n23562_ & ~new_n23563_;
  assign new_n23565_ = ~ys__n24463 & ~new_n23564_;
  assign new_n23566_ = ~new_n15124_ & ~new_n23565_;
  assign new_n23567_ = ~ys__n1120 & ~ys__n24461;
  assign new_n23568_ = ~new_n23566_ & new_n23567_;
  assign new_n23569_ = ~ys__n1120 & ~new_n23568_;
  assign new_n23570_ = ~ys__n1116 & ~ys__n1117;
  assign new_n23571_ = ~ys__n1119 & new_n23570_;
  assign new_n23572_ = ~new_n23569_ & new_n23571_;
  assign new_n23573_ = ys__n690 & ys__n692;
  assign new_n23574_ = ys__n694 & ys__n696;
  assign new_n23575_ = new_n23573_ & new_n23574_;
  assign new_n23576_ = ys__n606 & ys__n608;
  assign new_n23577_ = ys__n610 & ys__n688;
  assign new_n23578_ = new_n23576_ & new_n23577_;
  assign new_n23579_ = new_n23575_ & new_n23578_;
  assign new_n23580_ = ~ys__n38654 & ~new_n23579_;
  assign new_n23581_ = new_n17716_ & new_n23580_;
  assign new_n23582_ = ys__n140 & ys__n1119;
  assign new_n23583_ = new_n23581_ & new_n23582_;
  assign new_n23584_ = ~new_n23572_ & ~new_n23583_;
  assign new_n23585_ = new_n13631_ & ~new_n23584_;
  assign new_n23586_ = ~ys__n1110 & ~new_n23585_;
  assign new_n23587_ = ~ys__n1099 & ~ys__n1109;
  assign new_n23588_ = new_n13609_ & new_n23587_;
  assign new_n23589_ = ~new_n23586_ & new_n23588_;
  assign new_n23590_ = ys__n1099 & ys__n24506;
  assign new_n23591_ = ~new_n23589_ & ~new_n23590_;
  assign new_n23592_ = ~ys__n1106 & ~new_n23591_;
  assign new_n23593_ = ys__n1106 & ys__n33495;
  assign new_n23594_ = new_n17716_ & new_n23593_;
  assign new_n23595_ = ~ys__n4696 & new_n23594_;
  assign new_n23596_ = ys__n33481 & new_n23595_;
  assign new_n23597_ = ~ys__n33493 & ys__n4696;
  assign new_n23598_ = ys__n33495 & ~new_n23580_;
  assign new_n23599_ = ~ys__n33497 & ~new_n13606_;
  assign new_n23600_ = ys__n1106 & ys__n33491;
  assign new_n23601_ = ~new_n23599_ & new_n23600_;
  assign new_n23602_ = ~ys__n24567 & ~ys__n33495;
  assign new_n23603_ = ~ys__n33497 & ~ys__n33499;
  assign new_n23604_ = new_n23602_ & new_n23603_;
  assign new_n23605_ = new_n17716_ & ~new_n23604_;
  assign new_n23606_ = ~new_n23601_ & new_n23605_;
  assign new_n23607_ = ~ys__n4566 & new_n23606_;
  assign new_n23608_ = ~new_n23598_ & new_n23607_;
  assign new_n23609_ = ~new_n23597_ & new_n23608_;
  assign new_n23610_ = ~new_n23596_ & new_n23609_;
  assign new_n23611_ = ys__n1106 & ~new_n23610_;
  assign new_n23612_ = ~new_n23592_ & ~new_n23611_;
  assign ys__n24502 = ~ys__n1094 & ~new_n23612_;
  assign new_n23614_ = ys__n1106 & ~ys__n33493;
  assign new_n23615_ = ~new_n23580_ & new_n23614_;
  assign new_n23616_ = ~ys__n33493 & ys__n1088;
  assign new_n23617_ = ys__n1106 & ys__n33479;
  assign new_n23618_ = ~ys__n1119 & ~new_n23617_;
  assign new_n23619_ = ~new_n23616_ & new_n23618_;
  assign new_n23620_ = ~new_n23615_ & new_n23619_;
  assign new_n23621_ = ~ys__n33495 & ~ys__n33497;
  assign new_n23622_ = new_n17716_ & ~new_n23621_;
  assign new_n23623_ = ~new_n23620_ & new_n23622_;
  assign ys__n24271 = ~ys__n4696 & new_n23623_;
  assign new_n23625_ = ys__n1106 & ~new_n23601_;
  assign new_n23626_ = new_n23580_ & new_n23625_;
  assign new_n23627_ = ~ys__n4566 & new_n23626_;
  assign new_n23628_ = new_n23595_ & new_n23627_;
  assign ys__n33457 = ~ys__n24271 & new_n23628_;
  assign new_n23630_ = ys__n24502 & ys__n33457;
  assign ys__n33455 = ys__n24519 & ~new_n13610_;
  assign new_n23632_ = ys__n38631 & ~ys__n4696;
  assign ys__n38633 = ys__n33455 | new_n23632_;
  assign ys__n24258 = ys__n38624 | ~new_n17716_;
  assign new_n23635_ = ys__n24256 & ~ys__n24258;
  assign new_n23636_ = ys__n33497 & ys__n24258;
  assign new_n23637_ = ~ys__n4566 & new_n23636_;
  assign ys__n24259 = new_n23635_ | new_n23637_;
  assign new_n23639_ = ~ys__n1511 & ys__n30216;
  assign new_n23640_ = ~ys__n24258 & new_n23639_;
  assign new_n23641_ = ~ys__n4566 & new_n23640_;
  assign new_n23642_ = ys__n38670 & ys__n24258;
  assign new_n23643_ = ~ys__n4566 & new_n23642_;
  assign ys__n24265 = new_n23641_ | new_n23643_;
  assign new_n23645_ = ~ys__n24259 & ~ys__n24265;
  assign new_n23646_ = ~ys__n1106 & ~ys__n1119;
  assign new_n23647_ = ~ys__n1120 & ~ys__n24463;
  assign new_n23648_ = ~ys__n24464 & new_n23647_;
  assign new_n23649_ = new_n23646_ & new_n23648_;
  assign new_n23650_ = ~new_n23645_ & ~new_n23649_;
  assign new_n23651_ = ys__n38633 & new_n23650_;
  assign new_n23652_ = ~new_n23630_ & new_n23651_;
  assign new_n23653_ = ~ys__n33464 & ys__n33488;
  assign new_n23654_ = new_n13617_ & new_n23653_;
  assign ys__n38628 = ~ys__n33481 & new_n23595_;
  assign new_n23656_ = ~new_n13617_ & ys__n38628;
  assign new_n23657_ = ~new_n23654_ & ~new_n23656_;
  assign new_n23658_ = ~ys__n24271 & ~new_n23657_;
  assign new_n23659_ = ys__n24271 & new_n23654_;
  assign ys__n24272 = new_n23658_ | new_n23659_;
  assign new_n23661_ = ys__n33552 & ys__n24272;
  assign new_n23662_ = new_n23645_ & ~new_n23661_;
  assign new_n23663_ = ys__n38633 & ~new_n23649_;
  assign new_n23664_ = new_n23630_ & new_n23663_;
  assign new_n23665_ = ~new_n23662_ & new_n23664_;
  assign ys__n24255 = new_n23652_ | new_n23665_;
  assign ys__n24260 = ys__n30216 & ~ys__n4566;
  assign new_n23668_ = ~ys__n24258 & ys__n24260;
  assign new_n23669_ = ys__n33495 & ys__n24258;
  assign new_n23670_ = ~ys__n4566 & new_n23669_;
  assign ys__n24262 = new_n23668_ | new_n23670_;
  assign new_n23672_ = ~ys__n1511 & ys__n30219;
  assign new_n23673_ = ~ys__n24258 & new_n23672_;
  assign new_n23674_ = ~ys__n4566 & new_n23673_;
  assign new_n23675_ = ys__n33493 & ys__n24258;
  assign new_n23676_ = ~ys__n4566 & new_n23675_;
  assign ys__n24268 = new_n23674_ | new_n23676_;
  assign ys__n24274 = ~ys__n24107 & ys__n24279;
  assign new_n23679_ = ~ys__n454 & ~ys__n38693;
  assign new_n23680_ = ys__n454 & ys__n38693;
  assign new_n23681_ = ~new_n23679_ & ~new_n23680_;
  assign new_n23682_ = ~ys__n24112 & ~new_n23681_;
  assign new_n23683_ = ~ys__n452 & ys__n24112;
  assign new_n23684_ = ~new_n23682_ & ~new_n23683_;
  assign new_n23685_ = ~ys__n1088 & ys__n1089;
  assign new_n23686_ = ~new_n23684_ & new_n23685_;
  assign new_n23687_ = ys__n1088 & ys__n24274;
  assign ys__n24275 = new_n23686_ | new_n23687_;
  assign ys__n24277 = ~ys__n24107 & ys__n24280;
  assign new_n23690_ = ys__n454 & ~ys__n712;
  assign new_n23691_ = ~ys__n454 & ys__n712;
  assign ys__n35425 = new_n23690_ | new_n23691_;
  assign new_n23693_ = ~ys__n38694 & ys__n35425;
  assign new_n23694_ = ys__n38694 & ~ys__n35425;
  assign new_n23695_ = ~new_n23693_ & ~new_n23694_;
  assign new_n23696_ = ~ys__n24112 & ~new_n23695_;
  assign new_n23697_ = ys__n452 & ~ys__n35426;
  assign new_n23698_ = ~ys__n452 & ys__n35426;
  assign new_n23699_ = ~new_n23697_ & ~new_n23698_;
  assign new_n23700_ = ys__n24112 & ~new_n23699_;
  assign new_n23701_ = ~new_n23696_ & ~new_n23700_;
  assign new_n23702_ = new_n23685_ & ~new_n23701_;
  assign new_n23703_ = ys__n1088 & ys__n24277;
  assign ys__n24278 = new_n23702_ | new_n23703_;
  assign new_n23705_ = ~ys__n80 & ~ys__n82;
  assign new_n23706_ = ys__n84 & ys__n86;
  assign new_n23707_ = new_n23705_ & new_n23706_;
  assign new_n23708_ = ys__n84 & ~ys__n86;
  assign new_n23709_ = new_n23705_ & new_n23708_;
  assign new_n23710_ = ~new_n23707_ & ~new_n23709_;
  assign new_n23711_ = ~ys__n84 & ys__n86;
  assign new_n23712_ = new_n23705_ & new_n23711_;
  assign new_n23713_ = ~ys__n84 & ~ys__n86;
  assign new_n23714_ = new_n23705_ & new_n23713_;
  assign new_n23715_ = ~new_n23712_ & ~new_n23714_;
  assign new_n23716_ = new_n23710_ & new_n23715_;
  assign new_n23717_ = ys__n80 & ~ys__n82;
  assign new_n23718_ = new_n23708_ & new_n23717_;
  assign new_n23719_ = new_n23713_ & new_n23717_;
  assign new_n23720_ = ~new_n23718_ & ~new_n23719_;
  assign new_n23721_ = new_n23716_ & new_n23720_;
  assign new_n23722_ = ys__n80 & ys__n82;
  assign new_n23723_ = new_n23713_ & new_n23722_;
  assign new_n23724_ = new_n23721_ & ~new_n23723_;
  assign new_n23725_ = ~new_n23721_ & ~new_n23724_;
  assign new_n23726_ = ys__n47194 & ~new_n23725_;
  assign new_n23727_ = ~new_n23709_ & ~new_n23718_;
  assign new_n23728_ = ys__n47193 & ~new_n23727_;
  assign new_n23729_ = ~new_n23714_ & ~new_n23719_;
  assign new_n23730_ = ys__n47201 & ~new_n23729_;
  assign new_n23731_ = ys__n47009 & new_n23712_;
  assign new_n23732_ = ys__n47001 & new_n23707_;
  assign new_n23733_ = ~new_n23731_ & ~new_n23732_;
  assign new_n23734_ = ~new_n23730_ & new_n23733_;
  assign new_n23735_ = ~new_n23728_ & new_n23734_;
  assign new_n23736_ = ~new_n23707_ & ~new_n23712_;
  assign new_n23737_ = new_n23727_ & new_n23729_;
  assign new_n23738_ = new_n23736_ & new_n23737_;
  assign new_n23739_ = ys__n38898 & ~new_n23738_;
  assign new_n23740_ = ~new_n23735_ & new_n23739_;
  assign new_n23741_ = new_n23725_ & new_n23740_;
  assign new_n23742_ = ~new_n23726_ & ~new_n23741_;
  assign new_n23743_ = ys__n18149 & ys__n18137;
  assign new_n23744_ = new_n17355_ & new_n23743_;
  assign new_n23745_ = ~ys__n1154 & ~ys__n38805;
  assign new_n23746_ = ~new_n23744_ & new_n23745_;
  assign new_n23747_ = new_n11743_ & ~new_n23746_;
  assign new_n23748_ = ~new_n23742_ & ~new_n23747_;
  assign new_n23749_ = ~ys__n1106 & ~ys__n1109;
  assign new_n23750_ = ~ys__n1116 & new_n23749_;
  assign new_n23751_ = new_n23748_ & new_n23750_;
  assign new_n23752_ = ~ys__n4176 & new_n11743_;
  assign new_n23753_ = ys__n33407 & new_n23752_;
  assign new_n23754_ = ys__n28932 & new_n23753_;
  assign new_n23755_ = ys__n33409 & new_n23752_;
  assign new_n23756_ = ys__n29286 & new_n23755_;
  assign new_n23757_ = ys__n33411 & new_n23752_;
  assign new_n23758_ = ys__n29593 & new_n23757_;
  assign new_n23759_ = ys__n29594 & ~new_n23757_;
  assign new_n23760_ = ~new_n23758_ & ~new_n23759_;
  assign new_n23761_ = ~new_n23755_ & ~new_n23760_;
  assign new_n23762_ = ~new_n23756_ & ~new_n23761_;
  assign new_n23763_ = ~new_n23753_ & ~new_n23762_;
  assign new_n23764_ = ~new_n23754_ & ~new_n23763_;
  assign new_n23765_ = ~new_n23750_ & ~new_n23764_;
  assign ys__n24286 = new_n23751_ | new_n23765_;
  assign new_n23767_ = ys__n47195 & ~new_n23725_;
  assign new_n23768_ = ~new_n23741_ & ~new_n23767_;
  assign new_n23769_ = ~new_n23747_ & ~new_n23768_;
  assign new_n23770_ = new_n23750_ & new_n23769_;
  assign new_n23771_ = ys__n28935 & new_n23753_;
  assign new_n23772_ = ys__n29288 & new_n23755_;
  assign new_n23773_ = ys__n29595 & new_n23757_;
  assign new_n23774_ = ys__n29596 & ~new_n23757_;
  assign new_n23775_ = ~new_n23773_ & ~new_n23774_;
  assign new_n23776_ = ~new_n23755_ & ~new_n23775_;
  assign new_n23777_ = ~new_n23772_ & ~new_n23776_;
  assign new_n23778_ = ~new_n23753_ & ~new_n23777_;
  assign new_n23779_ = ~new_n23771_ & ~new_n23778_;
  assign new_n23780_ = ~new_n23750_ & ~new_n23779_;
  assign ys__n24289 = new_n23770_ | new_n23780_;
  assign new_n23782_ = ys__n47196 & ~new_n23725_;
  assign new_n23783_ = ~new_n23741_ & ~new_n23782_;
  assign new_n23784_ = ~new_n23747_ & ~new_n23783_;
  assign new_n23785_ = new_n23750_ & new_n23784_;
  assign new_n23786_ = ys__n28938 & new_n23753_;
  assign new_n23787_ = ys__n29290 & new_n23755_;
  assign new_n23788_ = ys__n29597 & new_n23757_;
  assign new_n23789_ = ys__n29598 & ~new_n23757_;
  assign new_n23790_ = ~new_n23788_ & ~new_n23789_;
  assign new_n23791_ = ~new_n23755_ & ~new_n23790_;
  assign new_n23792_ = ~new_n23787_ & ~new_n23791_;
  assign new_n23793_ = ~new_n23753_ & ~new_n23792_;
  assign new_n23794_ = ~new_n23786_ & ~new_n23793_;
  assign new_n23795_ = ~new_n23750_ & ~new_n23794_;
  assign ys__n24291 = new_n23785_ | new_n23795_;
  assign new_n23797_ = ys__n47197 & ~new_n23725_;
  assign new_n23798_ = ~new_n23741_ & ~new_n23797_;
  assign new_n23799_ = ~new_n23747_ & ~new_n23798_;
  assign new_n23800_ = new_n23750_ & new_n23799_;
  assign new_n23801_ = ys__n28941 & new_n23753_;
  assign new_n23802_ = ys__n29292 & new_n23755_;
  assign new_n23803_ = ys__n29599 & new_n23757_;
  assign new_n23804_ = ys__n29600 & ~new_n23757_;
  assign new_n23805_ = ~new_n23803_ & ~new_n23804_;
  assign new_n23806_ = ~new_n23755_ & ~new_n23805_;
  assign new_n23807_ = ~new_n23802_ & ~new_n23806_;
  assign new_n23808_ = ~new_n23753_ & ~new_n23807_;
  assign new_n23809_ = ~new_n23801_ & ~new_n23808_;
  assign new_n23810_ = ~new_n23750_ & ~new_n23809_;
  assign ys__n24293 = new_n23800_ | new_n23810_;
  assign new_n23812_ = ys__n47198 & ~new_n23725_;
  assign new_n23813_ = ~new_n23741_ & ~new_n23812_;
  assign new_n23814_ = ~new_n23747_ & ~new_n23813_;
  assign new_n23815_ = new_n23750_ & new_n23814_;
  assign new_n23816_ = ys__n28944 & new_n23753_;
  assign new_n23817_ = ys__n29294 & new_n23755_;
  assign new_n23818_ = ys__n29601 & new_n23757_;
  assign new_n23819_ = ys__n29602 & ~new_n23757_;
  assign new_n23820_ = ~new_n23818_ & ~new_n23819_;
  assign new_n23821_ = ~new_n23755_ & ~new_n23820_;
  assign new_n23822_ = ~new_n23817_ & ~new_n23821_;
  assign new_n23823_ = ~new_n23753_ & ~new_n23822_;
  assign new_n23824_ = ~new_n23816_ & ~new_n23823_;
  assign new_n23825_ = ~new_n23750_ & ~new_n23824_;
  assign ys__n24295 = new_n23815_ | new_n23825_;
  assign new_n23827_ = ys__n47199 & ~new_n23725_;
  assign new_n23828_ = ~new_n23741_ & ~new_n23827_;
  assign new_n23829_ = ~new_n23747_ & ~new_n23828_;
  assign new_n23830_ = new_n23750_ & new_n23829_;
  assign new_n23831_ = ys__n28947 & new_n23753_;
  assign new_n23832_ = ys__n29296 & new_n23755_;
  assign new_n23833_ = ys__n29603 & new_n23757_;
  assign new_n23834_ = ys__n29604 & ~new_n23757_;
  assign new_n23835_ = ~new_n23833_ & ~new_n23834_;
  assign new_n23836_ = ~new_n23755_ & ~new_n23835_;
  assign new_n23837_ = ~new_n23832_ & ~new_n23836_;
  assign new_n23838_ = ~new_n23753_ & ~new_n23837_;
  assign new_n23839_ = ~new_n23831_ & ~new_n23838_;
  assign new_n23840_ = ~new_n23750_ & ~new_n23839_;
  assign ys__n24297 = new_n23830_ | new_n23840_;
  assign new_n23842_ = ys__n47200 & ~new_n23725_;
  assign new_n23843_ = ~new_n23741_ & ~new_n23842_;
  assign new_n23844_ = ~new_n23747_ & ~new_n23843_;
  assign new_n23845_ = new_n23750_ & new_n23844_;
  assign new_n23846_ = ys__n28950 & new_n23753_;
  assign new_n23847_ = ys__n29298 & new_n23755_;
  assign new_n23848_ = ys__n29605 & new_n23757_;
  assign new_n23849_ = ys__n29606 & ~new_n23757_;
  assign new_n23850_ = ~new_n23848_ & ~new_n23849_;
  assign new_n23851_ = ~new_n23755_ & ~new_n23850_;
  assign new_n23852_ = ~new_n23847_ & ~new_n23851_;
  assign new_n23853_ = ~new_n23753_ & ~new_n23852_;
  assign new_n23854_ = ~new_n23846_ & ~new_n23853_;
  assign new_n23855_ = ~new_n23750_ & ~new_n23854_;
  assign ys__n24299 = new_n23845_ | new_n23855_;
  assign new_n23857_ = ys__n47201 & ~new_n23725_;
  assign new_n23858_ = ~new_n23741_ & ~new_n23857_;
  assign new_n23859_ = ~new_n23747_ & ~new_n23858_;
  assign new_n23860_ = new_n23750_ & new_n23859_;
  assign new_n23861_ = ys__n28953 & new_n23753_;
  assign new_n23862_ = ys__n29300 & new_n23755_;
  assign new_n23863_ = ys__n29607 & new_n23757_;
  assign new_n23864_ = ys__n29608 & ~new_n23757_;
  assign new_n23865_ = ~new_n23863_ & ~new_n23864_;
  assign new_n23866_ = ~new_n23755_ & ~new_n23865_;
  assign new_n23867_ = ~new_n23862_ & ~new_n23866_;
  assign new_n23868_ = ~new_n23753_ & ~new_n23867_;
  assign new_n23869_ = ~new_n23861_ & ~new_n23868_;
  assign new_n23870_ = ~new_n23750_ & ~new_n23869_;
  assign ys__n24301 = new_n23860_ | new_n23870_;
  assign new_n23872_ = ~ys__n33469 & new_n13607_;
  assign new_n23873_ = ys__n1107 & ys__n2693;
  assign new_n23874_ = new_n15121_ & new_n23873_;
  assign new_n23875_ = ~new_n23872_ & ~new_n23874_;
  assign new_n23876_ = ys__n24286 & new_n23875_;
  assign new_n23877_ = ys__n24303 & new_n23874_;
  assign ys__n24305 = new_n23876_ | new_n23877_;
  assign new_n23879_ = ys__n24289 & new_n23875_;
  assign new_n23880_ = ys__n24306 & new_n23874_;
  assign ys__n24307 = new_n23879_ | new_n23880_;
  assign new_n23882_ = ys__n24291 & new_n23875_;
  assign new_n23883_ = ys__n24308 & new_n23874_;
  assign ys__n24309 = new_n23882_ | new_n23883_;
  assign new_n23885_ = ys__n24293 & new_n23875_;
  assign new_n23886_ = ys__n24310 & new_n23874_;
  assign ys__n24311 = new_n23885_ | new_n23886_;
  assign new_n23888_ = ys__n24295 & new_n23875_;
  assign new_n23889_ = ys__n24312 & new_n23874_;
  assign ys__n24313 = new_n23888_ | new_n23889_;
  assign new_n23891_ = ys__n24297 & new_n23875_;
  assign new_n23892_ = ys__n24314 & new_n23874_;
  assign ys__n24315 = new_n23891_ | new_n23892_;
  assign new_n23894_ = ys__n24299 & new_n23875_;
  assign new_n23895_ = ys__n24316 & new_n23874_;
  assign ys__n24317 = new_n23894_ | new_n23895_;
  assign new_n23897_ = ys__n24301 & new_n23875_;
  assign new_n23898_ = ys__n24318 & new_n23874_;
  assign ys__n24319 = new_n23897_ | new_n23898_;
  assign new_n23900_ = ys__n47002 & ~new_n23725_;
  assign new_n23901_ = ~new_n23741_ & ~new_n23900_;
  assign new_n23902_ = ~new_n23747_ & ~new_n23901_;
  assign new_n23903_ = new_n23750_ & new_n23902_;
  assign new_n23904_ = ys__n28908 & new_n23753_;
  assign new_n23905_ = ys__n29270 & new_n23755_;
  assign new_n23906_ = ys__n29577 & new_n23757_;
  assign new_n23907_ = ys__n29578 & ~new_n23757_;
  assign new_n23908_ = ~new_n23906_ & ~new_n23907_;
  assign new_n23909_ = ~new_n23755_ & ~new_n23908_;
  assign new_n23910_ = ~new_n23905_ & ~new_n23909_;
  assign new_n23911_ = ~new_n23753_ & ~new_n23910_;
  assign new_n23912_ = ~new_n23904_ & ~new_n23911_;
  assign new_n23913_ = ~new_n23750_ & ~new_n23912_;
  assign ys__n24320 = new_n23903_ | new_n23913_;
  assign new_n23915_ = ys__n47003 & ~new_n23725_;
  assign new_n23916_ = ~new_n23741_ & ~new_n23915_;
  assign new_n23917_ = ~new_n23747_ & ~new_n23916_;
  assign new_n23918_ = new_n23750_ & new_n23917_;
  assign new_n23919_ = ys__n28911 & new_n23753_;
  assign new_n23920_ = ys__n29272 & new_n23755_;
  assign new_n23921_ = ys__n29579 & new_n23757_;
  assign new_n23922_ = ys__n29580 & ~new_n23757_;
  assign new_n23923_ = ~new_n23921_ & ~new_n23922_;
  assign new_n23924_ = ~new_n23755_ & ~new_n23923_;
  assign new_n23925_ = ~new_n23920_ & ~new_n23924_;
  assign new_n23926_ = ~new_n23753_ & ~new_n23925_;
  assign new_n23927_ = ~new_n23919_ & ~new_n23926_;
  assign new_n23928_ = ~new_n23750_ & ~new_n23927_;
  assign ys__n24323 = new_n23918_ | new_n23928_;
  assign new_n23930_ = ys__n47004 & ~new_n23725_;
  assign new_n23931_ = ~new_n23741_ & ~new_n23930_;
  assign new_n23932_ = ~new_n23747_ & ~new_n23931_;
  assign new_n23933_ = new_n23750_ & new_n23932_;
  assign new_n23934_ = ys__n28914 & new_n23753_;
  assign new_n23935_ = ys__n29274 & new_n23755_;
  assign new_n23936_ = ys__n29581 & new_n23757_;
  assign new_n23937_ = ys__n29582 & ~new_n23757_;
  assign new_n23938_ = ~new_n23936_ & ~new_n23937_;
  assign new_n23939_ = ~new_n23755_ & ~new_n23938_;
  assign new_n23940_ = ~new_n23935_ & ~new_n23939_;
  assign new_n23941_ = ~new_n23753_ & ~new_n23940_;
  assign new_n23942_ = ~new_n23934_ & ~new_n23941_;
  assign new_n23943_ = ~new_n23750_ & ~new_n23942_;
  assign ys__n24325 = new_n23933_ | new_n23943_;
  assign new_n23945_ = ys__n47005 & ~new_n23725_;
  assign new_n23946_ = ~new_n23741_ & ~new_n23945_;
  assign new_n23947_ = ~new_n23747_ & ~new_n23946_;
  assign new_n23948_ = new_n23750_ & new_n23947_;
  assign new_n23949_ = ys__n28917 & new_n23753_;
  assign new_n23950_ = ys__n29276 & new_n23755_;
  assign new_n23951_ = ys__n29583 & new_n23757_;
  assign new_n23952_ = ys__n29584 & ~new_n23757_;
  assign new_n23953_ = ~new_n23951_ & ~new_n23952_;
  assign new_n23954_ = ~new_n23755_ & ~new_n23953_;
  assign new_n23955_ = ~new_n23950_ & ~new_n23954_;
  assign new_n23956_ = ~new_n23753_ & ~new_n23955_;
  assign new_n23957_ = ~new_n23949_ & ~new_n23956_;
  assign new_n23958_ = ~new_n23750_ & ~new_n23957_;
  assign ys__n24327 = new_n23948_ | new_n23958_;
  assign new_n23960_ = ys__n47006 & ~new_n23725_;
  assign new_n23961_ = ~new_n23741_ & ~new_n23960_;
  assign new_n23962_ = ~new_n23747_ & ~new_n23961_;
  assign new_n23963_ = new_n23750_ & new_n23962_;
  assign new_n23964_ = ys__n28920 & new_n23753_;
  assign new_n23965_ = ys__n29278 & new_n23755_;
  assign new_n23966_ = ys__n29585 & new_n23757_;
  assign new_n23967_ = ys__n29586 & ~new_n23757_;
  assign new_n23968_ = ~new_n23966_ & ~new_n23967_;
  assign new_n23969_ = ~new_n23755_ & ~new_n23968_;
  assign new_n23970_ = ~new_n23965_ & ~new_n23969_;
  assign new_n23971_ = ~new_n23753_ & ~new_n23970_;
  assign new_n23972_ = ~new_n23964_ & ~new_n23971_;
  assign new_n23973_ = ~new_n23750_ & ~new_n23972_;
  assign ys__n24329 = new_n23963_ | new_n23973_;
  assign new_n23975_ = ys__n47007 & ~new_n23725_;
  assign new_n23976_ = ~new_n23741_ & ~new_n23975_;
  assign new_n23977_ = ~new_n23747_ & ~new_n23976_;
  assign new_n23978_ = new_n23750_ & new_n23977_;
  assign new_n23979_ = ys__n28923 & new_n23753_;
  assign new_n23980_ = ys__n29280 & new_n23755_;
  assign new_n23981_ = ys__n29587 & new_n23757_;
  assign new_n23982_ = ys__n29588 & ~new_n23757_;
  assign new_n23983_ = ~new_n23981_ & ~new_n23982_;
  assign new_n23984_ = ~new_n23755_ & ~new_n23983_;
  assign new_n23985_ = ~new_n23980_ & ~new_n23984_;
  assign new_n23986_ = ~new_n23753_ & ~new_n23985_;
  assign new_n23987_ = ~new_n23979_ & ~new_n23986_;
  assign new_n23988_ = ~new_n23750_ & ~new_n23987_;
  assign ys__n24331 = new_n23978_ | new_n23988_;
  assign new_n23990_ = ys__n47008 & ~new_n23725_;
  assign new_n23991_ = ~new_n23741_ & ~new_n23990_;
  assign new_n23992_ = ~new_n23747_ & ~new_n23991_;
  assign new_n23993_ = new_n23750_ & new_n23992_;
  assign new_n23994_ = ys__n28926 & new_n23753_;
  assign new_n23995_ = ys__n29282 & new_n23755_;
  assign new_n23996_ = ys__n29589 & new_n23757_;
  assign new_n23997_ = ys__n29590 & ~new_n23757_;
  assign new_n23998_ = ~new_n23996_ & ~new_n23997_;
  assign new_n23999_ = ~new_n23755_ & ~new_n23998_;
  assign new_n24000_ = ~new_n23995_ & ~new_n23999_;
  assign new_n24001_ = ~new_n23753_ & ~new_n24000_;
  assign new_n24002_ = ~new_n23994_ & ~new_n24001_;
  assign new_n24003_ = ~new_n23750_ & ~new_n24002_;
  assign ys__n24333 = new_n23993_ | new_n24003_;
  assign new_n24005_ = ys__n47009 & ~new_n23725_;
  assign new_n24006_ = ~new_n23741_ & ~new_n24005_;
  assign new_n24007_ = ~new_n23747_ & ~new_n24006_;
  assign new_n24008_ = new_n23750_ & new_n24007_;
  assign new_n24009_ = ys__n28929 & new_n23753_;
  assign new_n24010_ = ys__n29284 & new_n23755_;
  assign new_n24011_ = ys__n29591 & new_n23757_;
  assign new_n24012_ = ys__n29592 & ~new_n23757_;
  assign new_n24013_ = ~new_n24011_ & ~new_n24012_;
  assign new_n24014_ = ~new_n23755_ & ~new_n24013_;
  assign new_n24015_ = ~new_n24010_ & ~new_n24014_;
  assign new_n24016_ = ~new_n23753_ & ~new_n24015_;
  assign new_n24017_ = ~new_n24009_ & ~new_n24016_;
  assign new_n24018_ = ~new_n23750_ & ~new_n24017_;
  assign ys__n24335 = new_n24008_ | new_n24018_;
  assign new_n24020_ = ~ys__n33471 & new_n13607_;
  assign new_n24021_ = ys__n16 & ys__n1107;
  assign new_n24022_ = new_n15121_ & new_n24021_;
  assign new_n24023_ = ~new_n24020_ & ~new_n24022_;
  assign new_n24024_ = ys__n24320 & new_n24023_;
  assign new_n24025_ = ys__n24337 & new_n24022_;
  assign ys__n24339 = new_n24024_ | new_n24025_;
  assign new_n24027_ = ys__n24323 & new_n24023_;
  assign new_n24028_ = ys__n24340 & new_n24022_;
  assign ys__n24341 = new_n24027_ | new_n24028_;
  assign new_n24030_ = ys__n24325 & new_n24023_;
  assign new_n24031_ = ys__n24342 & new_n24022_;
  assign ys__n24343 = new_n24030_ | new_n24031_;
  assign new_n24033_ = ys__n24327 & new_n24023_;
  assign new_n24034_ = ys__n24344 & new_n24022_;
  assign ys__n24345 = new_n24033_ | new_n24034_;
  assign new_n24036_ = ys__n24329 & new_n24023_;
  assign new_n24037_ = ys__n24346 & new_n24022_;
  assign ys__n24347 = new_n24036_ | new_n24037_;
  assign new_n24039_ = ys__n24331 & new_n24023_;
  assign new_n24040_ = ys__n24348 & new_n24022_;
  assign ys__n24349 = new_n24039_ | new_n24040_;
  assign new_n24042_ = ys__n24333 & new_n24023_;
  assign new_n24043_ = ys__n24350 & new_n24022_;
  assign ys__n24351 = new_n24042_ | new_n24043_;
  assign new_n24045_ = ys__n24335 & new_n24023_;
  assign new_n24046_ = ys__n24352 & new_n24022_;
  assign ys__n24353 = new_n24045_ | new_n24046_;
  assign new_n24048_ = new_n23715_ & ~new_n23719_;
  assign new_n24049_ = ~new_n23718_ & ~new_n23723_;
  assign new_n24050_ = new_n23710_ & new_n24049_;
  assign new_n24051_ = new_n24048_ & new_n24050_;
  assign new_n24052_ = ~new_n24048_ & ~new_n24051_;
  assign new_n24053_ = ys__n47186 & ~new_n24052_;
  assign new_n24054_ = ys__n47194 & new_n24052_;
  assign new_n24055_ = ~new_n24053_ & ~new_n24054_;
  assign new_n24056_ = new_n23720_ & ~new_n23723_;
  assign new_n24057_ = new_n23716_ & new_n24056_;
  assign new_n24058_ = ~new_n23716_ & ~new_n24057_;
  assign new_n24059_ = ~new_n24055_ & ~new_n24058_;
  assign new_n24060_ = new_n23740_ & new_n24058_;
  assign new_n24061_ = ~new_n24059_ & ~new_n24060_;
  assign new_n24062_ = ~new_n23747_ & ~new_n24061_;
  assign new_n24063_ = new_n23750_ & new_n24062_;
  assign new_n24064_ = ys__n28884 & new_n23753_;
  assign new_n24065_ = ys__n29254 & new_n23755_;
  assign new_n24066_ = ys__n29561 & new_n23757_;
  assign new_n24067_ = ys__n29562 & ~new_n23757_;
  assign new_n24068_ = ~new_n24066_ & ~new_n24067_;
  assign new_n24069_ = ~new_n23755_ & ~new_n24068_;
  assign new_n24070_ = ~new_n24065_ & ~new_n24069_;
  assign new_n24071_ = ~new_n23753_ & ~new_n24070_;
  assign new_n24072_ = ~new_n24064_ & ~new_n24071_;
  assign new_n24073_ = ~new_n23750_ & ~new_n24072_;
  assign ys__n24354 = new_n24063_ | new_n24073_;
  assign new_n24075_ = ys__n47187 & ~new_n24052_;
  assign new_n24076_ = ys__n47195 & new_n24052_;
  assign new_n24077_ = ~new_n24075_ & ~new_n24076_;
  assign new_n24078_ = ~new_n24058_ & ~new_n24077_;
  assign new_n24079_ = ~new_n24060_ & ~new_n24078_;
  assign new_n24080_ = ~new_n23747_ & ~new_n24079_;
  assign new_n24081_ = new_n23750_ & new_n24080_;
  assign new_n24082_ = ys__n28887 & new_n23753_;
  assign new_n24083_ = ys__n29256 & new_n23755_;
  assign new_n24084_ = ys__n29563 & new_n23757_;
  assign new_n24085_ = ys__n29564 & ~new_n23757_;
  assign new_n24086_ = ~new_n24084_ & ~new_n24085_;
  assign new_n24087_ = ~new_n23755_ & ~new_n24086_;
  assign new_n24088_ = ~new_n24083_ & ~new_n24087_;
  assign new_n24089_ = ~new_n23753_ & ~new_n24088_;
  assign new_n24090_ = ~new_n24082_ & ~new_n24089_;
  assign new_n24091_ = ~new_n23750_ & ~new_n24090_;
  assign ys__n24357 = new_n24081_ | new_n24091_;
  assign new_n24093_ = ys__n47188 & ~new_n24052_;
  assign new_n24094_ = ys__n47196 & new_n24052_;
  assign new_n24095_ = ~new_n24093_ & ~new_n24094_;
  assign new_n24096_ = ~new_n24058_ & ~new_n24095_;
  assign new_n24097_ = ~new_n24060_ & ~new_n24096_;
  assign new_n24098_ = ~new_n23747_ & ~new_n24097_;
  assign new_n24099_ = new_n23750_ & new_n24098_;
  assign new_n24100_ = ys__n28890 & new_n23753_;
  assign new_n24101_ = ys__n29258 & new_n23755_;
  assign new_n24102_ = ys__n29565 & new_n23757_;
  assign new_n24103_ = ys__n29566 & ~new_n23757_;
  assign new_n24104_ = ~new_n24102_ & ~new_n24103_;
  assign new_n24105_ = ~new_n23755_ & ~new_n24104_;
  assign new_n24106_ = ~new_n24101_ & ~new_n24105_;
  assign new_n24107_ = ~new_n23753_ & ~new_n24106_;
  assign new_n24108_ = ~new_n24100_ & ~new_n24107_;
  assign new_n24109_ = ~new_n23750_ & ~new_n24108_;
  assign ys__n24359 = new_n24099_ | new_n24109_;
  assign new_n24111_ = ys__n47189 & ~new_n24052_;
  assign new_n24112_ = ys__n47197 & new_n24052_;
  assign new_n24113_ = ~new_n24111_ & ~new_n24112_;
  assign new_n24114_ = ~new_n24058_ & ~new_n24113_;
  assign new_n24115_ = ~new_n24060_ & ~new_n24114_;
  assign new_n24116_ = ~new_n23747_ & ~new_n24115_;
  assign new_n24117_ = new_n23750_ & new_n24116_;
  assign new_n24118_ = ys__n28893 & new_n23753_;
  assign new_n24119_ = ys__n29260 & new_n23755_;
  assign new_n24120_ = ys__n29567 & new_n23757_;
  assign new_n24121_ = ys__n29568 & ~new_n23757_;
  assign new_n24122_ = ~new_n24120_ & ~new_n24121_;
  assign new_n24123_ = ~new_n23755_ & ~new_n24122_;
  assign new_n24124_ = ~new_n24119_ & ~new_n24123_;
  assign new_n24125_ = ~new_n23753_ & ~new_n24124_;
  assign new_n24126_ = ~new_n24118_ & ~new_n24125_;
  assign new_n24127_ = ~new_n23750_ & ~new_n24126_;
  assign ys__n24361 = new_n24117_ | new_n24127_;
  assign new_n24129_ = ys__n47190 & ~new_n24052_;
  assign new_n24130_ = ys__n47198 & new_n24052_;
  assign new_n24131_ = ~new_n24129_ & ~new_n24130_;
  assign new_n24132_ = ~new_n24058_ & ~new_n24131_;
  assign new_n24133_ = ~new_n24060_ & ~new_n24132_;
  assign new_n24134_ = ~new_n23747_ & ~new_n24133_;
  assign new_n24135_ = new_n23750_ & new_n24134_;
  assign new_n24136_ = ys__n28896 & new_n23753_;
  assign new_n24137_ = ys__n29262 & new_n23755_;
  assign new_n24138_ = ys__n29569 & new_n23757_;
  assign new_n24139_ = ys__n29570 & ~new_n23757_;
  assign new_n24140_ = ~new_n24138_ & ~new_n24139_;
  assign new_n24141_ = ~new_n23755_ & ~new_n24140_;
  assign new_n24142_ = ~new_n24137_ & ~new_n24141_;
  assign new_n24143_ = ~new_n23753_ & ~new_n24142_;
  assign new_n24144_ = ~new_n24136_ & ~new_n24143_;
  assign new_n24145_ = ~new_n23750_ & ~new_n24144_;
  assign ys__n24363 = new_n24135_ | new_n24145_;
  assign new_n24147_ = ys__n47191 & ~new_n24052_;
  assign new_n24148_ = ys__n47199 & new_n24052_;
  assign new_n24149_ = ~new_n24147_ & ~new_n24148_;
  assign new_n24150_ = ~new_n24058_ & ~new_n24149_;
  assign new_n24151_ = ~new_n24060_ & ~new_n24150_;
  assign new_n24152_ = ~new_n23747_ & ~new_n24151_;
  assign new_n24153_ = new_n23750_ & new_n24152_;
  assign new_n24154_ = ys__n28899 & new_n23753_;
  assign new_n24155_ = ys__n29264 & new_n23755_;
  assign new_n24156_ = ys__n29571 & new_n23757_;
  assign new_n24157_ = ys__n29572 & ~new_n23757_;
  assign new_n24158_ = ~new_n24156_ & ~new_n24157_;
  assign new_n24159_ = ~new_n23755_ & ~new_n24158_;
  assign new_n24160_ = ~new_n24155_ & ~new_n24159_;
  assign new_n24161_ = ~new_n23753_ & ~new_n24160_;
  assign new_n24162_ = ~new_n24154_ & ~new_n24161_;
  assign new_n24163_ = ~new_n23750_ & ~new_n24162_;
  assign ys__n24365 = new_n24153_ | new_n24163_;
  assign new_n24165_ = ys__n47192 & ~new_n24052_;
  assign new_n24166_ = ys__n47200 & new_n24052_;
  assign new_n24167_ = ~new_n24165_ & ~new_n24166_;
  assign new_n24168_ = ~new_n24058_ & ~new_n24167_;
  assign new_n24169_ = ~new_n24060_ & ~new_n24168_;
  assign new_n24170_ = ~new_n23747_ & ~new_n24169_;
  assign new_n24171_ = new_n23750_ & new_n24170_;
  assign new_n24172_ = ys__n28902 & new_n23753_;
  assign new_n24173_ = ys__n29266 & new_n23755_;
  assign new_n24174_ = ys__n29573 & new_n23757_;
  assign new_n24175_ = ys__n29574 & ~new_n23757_;
  assign new_n24176_ = ~new_n24174_ & ~new_n24175_;
  assign new_n24177_ = ~new_n23755_ & ~new_n24176_;
  assign new_n24178_ = ~new_n24173_ & ~new_n24177_;
  assign new_n24179_ = ~new_n23753_ & ~new_n24178_;
  assign new_n24180_ = ~new_n24172_ & ~new_n24179_;
  assign new_n24181_ = ~new_n23750_ & ~new_n24180_;
  assign ys__n24367 = new_n24171_ | new_n24181_;
  assign new_n24183_ = ys__n47193 & ~new_n24052_;
  assign new_n24184_ = ys__n47201 & new_n24052_;
  assign new_n24185_ = ~new_n24183_ & ~new_n24184_;
  assign new_n24186_ = ~new_n24058_ & ~new_n24185_;
  assign new_n24187_ = ~new_n24060_ & ~new_n24186_;
  assign new_n24188_ = ~new_n23747_ & ~new_n24187_;
  assign new_n24189_ = new_n23750_ & new_n24188_;
  assign new_n24190_ = ys__n28905 & new_n23753_;
  assign new_n24191_ = ys__n29268 & new_n23755_;
  assign new_n24192_ = ys__n29575 & new_n23757_;
  assign new_n24193_ = ys__n29576 & ~new_n23757_;
  assign new_n24194_ = ~new_n24192_ & ~new_n24193_;
  assign new_n24195_ = ~new_n23755_ & ~new_n24194_;
  assign new_n24196_ = ~new_n24191_ & ~new_n24195_;
  assign new_n24197_ = ~new_n23753_ & ~new_n24196_;
  assign new_n24198_ = ~new_n24190_ & ~new_n24197_;
  assign new_n24199_ = ~new_n23750_ & ~new_n24198_;
  assign ys__n24369 = new_n24189_ | new_n24199_;
  assign new_n24201_ = ~ys__n33473 & new_n13607_;
  assign new_n24202_ = ys__n14 & ys__n1107;
  assign new_n24203_ = new_n15121_ & new_n24202_;
  assign new_n24204_ = ~new_n24201_ & ~new_n24203_;
  assign new_n24205_ = ys__n24354 & new_n24204_;
  assign new_n24206_ = ys__n24371 & new_n24203_;
  assign ys__n24373 = new_n24205_ | new_n24206_;
  assign new_n24208_ = ys__n24357 & new_n24204_;
  assign new_n24209_ = ys__n24374 & new_n24203_;
  assign ys__n24375 = new_n24208_ | new_n24209_;
  assign new_n24211_ = ys__n24359 & new_n24204_;
  assign new_n24212_ = ys__n24376 & new_n24203_;
  assign ys__n24377 = new_n24211_ | new_n24212_;
  assign new_n24214_ = ys__n24361 & new_n24204_;
  assign new_n24215_ = ys__n24378 & new_n24203_;
  assign ys__n24379 = new_n24214_ | new_n24215_;
  assign new_n24217_ = ys__n24363 & new_n24204_;
  assign new_n24218_ = ys__n24380 & new_n24203_;
  assign ys__n24381 = new_n24217_ | new_n24218_;
  assign new_n24220_ = ys__n24365 & new_n24204_;
  assign new_n24221_ = ys__n24382 & new_n24203_;
  assign ys__n24383 = new_n24220_ | new_n24221_;
  assign new_n24223_ = ys__n24367 & new_n24204_;
  assign new_n24224_ = ys__n24384 & new_n24203_;
  assign ys__n24385 = new_n24223_ | new_n24224_;
  assign new_n24226_ = ys__n24369 & new_n24204_;
  assign new_n24227_ = ys__n24386 & new_n24203_;
  assign ys__n24387 = new_n24226_ | new_n24227_;
  assign new_n24229_ = ~ys__n1154 & ys__n24575;
  assign new_n24230_ = ~ys__n90 & ~ys__n4736;
  assign new_n24231_ = ~ys__n88 & ~ys__n4736;
  assign new_n24232_ = ys__n1154 & ys__n47448;
  assign new_n24233_ = ~new_n24231_ & new_n24232_;
  assign new_n24234_ = ~new_n24230_ & new_n24233_;
  assign new_n24235_ = ~new_n24229_ & ~new_n24234_;
  assign new_n24236_ = new_n23747_ & ~new_n24235_;
  assign new_n24237_ = ys__n46994 & ~new_n24052_;
  assign new_n24238_ = ys__n47002 & new_n24052_;
  assign new_n24239_ = ~new_n24237_ & ~new_n24238_;
  assign new_n24240_ = ~new_n23709_ & ~new_n23714_;
  assign new_n24241_ = new_n23736_ & new_n24240_;
  assign new_n24242_ = new_n24056_ & new_n24241_;
  assign new_n24243_ = ~new_n24240_ & ~new_n24242_;
  assign new_n24244_ = ~new_n24239_ & ~new_n24243_;
  assign new_n24245_ = ~new_n24055_ & new_n24243_;
  assign new_n24246_ = ~new_n24244_ & ~new_n24245_;
  assign new_n24247_ = ~new_n23747_ & ~new_n24246_;
  assign new_n24248_ = ~new_n24236_ & ~new_n24247_;
  assign new_n24249_ = new_n23750_ & ~new_n24248_;
  assign new_n24250_ = ys__n28859 & new_n23753_;
  assign new_n24251_ = ys__n29237 & new_n23755_;
  assign new_n24252_ = ys__n29550 & new_n23757_;
  assign new_n24253_ = ys__n28462 & ~new_n23757_;
  assign new_n24254_ = ~new_n24252_ & ~new_n24253_;
  assign new_n24255_ = ~new_n23755_ & ~new_n24254_;
  assign new_n24256_ = ~new_n24251_ & ~new_n24255_;
  assign new_n24257_ = ~new_n23753_ & ~new_n24256_;
  assign new_n24258_ = ~new_n24250_ & ~new_n24257_;
  assign new_n24259_ = ~new_n23750_ & ~new_n24258_;
  assign ys__n24388 = new_n24249_ | new_n24259_;
  assign new_n24261_ = ys__n46995 & ~new_n24052_;
  assign new_n24262_ = ys__n47003 & new_n24052_;
  assign new_n24263_ = ~new_n24261_ & ~new_n24262_;
  assign new_n24264_ = ~new_n24243_ & ~new_n24263_;
  assign new_n24265_ = ~new_n24077_ & new_n24243_;
  assign new_n24266_ = ~new_n24264_ & ~new_n24265_;
  assign new_n24267_ = ~new_n23747_ & ~new_n24266_;
  assign new_n24268_ = new_n23750_ & new_n24267_;
  assign new_n24269_ = ys__n28863 & new_n23753_;
  assign new_n24270_ = ys__n29240 & new_n23755_;
  assign new_n24271_ = ys__n29552 & new_n23757_;
  assign new_n24272_ = ys__n28464 & ~new_n23757_;
  assign new_n24273_ = ~new_n24271_ & ~new_n24272_;
  assign new_n24274_ = ~new_n23755_ & ~new_n24273_;
  assign new_n24275_ = ~new_n24270_ & ~new_n24274_;
  assign new_n24276_ = ~new_n23753_ & ~new_n24275_;
  assign new_n24277_ = ~new_n24269_ & ~new_n24276_;
  assign new_n24278_ = ~new_n23750_ & ~new_n24277_;
  assign ys__n24392 = new_n24268_ | new_n24278_;
  assign new_n24280_ = ys__n46996 & ~new_n24052_;
  assign new_n24281_ = ys__n47004 & new_n24052_;
  assign new_n24282_ = ~new_n24280_ & ~new_n24281_;
  assign new_n24283_ = ~new_n24243_ & ~new_n24282_;
  assign new_n24284_ = ~new_n24095_ & new_n24243_;
  assign new_n24285_ = ~new_n24283_ & ~new_n24284_;
  assign new_n24286_ = ~new_n23747_ & ~new_n24285_;
  assign new_n24287_ = new_n23750_ & new_n24286_;
  assign new_n24288_ = ys__n28866 & new_n23753_;
  assign new_n24289_ = ys__n29242 & new_n23755_;
  assign new_n24290_ = ys__n29553 & new_n23757_;
  assign new_n24291_ = ys__n28466 & ~new_n23757_;
  assign new_n24292_ = ~new_n24290_ & ~new_n24291_;
  assign new_n24293_ = ~new_n23755_ & ~new_n24292_;
  assign new_n24294_ = ~new_n24289_ & ~new_n24293_;
  assign new_n24295_ = ~new_n23753_ & ~new_n24294_;
  assign new_n24296_ = ~new_n24288_ & ~new_n24295_;
  assign new_n24297_ = ~new_n23750_ & ~new_n24296_;
  assign ys__n24394 = new_n24287_ | new_n24297_;
  assign new_n24299_ = ys__n46997 & ~new_n24052_;
  assign new_n24300_ = ys__n47005 & new_n24052_;
  assign new_n24301_ = ~new_n24299_ & ~new_n24300_;
  assign new_n24302_ = ~new_n24243_ & ~new_n24301_;
  assign new_n24303_ = ~new_n24113_ & new_n24243_;
  assign new_n24304_ = ~new_n24302_ & ~new_n24303_;
  assign new_n24305_ = ~new_n23747_ & ~new_n24304_;
  assign new_n24306_ = new_n23750_ & new_n24305_;
  assign new_n24307_ = ys__n28869 & new_n23753_;
  assign new_n24308_ = ys__n29244 & new_n23755_;
  assign new_n24309_ = ys__n29554 & new_n23757_;
  assign new_n24310_ = ys__n28468 & ~new_n23757_;
  assign new_n24311_ = ~new_n24309_ & ~new_n24310_;
  assign new_n24312_ = ~new_n23755_ & ~new_n24311_;
  assign new_n24313_ = ~new_n24308_ & ~new_n24312_;
  assign new_n24314_ = ~new_n23753_ & ~new_n24313_;
  assign new_n24315_ = ~new_n24307_ & ~new_n24314_;
  assign new_n24316_ = ~new_n23750_ & ~new_n24315_;
  assign ys__n24396 = new_n24306_ | new_n24316_;
  assign new_n24318_ = ys__n46998 & ~new_n24052_;
  assign new_n24319_ = ys__n47006 & new_n24052_;
  assign new_n24320_ = ~new_n24318_ & ~new_n24319_;
  assign new_n24321_ = ~new_n24243_ & ~new_n24320_;
  assign new_n24322_ = ~new_n24131_ & new_n24243_;
  assign new_n24323_ = ~new_n24321_ & ~new_n24322_;
  assign new_n24324_ = ~new_n23747_ & ~new_n24323_;
  assign new_n24325_ = new_n23750_ & new_n24324_;
  assign new_n24326_ = ys__n28872 & new_n23753_;
  assign new_n24327_ = ys__n29246 & new_n23755_;
  assign new_n24328_ = ys__n29555 & new_n23757_;
  assign new_n24329_ = ys__n28470 & ~new_n23757_;
  assign new_n24330_ = ~new_n24328_ & ~new_n24329_;
  assign new_n24331_ = ~new_n23755_ & ~new_n24330_;
  assign new_n24332_ = ~new_n24327_ & ~new_n24331_;
  assign new_n24333_ = ~new_n23753_ & ~new_n24332_;
  assign new_n24334_ = ~new_n24326_ & ~new_n24333_;
  assign new_n24335_ = ~new_n23750_ & ~new_n24334_;
  assign ys__n24398 = new_n24325_ | new_n24335_;
  assign new_n24337_ = ys__n46999 & ~new_n24052_;
  assign new_n24338_ = ys__n47007 & new_n24052_;
  assign new_n24339_ = ~new_n24337_ & ~new_n24338_;
  assign new_n24340_ = ~new_n24243_ & ~new_n24339_;
  assign new_n24341_ = ~new_n24149_ & new_n24243_;
  assign new_n24342_ = ~new_n24340_ & ~new_n24341_;
  assign new_n24343_ = ~new_n23747_ & ~new_n24342_;
  assign new_n24344_ = new_n23750_ & new_n24343_;
  assign new_n24345_ = ys__n28875 & new_n23753_;
  assign new_n24346_ = ys__n29248 & new_n23755_;
  assign new_n24347_ = ys__n29556 & new_n23757_;
  assign new_n24348_ = ys__n28472 & ~new_n23757_;
  assign new_n24349_ = ~new_n24347_ & ~new_n24348_;
  assign new_n24350_ = ~new_n23755_ & ~new_n24349_;
  assign new_n24351_ = ~new_n24346_ & ~new_n24350_;
  assign new_n24352_ = ~new_n23753_ & ~new_n24351_;
  assign new_n24353_ = ~new_n24345_ & ~new_n24352_;
  assign new_n24354_ = ~new_n23750_ & ~new_n24353_;
  assign ys__n24400 = new_n24344_ | new_n24354_;
  assign new_n24356_ = ys__n47000 & ~new_n24052_;
  assign new_n24357_ = ys__n47008 & new_n24052_;
  assign new_n24358_ = ~new_n24356_ & ~new_n24357_;
  assign new_n24359_ = ~new_n24243_ & ~new_n24358_;
  assign new_n24360_ = ~new_n24167_ & new_n24243_;
  assign new_n24361_ = ~new_n24359_ & ~new_n24360_;
  assign new_n24362_ = ~new_n23747_ & ~new_n24361_;
  assign new_n24363_ = new_n23750_ & new_n24362_;
  assign new_n24364_ = ys__n28878 & new_n23753_;
  assign new_n24365_ = ys__n29250 & new_n23755_;
  assign new_n24366_ = ys__n29557 & new_n23757_;
  assign new_n24367_ = ys__n29558 & ~new_n23757_;
  assign new_n24368_ = ~new_n24366_ & ~new_n24367_;
  assign new_n24369_ = ~new_n23755_ & ~new_n24368_;
  assign new_n24370_ = ~new_n24365_ & ~new_n24369_;
  assign new_n24371_ = ~new_n23753_ & ~new_n24370_;
  assign new_n24372_ = ~new_n24364_ & ~new_n24371_;
  assign new_n24373_ = ~new_n23750_ & ~new_n24372_;
  assign ys__n24402 = new_n24363_ | new_n24373_;
  assign new_n24375_ = ys__n47001 & ~new_n24052_;
  assign new_n24376_ = ys__n47009 & new_n24052_;
  assign new_n24377_ = ~new_n24375_ & ~new_n24376_;
  assign new_n24378_ = ~new_n24243_ & ~new_n24377_;
  assign new_n24379_ = ~new_n24185_ & new_n24243_;
  assign new_n24380_ = ~new_n24378_ & ~new_n24379_;
  assign new_n24381_ = ~new_n23747_ & ~new_n24380_;
  assign new_n24382_ = new_n23750_ & new_n24381_;
  assign new_n24383_ = ys__n28881 & new_n23753_;
  assign new_n24384_ = ys__n29252 & new_n23755_;
  assign new_n24385_ = ys__n29559 & new_n23757_;
  assign new_n24386_ = ys__n29560 & ~new_n23757_;
  assign new_n24387_ = ~new_n24385_ & ~new_n24386_;
  assign new_n24388_ = ~new_n23755_ & ~new_n24387_;
  assign new_n24389_ = ~new_n24384_ & ~new_n24388_;
  assign new_n24390_ = ~new_n23753_ & ~new_n24389_;
  assign new_n24391_ = ~new_n24383_ & ~new_n24390_;
  assign new_n24392_ = ~new_n23750_ & ~new_n24391_;
  assign ys__n24404 = new_n24382_ | new_n24392_;
  assign new_n24394_ = ~ys__n33475 & new_n13607_;
  assign new_n24395_ = ys__n24388 & ~new_n24394_;
  assign new_n24396_ = ys__n24389 & new_n24394_;
  assign new_n24397_ = ~new_n24395_ & ~new_n24396_;
  assign new_n24398_ = ys__n1107 & ys__n4688;
  assign new_n24399_ = new_n15121_ & new_n24398_;
  assign new_n24400_ = ~new_n24397_ & ~new_n24399_;
  assign new_n24401_ = ys__n24406 & new_n24399_;
  assign ys__n24408 = new_n24400_ | new_n24401_;
  assign new_n24403_ = ~new_n24394_ & ~new_n24399_;
  assign new_n24404_ = ys__n24392 & new_n24403_;
  assign new_n24405_ = ys__n24409 & new_n24399_;
  assign ys__n24410 = new_n24404_ | new_n24405_;
  assign new_n24407_ = ys__n24394 & new_n24403_;
  assign new_n24408_ = ys__n24411 & new_n24399_;
  assign ys__n24412 = new_n24407_ | new_n24408_;
  assign new_n24410_ = ys__n24396 & new_n24403_;
  assign new_n24411_ = ys__n24413 & new_n24399_;
  assign ys__n24414 = new_n24410_ | new_n24411_;
  assign new_n24413_ = ys__n24398 & new_n24403_;
  assign new_n24414_ = ys__n24415 & new_n24399_;
  assign ys__n24416 = new_n24413_ | new_n24414_;
  assign new_n24416_ = ys__n24400 & new_n24403_;
  assign new_n24417_ = ys__n24417 & new_n24399_;
  assign ys__n24418 = new_n24416_ | new_n24417_;
  assign new_n24419_ = ys__n24402 & new_n24403_;
  assign new_n24420_ = ys__n24419 & new_n24399_;
  assign ys__n24420 = new_n24419_ | new_n24420_;
  assign new_n24422_ = ys__n24404 & new_n24403_;
  assign new_n24423_ = ys__n24421 & new_n24399_;
  assign ys__n24422 = new_n24422_ | new_n24423_;
  assign new_n24425_ = ~ys__n1116 & new_n13610_;
  assign new_n24426_ = ys__n24279 & new_n24425_;
  assign new_n24427_ = ys__n452 & ~new_n24425_;
  assign new_n24428_ = ~new_n24426_ & ~new_n24427_;
  assign new_n24429_ = ~ys__n1109 & ~ys__n1116;
  assign new_n24430_ = ~ys__n1117 & new_n24429_;
  assign new_n24431_ = ~new_n24428_ & new_n24430_;
  assign new_n24432_ = ys__n24427 & ~new_n24430_;
  assign new_n24433_ = ~new_n24431_ & ~new_n24432_;
  assign new_n24434_ = ys__n33495 & new_n23580_;
  assign new_n24435_ = ~ys__n24258 & ~new_n23649_;
  assign new_n24436_ = ~new_n24434_ & new_n24435_;
  assign new_n24437_ = ~new_n24433_ & ~new_n24436_;
  assign new_n24438_ = ys__n20008 & new_n24436_;
  assign ys__n24425 = new_n24437_ | new_n24438_;
  assign new_n24440_ = ys__n1094 & ~ys__n1147;
  assign new_n24441_ = ~ys__n24433 & ys__n24434;
  assign new_n24442_ = new_n24440_ & new_n24441_;
  assign new_n24443_ = ys__n1147 & ~ys__n18019;
  assign new_n24444_ = ~new_n24442_ & ~new_n24443_;
  assign new_n24445_ = ~ys__n140 & ~new_n24444_;
  assign ys__n24430 = ys__n140 | new_n24445_;
  assign new_n24447_ = ~ys__n1094 & ~ys__n24433;
  assign new_n24448_ = ys__n24434 & new_n24447_;
  assign ys__n24436 = ys__n24433 | new_n24448_;
  assign new_n24450_ = ys__n454 & ys__n712;
  assign ys__n24470 = ys__n24519 & new_n24450_;
  assign new_n24452_ = ~ys__n1098 & ~ys__n1099;
  assign new_n24453_ = ys__n1107 & new_n24452_;
  assign new_n24454_ = ~ys__n24470 & new_n24453_;
  assign new_n24455_ = ys__n1099 & ~ys__n24506;
  assign new_n24456_ = ys__n33488 & new_n24455_;
  assign ys__n24440 = new_n24454_ | new_n24456_;
  assign new_n24458_ = ys__n1098 & ~ys__n1099;
  assign new_n24459_ = ~ys__n24470 & new_n24458_;
  assign new_n24460_ = ~ys__n33488 & new_n24455_;
  assign ys__n24445 = new_n24459_ | new_n24460_;
  assign new_n24462_ = ~ys__n1107 & ~ys__n1110;
  assign new_n24463_ = new_n23749_ & new_n24462_;
  assign new_n24464_ = new_n24452_ & new_n24463_;
  assign new_n24465_ = ~ys__n1129 & ~ys__n24461;
  assign new_n24466_ = ~ys__n24463 & new_n24465_;
  assign new_n24467_ = new_n13634_ & new_n23570_;
  assign new_n24468_ = new_n24466_ & new_n24467_;
  assign new_n24469_ = new_n24464_ & new_n24468_;
  assign new_n24470_ = new_n17724_ & new_n24469_;
  assign new_n24471_ = ys__n33493 & new_n17716_;
  assign new_n24472_ = ys__n1106 & ~ys__n33491;
  assign new_n24473_ = new_n24471_ & new_n24472_;
  assign new_n24474_ = ~ys__n4566 & new_n24473_;
  assign new_n24475_ = ys__n4696 & new_n24474_;
  assign new_n24476_ = ~new_n24470_ & ~new_n24475_;
  assign ys__n24447 = ~ys__n1094 & ~new_n24476_;
  assign new_n24478_ = new_n13609_ & new_n13622_;
  assign new_n24479_ = new_n24467_ & new_n24478_;
  assign new_n24480_ = ~ys__n24483 & ys__n24485;
  assign new_n24481_ = ~ys__n24567 & new_n24480_;
  assign new_n24482_ = ~ys__n24463 & ~ys__n24464;
  assign new_n24483_ = new_n24465_ & new_n24482_;
  assign new_n24484_ = new_n24481_ & new_n24483_;
  assign new_n24485_ = new_n24479_ & new_n24484_;
  assign new_n24486_ = ys__n1098 & ys__n24470;
  assign new_n24487_ = ~new_n24485_ & ~new_n24486_;
  assign new_n24488_ = ~ys__n1099 & new_n13617_;
  assign new_n24489_ = ~new_n24487_ & new_n24488_;
  assign new_n24490_ = ys__n1094 & ys__n24433;
  assign ys__n24466 = new_n24489_ | new_n24490_;
  assign new_n24492_ = ys__n1119 & ~ys__n1129;
  assign new_n24493_ = new_n24462_ & new_n24492_;
  assign new_n24494_ = new_n23749_ & new_n24452_;
  assign new_n24495_ = new_n24493_ & new_n24494_;
  assign new_n24496_ = new_n17716_ & new_n24495_;
  assign new_n24497_ = ~new_n23580_ & new_n24496_;
  assign new_n24498_ = ys__n33481 & ys__n33497;
  assign new_n24499_ = new_n24472_ & new_n24498_;
  assign new_n24500_ = new_n17716_ & new_n24499_;
  assign new_n24501_ = ~new_n23580_ & new_n24500_;
  assign new_n24502_ = ~ys__n4566 & new_n24501_;
  assign new_n24503_ = ~ys__n4696 & new_n24502_;
  assign ys__n24488 = new_n24497_ | new_n24503_;
  assign new_n24505_ = ~ys__n1094 & ys__n1106;
  assign new_n24506_ = ys__n33499 & new_n23621_;
  assign new_n24507_ = new_n24505_ & new_n24506_;
  assign new_n24508_ = new_n17716_ & new_n24507_;
  assign new_n24509_ = ~ys__n4566 & new_n24508_;
  assign new_n24510_ = ys__n1094 & ~ys__n24433;
  assign ys__n24499 = new_n24509_ | new_n24510_;
  assign new_n24512_ = ~ys__n140 & ys__n1119;
  assign new_n24513_ = ~ys__n1129 & new_n24512_;
  assign new_n24514_ = new_n23581_ & new_n24513_;
  assign new_n24515_ = ys__n1129 & ~ys__n24470;
  assign ys__n24522 = new_n24514_ | new_n24515_;
  assign new_n24517_ = ~ys__n24461 & ys__n24463;
  assign new_n24518_ = ~ys__n24519 & new_n24517_;
  assign ys__n24532 = ys__n24461 | new_n24518_;
  assign new_n24520_ = ~ys__n1129 & new_n24462_;
  assign new_n24521_ = new_n24494_ & new_n24520_;
  assign new_n24522_ = new_n17717_ & new_n24521_;
  assign new_n24523_ = ~ys__n4696 & new_n24474_;
  assign new_n24524_ = ~new_n24522_ & ~new_n24523_;
  assign ys__n24541 = ~ys__n1094 & ~new_n24524_;
  assign ys__n38677 = ys__n24485 & ys__n24567;
  assign new_n24527_ = new_n24494_ & ys__n38677;
  assign new_n24528_ = ~ys__n24483 & new_n24482_;
  assign new_n24529_ = new_n13634_ & new_n24465_;
  assign new_n24530_ = new_n23570_ & new_n24462_;
  assign new_n24531_ = new_n24529_ & new_n24530_;
  assign new_n24532_ = new_n24528_ & new_n24531_;
  assign new_n24533_ = new_n24527_ & new_n24532_;
  assign new_n24534_ = ys__n1106 & ys__n24567;
  assign new_n24535_ = ~ys__n33499 & new_n23621_;
  assign new_n24536_ = new_n24534_ & new_n24535_;
  assign new_n24537_ = new_n17716_ & new_n24536_;
  assign new_n24538_ = ~new_n23601_ & new_n24537_;
  assign new_n24539_ = ~ys__n4566 & new_n24538_;
  assign ys__n24552 = new_n24533_ | new_n24539_;
  assign new_n24541_ = ~ys__n18227 & ys__n24260;
  assign new_n24542_ = ys__n18150 & ~ys__n4566;
  assign new_n24543_ = ys__n18227 & new_n24542_;
  assign ys__n24570 = new_n24541_ | new_n24543_;
  assign new_n24545_ = new_n17684_ & ys__n33521;
  assign new_n24546_ = ys__n18143 & ~ys__n4566;
  assign new_n24547_ = ys__n18227 & new_n24546_;
  assign ys__n24573 = new_n24545_ | new_n24547_;
  assign new_n24549_ = ~ys__n14 & ~ys__n4688;
  assign new_n24550_ = ys__n30011 & ~new_n24549_;
  assign new_n24551_ = ys__n30044 & new_n24549_;
  assign new_n24552_ = ~new_n24550_ & ~new_n24551_;
  assign new_n24553_ = ~ys__n16 & ~ys__n4688;
  assign new_n24554_ = ~new_n24552_ & ~new_n24553_;
  assign new_n24555_ = ys__n30028 & ~new_n24549_;
  assign new_n24556_ = ys__n30060 & new_n24549_;
  assign new_n24557_ = ~new_n24555_ & ~new_n24556_;
  assign new_n24558_ = new_n24553_ & ~new_n24557_;
  assign new_n24559_ = ~new_n24554_ & ~new_n24558_;
  assign new_n24560_ = ys__n33552 & ys__n38680;
  assign new_n24561_ = new_n23617_ & new_n24560_;
  assign new_n24562_ = ~new_n24559_ & ~new_n24561_;
  assign new_n24563_ = ys__n30011 & new_n24561_;
  assign new_n24564_ = ~new_n24562_ & ~new_n24563_;
  assign new_n24565_ = new_n13634_ & ~new_n24561_;
  assign new_n24566_ = ~new_n24564_ & ~new_n24565_;
  assign new_n24567_ = ys__n24389 & new_n24565_;
  assign new_n24568_ = ~new_n24566_ & ~new_n24567_;
  assign new_n24569_ = ~ys__n4176 & ~ys__n4696;
  assign new_n24570_ = new_n11743_ & ~new_n24569_;
  assign new_n24571_ = ys__n33497 & ys__n1088;
  assign new_n24572_ = ~ys__n1117 & ~ys__n1119;
  assign new_n24573_ = new_n15125_ & new_n24572_;
  assign new_n24574_ = ~new_n24561_ & new_n24573_;
  assign new_n24575_ = ~new_n24571_ & new_n24574_;
  assign new_n24576_ = ~new_n24570_ & ~new_n24575_;
  assign new_n24577_ = ~new_n24568_ & new_n24576_;
  assign new_n24578_ = ~new_n24258_ & ~new_n24576_;
  assign new_n24579_ = ~new_n24577_ & ~new_n24578_;
  assign new_n24580_ = ys__n1151 & ~ys__n33522;
  assign new_n24581_ = new_n17697_ & new_n24580_;
  assign new_n24582_ = ~new_n24579_ & ~new_n24581_;
  assign new_n24583_ = ys__n24575 & new_n24581_;
  assign ys__n24577 = new_n24582_ | new_n24583_;
  assign new_n24585_ = ys__n1151 & ys__n18143;
  assign new_n24586_ = new_n17689_ & new_n24585_;
  assign new_n24587_ = new_n17689_ & new_n17692_;
  assign new_n24588_ = new_n13651_ & ~ys__n18137;
  assign new_n24589_ = ~ys__n18227 & ~new_n24588_;
  assign new_n24590_ = ~new_n24587_ & new_n24589_;
  assign new_n24591_ = ~new_n24586_ & new_n24590_;
  assign new_n24592_ = ys__n24578 & ~new_n24591_;
  assign new_n24593_ = ys__n20008 & new_n24591_;
  assign ys__n24579 = new_n24592_ | new_n24593_;
  assign new_n24595_ = ~ys__n140 & ys__n1151;
  assign ys__n24581 = ~new_n17723_ & new_n24595_;
  assign new_n24597_ = ~ys__n1157 & new_n13651_;
  assign ys__n38801 = ys__n24590 & ys__n24591;
  assign new_n24599_ = ~ys__n18137 & ys__n38801;
  assign new_n24600_ = new_n24597_ & new_n24599_;
  assign new_n24601_ = ys__n1151 & new_n17727_;
  assign ys__n24585 = new_n24600_ | new_n24601_;
  assign new_n24603_ = ys__n1154 & ~ys__n18137;
  assign new_n24604_ = ~new_n17682_ & new_n24603_;
  assign new_n24605_ = ys__n1151 & ~new_n17726_;
  assign new_n24606_ = ~new_n24604_ & ~new_n24605_;
  assign ys__n24604 = ~ys__n140 & ~new_n24606_;
  assign ys__n24713 = new_n13261_ & ys__n19183;
  assign ys__n24714 = ~new_n13261_ & new_n18052_;
  assign new_n24610_ = ~ys__n44906 & ~ys__n44907;
  assign new_n24611_ = ~ys__n44908 & new_n24610_;
  assign new_n24612_ = ys__n30819 & ys__n31031;
  assign new_n24613_ = ~new_n24611_ & new_n24612_;
  assign new_n24614_ = ~ys__n2779 & ~new_n24613_;
  assign new_n24615_ = ys__n31031 & ys__n47026;
  assign new_n24616_ = new_n24614_ & new_n24615_;
  assign new_n24617_ = ys__n34762 & ys__n34764;
  assign new_n24618_ = ys__n34766 & new_n24617_;
  assign new_n24619_ = ~ys__n34762 & ~ys__n34764;
  assign new_n24620_ = ys__n34766 & new_n24619_;
  assign new_n24621_ = ~new_n24618_ & ~new_n24620_;
  assign new_n24622_ = ~ys__n34762 & ys__n34764;
  assign new_n24623_ = ~ys__n34766 & new_n24622_;
  assign new_n24624_ = ys__n34762 & ~ys__n34764;
  assign new_n24625_ = ~ys__n34766 & new_n24624_;
  assign new_n24626_ = ~new_n24623_ & ~new_n24625_;
  assign new_n24627_ = new_n24621_ & new_n24626_;
  assign new_n24628_ = ys__n34770 & ys__n34772;
  assign new_n24629_ = ys__n34768 & ys__n34770;
  assign new_n24630_ = ys__n34768 & ys__n34772;
  assign new_n24631_ = ~new_n24629_ & ~new_n24630_;
  assign new_n24632_ = ~new_n24628_ & new_n24631_;
  assign new_n24633_ = new_n24627_ & ~new_n24632_;
  assign new_n24634_ = ~new_n24627_ & new_n24632_;
  assign new_n24635_ = ~new_n24633_ & ~new_n24634_;
  assign new_n24636_ = ys__n34852 & ys__n34854;
  assign new_n24637_ = ys__n34856 & new_n24636_;
  assign new_n24638_ = ~ys__n34852 & ~ys__n34854;
  assign new_n24639_ = ys__n34856 & new_n24638_;
  assign new_n24640_ = ~new_n24637_ & ~new_n24639_;
  assign new_n24641_ = ~ys__n34852 & ys__n34854;
  assign new_n24642_ = ~ys__n34856 & new_n24641_;
  assign new_n24643_ = ys__n34852 & ~ys__n34854;
  assign new_n24644_ = ~ys__n34856 & new_n24643_;
  assign new_n24645_ = ~new_n24642_ & ~new_n24644_;
  assign new_n24646_ = new_n24640_ & new_n24645_;
  assign new_n24647_ = ys__n34860 & ys__n34862;
  assign new_n24648_ = ys__n34858 & ys__n34860;
  assign new_n24649_ = ys__n34858 & ys__n34862;
  assign new_n24650_ = ~new_n24648_ & ~new_n24649_;
  assign new_n24651_ = ~new_n24647_ & new_n24650_;
  assign new_n24652_ = ~new_n24646_ & ~new_n24651_;
  assign new_n24653_ = new_n24646_ & ~new_n24651_;
  assign new_n24654_ = ~new_n24646_ & new_n24651_;
  assign new_n24655_ = ~new_n24653_ & ~new_n24654_;
  assign new_n24656_ = ys__n34862 & new_n24648_;
  assign new_n24657_ = ~ys__n34858 & ~ys__n34860;
  assign new_n24658_ = ys__n34862 & new_n24657_;
  assign new_n24659_ = ~new_n24656_ & ~new_n24658_;
  assign new_n24660_ = ~ys__n34858 & ys__n34860;
  assign new_n24661_ = ~ys__n34862 & new_n24660_;
  assign new_n24662_ = ys__n34858 & ~ys__n34860;
  assign new_n24663_ = ~ys__n34862 & new_n24662_;
  assign new_n24664_ = ~new_n24661_ & ~new_n24663_;
  assign new_n24665_ = new_n24659_ & new_n24664_;
  assign new_n24666_ = ys__n34866 & ys__n34868;
  assign new_n24667_ = ys__n34864 & ys__n34866;
  assign new_n24668_ = ys__n34864 & ys__n34868;
  assign new_n24669_ = ~new_n24667_ & ~new_n24668_;
  assign new_n24670_ = ~new_n24666_ & new_n24669_;
  assign new_n24671_ = ~new_n24665_ & ~new_n24670_;
  assign new_n24672_ = ~new_n24655_ & new_n24671_;
  assign new_n24673_ = ~new_n24652_ & ~new_n24672_;
  assign new_n24674_ = ys__n34840 & ys__n34842;
  assign new_n24675_ = ys__n34844 & new_n24674_;
  assign new_n24676_ = ~ys__n34840 & ~ys__n34842;
  assign new_n24677_ = ys__n34844 & new_n24676_;
  assign new_n24678_ = ~new_n24675_ & ~new_n24677_;
  assign new_n24679_ = ~ys__n34840 & ys__n34842;
  assign new_n24680_ = ~ys__n34844 & new_n24679_;
  assign new_n24681_ = ys__n34840 & ~ys__n34842;
  assign new_n24682_ = ~ys__n34844 & new_n24681_;
  assign new_n24683_ = ~new_n24680_ & ~new_n24682_;
  assign new_n24684_ = new_n24678_ & new_n24683_;
  assign new_n24685_ = ys__n34848 & ys__n34850;
  assign new_n24686_ = ys__n34846 & ys__n34848;
  assign new_n24687_ = ys__n34846 & ys__n34850;
  assign new_n24688_ = ~new_n24686_ & ~new_n24687_;
  assign new_n24689_ = ~new_n24685_ & new_n24688_;
  assign new_n24690_ = new_n24684_ & ~new_n24689_;
  assign new_n24691_ = ~new_n24684_ & new_n24689_;
  assign new_n24692_ = ~new_n24690_ & ~new_n24691_;
  assign new_n24693_ = ys__n34850 & new_n24686_;
  assign new_n24694_ = ~ys__n34846 & ~ys__n34848;
  assign new_n24695_ = ys__n34850 & new_n24694_;
  assign new_n24696_ = ~new_n24693_ & ~new_n24695_;
  assign new_n24697_ = ~ys__n34846 & ys__n34848;
  assign new_n24698_ = ~ys__n34850 & new_n24697_;
  assign new_n24699_ = ys__n34846 & ~ys__n34848;
  assign new_n24700_ = ~ys__n34850 & new_n24699_;
  assign new_n24701_ = ~new_n24698_ & ~new_n24700_;
  assign new_n24702_ = new_n24696_ & new_n24701_;
  assign new_n24703_ = ys__n34854 & ys__n34856;
  assign new_n24704_ = ys__n34852 & ys__n34856;
  assign new_n24705_ = ~new_n24636_ & ~new_n24704_;
  assign new_n24706_ = ~new_n24703_ & new_n24705_;
  assign new_n24707_ = new_n24702_ & ~new_n24706_;
  assign new_n24708_ = ~new_n24702_ & new_n24706_;
  assign new_n24709_ = ~new_n24707_ & ~new_n24708_;
  assign new_n24710_ = ~new_n24692_ & ~new_n24709_;
  assign new_n24711_ = ~new_n24673_ & new_n24710_;
  assign new_n24712_ = ~new_n24684_ & ~new_n24689_;
  assign new_n24713_ = ~new_n24702_ & ~new_n24706_;
  assign new_n24714_ = ~new_n24692_ & new_n24713_;
  assign new_n24715_ = ~new_n24712_ & ~new_n24714_;
  assign new_n24716_ = ~new_n24711_ & new_n24715_;
  assign new_n24717_ = ys__n34816 & ys__n34818;
  assign new_n24718_ = ys__n34820 & new_n24717_;
  assign new_n24719_ = ~ys__n34816 & ~ys__n34818;
  assign new_n24720_ = ys__n34820 & new_n24719_;
  assign new_n24721_ = ~new_n24718_ & ~new_n24720_;
  assign new_n24722_ = ~ys__n34816 & ys__n34818;
  assign new_n24723_ = ~ys__n34820 & new_n24722_;
  assign new_n24724_ = ys__n34816 & ~ys__n34818;
  assign new_n24725_ = ~ys__n34820 & new_n24724_;
  assign new_n24726_ = ~new_n24723_ & ~new_n24725_;
  assign new_n24727_ = new_n24721_ & new_n24726_;
  assign new_n24728_ = ys__n34824 & ys__n34826;
  assign new_n24729_ = ys__n34822 & ys__n34824;
  assign new_n24730_ = ys__n34822 & ys__n34826;
  assign new_n24731_ = ~new_n24729_ & ~new_n24730_;
  assign new_n24732_ = ~new_n24728_ & new_n24731_;
  assign new_n24733_ = new_n24727_ & ~new_n24732_;
  assign new_n24734_ = ~new_n24727_ & new_n24732_;
  assign new_n24735_ = ~new_n24733_ & ~new_n24734_;
  assign new_n24736_ = ys__n34826 & new_n24729_;
  assign new_n24737_ = ~ys__n34822 & ~ys__n34824;
  assign new_n24738_ = ys__n34826 & new_n24737_;
  assign new_n24739_ = ~new_n24736_ & ~new_n24738_;
  assign new_n24740_ = ~ys__n34822 & ys__n34824;
  assign new_n24741_ = ~ys__n34826 & new_n24740_;
  assign new_n24742_ = ys__n34822 & ~ys__n34824;
  assign new_n24743_ = ~ys__n34826 & new_n24742_;
  assign new_n24744_ = ~new_n24741_ & ~new_n24743_;
  assign new_n24745_ = new_n24739_ & new_n24744_;
  assign new_n24746_ = ys__n34830 & ys__n34832;
  assign new_n24747_ = ys__n34828 & ys__n34830;
  assign new_n24748_ = ys__n34828 & ys__n34832;
  assign new_n24749_ = ~new_n24747_ & ~new_n24748_;
  assign new_n24750_ = ~new_n24746_ & new_n24749_;
  assign new_n24751_ = new_n24745_ & ~new_n24750_;
  assign new_n24752_ = ~new_n24745_ & new_n24750_;
  assign new_n24753_ = ~new_n24751_ & ~new_n24752_;
  assign new_n24754_ = ~new_n24735_ & ~new_n24753_;
  assign new_n24755_ = ys__n34832 & new_n24747_;
  assign new_n24756_ = ~ys__n34828 & ~ys__n34830;
  assign new_n24757_ = ys__n34832 & new_n24756_;
  assign new_n24758_ = ~new_n24755_ & ~new_n24757_;
  assign new_n24759_ = ~ys__n34828 & ys__n34830;
  assign new_n24760_ = ~ys__n34832 & new_n24759_;
  assign new_n24761_ = ys__n34828 & ~ys__n34830;
  assign new_n24762_ = ~ys__n34832 & new_n24761_;
  assign new_n24763_ = ~new_n24760_ & ~new_n24762_;
  assign new_n24764_ = new_n24758_ & new_n24763_;
  assign new_n24765_ = ys__n34836 & ys__n34838;
  assign new_n24766_ = ys__n34834 & ys__n34836;
  assign new_n24767_ = ys__n34834 & ys__n34838;
  assign new_n24768_ = ~new_n24766_ & ~new_n24767_;
  assign new_n24769_ = ~new_n24765_ & new_n24768_;
  assign new_n24770_ = new_n24764_ & ~new_n24769_;
  assign new_n24771_ = ~new_n24764_ & new_n24769_;
  assign new_n24772_ = ~new_n24770_ & ~new_n24771_;
  assign new_n24773_ = ys__n34838 & new_n24766_;
  assign new_n24774_ = ~ys__n34834 & ~ys__n34836;
  assign new_n24775_ = ys__n34838 & new_n24774_;
  assign new_n24776_ = ~new_n24773_ & ~new_n24775_;
  assign new_n24777_ = ~ys__n34834 & ys__n34836;
  assign new_n24778_ = ~ys__n34838 & new_n24777_;
  assign new_n24779_ = ys__n34834 & ~ys__n34836;
  assign new_n24780_ = ~ys__n34838 & new_n24779_;
  assign new_n24781_ = ~new_n24778_ & ~new_n24780_;
  assign new_n24782_ = new_n24776_ & new_n24781_;
  assign new_n24783_ = ys__n34842 & ys__n34844;
  assign new_n24784_ = ys__n34840 & ys__n34844;
  assign new_n24785_ = ~new_n24674_ & ~new_n24784_;
  assign new_n24786_ = ~new_n24783_ & new_n24785_;
  assign new_n24787_ = new_n24782_ & ~new_n24786_;
  assign new_n24788_ = ~new_n24782_ & new_n24786_;
  assign new_n24789_ = ~new_n24787_ & ~new_n24788_;
  assign new_n24790_ = ~new_n24772_ & ~new_n24789_;
  assign new_n24791_ = new_n24754_ & new_n24790_;
  assign new_n24792_ = ~new_n24716_ & new_n24791_;
  assign new_n24793_ = ~new_n24764_ & ~new_n24769_;
  assign new_n24794_ = ~new_n24782_ & ~new_n24786_;
  assign new_n24795_ = ~new_n24772_ & new_n24794_;
  assign new_n24796_ = ~new_n24793_ & ~new_n24795_;
  assign new_n24797_ = new_n24754_ & ~new_n24796_;
  assign new_n24798_ = ~new_n24727_ & ~new_n24732_;
  assign new_n24799_ = ~new_n24745_ & ~new_n24750_;
  assign new_n24800_ = ~new_n24735_ & new_n24799_;
  assign new_n24801_ = ~new_n24798_ & ~new_n24800_;
  assign new_n24802_ = ~new_n24797_ & new_n24801_;
  assign new_n24803_ = ~new_n24792_ & new_n24802_;
  assign new_n24804_ = ys__n34772 & new_n24629_;
  assign new_n24805_ = ~ys__n34768 & ~ys__n34770;
  assign new_n24806_ = ys__n34772 & new_n24805_;
  assign new_n24807_ = ~new_n24804_ & ~new_n24806_;
  assign new_n24808_ = ~ys__n34768 & ys__n34770;
  assign new_n24809_ = ~ys__n34772 & new_n24808_;
  assign new_n24810_ = ys__n34768 & ~ys__n34770;
  assign new_n24811_ = ~ys__n34772 & new_n24810_;
  assign new_n24812_ = ~new_n24809_ & ~new_n24811_;
  assign new_n24813_ = new_n24807_ & new_n24812_;
  assign new_n24814_ = ys__n34776 & ys__n34778;
  assign new_n24815_ = ys__n34774 & ys__n34776;
  assign new_n24816_ = ys__n34774 & ys__n34778;
  assign new_n24817_ = ~new_n24815_ & ~new_n24816_;
  assign new_n24818_ = ~new_n24814_ & new_n24817_;
  assign new_n24819_ = new_n24813_ & ~new_n24818_;
  assign new_n24820_ = ~new_n24813_ & new_n24818_;
  assign new_n24821_ = ~new_n24819_ & ~new_n24820_;
  assign new_n24822_ = ys__n34778 & new_n24815_;
  assign new_n24823_ = ~ys__n34774 & ~ys__n34776;
  assign new_n24824_ = ys__n34778 & new_n24823_;
  assign new_n24825_ = ~new_n24822_ & ~new_n24824_;
  assign new_n24826_ = ~ys__n34774 & ys__n34776;
  assign new_n24827_ = ~ys__n34778 & new_n24826_;
  assign new_n24828_ = ys__n34774 & ~ys__n34776;
  assign new_n24829_ = ~ys__n34778 & new_n24828_;
  assign new_n24830_ = ~new_n24827_ & ~new_n24829_;
  assign new_n24831_ = new_n24825_ & new_n24830_;
  assign new_n24832_ = ys__n34782 & ys__n34784;
  assign new_n24833_ = ys__n34780 & ys__n34782;
  assign new_n24834_ = ys__n34780 & ys__n34784;
  assign new_n24835_ = ~new_n24833_ & ~new_n24834_;
  assign new_n24836_ = ~new_n24832_ & new_n24835_;
  assign new_n24837_ = new_n24831_ & ~new_n24836_;
  assign new_n24838_ = ~new_n24831_ & new_n24836_;
  assign new_n24839_ = ~new_n24837_ & ~new_n24838_;
  assign new_n24840_ = ~new_n24821_ & ~new_n24839_;
  assign new_n24841_ = ys__n34784 & new_n24833_;
  assign new_n24842_ = ~ys__n34780 & ~ys__n34782;
  assign new_n24843_ = ys__n34784 & new_n24842_;
  assign new_n24844_ = ~new_n24841_ & ~new_n24843_;
  assign new_n24845_ = ~ys__n34780 & ys__n34782;
  assign new_n24846_ = ~ys__n34784 & new_n24845_;
  assign new_n24847_ = ys__n34780 & ~ys__n34782;
  assign new_n24848_ = ~ys__n34784 & new_n24847_;
  assign new_n24849_ = ~new_n24846_ & ~new_n24848_;
  assign new_n24850_ = new_n24844_ & new_n24849_;
  assign new_n24851_ = ys__n34788 & ys__n34790;
  assign new_n24852_ = ys__n34786 & ys__n34788;
  assign new_n24853_ = ys__n34786 & ys__n34790;
  assign new_n24854_ = ~new_n24852_ & ~new_n24853_;
  assign new_n24855_ = ~new_n24851_ & new_n24854_;
  assign new_n24856_ = new_n24850_ & ~new_n24855_;
  assign new_n24857_ = ~new_n24850_ & new_n24855_;
  assign new_n24858_ = ~new_n24856_ & ~new_n24857_;
  assign new_n24859_ = ys__n34790 & new_n24852_;
  assign new_n24860_ = ~ys__n34786 & ~ys__n34788;
  assign new_n24861_ = ys__n34790 & new_n24860_;
  assign new_n24862_ = ~new_n24859_ & ~new_n24861_;
  assign new_n24863_ = ~ys__n34786 & ys__n34788;
  assign new_n24864_ = ~ys__n34790 & new_n24863_;
  assign new_n24865_ = ys__n34786 & ~ys__n34788;
  assign new_n24866_ = ~ys__n34790 & new_n24865_;
  assign new_n24867_ = ~new_n24864_ & ~new_n24866_;
  assign new_n24868_ = new_n24862_ & new_n24867_;
  assign new_n24869_ = ys__n34794 & ys__n34796;
  assign new_n24870_ = ys__n34792 & ys__n34794;
  assign new_n24871_ = ys__n34792 & ys__n34796;
  assign new_n24872_ = ~new_n24870_ & ~new_n24871_;
  assign new_n24873_ = ~new_n24869_ & new_n24872_;
  assign new_n24874_ = new_n24868_ & ~new_n24873_;
  assign new_n24875_ = ~new_n24868_ & new_n24873_;
  assign new_n24876_ = ~new_n24874_ & ~new_n24875_;
  assign new_n24877_ = ~new_n24858_ & ~new_n24876_;
  assign new_n24878_ = new_n24840_ & new_n24877_;
  assign new_n24879_ = ys__n34796 & new_n24870_;
  assign new_n24880_ = ~ys__n34792 & ~ys__n34794;
  assign new_n24881_ = ys__n34796 & new_n24880_;
  assign new_n24882_ = ~new_n24879_ & ~new_n24881_;
  assign new_n24883_ = ~ys__n34792 & ys__n34794;
  assign new_n24884_ = ~ys__n34796 & new_n24883_;
  assign new_n24885_ = ys__n34792 & ~ys__n34794;
  assign new_n24886_ = ~ys__n34796 & new_n24885_;
  assign new_n24887_ = ~new_n24884_ & ~new_n24886_;
  assign new_n24888_ = new_n24882_ & new_n24887_;
  assign new_n24889_ = ys__n34800 & ys__n34802;
  assign new_n24890_ = ys__n34798 & ys__n34800;
  assign new_n24891_ = ys__n34798 & ys__n34802;
  assign new_n24892_ = ~new_n24890_ & ~new_n24891_;
  assign new_n24893_ = ~new_n24889_ & new_n24892_;
  assign new_n24894_ = new_n24888_ & ~new_n24893_;
  assign new_n24895_ = ~new_n24888_ & new_n24893_;
  assign new_n24896_ = ~new_n24894_ & ~new_n24895_;
  assign new_n24897_ = ys__n34802 & new_n24890_;
  assign new_n24898_ = ~ys__n34798 & ~ys__n34800;
  assign new_n24899_ = ys__n34802 & new_n24898_;
  assign new_n24900_ = ~new_n24897_ & ~new_n24899_;
  assign new_n24901_ = ~ys__n34798 & ys__n34800;
  assign new_n24902_ = ~ys__n34802 & new_n24901_;
  assign new_n24903_ = ys__n34798 & ~ys__n34800;
  assign new_n24904_ = ~ys__n34802 & new_n24903_;
  assign new_n24905_ = ~new_n24902_ & ~new_n24904_;
  assign new_n24906_ = new_n24900_ & new_n24905_;
  assign new_n24907_ = ys__n34806 & ys__n34808;
  assign new_n24908_ = ys__n34804 & ys__n34806;
  assign new_n24909_ = ys__n34804 & ys__n34808;
  assign new_n24910_ = ~new_n24908_ & ~new_n24909_;
  assign new_n24911_ = ~new_n24907_ & new_n24910_;
  assign new_n24912_ = new_n24906_ & ~new_n24911_;
  assign new_n24913_ = ~new_n24906_ & new_n24911_;
  assign new_n24914_ = ~new_n24912_ & ~new_n24913_;
  assign new_n24915_ = ~new_n24896_ & ~new_n24914_;
  assign new_n24916_ = ys__n34808 & new_n24908_;
  assign new_n24917_ = ~ys__n34804 & ~ys__n34806;
  assign new_n24918_ = ys__n34808 & new_n24917_;
  assign new_n24919_ = ~new_n24916_ & ~new_n24918_;
  assign new_n24920_ = ~ys__n34804 & ys__n34806;
  assign new_n24921_ = ~ys__n34808 & new_n24920_;
  assign new_n24922_ = ys__n34804 & ~ys__n34806;
  assign new_n24923_ = ~ys__n34808 & new_n24922_;
  assign new_n24924_ = ~new_n24921_ & ~new_n24923_;
  assign new_n24925_ = new_n24919_ & new_n24924_;
  assign new_n24926_ = ys__n34812 & ys__n34814;
  assign new_n24927_ = ys__n34810 & ys__n34812;
  assign new_n24928_ = ys__n34810 & ys__n34814;
  assign new_n24929_ = ~new_n24927_ & ~new_n24928_;
  assign new_n24930_ = ~new_n24926_ & new_n24929_;
  assign new_n24931_ = new_n24925_ & ~new_n24930_;
  assign new_n24932_ = ~new_n24925_ & new_n24930_;
  assign new_n24933_ = ~new_n24931_ & ~new_n24932_;
  assign new_n24934_ = ys__n34814 & new_n24927_;
  assign new_n24935_ = ~ys__n34810 & ~ys__n34812;
  assign new_n24936_ = ys__n34814 & new_n24935_;
  assign new_n24937_ = ~new_n24934_ & ~new_n24936_;
  assign new_n24938_ = ~ys__n34810 & ys__n34812;
  assign new_n24939_ = ~ys__n34814 & new_n24938_;
  assign new_n24940_ = ys__n34810 & ~ys__n34812;
  assign new_n24941_ = ~ys__n34814 & new_n24940_;
  assign new_n24942_ = ~new_n24939_ & ~new_n24941_;
  assign new_n24943_ = new_n24937_ & new_n24942_;
  assign new_n24944_ = ys__n34818 & ys__n34820;
  assign new_n24945_ = ys__n34816 & ys__n34820;
  assign new_n24946_ = ~new_n24717_ & ~new_n24945_;
  assign new_n24947_ = ~new_n24944_ & new_n24946_;
  assign new_n24948_ = new_n24943_ & ~new_n24947_;
  assign new_n24949_ = ~new_n24943_ & new_n24947_;
  assign new_n24950_ = ~new_n24948_ & ~new_n24949_;
  assign new_n24951_ = ~new_n24933_ & ~new_n24950_;
  assign new_n24952_ = new_n24915_ & new_n24951_;
  assign new_n24953_ = new_n24878_ & new_n24952_;
  assign new_n24954_ = ~new_n24803_ & new_n24953_;
  assign new_n24955_ = ~new_n24925_ & ~new_n24930_;
  assign new_n24956_ = ~new_n24943_ & ~new_n24947_;
  assign new_n24957_ = ~new_n24933_ & new_n24956_;
  assign new_n24958_ = ~new_n24955_ & ~new_n24957_;
  assign new_n24959_ = new_n24915_ & ~new_n24958_;
  assign new_n24960_ = ~new_n24888_ & ~new_n24893_;
  assign new_n24961_ = ~new_n24906_ & ~new_n24911_;
  assign new_n24962_ = ~new_n24896_ & new_n24961_;
  assign new_n24963_ = ~new_n24960_ & ~new_n24962_;
  assign new_n24964_ = ~new_n24959_ & new_n24963_;
  assign new_n24965_ = new_n24878_ & ~new_n24964_;
  assign new_n24966_ = ~new_n24850_ & ~new_n24855_;
  assign new_n24967_ = ~new_n24868_ & ~new_n24873_;
  assign new_n24968_ = ~new_n24858_ & new_n24967_;
  assign new_n24969_ = ~new_n24966_ & ~new_n24968_;
  assign new_n24970_ = new_n24840_ & ~new_n24969_;
  assign new_n24971_ = ~new_n24813_ & ~new_n24818_;
  assign new_n24972_ = ~new_n24831_ & ~new_n24836_;
  assign new_n24973_ = ~new_n24821_ & new_n24972_;
  assign new_n24974_ = ~new_n24971_ & ~new_n24973_;
  assign new_n24975_ = ~new_n24970_ & new_n24974_;
  assign new_n24976_ = ~new_n24965_ & new_n24975_;
  assign new_n24977_ = ~new_n24954_ & new_n24976_;
  assign new_n24978_ = ys__n34938 & ys__n34940;
  assign new_n24979_ = ys__n34942 & new_n24978_;
  assign new_n24980_ = ~ys__n34938 & ~ys__n34940;
  assign new_n24981_ = ys__n34942 & new_n24980_;
  assign new_n24982_ = ~new_n24979_ & ~new_n24981_;
  assign new_n24983_ = ~ys__n34938 & ys__n34940;
  assign new_n24984_ = ~ys__n34942 & new_n24983_;
  assign new_n24985_ = ys__n34938 & ~ys__n34940;
  assign new_n24986_ = ~ys__n34942 & new_n24985_;
  assign new_n24987_ = ~new_n24984_ & ~new_n24986_;
  assign new_n24988_ = new_n24982_ & new_n24987_;
  assign new_n24989_ = ys__n34944 & ys__n34946;
  assign new_n24990_ = new_n24988_ & new_n24989_;
  assign new_n24991_ = ~new_n24988_ & ~new_n24989_;
  assign new_n24992_ = ~new_n24990_ & ~new_n24991_;
  assign new_n24993_ = ~ys__n34934 & ys__n34936;
  assign new_n24994_ = ys__n34934 & ~ys__n34936;
  assign new_n24995_ = ~new_n24993_ & ~new_n24994_;
  assign new_n24996_ = ys__n34940 & ys__n34942;
  assign new_n24997_ = ys__n34938 & ys__n34942;
  assign new_n24998_ = ~new_n24978_ & ~new_n24997_;
  assign new_n24999_ = ~new_n24996_ & new_n24998_;
  assign new_n25000_ = new_n24995_ & ~new_n24999_;
  assign new_n25001_ = ~new_n24995_ & new_n24999_;
  assign new_n25002_ = ~new_n25000_ & ~new_n25001_;
  assign new_n25003_ = ~ys__n34944 & ys__n34946;
  assign new_n25004_ = ys__n34944 & ~ys__n34946;
  assign new_n25005_ = ~new_n25003_ & ~new_n25004_;
  assign new_n25006_ = ys__n34948 & ys__n34950;
  assign new_n25007_ = ~new_n25005_ & new_n25006_;
  assign new_n25008_ = ~new_n25002_ & new_n25007_;
  assign new_n25009_ = ~new_n24992_ & new_n25008_;
  assign new_n25010_ = ~new_n24995_ & ~new_n24999_;
  assign new_n25011_ = ~new_n24988_ & new_n24989_;
  assign new_n25012_ = ~new_n25002_ & new_n25011_;
  assign new_n25013_ = ~new_n25010_ & ~new_n25012_;
  assign new_n25014_ = ~new_n25009_ & new_n25013_;
  assign new_n25015_ = ys__n34912 & ys__n34914;
  assign new_n25016_ = ys__n34916 & new_n25015_;
  assign new_n25017_ = ~ys__n34912 & ~ys__n34914;
  assign new_n25018_ = ys__n34916 & new_n25017_;
  assign new_n25019_ = ~new_n25016_ & ~new_n25018_;
  assign new_n25020_ = ~ys__n34912 & ys__n34914;
  assign new_n25021_ = ~ys__n34916 & new_n25020_;
  assign new_n25022_ = ys__n34912 & ~ys__n34914;
  assign new_n25023_ = ~ys__n34916 & new_n25022_;
  assign new_n25024_ = ~new_n25021_ & ~new_n25023_;
  assign new_n25025_ = new_n25019_ & new_n25024_;
  assign new_n25026_ = ys__n34920 & ys__n34922;
  assign new_n25027_ = ys__n34918 & ys__n34920;
  assign new_n25028_ = ys__n34918 & ys__n34922;
  assign new_n25029_ = ~new_n25027_ & ~new_n25028_;
  assign new_n25030_ = ~new_n25026_ & new_n25029_;
  assign new_n25031_ = new_n25025_ & ~new_n25030_;
  assign new_n25032_ = ~new_n25025_ & new_n25030_;
  assign new_n25033_ = ~new_n25031_ & ~new_n25032_;
  assign new_n25034_ = ys__n34922 & new_n25027_;
  assign new_n25035_ = ~ys__n34918 & ~ys__n34920;
  assign new_n25036_ = ys__n34922 & new_n25035_;
  assign new_n25037_ = ~new_n25034_ & ~new_n25036_;
  assign new_n25038_ = ~ys__n34918 & ys__n34920;
  assign new_n25039_ = ~ys__n34922 & new_n25038_;
  assign new_n25040_ = ys__n34918 & ~ys__n34920;
  assign new_n25041_ = ~ys__n34922 & new_n25040_;
  assign new_n25042_ = ~new_n25039_ & ~new_n25041_;
  assign new_n25043_ = new_n25037_ & new_n25042_;
  assign new_n25044_ = ys__n34926 & ys__n34928;
  assign new_n25045_ = ys__n34924 & ys__n34926;
  assign new_n25046_ = ys__n34924 & ys__n34928;
  assign new_n25047_ = ~new_n25045_ & ~new_n25046_;
  assign new_n25048_ = ~new_n25044_ & new_n25047_;
  assign new_n25049_ = new_n25043_ & ~new_n25048_;
  assign new_n25050_ = ~new_n25043_ & new_n25048_;
  assign new_n25051_ = ~new_n25049_ & ~new_n25050_;
  assign new_n25052_ = ~new_n25033_ & ~new_n25051_;
  assign new_n25053_ = ys__n34928 & new_n25045_;
  assign new_n25054_ = ~ys__n34924 & ~ys__n34926;
  assign new_n25055_ = ys__n34928 & new_n25054_;
  assign new_n25056_ = ~new_n25053_ & ~new_n25055_;
  assign new_n25057_ = ~ys__n34924 & ys__n34926;
  assign new_n25058_ = ~ys__n34928 & new_n25057_;
  assign new_n25059_ = ys__n34924 & ~ys__n34926;
  assign new_n25060_ = ~ys__n34928 & new_n25059_;
  assign new_n25061_ = ~new_n25058_ & ~new_n25060_;
  assign new_n25062_ = new_n25056_ & new_n25061_;
  assign new_n25063_ = ys__n34930 & ys__n34932;
  assign new_n25064_ = new_n25062_ & new_n25063_;
  assign new_n25065_ = ~new_n25062_ & ~new_n25063_;
  assign new_n25066_ = ~new_n25064_ & ~new_n25065_;
  assign new_n25067_ = ~ys__n34930 & ys__n34932;
  assign new_n25068_ = ys__n34930 & ~ys__n34932;
  assign new_n25069_ = ~new_n25067_ & ~new_n25068_;
  assign new_n25070_ = ys__n34934 & ys__n34936;
  assign new_n25071_ = new_n25069_ & new_n25070_;
  assign new_n25072_ = ~new_n25069_ & ~new_n25070_;
  assign new_n25073_ = ~new_n25071_ & ~new_n25072_;
  assign new_n25074_ = ~new_n25066_ & ~new_n25073_;
  assign new_n25075_ = new_n25052_ & new_n25074_;
  assign new_n25076_ = ~new_n25014_ & new_n25075_;
  assign new_n25077_ = ~new_n25062_ & new_n25063_;
  assign new_n25078_ = ~new_n25069_ & new_n25070_;
  assign new_n25079_ = ~new_n25066_ & new_n25078_;
  assign new_n25080_ = ~new_n25077_ & ~new_n25079_;
  assign new_n25081_ = new_n25052_ & ~new_n25080_;
  assign new_n25082_ = ~new_n25025_ & ~new_n25030_;
  assign new_n25083_ = ~new_n25043_ & ~new_n25048_;
  assign new_n25084_ = ~new_n25033_ & new_n25083_;
  assign new_n25085_ = ~new_n25082_ & ~new_n25084_;
  assign new_n25086_ = ~new_n25081_ & new_n25085_;
  assign new_n25087_ = ~new_n25076_ & new_n25086_;
  assign new_n25088_ = ys__n34868 & new_n24667_;
  assign new_n25089_ = ~ys__n34864 & ~ys__n34866;
  assign new_n25090_ = ys__n34868 & new_n25089_;
  assign new_n25091_ = ~new_n25088_ & ~new_n25090_;
  assign new_n25092_ = ~ys__n34864 & ys__n34866;
  assign new_n25093_ = ~ys__n34868 & new_n25092_;
  assign new_n25094_ = ys__n34864 & ~ys__n34866;
  assign new_n25095_ = ~ys__n34868 & new_n25094_;
  assign new_n25096_ = ~new_n25093_ & ~new_n25095_;
  assign new_n25097_ = new_n25091_ & new_n25096_;
  assign new_n25098_ = ys__n34872 & ys__n34874;
  assign new_n25099_ = ys__n34870 & ys__n34872;
  assign new_n25100_ = ys__n34870 & ys__n34874;
  assign new_n25101_ = ~new_n25099_ & ~new_n25100_;
  assign new_n25102_ = ~new_n25098_ & new_n25101_;
  assign new_n25103_ = new_n25097_ & ~new_n25102_;
  assign new_n25104_ = ~new_n25097_ & new_n25102_;
  assign new_n25105_ = ~new_n25103_ & ~new_n25104_;
  assign new_n25106_ = ys__n34874 & new_n25099_;
  assign new_n25107_ = ~ys__n34870 & ~ys__n34872;
  assign new_n25108_ = ys__n34874 & new_n25107_;
  assign new_n25109_ = ~new_n25106_ & ~new_n25108_;
  assign new_n25110_ = ~ys__n34870 & ys__n34872;
  assign new_n25111_ = ~ys__n34874 & new_n25110_;
  assign new_n25112_ = ys__n34870 & ~ys__n34872;
  assign new_n25113_ = ~ys__n34874 & new_n25112_;
  assign new_n25114_ = ~new_n25111_ & ~new_n25113_;
  assign new_n25115_ = new_n25109_ & new_n25114_;
  assign new_n25116_ = ys__n34878 & ys__n34880;
  assign new_n25117_ = ys__n34876 & ys__n34878;
  assign new_n25118_ = ys__n34876 & ys__n34880;
  assign new_n25119_ = ~new_n25117_ & ~new_n25118_;
  assign new_n25120_ = ~new_n25116_ & new_n25119_;
  assign new_n25121_ = new_n25115_ & ~new_n25120_;
  assign new_n25122_ = ~new_n25115_ & new_n25120_;
  assign new_n25123_ = ~new_n25121_ & ~new_n25122_;
  assign new_n25124_ = ~new_n25105_ & ~new_n25123_;
  assign new_n25125_ = ys__n34880 & new_n25117_;
  assign new_n25126_ = ~ys__n34876 & ~ys__n34878;
  assign new_n25127_ = ys__n34880 & new_n25126_;
  assign new_n25128_ = ~new_n25125_ & ~new_n25127_;
  assign new_n25129_ = ~ys__n34876 & ys__n34878;
  assign new_n25130_ = ~ys__n34880 & new_n25129_;
  assign new_n25131_ = ys__n34876 & ~ys__n34878;
  assign new_n25132_ = ~ys__n34880 & new_n25131_;
  assign new_n25133_ = ~new_n25130_ & ~new_n25132_;
  assign new_n25134_ = new_n25128_ & new_n25133_;
  assign new_n25135_ = ys__n34884 & ys__n34886;
  assign new_n25136_ = ys__n34882 & ys__n34884;
  assign new_n25137_ = ys__n34882 & ys__n34886;
  assign new_n25138_ = ~new_n25136_ & ~new_n25137_;
  assign new_n25139_ = ~new_n25135_ & new_n25138_;
  assign new_n25140_ = new_n25134_ & ~new_n25139_;
  assign new_n25141_ = ~new_n25134_ & new_n25139_;
  assign new_n25142_ = ~new_n25140_ & ~new_n25141_;
  assign new_n25143_ = ys__n34886 & new_n25136_;
  assign new_n25144_ = ~ys__n34882 & ~ys__n34884;
  assign new_n25145_ = ys__n34886 & new_n25144_;
  assign new_n25146_ = ~new_n25143_ & ~new_n25145_;
  assign new_n25147_ = ~ys__n34882 & ys__n34884;
  assign new_n25148_ = ~ys__n34886 & new_n25147_;
  assign new_n25149_ = ys__n34882 & ~ys__n34884;
  assign new_n25150_ = ~ys__n34886 & new_n25149_;
  assign new_n25151_ = ~new_n25148_ & ~new_n25150_;
  assign new_n25152_ = new_n25146_ & new_n25151_;
  assign new_n25153_ = ys__n34890 & ys__n34892;
  assign new_n25154_ = ys__n34888 & ys__n34890;
  assign new_n25155_ = ys__n34888 & ys__n34892;
  assign new_n25156_ = ~new_n25154_ & ~new_n25155_;
  assign new_n25157_ = ~new_n25153_ & new_n25156_;
  assign new_n25158_ = new_n25152_ & ~new_n25157_;
  assign new_n25159_ = ~new_n25152_ & new_n25157_;
  assign new_n25160_ = ~new_n25158_ & ~new_n25159_;
  assign new_n25161_ = ~new_n25142_ & ~new_n25160_;
  assign new_n25162_ = new_n25124_ & new_n25161_;
  assign new_n25163_ = ys__n34892 & new_n25154_;
  assign new_n25164_ = ~ys__n34888 & ~ys__n34890;
  assign new_n25165_ = ys__n34892 & new_n25164_;
  assign new_n25166_ = ~new_n25163_ & ~new_n25165_;
  assign new_n25167_ = ~ys__n34888 & ys__n34890;
  assign new_n25168_ = ~ys__n34892 & new_n25167_;
  assign new_n25169_ = ys__n34888 & ~ys__n34890;
  assign new_n25170_ = ~ys__n34892 & new_n25169_;
  assign new_n25171_ = ~new_n25168_ & ~new_n25170_;
  assign new_n25172_ = new_n25166_ & new_n25171_;
  assign new_n25173_ = ys__n34896 & ys__n34898;
  assign new_n25174_ = ys__n34894 & ys__n34896;
  assign new_n25175_ = ys__n34894 & ys__n34898;
  assign new_n25176_ = ~new_n25174_ & ~new_n25175_;
  assign new_n25177_ = ~new_n25173_ & new_n25176_;
  assign new_n25178_ = new_n25172_ & ~new_n25177_;
  assign new_n25179_ = ~new_n25172_ & new_n25177_;
  assign new_n25180_ = ~new_n25178_ & ~new_n25179_;
  assign new_n25181_ = ys__n34898 & new_n25174_;
  assign new_n25182_ = ~ys__n34894 & ~ys__n34896;
  assign new_n25183_ = ys__n34898 & new_n25182_;
  assign new_n25184_ = ~new_n25181_ & ~new_n25183_;
  assign new_n25185_ = ~ys__n34894 & ys__n34896;
  assign new_n25186_ = ~ys__n34898 & new_n25185_;
  assign new_n25187_ = ys__n34894 & ~ys__n34896;
  assign new_n25188_ = ~ys__n34898 & new_n25187_;
  assign new_n25189_ = ~new_n25186_ & ~new_n25188_;
  assign new_n25190_ = new_n25184_ & new_n25189_;
  assign new_n25191_ = ys__n34902 & ys__n34904;
  assign new_n25192_ = ys__n34900 & ys__n34902;
  assign new_n25193_ = ys__n34900 & ys__n34904;
  assign new_n25194_ = ~new_n25192_ & ~new_n25193_;
  assign new_n25195_ = ~new_n25191_ & new_n25194_;
  assign new_n25196_ = new_n25190_ & ~new_n25195_;
  assign new_n25197_ = ~new_n25190_ & new_n25195_;
  assign new_n25198_ = ~new_n25196_ & ~new_n25197_;
  assign new_n25199_ = ~new_n25180_ & ~new_n25198_;
  assign new_n25200_ = ys__n34904 & new_n25192_;
  assign new_n25201_ = ~ys__n34900 & ~ys__n34902;
  assign new_n25202_ = ys__n34904 & new_n25201_;
  assign new_n25203_ = ~new_n25200_ & ~new_n25202_;
  assign new_n25204_ = ~ys__n34900 & ys__n34902;
  assign new_n25205_ = ~ys__n34904 & new_n25204_;
  assign new_n25206_ = ys__n34900 & ~ys__n34902;
  assign new_n25207_ = ~ys__n34904 & new_n25206_;
  assign new_n25208_ = ~new_n25205_ & ~new_n25207_;
  assign new_n25209_ = new_n25203_ & new_n25208_;
  assign new_n25210_ = ys__n34908 & ys__n34910;
  assign new_n25211_ = ys__n34906 & ys__n34908;
  assign new_n25212_ = ys__n34906 & ys__n34910;
  assign new_n25213_ = ~new_n25211_ & ~new_n25212_;
  assign new_n25214_ = ~new_n25210_ & new_n25213_;
  assign new_n25215_ = new_n25209_ & ~new_n25214_;
  assign new_n25216_ = ~new_n25209_ & new_n25214_;
  assign new_n25217_ = ~new_n25215_ & ~new_n25216_;
  assign new_n25218_ = ys__n34910 & new_n25211_;
  assign new_n25219_ = ~ys__n34906 & ~ys__n34908;
  assign new_n25220_ = ys__n34910 & new_n25219_;
  assign new_n25221_ = ~new_n25218_ & ~new_n25220_;
  assign new_n25222_ = ~ys__n34906 & ys__n34908;
  assign new_n25223_ = ~ys__n34910 & new_n25222_;
  assign new_n25224_ = ys__n34906 & ~ys__n34908;
  assign new_n25225_ = ~ys__n34910 & new_n25224_;
  assign new_n25226_ = ~new_n25223_ & ~new_n25225_;
  assign new_n25227_ = new_n25221_ & new_n25226_;
  assign new_n25228_ = ys__n34914 & ys__n34916;
  assign new_n25229_ = ys__n34912 & ys__n34916;
  assign new_n25230_ = ~new_n25015_ & ~new_n25229_;
  assign new_n25231_ = ~new_n25228_ & new_n25230_;
  assign new_n25232_ = new_n25227_ & ~new_n25231_;
  assign new_n25233_ = ~new_n25227_ & new_n25231_;
  assign new_n25234_ = ~new_n25232_ & ~new_n25233_;
  assign new_n25235_ = ~new_n25217_ & ~new_n25234_;
  assign new_n25236_ = new_n25199_ & new_n25235_;
  assign new_n25237_ = new_n25162_ & new_n25236_;
  assign new_n25238_ = ~new_n25087_ & new_n25237_;
  assign new_n25239_ = ~new_n25209_ & ~new_n25214_;
  assign new_n25240_ = ~new_n25227_ & ~new_n25231_;
  assign new_n25241_ = ~new_n25217_ & new_n25240_;
  assign new_n25242_ = ~new_n25239_ & ~new_n25241_;
  assign new_n25243_ = new_n25199_ & ~new_n25242_;
  assign new_n25244_ = ~new_n25172_ & ~new_n25177_;
  assign new_n25245_ = ~new_n25190_ & ~new_n25195_;
  assign new_n25246_ = ~new_n25180_ & new_n25245_;
  assign new_n25247_ = ~new_n25244_ & ~new_n25246_;
  assign new_n25248_ = ~new_n25243_ & new_n25247_;
  assign new_n25249_ = new_n25162_ & ~new_n25248_;
  assign new_n25250_ = ~new_n25134_ & ~new_n25139_;
  assign new_n25251_ = ~new_n25152_ & ~new_n25157_;
  assign new_n25252_ = ~new_n25142_ & new_n25251_;
  assign new_n25253_ = ~new_n25250_ & ~new_n25252_;
  assign new_n25254_ = new_n25124_ & ~new_n25253_;
  assign new_n25255_ = ~new_n25097_ & ~new_n25102_;
  assign new_n25256_ = ~new_n25115_ & ~new_n25120_;
  assign new_n25257_ = ~new_n25105_ & new_n25256_;
  assign new_n25258_ = ~new_n25255_ & ~new_n25257_;
  assign new_n25259_ = ~new_n25254_ & new_n25258_;
  assign new_n25260_ = ~new_n25249_ & new_n25259_;
  assign new_n25261_ = ~new_n25238_ & new_n25260_;
  assign new_n25262_ = ~new_n24977_ & new_n25261_;
  assign new_n25263_ = ~new_n24803_ & new_n24952_;
  assign new_n25264_ = new_n24964_ & ~new_n25263_;
  assign new_n25265_ = new_n24877_ & ~new_n25264_;
  assign new_n25266_ = new_n24969_ & ~new_n25265_;
  assign new_n25267_ = ~new_n24839_ & ~new_n25266_;
  assign new_n25268_ = ~new_n24972_ & ~new_n25267_;
  assign new_n25269_ = new_n24821_ & ~new_n25268_;
  assign new_n25270_ = ~new_n24821_ & new_n25268_;
  assign new_n25271_ = ~new_n25269_ & ~new_n25270_;
  assign new_n25272_ = ~new_n24803_ & new_n24951_;
  assign new_n25273_ = new_n24958_ & ~new_n25272_;
  assign new_n25274_ = ~new_n24914_ & ~new_n25273_;
  assign new_n25275_ = ~new_n24961_ & ~new_n25274_;
  assign new_n25276_ = new_n24896_ & ~new_n25275_;
  assign new_n25277_ = ~new_n24896_ & new_n25275_;
  assign new_n25278_ = ~new_n25276_ & ~new_n25277_;
  assign new_n25279_ = new_n24914_ & ~new_n25273_;
  assign new_n25280_ = ~new_n24914_ & new_n25273_;
  assign new_n25281_ = ~new_n25279_ & ~new_n25280_;
  assign new_n25282_ = ~new_n24803_ & ~new_n24950_;
  assign new_n25283_ = ~new_n24956_ & ~new_n25282_;
  assign new_n25284_ = new_n24933_ & ~new_n25283_;
  assign new_n25285_ = ~new_n24933_ & new_n25283_;
  assign new_n25286_ = ~new_n25284_ & ~new_n25285_;
  assign new_n25287_ = ~new_n24803_ & new_n24950_;
  assign new_n25288_ = new_n24803_ & ~new_n24950_;
  assign new_n25289_ = ~new_n25287_ & ~new_n25288_;
  assign new_n25290_ = ~new_n25286_ & ~new_n25289_;
  assign new_n25291_ = ~new_n25281_ & new_n25290_;
  assign new_n25292_ = ~new_n25278_ & new_n25291_;
  assign new_n25293_ = ~new_n24876_ & ~new_n25264_;
  assign new_n25294_ = ~new_n24967_ & ~new_n25293_;
  assign new_n25295_ = new_n24858_ & ~new_n25294_;
  assign new_n25296_ = ~new_n24858_ & new_n25294_;
  assign new_n25297_ = ~new_n25295_ & ~new_n25296_;
  assign new_n25298_ = new_n24876_ & ~new_n25264_;
  assign new_n25299_ = ~new_n24876_ & new_n25264_;
  assign new_n25300_ = ~new_n25298_ & ~new_n25299_;
  assign new_n25301_ = ~new_n25297_ & ~new_n25300_;
  assign new_n25302_ = new_n24839_ & ~new_n25266_;
  assign new_n25303_ = ~new_n24839_ & new_n25266_;
  assign new_n25304_ = ~new_n25302_ & ~new_n25303_;
  assign new_n25305_ = ~new_n24716_ & new_n24790_;
  assign new_n25306_ = new_n24796_ & ~new_n25305_;
  assign new_n25307_ = ~new_n24753_ & ~new_n25306_;
  assign new_n25308_ = ~new_n24799_ & ~new_n25307_;
  assign new_n25309_ = new_n24735_ & ~new_n25308_;
  assign new_n25310_ = ~new_n24735_ & new_n25308_;
  assign new_n25311_ = ~new_n25309_ & ~new_n25310_;
  assign new_n25312_ = ~new_n24716_ & ~new_n24789_;
  assign new_n25313_ = ~new_n24794_ & ~new_n25312_;
  assign new_n25314_ = new_n24772_ & ~new_n25313_;
  assign new_n25315_ = ~new_n24772_ & new_n25313_;
  assign new_n25316_ = ~new_n25314_ & ~new_n25315_;
  assign new_n25317_ = ~new_n24716_ & new_n24789_;
  assign new_n25318_ = new_n24716_ & ~new_n24789_;
  assign new_n25319_ = ~new_n25317_ & ~new_n25318_;
  assign new_n25320_ = ~new_n25316_ & ~new_n25319_;
  assign new_n25321_ = new_n24753_ & ~new_n25306_;
  assign new_n25322_ = ~new_n24753_ & new_n25306_;
  assign new_n25323_ = ~new_n25321_ & ~new_n25322_;
  assign new_n25324_ = ~new_n24673_ & ~new_n24709_;
  assign new_n25325_ = ~new_n24713_ & ~new_n25324_;
  assign new_n25326_ = new_n24692_ & ~new_n25325_;
  assign new_n25327_ = ~new_n24692_ & new_n25325_;
  assign new_n25328_ = ~new_n25326_ & ~new_n25327_;
  assign new_n25329_ = ~new_n24673_ & new_n24709_;
  assign new_n25330_ = new_n24673_ & ~new_n24709_;
  assign new_n25331_ = ~new_n25329_ & ~new_n25330_;
  assign new_n25332_ = new_n24655_ & new_n24671_;
  assign new_n25333_ = ~new_n24655_ & ~new_n24671_;
  assign new_n25334_ = ~new_n25332_ & ~new_n25333_;
  assign new_n25335_ = new_n24665_ & ~new_n24670_;
  assign new_n25336_ = ~new_n24665_ & new_n24670_;
  assign new_n25337_ = ~new_n25335_ & ~new_n25336_;
  assign new_n25338_ = ~new_n25334_ & ~new_n25337_;
  assign new_n25339_ = ~new_n25331_ & new_n25338_;
  assign new_n25340_ = ~new_n25328_ & new_n25339_;
  assign new_n25341_ = ~new_n25323_ & new_n25340_;
  assign new_n25342_ = new_n25320_ & new_n25341_;
  assign new_n25343_ = ~new_n25311_ & new_n25342_;
  assign new_n25344_ = ~new_n25304_ & new_n25343_;
  assign new_n25345_ = new_n25301_ & new_n25344_;
  assign new_n25346_ = new_n25292_ & new_n25345_;
  assign new_n25347_ = ~new_n25271_ & new_n25346_;
  assign new_n25348_ = new_n24977_ & new_n25347_;
  assign new_n25349_ = ~new_n24977_ & ~new_n25347_;
  assign new_n25350_ = ~new_n25348_ & ~new_n25349_;
  assign new_n25351_ = ~new_n25261_ & ~new_n25350_;
  assign new_n25352_ = ~new_n25262_ & ~new_n25351_;
  assign new_n25353_ = ~ys__n33749 & ~new_n25352_;
  assign new_n25354_ = ~ys__n33749 & ~new_n25353_;
  assign new_n25355_ = ~new_n24635_ & new_n25354_;
  assign new_n25356_ = new_n24635_ & ~new_n25354_;
  assign new_n25357_ = ~new_n25355_ & ~new_n25356_;
  assign new_n25358_ = ys__n33749 & ~new_n25352_;
  assign new_n25359_ = ~new_n25357_ & ~new_n25358_;
  assign new_n25360_ = ~new_n24635_ & new_n25358_;
  assign new_n25361_ = ~new_n25359_ & ~new_n25360_;
  assign new_n25362_ = ~new_n24614_ & ~new_n25361_;
  assign new_n25363_ = ~new_n24616_ & ~new_n25362_;
  assign new_n25364_ = ys__n31031 & new_n13350_;
  assign new_n25365_ = ~new_n25363_ & ~new_n25364_;
  assign new_n25366_ = ~ys__n34948 & ys__n34950;
  assign new_n25367_ = ys__n34948 & ~ys__n34950;
  assign new_n25368_ = ~new_n25366_ & ~new_n25367_;
  assign new_n25369_ = new_n25364_ & ~new_n25368_;
  assign new_n25370_ = ~new_n25365_ & ~new_n25369_;
  assign new_n25371_ = ys__n2779 & ~ys__n2535;
  assign new_n25372_ = ~new_n25370_ & new_n25371_;
  assign new_n25373_ = ys__n2535 & ~new_n25370_;
  assign new_n25374_ = ~new_n25372_ & ~new_n25373_;
  assign new_n25375_ = ~new_n13708_ & ~new_n25374_;
  assign new_n25376_ = ys__n166 & ys__n30819;
  assign new_n25377_ = ~new_n24611_ & new_n25376_;
  assign new_n25378_ = ys__n168 & ys__n30816;
  assign new_n25379_ = ys__n30818 & new_n25378_;
  assign new_n25380_ = ys__n168 & ys__n30820;
  assign new_n25381_ = ~new_n24611_ & new_n25380_;
  assign new_n25382_ = ~new_n25379_ & ~new_n25381_;
  assign new_n25383_ = ~new_n25377_ & new_n25382_;
  assign new_n25384_ = ~ys__n166 & ys__n168;
  assign new_n25385_ = ys__n47074 & new_n25384_;
  assign new_n25386_ = ys__n166 & ~ys__n168;
  assign new_n25387_ = ys__n47010 & new_n25386_;
  assign new_n25388_ = ~new_n25385_ & ~new_n25387_;
  assign new_n25389_ = ~new_n25384_ & ~new_n25386_;
  assign new_n25390_ = ~new_n25388_ & ~new_n25389_;
  assign new_n25391_ = new_n25383_ & new_n25390_;
  assign new_n25392_ = new_n25261_ & ~new_n25337_;
  assign new_n25393_ = ~new_n25261_ & new_n25337_;
  assign new_n25394_ = ~new_n25392_ & ~new_n25393_;
  assign new_n25395_ = ~new_n25383_ & ~new_n25394_;
  assign new_n25396_ = ~new_n25391_ & ~new_n25395_;
  assign new_n25397_ = ys__n166 & ys__n30815;
  assign new_n25398_ = ys__n30816 & new_n25397_;
  assign new_n25399_ = ~ys__n2779 & ~new_n25398_;
  assign new_n25400_ = ~new_n25396_ & new_n25399_;
  assign new_n25401_ = ys__n314 & ~new_n25399_;
  assign new_n25402_ = ~new_n25400_ & ~new_n25401_;
  assign new_n25403_ = new_n13708_ & ~new_n25402_;
  assign new_n25404_ = ~new_n25375_ & ~new_n25403_;
  assign new_n25405_ = ~ys__n1598 & ~new_n25404_;
  assign new_n25406_ = ys__n24741 & ys__n1598;
  assign ys__n24742 = new_n25405_ | new_n25406_;
  assign new_n25408_ = ys__n31031 & ys__n47027;
  assign new_n25409_ = new_n24614_ & new_n25408_;
  assign new_n25410_ = ys__n34756 & ys__n34758;
  assign new_n25411_ = ys__n34760 & new_n25410_;
  assign new_n25412_ = ~ys__n34756 & ~ys__n34758;
  assign new_n25413_ = ys__n34760 & new_n25412_;
  assign new_n25414_ = ~new_n25411_ & ~new_n25413_;
  assign new_n25415_ = ~ys__n34756 & ys__n34758;
  assign new_n25416_ = ~ys__n34760 & new_n25415_;
  assign new_n25417_ = ys__n34756 & ~ys__n34758;
  assign new_n25418_ = ~ys__n34760 & new_n25417_;
  assign new_n25419_ = ~new_n25416_ & ~new_n25418_;
  assign new_n25420_ = new_n25414_ & new_n25419_;
  assign new_n25421_ = ys__n34764 & ys__n34766;
  assign new_n25422_ = ys__n34762 & ys__n34766;
  assign new_n25423_ = ~new_n24617_ & ~new_n25422_;
  assign new_n25424_ = ~new_n25421_ & new_n25423_;
  assign new_n25425_ = new_n25420_ & ~new_n25424_;
  assign new_n25426_ = ~new_n25420_ & new_n25424_;
  assign new_n25427_ = ~new_n25425_ & ~new_n25426_;
  assign new_n25428_ = ~new_n24627_ & ~new_n24632_;
  assign new_n25429_ = new_n25427_ & new_n25428_;
  assign new_n25430_ = ~new_n25427_ & ~new_n25428_;
  assign new_n25431_ = ~new_n25429_ & ~new_n25430_;
  assign new_n25432_ = new_n25354_ & ~new_n25431_;
  assign new_n25433_ = ~new_n24635_ & new_n25431_;
  assign new_n25434_ = new_n24635_ & ~new_n25431_;
  assign new_n25435_ = ~new_n25433_ & ~new_n25434_;
  assign new_n25436_ = ~new_n25354_ & ~new_n25435_;
  assign new_n25437_ = ~new_n25432_ & ~new_n25436_;
  assign new_n25438_ = ~new_n25358_ & ~new_n25437_;
  assign new_n25439_ = new_n25358_ & new_n25431_;
  assign new_n25440_ = ~new_n25438_ & ~new_n25439_;
  assign new_n25441_ = ~new_n24614_ & ~new_n25440_;
  assign new_n25442_ = ~new_n25409_ & ~new_n25441_;
  assign new_n25443_ = ~new_n25364_ & ~new_n25442_;
  assign new_n25444_ = new_n25005_ & new_n25006_;
  assign new_n25445_ = ~new_n25005_ & ~new_n25006_;
  assign new_n25446_ = ~new_n25444_ & ~new_n25445_;
  assign new_n25447_ = new_n25364_ & ~new_n25446_;
  assign new_n25448_ = ~new_n25443_ & ~new_n25447_;
  assign new_n25449_ = new_n25371_ & ~new_n25448_;
  assign new_n25450_ = ys__n2535 & ~new_n25448_;
  assign new_n25451_ = ~new_n25449_ & ~new_n25450_;
  assign new_n25452_ = ~new_n13708_ & ~new_n25451_;
  assign new_n25453_ = ys__n47075 & new_n25384_;
  assign new_n25454_ = ys__n47011 & new_n25386_;
  assign new_n25455_ = ~new_n25453_ & ~new_n25454_;
  assign new_n25456_ = ~new_n25389_ & ~new_n25455_;
  assign new_n25457_ = new_n25383_ & new_n25456_;
  assign new_n25458_ = new_n25261_ & ~new_n25334_;
  assign new_n25459_ = new_n25334_ & ~new_n25337_;
  assign new_n25460_ = ~new_n25334_ & new_n25337_;
  assign new_n25461_ = ~new_n25459_ & ~new_n25460_;
  assign new_n25462_ = ~new_n25261_ & ~new_n25461_;
  assign new_n25463_ = ~new_n25458_ & ~new_n25462_;
  assign new_n25464_ = ~new_n25383_ & ~new_n25463_;
  assign new_n25465_ = ~new_n25457_ & ~new_n25464_;
  assign new_n25466_ = new_n25399_ & ~new_n25465_;
  assign new_n25467_ = ys__n170 & ~new_n25399_;
  assign new_n25468_ = ~new_n25466_ & ~new_n25467_;
  assign new_n25469_ = new_n13708_ & ~new_n25468_;
  assign new_n25470_ = ~new_n25452_ & ~new_n25469_;
  assign new_n25471_ = ~ys__n1598 & ~new_n25470_;
  assign new_n25472_ = ys__n24744 & ys__n1598;
  assign ys__n24745 = new_n25471_ | new_n25472_;
  assign new_n25474_ = ys__n31031 & ys__n47028;
  assign new_n25475_ = new_n24614_ & new_n25474_;
  assign new_n25476_ = ys__n34750 & ys__n34752;
  assign new_n25477_ = ys__n34754 & new_n25476_;
  assign new_n25478_ = ~ys__n34750 & ~ys__n34752;
  assign new_n25479_ = ys__n34754 & new_n25478_;
  assign new_n25480_ = ~new_n25477_ & ~new_n25479_;
  assign new_n25481_ = ~ys__n34750 & ys__n34752;
  assign new_n25482_ = ~ys__n34754 & new_n25481_;
  assign new_n25483_ = ys__n34750 & ~ys__n34752;
  assign new_n25484_ = ~ys__n34754 & new_n25483_;
  assign new_n25485_ = ~new_n25482_ & ~new_n25484_;
  assign new_n25486_ = new_n25480_ & new_n25485_;
  assign new_n25487_ = ys__n34758 & ys__n34760;
  assign new_n25488_ = ys__n34756 & ys__n34760;
  assign new_n25489_ = ~new_n25410_ & ~new_n25488_;
  assign new_n25490_ = ~new_n25487_ & new_n25489_;
  assign new_n25491_ = new_n25486_ & ~new_n25490_;
  assign new_n25492_ = ~new_n25486_ & new_n25490_;
  assign new_n25493_ = ~new_n25491_ & ~new_n25492_;
  assign new_n25494_ = ~new_n25420_ & ~new_n25424_;
  assign new_n25495_ = ~new_n25427_ & new_n25428_;
  assign new_n25496_ = ~new_n25494_ & ~new_n25495_;
  assign new_n25497_ = new_n25493_ & ~new_n25496_;
  assign new_n25498_ = ~new_n25493_ & new_n25496_;
  assign new_n25499_ = ~new_n25497_ & ~new_n25498_;
  assign new_n25500_ = new_n25354_ & ~new_n25499_;
  assign new_n25501_ = ~new_n24635_ & ~new_n25431_;
  assign new_n25502_ = new_n25499_ & new_n25501_;
  assign new_n25503_ = ~new_n25499_ & ~new_n25501_;
  assign new_n25504_ = ~new_n25502_ & ~new_n25503_;
  assign new_n25505_ = ~new_n25354_ & ~new_n25504_;
  assign new_n25506_ = ~new_n25500_ & ~new_n25505_;
  assign new_n25507_ = ~new_n25358_ & ~new_n25506_;
  assign new_n25508_ = ~new_n25431_ & new_n25499_;
  assign new_n25509_ = new_n25431_ & ~new_n25499_;
  assign new_n25510_ = ~new_n25508_ & ~new_n25509_;
  assign new_n25511_ = new_n25358_ & ~new_n25510_;
  assign new_n25512_ = ~new_n25507_ & ~new_n25511_;
  assign new_n25513_ = ~new_n24614_ & ~new_n25512_;
  assign new_n25514_ = ~new_n25475_ & ~new_n25513_;
  assign new_n25515_ = ~new_n25364_ & ~new_n25514_;
  assign new_n25516_ = new_n24992_ & new_n25007_;
  assign new_n25517_ = ~new_n24992_ & ~new_n25007_;
  assign new_n25518_ = ~new_n25516_ & ~new_n25517_;
  assign new_n25519_ = new_n25364_ & ~new_n25518_;
  assign new_n25520_ = ~new_n25515_ & ~new_n25519_;
  assign new_n25521_ = new_n25371_ & ~new_n25520_;
  assign new_n25522_ = ys__n2535 & ~new_n25520_;
  assign new_n25523_ = ~new_n25521_ & ~new_n25522_;
  assign new_n25524_ = ~new_n13708_ & ~new_n25523_;
  assign new_n25525_ = ys__n47076 & new_n25384_;
  assign new_n25526_ = ys__n47012 & new_n25386_;
  assign new_n25527_ = ~new_n25525_ & ~new_n25526_;
  assign new_n25528_ = ~new_n25389_ & ~new_n25527_;
  assign new_n25529_ = new_n25383_ & new_n25528_;
  assign new_n25530_ = new_n25261_ & ~new_n25331_;
  assign new_n25531_ = new_n25331_ & new_n25338_;
  assign new_n25532_ = ~new_n25331_ & ~new_n25338_;
  assign new_n25533_ = ~new_n25531_ & ~new_n25532_;
  assign new_n25534_ = ~new_n25261_ & ~new_n25533_;
  assign new_n25535_ = ~new_n25530_ & ~new_n25534_;
  assign new_n25536_ = ~new_n25383_ & ~new_n25535_;
  assign new_n25537_ = ~new_n25529_ & ~new_n25536_;
  assign new_n25538_ = new_n25399_ & ~new_n25537_;
  assign new_n25539_ = ys__n380 & ~new_n25399_;
  assign new_n25540_ = ~new_n25538_ & ~new_n25539_;
  assign new_n25541_ = new_n13708_ & ~new_n25540_;
  assign new_n25542_ = ~new_n25524_ & ~new_n25541_;
  assign new_n25543_ = ~ys__n1598 & ~new_n25542_;
  assign new_n25544_ = ys__n24747 & ys__n1598;
  assign ys__n24748 = new_n25543_ | new_n25544_;
  assign new_n25546_ = ys__n31031 & ys__n47029;
  assign new_n25547_ = new_n24614_ & new_n25546_;
  assign new_n25548_ = ys__n34744 & ys__n34746;
  assign new_n25549_ = ys__n34748 & new_n25548_;
  assign new_n25550_ = ~ys__n34744 & ~ys__n34746;
  assign new_n25551_ = ys__n34748 & new_n25550_;
  assign new_n25552_ = ~new_n25549_ & ~new_n25551_;
  assign new_n25553_ = ~ys__n34744 & ys__n34746;
  assign new_n25554_ = ~ys__n34748 & new_n25553_;
  assign new_n25555_ = ys__n34744 & ~ys__n34746;
  assign new_n25556_ = ~ys__n34748 & new_n25555_;
  assign new_n25557_ = ~new_n25554_ & ~new_n25556_;
  assign new_n25558_ = new_n25552_ & new_n25557_;
  assign new_n25559_ = ys__n34752 & ys__n34754;
  assign new_n25560_ = ys__n34750 & ys__n34754;
  assign new_n25561_ = ~new_n25476_ & ~new_n25560_;
  assign new_n25562_ = ~new_n25559_ & new_n25561_;
  assign new_n25563_ = new_n25558_ & ~new_n25562_;
  assign new_n25564_ = ~new_n25558_ & new_n25562_;
  assign new_n25565_ = ~new_n25563_ & ~new_n25564_;
  assign new_n25566_ = ~new_n25486_ & ~new_n25490_;
  assign new_n25567_ = ~new_n25493_ & ~new_n25496_;
  assign new_n25568_ = ~new_n25566_ & ~new_n25567_;
  assign new_n25569_ = new_n25565_ & ~new_n25568_;
  assign new_n25570_ = ~new_n25565_ & new_n25568_;
  assign new_n25571_ = ~new_n25569_ & ~new_n25570_;
  assign new_n25572_ = new_n25354_ & ~new_n25571_;
  assign new_n25573_ = ~new_n25499_ & new_n25501_;
  assign new_n25574_ = new_n25571_ & new_n25573_;
  assign new_n25575_ = ~new_n25571_ & ~new_n25573_;
  assign new_n25576_ = ~new_n25574_ & ~new_n25575_;
  assign new_n25577_ = ~new_n25354_ & ~new_n25576_;
  assign new_n25578_ = ~new_n25572_ & ~new_n25577_;
  assign new_n25579_ = ~new_n25358_ & ~new_n25578_;
  assign new_n25580_ = ~new_n25431_ & ~new_n25499_;
  assign new_n25581_ = new_n25571_ & new_n25580_;
  assign new_n25582_ = ~new_n25571_ & ~new_n25580_;
  assign new_n25583_ = ~new_n25581_ & ~new_n25582_;
  assign new_n25584_ = new_n25358_ & ~new_n25583_;
  assign new_n25585_ = ~new_n25579_ & ~new_n25584_;
  assign new_n25586_ = ~new_n24614_ & ~new_n25585_;
  assign new_n25587_ = ~new_n25547_ & ~new_n25586_;
  assign new_n25588_ = ~new_n25364_ & ~new_n25587_;
  assign new_n25589_ = ~new_n24992_ & new_n25007_;
  assign new_n25590_ = ~new_n25011_ & ~new_n25589_;
  assign new_n25591_ = new_n25002_ & ~new_n25590_;
  assign new_n25592_ = ~new_n25002_ & new_n25590_;
  assign new_n25593_ = ~new_n25591_ & ~new_n25592_;
  assign new_n25594_ = new_n25364_ & ~new_n25593_;
  assign new_n25595_ = ~new_n25588_ & ~new_n25594_;
  assign new_n25596_ = new_n25371_ & ~new_n25595_;
  assign new_n25597_ = ys__n2535 & ~new_n25595_;
  assign new_n25598_ = ~new_n25596_ & ~new_n25597_;
  assign new_n25599_ = ~new_n13708_ & ~new_n25598_;
  assign new_n25600_ = ys__n47077 & new_n25384_;
  assign new_n25601_ = ys__n47013 & new_n25386_;
  assign new_n25602_ = ~new_n25600_ & ~new_n25601_;
  assign new_n25603_ = ~new_n25389_ & ~new_n25602_;
  assign new_n25604_ = new_n25383_ & new_n25603_;
  assign new_n25605_ = new_n25261_ & ~new_n25328_;
  assign new_n25606_ = new_n25328_ & new_n25339_;
  assign new_n25607_ = ~new_n25328_ & ~new_n25339_;
  assign new_n25608_ = ~new_n25606_ & ~new_n25607_;
  assign new_n25609_ = ~new_n25261_ & ~new_n25608_;
  assign new_n25610_ = ~new_n25605_ & ~new_n25609_;
  assign new_n25611_ = ~new_n25383_ & ~new_n25610_;
  assign new_n25612_ = ~new_n25604_ & ~new_n25611_;
  assign new_n25613_ = new_n25399_ & ~new_n25612_;
  assign new_n25614_ = ys__n378 & ~new_n25399_;
  assign new_n25615_ = ~new_n25613_ & ~new_n25614_;
  assign new_n25616_ = new_n13708_ & ~new_n25615_;
  assign new_n25617_ = ~new_n25599_ & ~new_n25616_;
  assign new_n25618_ = ~ys__n1598 & ~new_n25617_;
  assign new_n25619_ = ys__n24750 & ys__n1598;
  assign ys__n24751 = new_n25618_ | new_n25619_;
  assign new_n25621_ = ys__n31031 & ys__n47030;
  assign new_n25622_ = new_n24614_ & new_n25621_;
  assign new_n25623_ = ys__n34738 & ys__n34740;
  assign new_n25624_ = ys__n34742 & new_n25623_;
  assign new_n25625_ = ~ys__n34738 & ~ys__n34740;
  assign new_n25626_ = ys__n34742 & new_n25625_;
  assign new_n25627_ = ~new_n25624_ & ~new_n25626_;
  assign new_n25628_ = ~ys__n34738 & ys__n34740;
  assign new_n25629_ = ~ys__n34742 & new_n25628_;
  assign new_n25630_ = ys__n34738 & ~ys__n34740;
  assign new_n25631_ = ~ys__n34742 & new_n25630_;
  assign new_n25632_ = ~new_n25629_ & ~new_n25631_;
  assign new_n25633_ = new_n25627_ & new_n25632_;
  assign new_n25634_ = ys__n34746 & ys__n34748;
  assign new_n25635_ = ys__n34744 & ys__n34748;
  assign new_n25636_ = ~new_n25548_ & ~new_n25635_;
  assign new_n25637_ = ~new_n25634_ & new_n25636_;
  assign new_n25638_ = new_n25633_ & ~new_n25637_;
  assign new_n25639_ = ~new_n25633_ & new_n25637_;
  assign new_n25640_ = ~new_n25638_ & ~new_n25639_;
  assign new_n25641_ = ~new_n25493_ & ~new_n25565_;
  assign new_n25642_ = ~new_n25496_ & new_n25641_;
  assign new_n25643_ = ~new_n25558_ & ~new_n25562_;
  assign new_n25644_ = ~new_n25565_ & new_n25566_;
  assign new_n25645_ = ~new_n25643_ & ~new_n25644_;
  assign new_n25646_ = ~new_n25642_ & new_n25645_;
  assign new_n25647_ = new_n25640_ & ~new_n25646_;
  assign new_n25648_ = ~new_n25640_ & new_n25646_;
  assign new_n25649_ = ~new_n25647_ & ~new_n25648_;
  assign new_n25650_ = new_n25354_ & ~new_n25649_;
  assign new_n25651_ = ~new_n25499_ & ~new_n25571_;
  assign new_n25652_ = new_n25501_ & new_n25651_;
  assign new_n25653_ = new_n25649_ & new_n25652_;
  assign new_n25654_ = ~new_n25649_ & ~new_n25652_;
  assign new_n25655_ = ~new_n25653_ & ~new_n25654_;
  assign new_n25656_ = ~new_n25354_ & ~new_n25655_;
  assign new_n25657_ = ~new_n25650_ & ~new_n25656_;
  assign new_n25658_ = ~new_n25358_ & ~new_n25657_;
  assign new_n25659_ = ~new_n25431_ & new_n25651_;
  assign new_n25660_ = new_n25649_ & new_n25659_;
  assign new_n25661_ = ~new_n25649_ & ~new_n25659_;
  assign new_n25662_ = ~new_n25660_ & ~new_n25661_;
  assign new_n25663_ = new_n25358_ & ~new_n25662_;
  assign new_n25664_ = ~new_n25658_ & ~new_n25663_;
  assign new_n25665_ = ~new_n24614_ & ~new_n25664_;
  assign new_n25666_ = ~new_n25622_ & ~new_n25665_;
  assign new_n25667_ = ~new_n25364_ & ~new_n25666_;
  assign new_n25668_ = ~new_n25014_ & new_n25073_;
  assign new_n25669_ = new_n25014_ & ~new_n25073_;
  assign new_n25670_ = ~new_n25668_ & ~new_n25669_;
  assign new_n25671_ = new_n25364_ & ~new_n25670_;
  assign new_n25672_ = ~new_n25667_ & ~new_n25671_;
  assign new_n25673_ = new_n25371_ & ~new_n25672_;
  assign new_n25674_ = ys__n2535 & ~new_n25672_;
  assign new_n25675_ = ~new_n25673_ & ~new_n25674_;
  assign new_n25676_ = ~new_n13708_ & ~new_n25675_;
  assign new_n25677_ = ys__n47078 & new_n25384_;
  assign new_n25678_ = ys__n47014 & new_n25386_;
  assign new_n25679_ = ~new_n25677_ & ~new_n25678_;
  assign new_n25680_ = ~new_n25389_ & ~new_n25679_;
  assign new_n25681_ = new_n25383_ & new_n25680_;
  assign new_n25682_ = new_n25261_ & ~new_n25319_;
  assign new_n25683_ = new_n25319_ & new_n25340_;
  assign new_n25684_ = ~new_n25319_ & ~new_n25340_;
  assign new_n25685_ = ~new_n25683_ & ~new_n25684_;
  assign new_n25686_ = ~new_n25261_ & ~new_n25685_;
  assign new_n25687_ = ~new_n25682_ & ~new_n25686_;
  assign new_n25688_ = ~new_n25383_ & ~new_n25687_;
  assign new_n25689_ = ~new_n25681_ & ~new_n25688_;
  assign new_n25690_ = new_n25399_ & ~new_n25689_;
  assign new_n25691_ = ys__n382 & ~new_n25399_;
  assign new_n25692_ = ~new_n25690_ & ~new_n25691_;
  assign new_n25693_ = new_n13708_ & ~new_n25692_;
  assign new_n25694_ = ~new_n25676_ & ~new_n25693_;
  assign new_n25695_ = ~ys__n1598 & ~new_n25694_;
  assign new_n25696_ = ys__n24753 & ys__n1598;
  assign ys__n24754 = new_n25695_ | new_n25696_;
  assign new_n25698_ = ys__n31031 & ys__n47031;
  assign new_n25699_ = new_n24614_ & new_n25698_;
  assign new_n25700_ = ys__n34732 & ys__n34734;
  assign new_n25701_ = ys__n34736 & new_n25700_;
  assign new_n25702_ = ~ys__n34732 & ~ys__n34734;
  assign new_n25703_ = ys__n34736 & new_n25702_;
  assign new_n25704_ = ~new_n25701_ & ~new_n25703_;
  assign new_n25705_ = ~ys__n34732 & ys__n34734;
  assign new_n25706_ = ~ys__n34736 & new_n25705_;
  assign new_n25707_ = ys__n34732 & ~ys__n34734;
  assign new_n25708_ = ~ys__n34736 & new_n25707_;
  assign new_n25709_ = ~new_n25706_ & ~new_n25708_;
  assign new_n25710_ = new_n25704_ & new_n25709_;
  assign new_n25711_ = ys__n34740 & ys__n34742;
  assign new_n25712_ = ys__n34738 & ys__n34742;
  assign new_n25713_ = ~new_n25623_ & ~new_n25712_;
  assign new_n25714_ = ~new_n25711_ & new_n25713_;
  assign new_n25715_ = new_n25710_ & ~new_n25714_;
  assign new_n25716_ = ~new_n25710_ & new_n25714_;
  assign new_n25717_ = ~new_n25715_ & ~new_n25716_;
  assign new_n25718_ = ~new_n25633_ & ~new_n25637_;
  assign new_n25719_ = ~new_n25640_ & ~new_n25646_;
  assign new_n25720_ = ~new_n25718_ & ~new_n25719_;
  assign new_n25721_ = new_n25717_ & ~new_n25720_;
  assign new_n25722_ = ~new_n25717_ & new_n25720_;
  assign new_n25723_ = ~new_n25721_ & ~new_n25722_;
  assign new_n25724_ = new_n25354_ & ~new_n25723_;
  assign new_n25725_ = ~new_n25649_ & new_n25652_;
  assign new_n25726_ = new_n25723_ & new_n25725_;
  assign new_n25727_ = ~new_n25723_ & ~new_n25725_;
  assign new_n25728_ = ~new_n25726_ & ~new_n25727_;
  assign new_n25729_ = ~new_n25354_ & ~new_n25728_;
  assign new_n25730_ = ~new_n25724_ & ~new_n25729_;
  assign new_n25731_ = ~new_n25358_ & ~new_n25730_;
  assign new_n25732_ = ~new_n25649_ & new_n25659_;
  assign new_n25733_ = new_n25723_ & new_n25732_;
  assign new_n25734_ = ~new_n25723_ & ~new_n25732_;
  assign new_n25735_ = ~new_n25733_ & ~new_n25734_;
  assign new_n25736_ = new_n25358_ & ~new_n25735_;
  assign new_n25737_ = ~new_n25731_ & ~new_n25736_;
  assign new_n25738_ = ~new_n24614_ & ~new_n25737_;
  assign new_n25739_ = ~new_n25699_ & ~new_n25738_;
  assign new_n25740_ = ~new_n25364_ & ~new_n25739_;
  assign new_n25741_ = ~new_n25014_ & ~new_n25073_;
  assign new_n25742_ = ~new_n25078_ & ~new_n25741_;
  assign new_n25743_ = new_n25066_ & ~new_n25742_;
  assign new_n25744_ = ~new_n25066_ & new_n25742_;
  assign new_n25745_ = ~new_n25743_ & ~new_n25744_;
  assign new_n25746_ = new_n25364_ & ~new_n25745_;
  assign new_n25747_ = ~new_n25740_ & ~new_n25746_;
  assign new_n25748_ = new_n25371_ & ~new_n25747_;
  assign new_n25749_ = ys__n2535 & ~new_n25747_;
  assign new_n25750_ = ~new_n25748_ & ~new_n25749_;
  assign new_n25751_ = ~new_n13708_ & ~new_n25750_;
  assign new_n25752_ = ys__n47079 & new_n25384_;
  assign new_n25753_ = ys__n47015 & new_n25386_;
  assign new_n25754_ = ~new_n25752_ & ~new_n25753_;
  assign new_n25755_ = ~new_n25389_ & ~new_n25754_;
  assign new_n25756_ = new_n25383_ & new_n25755_;
  assign new_n25757_ = new_n25261_ & ~new_n25316_;
  assign new_n25758_ = ~new_n25319_ & new_n25340_;
  assign new_n25759_ = new_n25316_ & new_n25758_;
  assign new_n25760_ = ~new_n25316_ & ~new_n25758_;
  assign new_n25761_ = ~new_n25759_ & ~new_n25760_;
  assign new_n25762_ = ~new_n25261_ & ~new_n25761_;
  assign new_n25763_ = ~new_n25757_ & ~new_n25762_;
  assign new_n25764_ = ~new_n25383_ & ~new_n25763_;
  assign new_n25765_ = ~new_n25756_ & ~new_n25764_;
  assign new_n25766_ = new_n25399_ & ~new_n25765_;
  assign new_n25767_ = ys__n374 & ~new_n25399_;
  assign new_n25768_ = ~new_n25766_ & ~new_n25767_;
  assign new_n25769_ = new_n13708_ & ~new_n25768_;
  assign new_n25770_ = ~new_n25751_ & ~new_n25769_;
  assign new_n25771_ = ~ys__n1598 & ~new_n25770_;
  assign new_n25772_ = ys__n24756 & ys__n1598;
  assign ys__n24757 = new_n25771_ | new_n25772_;
  assign new_n25774_ = ys__n31031 & ys__n47032;
  assign new_n25775_ = new_n24614_ & new_n25774_;
  assign new_n25776_ = ys__n34726 & ys__n34728;
  assign new_n25777_ = ys__n34730 & new_n25776_;
  assign new_n25778_ = ~ys__n34726 & ~ys__n34728;
  assign new_n25779_ = ys__n34730 & new_n25778_;
  assign new_n25780_ = ~new_n25777_ & ~new_n25779_;
  assign new_n25781_ = ~ys__n34726 & ys__n34728;
  assign new_n25782_ = ~ys__n34730 & new_n25781_;
  assign new_n25783_ = ys__n34726 & ~ys__n34728;
  assign new_n25784_ = ~ys__n34730 & new_n25783_;
  assign new_n25785_ = ~new_n25782_ & ~new_n25784_;
  assign new_n25786_ = new_n25780_ & new_n25785_;
  assign new_n25787_ = ys__n34734 & ys__n34736;
  assign new_n25788_ = ys__n34732 & ys__n34736;
  assign new_n25789_ = ~new_n25700_ & ~new_n25788_;
  assign new_n25790_ = ~new_n25787_ & new_n25789_;
  assign new_n25791_ = new_n25786_ & ~new_n25790_;
  assign new_n25792_ = ~new_n25786_ & new_n25790_;
  assign new_n25793_ = ~new_n25791_ & ~new_n25792_;
  assign new_n25794_ = ~new_n25710_ & ~new_n25714_;
  assign new_n25795_ = ~new_n25717_ & new_n25718_;
  assign new_n25796_ = ~new_n25794_ & ~new_n25795_;
  assign new_n25797_ = ~new_n25640_ & ~new_n25717_;
  assign new_n25798_ = ~new_n25646_ & new_n25797_;
  assign new_n25799_ = new_n25796_ & ~new_n25798_;
  assign new_n25800_ = new_n25793_ & ~new_n25799_;
  assign new_n25801_ = ~new_n25793_ & new_n25799_;
  assign new_n25802_ = ~new_n25800_ & ~new_n25801_;
  assign new_n25803_ = new_n25354_ & ~new_n25802_;
  assign new_n25804_ = ~new_n25649_ & ~new_n25723_;
  assign new_n25805_ = new_n25652_ & new_n25804_;
  assign new_n25806_ = new_n25802_ & new_n25805_;
  assign new_n25807_ = ~new_n25802_ & ~new_n25805_;
  assign new_n25808_ = ~new_n25806_ & ~new_n25807_;
  assign new_n25809_ = ~new_n25354_ & ~new_n25808_;
  assign new_n25810_ = ~new_n25803_ & ~new_n25809_;
  assign new_n25811_ = ~new_n25358_ & ~new_n25810_;
  assign new_n25812_ = new_n25659_ & new_n25804_;
  assign new_n25813_ = new_n25802_ & new_n25812_;
  assign new_n25814_ = ~new_n25802_ & ~new_n25812_;
  assign new_n25815_ = ~new_n25813_ & ~new_n25814_;
  assign new_n25816_ = new_n25358_ & ~new_n25815_;
  assign new_n25817_ = ~new_n25811_ & ~new_n25816_;
  assign new_n25818_ = ~new_n24614_ & ~new_n25817_;
  assign new_n25819_ = ~new_n25775_ & ~new_n25818_;
  assign new_n25820_ = ~new_n25364_ & ~new_n25819_;
  assign new_n25821_ = ~new_n25014_ & new_n25074_;
  assign new_n25822_ = new_n25080_ & ~new_n25821_;
  assign new_n25823_ = new_n25051_ & ~new_n25822_;
  assign new_n25824_ = ~new_n25051_ & new_n25822_;
  assign new_n25825_ = ~new_n25823_ & ~new_n25824_;
  assign new_n25826_ = new_n25364_ & ~new_n25825_;
  assign new_n25827_ = ~new_n25820_ & ~new_n25826_;
  assign new_n25828_ = new_n25371_ & ~new_n25827_;
  assign new_n25829_ = ys__n2535 & ~new_n25827_;
  assign new_n25830_ = ~new_n25828_ & ~new_n25829_;
  assign new_n25831_ = ~new_n13708_ & ~new_n25830_;
  assign new_n25832_ = ys__n47080 & new_n25384_;
  assign new_n25833_ = ys__n47016 & new_n25386_;
  assign new_n25834_ = ~new_n25832_ & ~new_n25833_;
  assign new_n25835_ = ~new_n25389_ & ~new_n25834_;
  assign new_n25836_ = new_n25383_ & new_n25835_;
  assign new_n25837_ = new_n25261_ & ~new_n25323_;
  assign new_n25838_ = new_n25320_ & new_n25340_;
  assign new_n25839_ = new_n25323_ & new_n25838_;
  assign new_n25840_ = ~new_n25323_ & ~new_n25838_;
  assign new_n25841_ = ~new_n25839_ & ~new_n25840_;
  assign new_n25842_ = ~new_n25261_ & ~new_n25841_;
  assign new_n25843_ = ~new_n25837_ & ~new_n25842_;
  assign new_n25844_ = ~new_n25383_ & ~new_n25843_;
  assign new_n25845_ = ~new_n25836_ & ~new_n25844_;
  assign new_n25846_ = new_n25399_ & ~new_n25845_;
  assign new_n25847_ = ys__n376 & ~new_n25399_;
  assign new_n25848_ = ~new_n25846_ & ~new_n25847_;
  assign new_n25849_ = new_n13708_ & ~new_n25848_;
  assign new_n25850_ = ~new_n25831_ & ~new_n25849_;
  assign new_n25851_ = ~ys__n1598 & ~new_n25850_;
  assign new_n25852_ = ys__n24759 & ys__n1598;
  assign ys__n24760 = new_n25851_ | new_n25852_;
  assign new_n25854_ = ys__n31031 & ys__n47033;
  assign new_n25855_ = new_n24614_ & new_n25854_;
  assign new_n25856_ = ys__n34720 & ys__n34722;
  assign new_n25857_ = ys__n34724 & new_n25856_;
  assign new_n25858_ = ~ys__n34720 & ~ys__n34722;
  assign new_n25859_ = ys__n34724 & new_n25858_;
  assign new_n25860_ = ~new_n25857_ & ~new_n25859_;
  assign new_n25861_ = ~ys__n34720 & ys__n34722;
  assign new_n25862_ = ~ys__n34724 & new_n25861_;
  assign new_n25863_ = ys__n34720 & ~ys__n34722;
  assign new_n25864_ = ~ys__n34724 & new_n25863_;
  assign new_n25865_ = ~new_n25862_ & ~new_n25864_;
  assign new_n25866_ = new_n25860_ & new_n25865_;
  assign new_n25867_ = ys__n34728 & ys__n34730;
  assign new_n25868_ = ys__n34726 & ys__n34730;
  assign new_n25869_ = ~new_n25776_ & ~new_n25868_;
  assign new_n25870_ = ~new_n25867_ & new_n25869_;
  assign new_n25871_ = new_n25866_ & ~new_n25870_;
  assign new_n25872_ = ~new_n25866_ & new_n25870_;
  assign new_n25873_ = ~new_n25871_ & ~new_n25872_;
  assign new_n25874_ = ~new_n25786_ & ~new_n25790_;
  assign new_n25875_ = ~new_n25793_ & ~new_n25799_;
  assign new_n25876_ = ~new_n25874_ & ~new_n25875_;
  assign new_n25877_ = new_n25873_ & ~new_n25876_;
  assign new_n25878_ = ~new_n25873_ & new_n25876_;
  assign new_n25879_ = ~new_n25877_ & ~new_n25878_;
  assign new_n25880_ = new_n25354_ & ~new_n25879_;
  assign new_n25881_ = ~new_n25802_ & new_n25805_;
  assign new_n25882_ = new_n25879_ & new_n25881_;
  assign new_n25883_ = ~new_n25879_ & ~new_n25881_;
  assign new_n25884_ = ~new_n25882_ & ~new_n25883_;
  assign new_n25885_ = ~new_n25354_ & ~new_n25884_;
  assign new_n25886_ = ~new_n25880_ & ~new_n25885_;
  assign new_n25887_ = ~new_n25358_ & ~new_n25886_;
  assign new_n25888_ = ~new_n25802_ & new_n25812_;
  assign new_n25889_ = new_n25879_ & new_n25888_;
  assign new_n25890_ = ~new_n25879_ & ~new_n25888_;
  assign new_n25891_ = ~new_n25889_ & ~new_n25890_;
  assign new_n25892_ = new_n25358_ & ~new_n25891_;
  assign new_n25893_ = ~new_n25887_ & ~new_n25892_;
  assign new_n25894_ = ~new_n24614_ & ~new_n25893_;
  assign new_n25895_ = ~new_n25855_ & ~new_n25894_;
  assign new_n25896_ = ~new_n25364_ & ~new_n25895_;
  assign new_n25897_ = ~new_n25051_ & ~new_n25822_;
  assign new_n25898_ = ~new_n25083_ & ~new_n25897_;
  assign new_n25899_ = new_n25033_ & ~new_n25898_;
  assign new_n25900_ = ~new_n25033_ & new_n25898_;
  assign new_n25901_ = ~new_n25899_ & ~new_n25900_;
  assign new_n25902_ = new_n25364_ & ~new_n25901_;
  assign new_n25903_ = ~new_n25896_ & ~new_n25902_;
  assign new_n25904_ = new_n25371_ & ~new_n25903_;
  assign new_n25905_ = ys__n2535 & ~new_n25903_;
  assign new_n25906_ = ~new_n25904_ & ~new_n25905_;
  assign new_n25907_ = ~new_n13708_ & ~new_n25906_;
  assign new_n25908_ = ys__n47081 & new_n25384_;
  assign new_n25909_ = ys__n47017 & new_n25386_;
  assign new_n25910_ = ~new_n25908_ & ~new_n25909_;
  assign new_n25911_ = ~new_n25389_ & ~new_n25910_;
  assign new_n25912_ = new_n25383_ & new_n25911_;
  assign new_n25913_ = new_n25261_ & ~new_n25311_;
  assign new_n25914_ = ~new_n25323_ & new_n25838_;
  assign new_n25915_ = new_n25311_ & new_n25914_;
  assign new_n25916_ = ~new_n25311_ & ~new_n25914_;
  assign new_n25917_ = ~new_n25915_ & ~new_n25916_;
  assign new_n25918_ = ~new_n25261_ & ~new_n25917_;
  assign new_n25919_ = ~new_n25913_ & ~new_n25918_;
  assign new_n25920_ = ~new_n25383_ & ~new_n25919_;
  assign new_n25921_ = ~new_n25912_ & ~new_n25920_;
  assign new_n25922_ = new_n25399_ & ~new_n25921_;
  assign new_n25923_ = ys__n372 & ~new_n25399_;
  assign new_n25924_ = ~new_n25922_ & ~new_n25923_;
  assign new_n25925_ = new_n13708_ & ~new_n25924_;
  assign new_n25926_ = ~new_n25907_ & ~new_n25925_;
  assign new_n25927_ = ~ys__n1598 & ~new_n25926_;
  assign new_n25928_ = ys__n24762 & ys__n1598;
  assign ys__n24763 = new_n25927_ | new_n25928_;
  assign new_n25930_ = ys__n31031 & ys__n47034;
  assign new_n25931_ = new_n24614_ & new_n25930_;
  assign new_n25932_ = ys__n34714 & ys__n34716;
  assign new_n25933_ = ys__n34718 & new_n25932_;
  assign new_n25934_ = ~ys__n34714 & ~ys__n34716;
  assign new_n25935_ = ys__n34718 & new_n25934_;
  assign new_n25936_ = ~new_n25933_ & ~new_n25935_;
  assign new_n25937_ = ~ys__n34714 & ys__n34716;
  assign new_n25938_ = ~ys__n34718 & new_n25937_;
  assign new_n25939_ = ys__n34714 & ~ys__n34716;
  assign new_n25940_ = ~ys__n34718 & new_n25939_;
  assign new_n25941_ = ~new_n25938_ & ~new_n25940_;
  assign new_n25942_ = new_n25936_ & new_n25941_;
  assign new_n25943_ = ys__n34722 & ys__n34724;
  assign new_n25944_ = ys__n34720 & ys__n34724;
  assign new_n25945_ = ~new_n25856_ & ~new_n25944_;
  assign new_n25946_ = ~new_n25943_ & new_n25945_;
  assign new_n25947_ = new_n25942_ & ~new_n25946_;
  assign new_n25948_ = ~new_n25942_ & new_n25946_;
  assign new_n25949_ = ~new_n25947_ & ~new_n25948_;
  assign new_n25950_ = ~new_n25793_ & ~new_n25873_;
  assign new_n25951_ = new_n25797_ & new_n25950_;
  assign new_n25952_ = ~new_n25646_ & new_n25951_;
  assign new_n25953_ = ~new_n25796_ & new_n25950_;
  assign new_n25954_ = ~new_n25866_ & ~new_n25870_;
  assign new_n25955_ = ~new_n25873_ & new_n25874_;
  assign new_n25956_ = ~new_n25954_ & ~new_n25955_;
  assign new_n25957_ = ~new_n25953_ & new_n25956_;
  assign new_n25958_ = ~new_n25952_ & new_n25957_;
  assign new_n25959_ = new_n25949_ & ~new_n25958_;
  assign new_n25960_ = ~new_n25949_ & new_n25958_;
  assign new_n25961_ = ~new_n25959_ & ~new_n25960_;
  assign new_n25962_ = new_n25354_ & ~new_n25961_;
  assign new_n25963_ = ~new_n25802_ & new_n25804_;
  assign new_n25964_ = ~new_n25879_ & new_n25963_;
  assign new_n25965_ = new_n25652_ & new_n25964_;
  assign new_n25966_ = new_n25961_ & new_n25965_;
  assign new_n25967_ = ~new_n25961_ & ~new_n25965_;
  assign new_n25968_ = ~new_n25966_ & ~new_n25967_;
  assign new_n25969_ = ~new_n25354_ & ~new_n25968_;
  assign new_n25970_ = ~new_n25962_ & ~new_n25969_;
  assign new_n25971_ = ~new_n25358_ & ~new_n25970_;
  assign new_n25972_ = new_n25659_ & new_n25964_;
  assign new_n25973_ = new_n25961_ & new_n25972_;
  assign new_n25974_ = ~new_n25961_ & ~new_n25972_;
  assign new_n25975_ = ~new_n25973_ & ~new_n25974_;
  assign new_n25976_ = new_n25358_ & ~new_n25975_;
  assign new_n25977_ = ~new_n25971_ & ~new_n25976_;
  assign new_n25978_ = ~new_n24614_ & ~new_n25977_;
  assign new_n25979_ = ~new_n25931_ & ~new_n25978_;
  assign new_n25980_ = ~new_n25364_ & ~new_n25979_;
  assign new_n25981_ = ~new_n25087_ & new_n25234_;
  assign new_n25982_ = new_n25087_ & ~new_n25234_;
  assign new_n25983_ = ~new_n25981_ & ~new_n25982_;
  assign new_n25984_ = new_n25364_ & ~new_n25983_;
  assign new_n25985_ = ~new_n25980_ & ~new_n25984_;
  assign new_n25986_ = new_n25371_ & ~new_n25985_;
  assign new_n25987_ = ys__n2535 & ~new_n25985_;
  assign new_n25988_ = ~new_n25986_ & ~new_n25987_;
  assign new_n25989_ = ~new_n13708_ & ~new_n25988_;
  assign new_n25990_ = ys__n47082 & new_n25384_;
  assign new_n25991_ = ys__n47018 & new_n25386_;
  assign new_n25992_ = ~new_n25990_ & ~new_n25991_;
  assign new_n25993_ = ~new_n25389_ & ~new_n25992_;
  assign new_n25994_ = new_n25383_ & new_n25993_;
  assign new_n25995_ = new_n25261_ & ~new_n25289_;
  assign new_n25996_ = new_n25289_ & new_n25343_;
  assign new_n25997_ = ~new_n25289_ & ~new_n25343_;
  assign new_n25998_ = ~new_n25996_ & ~new_n25997_;
  assign new_n25999_ = ~new_n25261_ & ~new_n25998_;
  assign new_n26000_ = ~new_n25995_ & ~new_n25999_;
  assign new_n26001_ = ~new_n25383_ & ~new_n26000_;
  assign new_n26002_ = ~new_n25994_ & ~new_n26001_;
  assign new_n26003_ = new_n25399_ & ~new_n26002_;
  assign new_n26004_ = ys__n384 & ~new_n25399_;
  assign new_n26005_ = ~new_n26003_ & ~new_n26004_;
  assign new_n26006_ = new_n13708_ & ~new_n26005_;
  assign new_n26007_ = ~new_n25989_ & ~new_n26006_;
  assign new_n26008_ = ~ys__n1598 & ~new_n26007_;
  assign new_n26009_ = ys__n24765 & ys__n1598;
  assign ys__n24766 = new_n26008_ | new_n26009_;
  assign new_n26011_ = ys__n31031 & ys__n47035;
  assign new_n26012_ = new_n24614_ & new_n26011_;
  assign new_n26013_ = ys__n34708 & ys__n34710;
  assign new_n26014_ = ys__n34712 & new_n26013_;
  assign new_n26015_ = ~ys__n34708 & ~ys__n34710;
  assign new_n26016_ = ys__n34712 & new_n26015_;
  assign new_n26017_ = ~new_n26014_ & ~new_n26016_;
  assign new_n26018_ = ~ys__n34708 & ys__n34710;
  assign new_n26019_ = ~ys__n34712 & new_n26018_;
  assign new_n26020_ = ys__n34708 & ~ys__n34710;
  assign new_n26021_ = ~ys__n34712 & new_n26020_;
  assign new_n26022_ = ~new_n26019_ & ~new_n26021_;
  assign new_n26023_ = new_n26017_ & new_n26022_;
  assign new_n26024_ = ys__n34716 & ys__n34718;
  assign new_n26025_ = ys__n34714 & ys__n34718;
  assign new_n26026_ = ~new_n25932_ & ~new_n26025_;
  assign new_n26027_ = ~new_n26024_ & new_n26026_;
  assign new_n26028_ = new_n26023_ & ~new_n26027_;
  assign new_n26029_ = ~new_n26023_ & new_n26027_;
  assign new_n26030_ = ~new_n26028_ & ~new_n26029_;
  assign new_n26031_ = ~new_n25942_ & ~new_n25946_;
  assign new_n26032_ = ~new_n25949_ & ~new_n25958_;
  assign new_n26033_ = ~new_n26031_ & ~new_n26032_;
  assign new_n26034_ = new_n26030_ & ~new_n26033_;
  assign new_n26035_ = ~new_n26030_ & new_n26033_;
  assign new_n26036_ = ~new_n26034_ & ~new_n26035_;
  assign new_n26037_ = new_n25354_ & ~new_n26036_;
  assign new_n26038_ = ~new_n25961_ & new_n25965_;
  assign new_n26039_ = new_n26036_ & new_n26038_;
  assign new_n26040_ = ~new_n26036_ & ~new_n26038_;
  assign new_n26041_ = ~new_n26039_ & ~new_n26040_;
  assign new_n26042_ = ~new_n25354_ & ~new_n26041_;
  assign new_n26043_ = ~new_n26037_ & ~new_n26042_;
  assign new_n26044_ = ~new_n25358_ & ~new_n26043_;
  assign new_n26045_ = ~new_n25961_ & new_n25972_;
  assign new_n26046_ = new_n26036_ & new_n26045_;
  assign new_n26047_ = ~new_n26036_ & ~new_n26045_;
  assign new_n26048_ = ~new_n26046_ & ~new_n26047_;
  assign new_n26049_ = new_n25358_ & ~new_n26048_;
  assign new_n26050_ = ~new_n26044_ & ~new_n26049_;
  assign new_n26051_ = ~new_n24614_ & ~new_n26050_;
  assign new_n26052_ = ~new_n26012_ & ~new_n26051_;
  assign new_n26053_ = ~new_n25364_ & ~new_n26052_;
  assign new_n26054_ = ~new_n25087_ & ~new_n25234_;
  assign new_n26055_ = ~new_n25240_ & ~new_n26054_;
  assign new_n26056_ = new_n25217_ & ~new_n26055_;
  assign new_n26057_ = ~new_n25217_ & new_n26055_;
  assign new_n26058_ = ~new_n26056_ & ~new_n26057_;
  assign new_n26059_ = new_n25364_ & ~new_n26058_;
  assign new_n26060_ = ~new_n26053_ & ~new_n26059_;
  assign new_n26061_ = new_n25371_ & ~new_n26060_;
  assign new_n26062_ = ys__n2535 & ~new_n26060_;
  assign new_n26063_ = ~new_n26061_ & ~new_n26062_;
  assign new_n26064_ = ~new_n13708_ & ~new_n26063_;
  assign new_n26065_ = ys__n47083 & new_n25384_;
  assign new_n26066_ = ys__n47019 & new_n25386_;
  assign new_n26067_ = ~new_n26065_ & ~new_n26066_;
  assign new_n26068_ = ~new_n25389_ & ~new_n26067_;
  assign new_n26069_ = new_n25383_ & new_n26068_;
  assign new_n26070_ = new_n25261_ & ~new_n25286_;
  assign new_n26071_ = ~new_n25289_ & new_n25343_;
  assign new_n26072_ = new_n25286_ & new_n26071_;
  assign new_n26073_ = ~new_n25286_ & ~new_n26071_;
  assign new_n26074_ = ~new_n26072_ & ~new_n26073_;
  assign new_n26075_ = ~new_n25261_ & ~new_n26074_;
  assign new_n26076_ = ~new_n26070_ & ~new_n26075_;
  assign new_n26077_ = ~new_n25383_ & ~new_n26076_;
  assign new_n26078_ = ~new_n26069_ & ~new_n26077_;
  assign new_n26079_ = new_n25399_ & ~new_n26078_;
  assign new_n26080_ = ys__n366 & ~new_n25399_;
  assign new_n26081_ = ~new_n26079_ & ~new_n26080_;
  assign new_n26082_ = new_n13708_ & ~new_n26081_;
  assign new_n26083_ = ~new_n26064_ & ~new_n26082_;
  assign new_n26084_ = ~ys__n1598 & ~new_n26083_;
  assign new_n26085_ = ys__n24768 & ys__n1598;
  assign ys__n24769 = new_n26084_ | new_n26085_;
  assign new_n26087_ = ys__n31031 & ys__n47036;
  assign new_n26088_ = new_n24614_ & new_n26087_;
  assign new_n26089_ = ys__n34702 & ys__n34704;
  assign new_n26090_ = ys__n34706 & new_n26089_;
  assign new_n26091_ = ~ys__n34702 & ~ys__n34704;
  assign new_n26092_ = ys__n34706 & new_n26091_;
  assign new_n26093_ = ~new_n26090_ & ~new_n26092_;
  assign new_n26094_ = ~ys__n34702 & ys__n34704;
  assign new_n26095_ = ~ys__n34706 & new_n26094_;
  assign new_n26096_ = ys__n34702 & ~ys__n34704;
  assign new_n26097_ = ~ys__n34706 & new_n26096_;
  assign new_n26098_ = ~new_n26095_ & ~new_n26097_;
  assign new_n26099_ = new_n26093_ & new_n26098_;
  assign new_n26100_ = ys__n34710 & ys__n34712;
  assign new_n26101_ = ys__n34708 & ys__n34712;
  assign new_n26102_ = ~new_n26013_ & ~new_n26101_;
  assign new_n26103_ = ~new_n26100_ & new_n26102_;
  assign new_n26104_ = new_n26099_ & ~new_n26103_;
  assign new_n26105_ = ~new_n26099_ & new_n26103_;
  assign new_n26106_ = ~new_n26104_ & ~new_n26105_;
  assign new_n26107_ = ~new_n26023_ & ~new_n26027_;
  assign new_n26108_ = ~new_n26030_ & new_n26031_;
  assign new_n26109_ = ~new_n26107_ & ~new_n26108_;
  assign new_n26110_ = ~new_n25949_ & ~new_n26030_;
  assign new_n26111_ = ~new_n25958_ & new_n26110_;
  assign new_n26112_ = new_n26109_ & ~new_n26111_;
  assign new_n26113_ = new_n26106_ & ~new_n26112_;
  assign new_n26114_ = ~new_n26106_ & new_n26112_;
  assign new_n26115_ = ~new_n26113_ & ~new_n26114_;
  assign new_n26116_ = new_n25354_ & ~new_n26115_;
  assign new_n26117_ = ~new_n25961_ & ~new_n26036_;
  assign new_n26118_ = new_n25965_ & new_n26117_;
  assign new_n26119_ = new_n26115_ & new_n26118_;
  assign new_n26120_ = ~new_n26115_ & ~new_n26118_;
  assign new_n26121_ = ~new_n26119_ & ~new_n26120_;
  assign new_n26122_ = ~new_n25354_ & ~new_n26121_;
  assign new_n26123_ = ~new_n26116_ & ~new_n26122_;
  assign new_n26124_ = ~new_n25358_ & ~new_n26123_;
  assign new_n26125_ = new_n25972_ & new_n26117_;
  assign new_n26126_ = new_n26115_ & new_n26125_;
  assign new_n26127_ = ~new_n26115_ & ~new_n26125_;
  assign new_n26128_ = ~new_n26126_ & ~new_n26127_;
  assign new_n26129_ = new_n25358_ & ~new_n26128_;
  assign new_n26130_ = ~new_n26124_ & ~new_n26129_;
  assign new_n26131_ = ~new_n24614_ & ~new_n26130_;
  assign new_n26132_ = ~new_n26088_ & ~new_n26131_;
  assign new_n26133_ = ~new_n25364_ & ~new_n26132_;
  assign new_n26134_ = ~new_n25087_ & new_n25235_;
  assign new_n26135_ = new_n25242_ & ~new_n26134_;
  assign new_n26136_ = new_n25198_ & ~new_n26135_;
  assign new_n26137_ = ~new_n25198_ & new_n26135_;
  assign new_n26138_ = ~new_n26136_ & ~new_n26137_;
  assign new_n26139_ = new_n25364_ & ~new_n26138_;
  assign new_n26140_ = ~new_n26133_ & ~new_n26139_;
  assign new_n26141_ = new_n25371_ & ~new_n26140_;
  assign new_n26142_ = ys__n2535 & ~new_n26140_;
  assign new_n26143_ = ~new_n26141_ & ~new_n26142_;
  assign new_n26144_ = ~new_n13708_ & ~new_n26143_;
  assign new_n26145_ = ys__n47084 & new_n25384_;
  assign new_n26146_ = ys__n47020 & new_n25386_;
  assign new_n26147_ = ~new_n26145_ & ~new_n26146_;
  assign new_n26148_ = ~new_n25389_ & ~new_n26147_;
  assign new_n26149_ = new_n25383_ & new_n26148_;
  assign new_n26150_ = new_n25261_ & ~new_n25281_;
  assign new_n26151_ = new_n25290_ & new_n25343_;
  assign new_n26152_ = new_n25281_ & new_n26151_;
  assign new_n26153_ = ~new_n25281_ & ~new_n26151_;
  assign new_n26154_ = ~new_n26152_ & ~new_n26153_;
  assign new_n26155_ = ~new_n25261_ & ~new_n26154_;
  assign new_n26156_ = ~new_n26150_ & ~new_n26155_;
  assign new_n26157_ = ~new_n25383_ & ~new_n26156_;
  assign new_n26158_ = ~new_n26149_ & ~new_n26157_;
  assign new_n26159_ = new_n25399_ & ~new_n26158_;
  assign new_n26160_ = ys__n368 & ~new_n25399_;
  assign new_n26161_ = ~new_n26159_ & ~new_n26160_;
  assign new_n26162_ = new_n13708_ & ~new_n26161_;
  assign new_n26163_ = ~new_n26144_ & ~new_n26162_;
  assign new_n26164_ = ~ys__n1598 & ~new_n26163_;
  assign new_n26165_ = ys__n24771 & ys__n1598;
  assign ys__n24772 = new_n26164_ | new_n26165_;
  assign new_n26167_ = ys__n31031 & ys__n47037;
  assign new_n26168_ = new_n24614_ & new_n26167_;
  assign new_n26169_ = ys__n34696 & ys__n34698;
  assign new_n26170_ = ys__n34700 & new_n26169_;
  assign new_n26171_ = ~ys__n34696 & ~ys__n34698;
  assign new_n26172_ = ys__n34700 & new_n26171_;
  assign new_n26173_ = ~new_n26170_ & ~new_n26172_;
  assign new_n26174_ = ~ys__n34696 & ys__n34698;
  assign new_n26175_ = ~ys__n34700 & new_n26174_;
  assign new_n26176_ = ys__n34696 & ~ys__n34698;
  assign new_n26177_ = ~ys__n34700 & new_n26176_;
  assign new_n26178_ = ~new_n26175_ & ~new_n26177_;
  assign new_n26179_ = new_n26173_ & new_n26178_;
  assign new_n26180_ = ys__n34704 & ys__n34706;
  assign new_n26181_ = ys__n34702 & ys__n34706;
  assign new_n26182_ = ~new_n26089_ & ~new_n26181_;
  assign new_n26183_ = ~new_n26180_ & new_n26182_;
  assign new_n26184_ = new_n26179_ & ~new_n26183_;
  assign new_n26185_ = ~new_n26179_ & new_n26183_;
  assign new_n26186_ = ~new_n26184_ & ~new_n26185_;
  assign new_n26187_ = ~new_n26099_ & ~new_n26103_;
  assign new_n26188_ = ~new_n26106_ & ~new_n26112_;
  assign new_n26189_ = ~new_n26187_ & ~new_n26188_;
  assign new_n26190_ = new_n26186_ & ~new_n26189_;
  assign new_n26191_ = ~new_n26186_ & new_n26189_;
  assign new_n26192_ = ~new_n26190_ & ~new_n26191_;
  assign new_n26193_ = new_n25354_ & ~new_n26192_;
  assign new_n26194_ = ~new_n26115_ & new_n26118_;
  assign new_n26195_ = new_n26192_ & new_n26194_;
  assign new_n26196_ = ~new_n26192_ & ~new_n26194_;
  assign new_n26197_ = ~new_n26195_ & ~new_n26196_;
  assign new_n26198_ = ~new_n25354_ & ~new_n26197_;
  assign new_n26199_ = ~new_n26193_ & ~new_n26198_;
  assign new_n26200_ = ~new_n25358_ & ~new_n26199_;
  assign new_n26201_ = ~new_n26115_ & new_n26125_;
  assign new_n26202_ = new_n26192_ & new_n26201_;
  assign new_n26203_ = ~new_n26192_ & ~new_n26201_;
  assign new_n26204_ = ~new_n26202_ & ~new_n26203_;
  assign new_n26205_ = new_n25358_ & ~new_n26204_;
  assign new_n26206_ = ~new_n26200_ & ~new_n26205_;
  assign new_n26207_ = ~new_n24614_ & ~new_n26206_;
  assign new_n26208_ = ~new_n26168_ & ~new_n26207_;
  assign new_n26209_ = ~new_n25364_ & ~new_n26208_;
  assign new_n26210_ = ~new_n25198_ & ~new_n26135_;
  assign new_n26211_ = ~new_n25245_ & ~new_n26210_;
  assign new_n26212_ = new_n25180_ & ~new_n26211_;
  assign new_n26213_ = ~new_n25180_ & new_n26211_;
  assign new_n26214_ = ~new_n26212_ & ~new_n26213_;
  assign new_n26215_ = new_n25364_ & ~new_n26214_;
  assign new_n26216_ = ~new_n26209_ & ~new_n26215_;
  assign new_n26217_ = new_n25371_ & ~new_n26216_;
  assign new_n26218_ = ys__n2535 & ~new_n26216_;
  assign new_n26219_ = ~new_n26217_ & ~new_n26218_;
  assign new_n26220_ = ~new_n13708_ & ~new_n26219_;
  assign new_n26221_ = ys__n47085 & new_n25384_;
  assign new_n26222_ = ys__n47021 & new_n25386_;
  assign new_n26223_ = ~new_n26221_ & ~new_n26222_;
  assign new_n26224_ = ~new_n25389_ & ~new_n26223_;
  assign new_n26225_ = new_n25383_ & new_n26224_;
  assign new_n26226_ = new_n25261_ & ~new_n25278_;
  assign new_n26227_ = ~new_n25281_ & new_n26151_;
  assign new_n26228_ = new_n25278_ & new_n26227_;
  assign new_n26229_ = ~new_n25278_ & ~new_n26227_;
  assign new_n26230_ = ~new_n26228_ & ~new_n26229_;
  assign new_n26231_ = ~new_n25261_ & ~new_n26230_;
  assign new_n26232_ = ~new_n26226_ & ~new_n26231_;
  assign new_n26233_ = ~new_n25383_ & ~new_n26232_;
  assign new_n26234_ = ~new_n26225_ & ~new_n26233_;
  assign new_n26235_ = new_n25399_ & ~new_n26234_;
  assign new_n26236_ = ys__n364 & ~new_n25399_;
  assign new_n26237_ = ~new_n26235_ & ~new_n26236_;
  assign new_n26238_ = new_n13708_ & ~new_n26237_;
  assign new_n26239_ = ~new_n26220_ & ~new_n26238_;
  assign new_n26240_ = ~ys__n1598 & ~new_n26239_;
  assign new_n26241_ = ys__n24774 & ys__n1598;
  assign ys__n24775 = new_n26240_ | new_n26241_;
  assign new_n26243_ = ys__n31031 & ys__n47038;
  assign new_n26244_ = new_n24614_ & new_n26243_;
  assign new_n26245_ = ys__n34690 & ys__n34692;
  assign new_n26246_ = ys__n34694 & new_n26245_;
  assign new_n26247_ = ~ys__n34690 & ~ys__n34692;
  assign new_n26248_ = ys__n34694 & new_n26247_;
  assign new_n26249_ = ~new_n26246_ & ~new_n26248_;
  assign new_n26250_ = ~ys__n34690 & ys__n34692;
  assign new_n26251_ = ~ys__n34694 & new_n26250_;
  assign new_n26252_ = ys__n34690 & ~ys__n34692;
  assign new_n26253_ = ~ys__n34694 & new_n26252_;
  assign new_n26254_ = ~new_n26251_ & ~new_n26253_;
  assign new_n26255_ = new_n26249_ & new_n26254_;
  assign new_n26256_ = ys__n34698 & ys__n34700;
  assign new_n26257_ = ys__n34696 & ys__n34700;
  assign new_n26258_ = ~new_n26169_ & ~new_n26257_;
  assign new_n26259_ = ~new_n26256_ & new_n26258_;
  assign new_n26260_ = new_n26255_ & ~new_n26259_;
  assign new_n26261_ = ~new_n26255_ & new_n26259_;
  assign new_n26262_ = ~new_n26260_ & ~new_n26261_;
  assign new_n26263_ = ~new_n26106_ & ~new_n26186_;
  assign new_n26264_ = new_n26110_ & new_n26263_;
  assign new_n26265_ = ~new_n25958_ & new_n26264_;
  assign new_n26266_ = ~new_n26109_ & new_n26263_;
  assign new_n26267_ = ~new_n26179_ & ~new_n26183_;
  assign new_n26268_ = ~new_n26186_ & new_n26187_;
  assign new_n26269_ = ~new_n26267_ & ~new_n26268_;
  assign new_n26270_ = ~new_n26266_ & new_n26269_;
  assign new_n26271_ = ~new_n26265_ & new_n26270_;
  assign new_n26272_ = new_n26262_ & ~new_n26271_;
  assign new_n26273_ = ~new_n26262_ & new_n26271_;
  assign new_n26274_ = ~new_n26272_ & ~new_n26273_;
  assign new_n26275_ = new_n25354_ & ~new_n26274_;
  assign new_n26276_ = ~new_n26115_ & new_n26117_;
  assign new_n26277_ = ~new_n26192_ & new_n26276_;
  assign new_n26278_ = new_n25965_ & new_n26277_;
  assign new_n26279_ = new_n26274_ & new_n26278_;
  assign new_n26280_ = ~new_n26274_ & ~new_n26278_;
  assign new_n26281_ = ~new_n26279_ & ~new_n26280_;
  assign new_n26282_ = ~new_n25354_ & ~new_n26281_;
  assign new_n26283_ = ~new_n26275_ & ~new_n26282_;
  assign new_n26284_ = ~new_n25358_ & ~new_n26283_;
  assign new_n26285_ = new_n25972_ & new_n26277_;
  assign new_n26286_ = new_n26274_ & new_n26285_;
  assign new_n26287_ = ~new_n26274_ & ~new_n26285_;
  assign new_n26288_ = ~new_n26286_ & ~new_n26287_;
  assign new_n26289_ = new_n25358_ & ~new_n26288_;
  assign new_n26290_ = ~new_n26284_ & ~new_n26289_;
  assign new_n26291_ = ~new_n24614_ & ~new_n26290_;
  assign new_n26292_ = ~new_n26244_ & ~new_n26291_;
  assign new_n26293_ = ~new_n25364_ & ~new_n26292_;
  assign new_n26294_ = ~new_n25087_ & new_n25236_;
  assign new_n26295_ = new_n25248_ & ~new_n26294_;
  assign new_n26296_ = new_n25160_ & ~new_n26295_;
  assign new_n26297_ = ~new_n25160_ & new_n26295_;
  assign new_n26298_ = ~new_n26296_ & ~new_n26297_;
  assign new_n26299_ = new_n25364_ & ~new_n26298_;
  assign new_n26300_ = ~new_n26293_ & ~new_n26299_;
  assign new_n26301_ = new_n25371_ & ~new_n26300_;
  assign new_n26302_ = ys__n2535 & ~new_n26300_;
  assign new_n26303_ = ~new_n26301_ & ~new_n26302_;
  assign new_n26304_ = ~new_n13708_ & ~new_n26303_;
  assign new_n26305_ = ys__n47086 & new_n25384_;
  assign new_n26306_ = ys__n47022 & new_n25386_;
  assign new_n26307_ = ~new_n26305_ & ~new_n26306_;
  assign new_n26308_ = ~new_n25389_ & ~new_n26307_;
  assign new_n26309_ = new_n25383_ & new_n26308_;
  assign new_n26310_ = new_n25261_ & ~new_n25300_;
  assign new_n26311_ = new_n25292_ & new_n25343_;
  assign new_n26312_ = new_n25300_ & new_n26311_;
  assign new_n26313_ = ~new_n25300_ & ~new_n26311_;
  assign new_n26314_ = ~new_n26312_ & ~new_n26313_;
  assign new_n26315_ = ~new_n25261_ & ~new_n26314_;
  assign new_n26316_ = ~new_n26310_ & ~new_n26315_;
  assign new_n26317_ = ~new_n25383_ & ~new_n26316_;
  assign new_n26318_ = ~new_n26309_ & ~new_n26317_;
  assign new_n26319_ = new_n25399_ & ~new_n26318_;
  assign new_n26320_ = ys__n370 & ~new_n25399_;
  assign new_n26321_ = ~new_n26319_ & ~new_n26320_;
  assign new_n26322_ = new_n13708_ & ~new_n26321_;
  assign new_n26323_ = ~new_n26304_ & ~new_n26322_;
  assign new_n26324_ = ~ys__n1598 & ~new_n26323_;
  assign new_n26325_ = ys__n24777 & ys__n1598;
  assign ys__n24778 = new_n26324_ | new_n26325_;
  assign new_n26327_ = ys__n31031 & ys__n47039;
  assign new_n26328_ = new_n24614_ & new_n26327_;
  assign new_n26329_ = ys__n34684 & ys__n34686;
  assign new_n26330_ = ys__n34688 & new_n26329_;
  assign new_n26331_ = ~ys__n34684 & ~ys__n34686;
  assign new_n26332_ = ys__n34688 & new_n26331_;
  assign new_n26333_ = ~new_n26330_ & ~new_n26332_;
  assign new_n26334_ = ~ys__n34684 & ys__n34686;
  assign new_n26335_ = ~ys__n34688 & new_n26334_;
  assign new_n26336_ = ys__n34684 & ~ys__n34686;
  assign new_n26337_ = ~ys__n34688 & new_n26336_;
  assign new_n26338_ = ~new_n26335_ & ~new_n26337_;
  assign new_n26339_ = new_n26333_ & new_n26338_;
  assign new_n26340_ = ys__n34692 & ys__n34694;
  assign new_n26341_ = ys__n34690 & ys__n34694;
  assign new_n26342_ = ~new_n26245_ & ~new_n26341_;
  assign new_n26343_ = ~new_n26340_ & new_n26342_;
  assign new_n26344_ = new_n26339_ & ~new_n26343_;
  assign new_n26345_ = ~new_n26339_ & new_n26343_;
  assign new_n26346_ = ~new_n26344_ & ~new_n26345_;
  assign new_n26347_ = ~new_n26255_ & ~new_n26259_;
  assign new_n26348_ = ~new_n26262_ & ~new_n26271_;
  assign new_n26349_ = ~new_n26347_ & ~new_n26348_;
  assign new_n26350_ = new_n26346_ & ~new_n26349_;
  assign new_n26351_ = ~new_n26346_ & new_n26349_;
  assign new_n26352_ = ~new_n26350_ & ~new_n26351_;
  assign new_n26353_ = new_n25354_ & ~new_n26352_;
  assign new_n26354_ = ~new_n26274_ & new_n26278_;
  assign new_n26355_ = new_n26352_ & new_n26354_;
  assign new_n26356_ = ~new_n26352_ & ~new_n26354_;
  assign new_n26357_ = ~new_n26355_ & ~new_n26356_;
  assign new_n26358_ = ~new_n25354_ & ~new_n26357_;
  assign new_n26359_ = ~new_n26353_ & ~new_n26358_;
  assign new_n26360_ = ~new_n25358_ & ~new_n26359_;
  assign new_n26361_ = ~new_n26274_ & new_n26285_;
  assign new_n26362_ = new_n26352_ & new_n26361_;
  assign new_n26363_ = ~new_n26352_ & ~new_n26361_;
  assign new_n26364_ = ~new_n26362_ & ~new_n26363_;
  assign new_n26365_ = new_n25358_ & ~new_n26364_;
  assign new_n26366_ = ~new_n26360_ & ~new_n26365_;
  assign new_n26367_ = ~new_n24614_ & ~new_n26366_;
  assign new_n26368_ = ~new_n26328_ & ~new_n26367_;
  assign new_n26369_ = ~new_n25364_ & ~new_n26368_;
  assign new_n26370_ = ~new_n25160_ & ~new_n26295_;
  assign new_n26371_ = ~new_n25251_ & ~new_n26370_;
  assign new_n26372_ = new_n25142_ & ~new_n26371_;
  assign new_n26373_ = ~new_n25142_ & new_n26371_;
  assign new_n26374_ = ~new_n26372_ & ~new_n26373_;
  assign new_n26375_ = new_n25364_ & ~new_n26374_;
  assign new_n26376_ = ~new_n26369_ & ~new_n26375_;
  assign new_n26377_ = new_n25371_ & ~new_n26376_;
  assign new_n26378_ = ys__n2535 & ~new_n26376_;
  assign new_n26379_ = ~new_n26377_ & ~new_n26378_;
  assign new_n26380_ = ~new_n13708_ & ~new_n26379_;
  assign new_n26381_ = ys__n47087 & new_n25384_;
  assign new_n26382_ = ys__n47023 & new_n25386_;
  assign new_n26383_ = ~new_n26381_ & ~new_n26382_;
  assign new_n26384_ = ~new_n25389_ & ~new_n26383_;
  assign new_n26385_ = new_n25383_ & new_n26384_;
  assign new_n26386_ = new_n25261_ & ~new_n25297_;
  assign new_n26387_ = ~new_n25300_ & new_n26311_;
  assign new_n26388_ = new_n25297_ & new_n26387_;
  assign new_n26389_ = ~new_n25297_ & ~new_n26387_;
  assign new_n26390_ = ~new_n26388_ & ~new_n26389_;
  assign new_n26391_ = ~new_n25261_ & ~new_n26390_;
  assign new_n26392_ = ~new_n26386_ & ~new_n26391_;
  assign new_n26393_ = ~new_n25383_ & ~new_n26392_;
  assign new_n26394_ = ~new_n26385_ & ~new_n26393_;
  assign new_n26395_ = new_n25399_ & ~new_n26394_;
  assign new_n26396_ = ys__n360 & ~new_n25399_;
  assign new_n26397_ = ~new_n26395_ & ~new_n26396_;
  assign new_n26398_ = new_n13708_ & ~new_n26397_;
  assign new_n26399_ = ~new_n26380_ & ~new_n26398_;
  assign new_n26400_ = ~ys__n1598 & ~new_n26399_;
  assign new_n26401_ = ys__n24780 & ys__n1598;
  assign ys__n24781 = new_n26400_ | new_n26401_;
  assign new_n26403_ = ys__n31031 & ys__n47040;
  assign new_n26404_ = new_n24614_ & new_n26403_;
  assign new_n26405_ = ys__n34678 & ys__n34680;
  assign new_n26406_ = ys__n34682 & new_n26405_;
  assign new_n26407_ = ~ys__n34678 & ~ys__n34680;
  assign new_n26408_ = ys__n34682 & new_n26407_;
  assign new_n26409_ = ~new_n26406_ & ~new_n26408_;
  assign new_n26410_ = ~ys__n34678 & ys__n34680;
  assign new_n26411_ = ~ys__n34682 & new_n26410_;
  assign new_n26412_ = ys__n34678 & ~ys__n34680;
  assign new_n26413_ = ~ys__n34682 & new_n26412_;
  assign new_n26414_ = ~new_n26411_ & ~new_n26413_;
  assign new_n26415_ = new_n26409_ & new_n26414_;
  assign new_n26416_ = ys__n34686 & ys__n34688;
  assign new_n26417_ = ys__n34684 & ys__n34688;
  assign new_n26418_ = ~new_n26329_ & ~new_n26417_;
  assign new_n26419_ = ~new_n26416_ & new_n26418_;
  assign new_n26420_ = new_n26415_ & ~new_n26419_;
  assign new_n26421_ = ~new_n26415_ & new_n26419_;
  assign new_n26422_ = ~new_n26420_ & ~new_n26421_;
  assign new_n26423_ = ~new_n26262_ & ~new_n26346_;
  assign new_n26424_ = ~new_n26271_ & new_n26423_;
  assign new_n26425_ = ~new_n26339_ & ~new_n26343_;
  assign new_n26426_ = ~new_n26346_ & new_n26347_;
  assign new_n26427_ = ~new_n26425_ & ~new_n26426_;
  assign new_n26428_ = ~new_n26424_ & new_n26427_;
  assign new_n26429_ = new_n26422_ & ~new_n26428_;
  assign new_n26430_ = ~new_n26422_ & new_n26428_;
  assign new_n26431_ = ~new_n26429_ & ~new_n26430_;
  assign new_n26432_ = new_n25354_ & ~new_n26431_;
  assign new_n26433_ = ~new_n26274_ & ~new_n26352_;
  assign new_n26434_ = new_n26278_ & new_n26433_;
  assign new_n26435_ = new_n26431_ & new_n26434_;
  assign new_n26436_ = ~new_n26431_ & ~new_n26434_;
  assign new_n26437_ = ~new_n26435_ & ~new_n26436_;
  assign new_n26438_ = ~new_n25354_ & ~new_n26437_;
  assign new_n26439_ = ~new_n26432_ & ~new_n26438_;
  assign new_n26440_ = ~new_n25358_ & ~new_n26439_;
  assign new_n26441_ = new_n26285_ & new_n26433_;
  assign new_n26442_ = new_n26431_ & new_n26441_;
  assign new_n26443_ = ~new_n26431_ & ~new_n26441_;
  assign new_n26444_ = ~new_n26442_ & ~new_n26443_;
  assign new_n26445_ = new_n25358_ & ~new_n26444_;
  assign new_n26446_ = ~new_n26440_ & ~new_n26445_;
  assign new_n26447_ = ~new_n24614_ & ~new_n26446_;
  assign new_n26448_ = ~new_n26404_ & ~new_n26447_;
  assign new_n26449_ = ~new_n25364_ & ~new_n26448_;
  assign new_n26450_ = new_n25161_ & ~new_n26295_;
  assign new_n26451_ = new_n25253_ & ~new_n26450_;
  assign new_n26452_ = new_n25123_ & ~new_n26451_;
  assign new_n26453_ = ~new_n25123_ & new_n26451_;
  assign new_n26454_ = ~new_n26452_ & ~new_n26453_;
  assign new_n26455_ = new_n25364_ & ~new_n26454_;
  assign new_n26456_ = ~new_n26449_ & ~new_n26455_;
  assign new_n26457_ = new_n25371_ & ~new_n26456_;
  assign new_n26458_ = ys__n2535 & ~new_n26456_;
  assign new_n26459_ = ~new_n26457_ & ~new_n26458_;
  assign new_n26460_ = ~new_n13708_ & ~new_n26459_;
  assign new_n26461_ = ys__n47088 & new_n25384_;
  assign new_n26462_ = ys__n47024 & new_n25386_;
  assign new_n26463_ = ~new_n26461_ & ~new_n26462_;
  assign new_n26464_ = ~new_n25389_ & ~new_n26463_;
  assign new_n26465_ = new_n25383_ & new_n26464_;
  assign new_n26466_ = new_n25261_ & ~new_n25304_;
  assign new_n26467_ = new_n25301_ & new_n26311_;
  assign new_n26468_ = new_n25304_ & new_n26467_;
  assign new_n26469_ = ~new_n25304_ & ~new_n26467_;
  assign new_n26470_ = ~new_n26468_ & ~new_n26469_;
  assign new_n26471_ = ~new_n25261_ & ~new_n26470_;
  assign new_n26472_ = ~new_n26466_ & ~new_n26471_;
  assign new_n26473_ = ~new_n25383_ & ~new_n26472_;
  assign new_n26474_ = ~new_n26465_ & ~new_n26473_;
  assign new_n26475_ = new_n25399_ & ~new_n26474_;
  assign new_n26476_ = ys__n362 & ~new_n25399_;
  assign new_n26477_ = ~new_n26475_ & ~new_n26476_;
  assign new_n26478_ = new_n13708_ & ~new_n26477_;
  assign new_n26479_ = ~new_n26460_ & ~new_n26478_;
  assign new_n26480_ = ~ys__n1598 & ~new_n26479_;
  assign new_n26481_ = ys__n24783 & ys__n1598;
  assign ys__n24784 = new_n26480_ | new_n26481_;
  assign new_n26483_ = ys__n31031 & ys__n47041;
  assign new_n26484_ = new_n24614_ & new_n26483_;
  assign new_n26485_ = ~ys__n34674 & ys__n34676;
  assign new_n26486_ = ys__n34674 & ~ys__n34676;
  assign new_n26487_ = ~new_n26485_ & ~new_n26486_;
  assign new_n26488_ = ys__n34680 & ys__n34682;
  assign new_n26489_ = ys__n34678 & ys__n34682;
  assign new_n26490_ = ~new_n26405_ & ~new_n26489_;
  assign new_n26491_ = ~new_n26488_ & new_n26490_;
  assign new_n26492_ = new_n26487_ & ~new_n26491_;
  assign new_n26493_ = ~new_n26487_ & new_n26491_;
  assign new_n26494_ = ~new_n26492_ & ~new_n26493_;
  assign new_n26495_ = ~ys__n48324 & ~new_n26494_;
  assign new_n26496_ = ys__n48324 & new_n26494_;
  assign new_n26497_ = ~new_n26495_ & ~new_n26496_;
  assign new_n26498_ = ~new_n26415_ & ~new_n26419_;
  assign new_n26499_ = ~new_n26422_ & ~new_n26428_;
  assign new_n26500_ = ~new_n26498_ & ~new_n26499_;
  assign new_n26501_ = new_n25354_ & ~new_n26500_;
  assign new_n26502_ = ~new_n26431_ & new_n26434_;
  assign new_n26503_ = new_n26500_ & new_n26502_;
  assign new_n26504_ = ~new_n26500_ & ~new_n26502_;
  assign new_n26505_ = ~new_n26503_ & ~new_n26504_;
  assign new_n26506_ = ~new_n25354_ & ~new_n26505_;
  assign new_n26507_ = ~new_n26501_ & ~new_n26506_;
  assign new_n26508_ = ~new_n25358_ & ~new_n26507_;
  assign new_n26509_ = ~new_n26431_ & new_n26441_;
  assign new_n26510_ = new_n26500_ & new_n26509_;
  assign new_n26511_ = ~new_n26500_ & ~new_n26509_;
  assign new_n26512_ = ~new_n26510_ & ~new_n26511_;
  assign new_n26513_ = new_n25358_ & ~new_n26512_;
  assign new_n26514_ = ~new_n26508_ & ~new_n26513_;
  assign new_n26515_ = ~new_n26497_ & new_n26514_;
  assign new_n26516_ = ~ys__n48324 & new_n26494_;
  assign new_n26517_ = ys__n48324 & ~new_n26494_;
  assign new_n26518_ = ~new_n26516_ & ~new_n26517_;
  assign new_n26519_ = ~new_n26514_ & ~new_n26518_;
  assign new_n26520_ = ~new_n26515_ & ~new_n26519_;
  assign new_n26521_ = ~new_n24614_ & ~new_n26520_;
  assign new_n26522_ = ~new_n26484_ & ~new_n26521_;
  assign new_n26523_ = ~new_n25364_ & ~new_n26522_;
  assign new_n26524_ = ~new_n25123_ & ~new_n26451_;
  assign new_n26525_ = ~new_n25256_ & ~new_n26524_;
  assign new_n26526_ = new_n25105_ & ~new_n26525_;
  assign new_n26527_ = ~new_n25105_ & new_n26525_;
  assign new_n26528_ = ~new_n26526_ & ~new_n26527_;
  assign new_n26529_ = new_n25364_ & ~new_n26528_;
  assign new_n26530_ = ~new_n26523_ & ~new_n26529_;
  assign new_n26531_ = new_n25371_ & ~new_n26530_;
  assign new_n26532_ = ys__n2535 & ~new_n26530_;
  assign new_n26533_ = ~new_n26531_ & ~new_n26532_;
  assign new_n26534_ = ~new_n13708_ & ~new_n26533_;
  assign new_n26535_ = ys__n47089 & new_n25384_;
  assign new_n26536_ = ys__n47025 & new_n25386_;
  assign new_n26537_ = ~new_n26535_ & ~new_n26536_;
  assign new_n26538_ = ~new_n25389_ & ~new_n26537_;
  assign new_n26539_ = new_n25383_ & new_n26538_;
  assign new_n26540_ = new_n25261_ & ~new_n25271_;
  assign new_n26541_ = ~new_n25304_ & new_n26467_;
  assign new_n26542_ = new_n25271_ & new_n26541_;
  assign new_n26543_ = ~new_n25271_ & ~new_n26541_;
  assign new_n26544_ = ~new_n26542_ & ~new_n26543_;
  assign new_n26545_ = ~new_n25261_ & ~new_n26544_;
  assign new_n26546_ = ~new_n26540_ & ~new_n26545_;
  assign new_n26547_ = ~new_n25383_ & ~new_n26546_;
  assign new_n26548_ = ~new_n26539_ & ~new_n26547_;
  assign new_n26549_ = new_n25399_ & ~new_n26548_;
  assign new_n26550_ = ys__n358 & ~new_n25399_;
  assign new_n26551_ = ~new_n26549_ & ~new_n26550_;
  assign new_n26552_ = new_n13708_ & ~new_n26551_;
  assign new_n26553_ = ~new_n26534_ & ~new_n26552_;
  assign new_n26554_ = ~ys__n1598 & ~new_n26553_;
  assign new_n26555_ = ys__n24786 & ys__n1598;
  assign ys__n24787 = new_n26554_ | new_n26555_;
  assign new_n26557_ = ~ys__n34670 & ys__n34672;
  assign new_n26558_ = ys__n34670 & ~ys__n34672;
  assign new_n26559_ = ~new_n26557_ & ~new_n26558_;
  assign new_n26560_ = ys__n34674 & ys__n34676;
  assign new_n26561_ = new_n26559_ & new_n26560_;
  assign new_n26562_ = ~new_n26559_ & ~new_n26560_;
  assign new_n26563_ = ~new_n26561_ & ~new_n26562_;
  assign new_n26564_ = ~new_n26487_ & ~new_n26491_;
  assign new_n26565_ = new_n26563_ & new_n26564_;
  assign new_n26566_ = ~new_n26563_ & ~new_n26564_;
  assign new_n26567_ = ~new_n26565_ & ~new_n26566_;
  assign new_n26568_ = ~ys__n48325 & ~new_n26567_;
  assign new_n26569_ = ys__n48325 & new_n26567_;
  assign new_n26570_ = ~new_n26568_ & ~new_n26569_;
  assign new_n26571_ = new_n26517_ & new_n26570_;
  assign new_n26572_ = ~new_n26517_ & ~new_n26570_;
  assign new_n26573_ = ~new_n26571_ & ~new_n26572_;
  assign new_n26574_ = new_n26514_ & ~new_n26573_;
  assign new_n26575_ = ~new_n26494_ & new_n26567_;
  assign new_n26576_ = new_n26494_ & ~new_n26567_;
  assign new_n26577_ = ~new_n26575_ & ~new_n26576_;
  assign new_n26578_ = ~ys__n48325 & ~new_n26577_;
  assign new_n26579_ = ys__n48325 & new_n26577_;
  assign new_n26580_ = ~new_n26578_ & ~new_n26579_;
  assign new_n26581_ = new_n26496_ & new_n26580_;
  assign new_n26582_ = ~new_n26496_ & ~new_n26580_;
  assign new_n26583_ = ~new_n26581_ & ~new_n26582_;
  assign new_n26584_ = ~new_n26514_ & ~new_n26583_;
  assign new_n26585_ = ~new_n26574_ & ~new_n26584_;
  assign new_n26586_ = ys__n2779 & ~new_n26585_;
  assign new_n26587_ = ~ys__n34666 & ys__n34668;
  assign new_n26588_ = ys__n34666 & ~ys__n34668;
  assign new_n26589_ = ~new_n26587_ & ~new_n26588_;
  assign new_n26590_ = ys__n34670 & ys__n34672;
  assign new_n26591_ = new_n26589_ & new_n26590_;
  assign new_n26592_ = ~new_n26589_ & ~new_n26590_;
  assign new_n26593_ = ~new_n26591_ & ~new_n26592_;
  assign new_n26594_ = ~new_n26559_ & new_n26560_;
  assign new_n26595_ = ~new_n26563_ & new_n26564_;
  assign new_n26596_ = ~new_n26594_ & ~new_n26595_;
  assign new_n26597_ = new_n26593_ & ~new_n26596_;
  assign new_n26598_ = ~new_n26593_ & new_n26596_;
  assign new_n26599_ = ~new_n26597_ & ~new_n26598_;
  assign new_n26600_ = ~ys__n48327 & ~new_n26599_;
  assign new_n26601_ = ys__n48327 & new_n26599_;
  assign new_n26602_ = ~new_n26600_ & ~new_n26601_;
  assign new_n26603_ = ys__n48325 & ~new_n26567_;
  assign new_n26604_ = new_n26517_ & ~new_n26570_;
  assign new_n26605_ = ~new_n26603_ & ~new_n26604_;
  assign new_n26606_ = new_n26602_ & ~new_n26605_;
  assign new_n26607_ = ~new_n26602_ & new_n26605_;
  assign new_n26608_ = ~new_n26606_ & ~new_n26607_;
  assign new_n26609_ = new_n26514_ & ~new_n26608_;
  assign new_n26610_ = ~new_n26494_ & ~new_n26567_;
  assign new_n26611_ = new_n26599_ & new_n26610_;
  assign new_n26612_ = ~new_n26599_ & ~new_n26610_;
  assign new_n26613_ = ~new_n26611_ & ~new_n26612_;
  assign new_n26614_ = ~ys__n48327 & ~new_n26613_;
  assign new_n26615_ = ys__n48327 & new_n26613_;
  assign new_n26616_ = ~new_n26614_ & ~new_n26615_;
  assign new_n26617_ = ys__n48325 & ~new_n26577_;
  assign new_n26618_ = new_n26496_ & ~new_n26580_;
  assign new_n26619_ = ~new_n26617_ & ~new_n26618_;
  assign new_n26620_ = new_n26616_ & ~new_n26619_;
  assign new_n26621_ = ~new_n26616_ & new_n26619_;
  assign new_n26622_ = ~new_n26620_ & ~new_n26621_;
  assign new_n26623_ = ~new_n26514_ & ~new_n26622_;
  assign new_n26624_ = ~new_n26609_ & ~new_n26623_;
  assign new_n26625_ = new_n26586_ & ~new_n26624_;
  assign new_n26626_ = ys__n314 & ~new_n26625_;
  assign new_n26627_ = ~ys__n314 & new_n26625_;
  assign new_n26628_ = ~new_n26626_ & ~new_n26627_;
  assign new_n26629_ = new_n25371_ & ~new_n26628_;
  assign new_n26630_ = ys__n2535 & ~new_n25402_;
  assign new_n26631_ = ~new_n26629_ & ~new_n26630_;
  assign new_n26632_ = ~new_n13708_ & ~new_n26631_;
  assign new_n26633_ = ys__n47090 & new_n25384_;
  assign new_n26634_ = ys__n47026 & new_n25386_;
  assign new_n26635_ = ~new_n26633_ & ~new_n26634_;
  assign new_n26636_ = ~new_n25389_ & ~new_n26635_;
  assign new_n26637_ = new_n25383_ & new_n26636_;
  assign new_n26638_ = ~new_n25361_ & ~new_n25383_;
  assign new_n26639_ = ~new_n26637_ & ~new_n26638_;
  assign new_n26640_ = new_n25399_ & ~new_n26639_;
  assign new_n26641_ = ~new_n25368_ & ~new_n25399_;
  assign new_n26642_ = ~new_n26640_ & ~new_n26641_;
  assign new_n26643_ = new_n13708_ & ~new_n26642_;
  assign new_n26644_ = ~new_n26632_ & ~new_n26643_;
  assign new_n26645_ = ~ys__n1598 & ~new_n26644_;
  assign new_n26646_ = ys__n24789 & ys__n1598;
  assign ys__n24790 = new_n26645_ | new_n26646_;
  assign new_n26648_ = ys__n170 & ~new_n26625_;
  assign new_n26649_ = ys__n170 & ys__n314;
  assign new_n26650_ = ~ys__n170 & ~ys__n314;
  assign new_n26651_ = ~new_n26649_ & ~new_n26650_;
  assign new_n26652_ = new_n26625_ & ~new_n26651_;
  assign new_n26653_ = ~new_n26648_ & ~new_n26652_;
  assign new_n26654_ = new_n25371_ & ~new_n26653_;
  assign new_n26655_ = ys__n2535 & ~new_n25468_;
  assign new_n26656_ = ~new_n26654_ & ~new_n26655_;
  assign new_n26657_ = ~new_n13708_ & ~new_n26656_;
  assign new_n26658_ = ys__n47091 & new_n25384_;
  assign new_n26659_ = ys__n47027 & new_n25386_;
  assign new_n26660_ = ~new_n26658_ & ~new_n26659_;
  assign new_n26661_ = ~new_n25389_ & ~new_n26660_;
  assign new_n26662_ = new_n25383_ & new_n26661_;
  assign new_n26663_ = ~new_n25383_ & ~new_n25440_;
  assign new_n26664_ = ~new_n26662_ & ~new_n26663_;
  assign new_n26665_ = new_n25399_ & ~new_n26664_;
  assign new_n26666_ = ~new_n25399_ & ~new_n25446_;
  assign new_n26667_ = ~new_n26665_ & ~new_n26666_;
  assign new_n26668_ = new_n13708_ & ~new_n26667_;
  assign new_n26669_ = ~new_n26657_ & ~new_n26668_;
  assign new_n26670_ = ~ys__n1598 & ~new_n26669_;
  assign new_n26671_ = ys__n24792 & ys__n1598;
  assign ys__n24793 = new_n26670_ | new_n26671_;
  assign new_n26673_ = ys__n380 & ~new_n26625_;
  assign new_n26674_ = ~ys__n170 & ys__n314;
  assign new_n26675_ = ~ys__n170 & ~new_n26674_;
  assign new_n26676_ = ys__n380 & ~new_n26675_;
  assign new_n26677_ = ~ys__n380 & new_n26675_;
  assign new_n26678_ = ~new_n26676_ & ~new_n26677_;
  assign new_n26679_ = new_n26625_ & ~new_n26678_;
  assign new_n26680_ = ~new_n26673_ & ~new_n26679_;
  assign new_n26681_ = new_n25371_ & ~new_n26680_;
  assign new_n26682_ = ys__n2535 & ~new_n25540_;
  assign new_n26683_ = ~new_n26681_ & ~new_n26682_;
  assign new_n26684_ = ~new_n13708_ & ~new_n26683_;
  assign new_n26685_ = ys__n47092 & new_n25384_;
  assign new_n26686_ = ys__n47028 & new_n25386_;
  assign new_n26687_ = ~new_n26685_ & ~new_n26686_;
  assign new_n26688_ = ~new_n25389_ & ~new_n26687_;
  assign new_n26689_ = new_n25383_ & new_n26688_;
  assign new_n26690_ = ~new_n25383_ & ~new_n25512_;
  assign new_n26691_ = ~new_n26689_ & ~new_n26690_;
  assign new_n26692_ = new_n25399_ & ~new_n26691_;
  assign new_n26693_ = ~new_n25399_ & ~new_n25518_;
  assign new_n26694_ = ~new_n26692_ & ~new_n26693_;
  assign new_n26695_ = new_n13708_ & ~new_n26694_;
  assign new_n26696_ = ~new_n26684_ & ~new_n26695_;
  assign new_n26697_ = ~ys__n1598 & ~new_n26696_;
  assign new_n26698_ = ys__n24795 & ys__n1598;
  assign ys__n24796 = new_n26697_ | new_n26698_;
  assign new_n26700_ = ys__n378 & ~new_n26625_;
  assign new_n26701_ = ~ys__n380 & ~new_n26675_;
  assign new_n26702_ = ~ys__n380 & ~new_n26701_;
  assign new_n26703_ = ys__n378 & ~new_n26702_;
  assign new_n26704_ = ~ys__n378 & new_n26702_;
  assign new_n26705_ = ~new_n26703_ & ~new_n26704_;
  assign new_n26706_ = new_n26625_ & ~new_n26705_;
  assign new_n26707_ = ~new_n26700_ & ~new_n26706_;
  assign new_n26708_ = new_n25371_ & ~new_n26707_;
  assign new_n26709_ = ys__n2535 & ~new_n25615_;
  assign new_n26710_ = ~new_n26708_ & ~new_n26709_;
  assign new_n26711_ = ~new_n13708_ & ~new_n26710_;
  assign new_n26712_ = ys__n47093 & new_n25384_;
  assign new_n26713_ = ys__n47029 & new_n25386_;
  assign new_n26714_ = ~new_n26712_ & ~new_n26713_;
  assign new_n26715_ = ~new_n25389_ & ~new_n26714_;
  assign new_n26716_ = new_n25383_ & new_n26715_;
  assign new_n26717_ = ~new_n25383_ & ~new_n25585_;
  assign new_n26718_ = ~new_n26716_ & ~new_n26717_;
  assign new_n26719_ = new_n25399_ & ~new_n26718_;
  assign new_n26720_ = ~new_n25399_ & ~new_n25593_;
  assign new_n26721_ = ~new_n26719_ & ~new_n26720_;
  assign new_n26722_ = new_n13708_ & ~new_n26721_;
  assign new_n26723_ = ~new_n26711_ & ~new_n26722_;
  assign new_n26724_ = ~ys__n1598 & ~new_n26723_;
  assign new_n26725_ = ys__n24798 & ys__n1598;
  assign ys__n24799 = new_n26724_ | new_n26725_;
  assign new_n26727_ = ys__n382 & ~new_n26625_;
  assign new_n26728_ = ~ys__n378 & ~ys__n380;
  assign new_n26729_ = ~new_n26675_ & new_n26728_;
  assign new_n26730_ = ~ys__n378 & ys__n380;
  assign new_n26731_ = ~ys__n378 & ~new_n26730_;
  assign new_n26732_ = ~new_n26729_ & new_n26731_;
  assign new_n26733_ = ys__n382 & ~new_n26732_;
  assign new_n26734_ = ~ys__n382 & new_n26732_;
  assign new_n26735_ = ~new_n26733_ & ~new_n26734_;
  assign new_n26736_ = new_n26625_ & ~new_n26735_;
  assign new_n26737_ = ~new_n26727_ & ~new_n26736_;
  assign new_n26738_ = new_n25371_ & ~new_n26737_;
  assign new_n26739_ = ys__n2535 & ~new_n25692_;
  assign new_n26740_ = ~new_n26738_ & ~new_n26739_;
  assign new_n26741_ = ~new_n13708_ & ~new_n26740_;
  assign new_n26742_ = ys__n47094 & new_n25384_;
  assign new_n26743_ = ys__n47030 & new_n25386_;
  assign new_n26744_ = ~new_n26742_ & ~new_n26743_;
  assign new_n26745_ = ~new_n25389_ & ~new_n26744_;
  assign new_n26746_ = new_n25383_ & new_n26745_;
  assign new_n26747_ = ~new_n25383_ & ~new_n25664_;
  assign new_n26748_ = ~new_n26746_ & ~new_n26747_;
  assign new_n26749_ = new_n25399_ & ~new_n26748_;
  assign new_n26750_ = ~new_n25399_ & ~new_n25670_;
  assign new_n26751_ = ~new_n26749_ & ~new_n26750_;
  assign new_n26752_ = new_n13708_ & ~new_n26751_;
  assign new_n26753_ = ~new_n26741_ & ~new_n26752_;
  assign new_n26754_ = ~ys__n1598 & ~new_n26753_;
  assign new_n26755_ = ys__n24801 & ys__n1598;
  assign ys__n24802 = new_n26754_ | new_n26755_;
  assign new_n26757_ = ys__n374 & ~new_n26625_;
  assign new_n26758_ = ~ys__n382 & ~new_n26732_;
  assign new_n26759_ = ~ys__n382 & ~new_n26758_;
  assign new_n26760_ = ys__n374 & ~new_n26759_;
  assign new_n26761_ = ~ys__n374 & new_n26759_;
  assign new_n26762_ = ~new_n26760_ & ~new_n26761_;
  assign new_n26763_ = new_n26625_ & ~new_n26762_;
  assign new_n26764_ = ~new_n26757_ & ~new_n26763_;
  assign new_n26765_ = new_n25371_ & ~new_n26764_;
  assign new_n26766_ = ys__n2535 & ~new_n25768_;
  assign new_n26767_ = ~new_n26765_ & ~new_n26766_;
  assign new_n26768_ = ~new_n13708_ & ~new_n26767_;
  assign new_n26769_ = ys__n47095 & new_n25384_;
  assign new_n26770_ = ys__n47031 & new_n25386_;
  assign new_n26771_ = ~new_n26769_ & ~new_n26770_;
  assign new_n26772_ = ~new_n25389_ & ~new_n26771_;
  assign new_n26773_ = new_n25383_ & new_n26772_;
  assign new_n26774_ = ~new_n25383_ & ~new_n25737_;
  assign new_n26775_ = ~new_n26773_ & ~new_n26774_;
  assign new_n26776_ = new_n25399_ & ~new_n26775_;
  assign new_n26777_ = ~new_n25399_ & ~new_n25745_;
  assign new_n26778_ = ~new_n26776_ & ~new_n26777_;
  assign new_n26779_ = new_n13708_ & ~new_n26778_;
  assign new_n26780_ = ~new_n26768_ & ~new_n26779_;
  assign new_n26781_ = ~ys__n1598 & ~new_n26780_;
  assign new_n26782_ = ys__n24804 & ys__n1598;
  assign ys__n24805 = new_n26781_ | new_n26782_;
  assign new_n26784_ = ys__n376 & ~new_n26625_;
  assign new_n26785_ = ~ys__n374 & ys__n382;
  assign new_n26786_ = ~ys__n374 & ~new_n26785_;
  assign new_n26787_ = ~ys__n374 & ~ys__n382;
  assign new_n26788_ = ~new_n26732_ & new_n26787_;
  assign new_n26789_ = new_n26786_ & ~new_n26788_;
  assign new_n26790_ = ys__n376 & ~new_n26789_;
  assign new_n26791_ = ~ys__n376 & new_n26789_;
  assign new_n26792_ = ~new_n26790_ & ~new_n26791_;
  assign new_n26793_ = new_n26625_ & ~new_n26792_;
  assign new_n26794_ = ~new_n26784_ & ~new_n26793_;
  assign new_n26795_ = new_n25371_ & ~new_n26794_;
  assign new_n26796_ = ys__n2535 & ~new_n25848_;
  assign new_n26797_ = ~new_n26795_ & ~new_n26796_;
  assign new_n26798_ = ~new_n13708_ & ~new_n26797_;
  assign new_n26799_ = ys__n47096 & new_n25384_;
  assign new_n26800_ = ys__n47032 & new_n25386_;
  assign new_n26801_ = ~new_n26799_ & ~new_n26800_;
  assign new_n26802_ = ~new_n25389_ & ~new_n26801_;
  assign new_n26803_ = new_n25383_ & new_n26802_;
  assign new_n26804_ = ~new_n25383_ & ~new_n25817_;
  assign new_n26805_ = ~new_n26803_ & ~new_n26804_;
  assign new_n26806_ = new_n25399_ & ~new_n26805_;
  assign new_n26807_ = ~new_n25399_ & ~new_n25825_;
  assign new_n26808_ = ~new_n26806_ & ~new_n26807_;
  assign new_n26809_ = new_n13708_ & ~new_n26808_;
  assign new_n26810_ = ~new_n26798_ & ~new_n26809_;
  assign new_n26811_ = ~ys__n1598 & ~new_n26810_;
  assign new_n26812_ = ys__n24807 & ys__n1598;
  assign ys__n24808 = new_n26811_ | new_n26812_;
  assign new_n26814_ = ys__n372 & ~new_n26625_;
  assign new_n26815_ = ~ys__n376 & ~new_n26789_;
  assign new_n26816_ = ~ys__n376 & ~new_n26815_;
  assign new_n26817_ = ys__n372 & ~new_n26816_;
  assign new_n26818_ = ~ys__n372 & new_n26816_;
  assign new_n26819_ = ~new_n26817_ & ~new_n26818_;
  assign new_n26820_ = new_n26625_ & ~new_n26819_;
  assign new_n26821_ = ~new_n26814_ & ~new_n26820_;
  assign new_n26822_ = new_n25371_ & ~new_n26821_;
  assign new_n26823_ = ys__n2535 & ~new_n25924_;
  assign new_n26824_ = ~new_n26822_ & ~new_n26823_;
  assign new_n26825_ = ~new_n13708_ & ~new_n26824_;
  assign new_n26826_ = ys__n47097 & new_n25384_;
  assign new_n26827_ = ys__n47033 & new_n25386_;
  assign new_n26828_ = ~new_n26826_ & ~new_n26827_;
  assign new_n26829_ = ~new_n25389_ & ~new_n26828_;
  assign new_n26830_ = new_n25383_ & new_n26829_;
  assign new_n26831_ = ~new_n25383_ & ~new_n25893_;
  assign new_n26832_ = ~new_n26830_ & ~new_n26831_;
  assign new_n26833_ = new_n25399_ & ~new_n26832_;
  assign new_n26834_ = ~new_n25399_ & ~new_n25901_;
  assign new_n26835_ = ~new_n26833_ & ~new_n26834_;
  assign new_n26836_ = new_n13708_ & ~new_n26835_;
  assign new_n26837_ = ~new_n26825_ & ~new_n26836_;
  assign new_n26838_ = ~ys__n1598 & ~new_n26837_;
  assign new_n26839_ = ys__n24810 & ys__n1598;
  assign ys__n24811 = new_n26838_ | new_n26839_;
  assign new_n26841_ = ys__n384 & ~new_n26625_;
  assign new_n26842_ = ~ys__n372 & ~ys__n376;
  assign new_n26843_ = new_n26787_ & new_n26842_;
  assign new_n26844_ = ~new_n26732_ & new_n26843_;
  assign new_n26845_ = ~new_n26786_ & new_n26842_;
  assign new_n26846_ = ~ys__n372 & ys__n376;
  assign new_n26847_ = ~ys__n372 & ~new_n26846_;
  assign new_n26848_ = ~new_n26845_ & new_n26847_;
  assign new_n26849_ = ~new_n26844_ & new_n26848_;
  assign new_n26850_ = ys__n384 & ~new_n26849_;
  assign new_n26851_ = ~ys__n384 & new_n26849_;
  assign new_n26852_ = ~new_n26850_ & ~new_n26851_;
  assign new_n26853_ = new_n26625_ & ~new_n26852_;
  assign new_n26854_ = ~new_n26841_ & ~new_n26853_;
  assign new_n26855_ = new_n25371_ & ~new_n26854_;
  assign new_n26856_ = ys__n2535 & ~new_n26005_;
  assign new_n26857_ = ~new_n26855_ & ~new_n26856_;
  assign new_n26858_ = ~new_n13708_ & ~new_n26857_;
  assign new_n26859_ = ys__n47098 & new_n25384_;
  assign new_n26860_ = ys__n47034 & new_n25386_;
  assign new_n26861_ = ~new_n26859_ & ~new_n26860_;
  assign new_n26862_ = ~new_n25389_ & ~new_n26861_;
  assign new_n26863_ = new_n25383_ & new_n26862_;
  assign new_n26864_ = ~new_n25383_ & ~new_n25977_;
  assign new_n26865_ = ~new_n26863_ & ~new_n26864_;
  assign new_n26866_ = new_n25399_ & ~new_n26865_;
  assign new_n26867_ = ~new_n25399_ & ~new_n25983_;
  assign new_n26868_ = ~new_n26866_ & ~new_n26867_;
  assign new_n26869_ = new_n13708_ & ~new_n26868_;
  assign new_n26870_ = ~new_n26858_ & ~new_n26869_;
  assign new_n26871_ = ~ys__n1598 & ~new_n26870_;
  assign new_n26872_ = ys__n24813 & ys__n1598;
  assign ys__n24814 = new_n26871_ | new_n26872_;
  assign new_n26874_ = ys__n366 & ~new_n26625_;
  assign new_n26875_ = ~ys__n384 & ~new_n26849_;
  assign new_n26876_ = ~ys__n384 & ~new_n26875_;
  assign new_n26877_ = ys__n366 & ~new_n26876_;
  assign new_n26878_ = ~ys__n366 & new_n26876_;
  assign new_n26879_ = ~new_n26877_ & ~new_n26878_;
  assign new_n26880_ = new_n26625_ & ~new_n26879_;
  assign new_n26881_ = ~new_n26874_ & ~new_n26880_;
  assign new_n26882_ = new_n25371_ & ~new_n26881_;
  assign new_n26883_ = ys__n2535 & ~new_n26081_;
  assign new_n26884_ = ~new_n26882_ & ~new_n26883_;
  assign new_n26885_ = ~new_n13708_ & ~new_n26884_;
  assign new_n26886_ = ys__n47099 & new_n25384_;
  assign new_n26887_ = ys__n47035 & new_n25386_;
  assign new_n26888_ = ~new_n26886_ & ~new_n26887_;
  assign new_n26889_ = ~new_n25389_ & ~new_n26888_;
  assign new_n26890_ = new_n25383_ & new_n26889_;
  assign new_n26891_ = ~new_n25383_ & ~new_n26050_;
  assign new_n26892_ = ~new_n26890_ & ~new_n26891_;
  assign new_n26893_ = new_n25399_ & ~new_n26892_;
  assign new_n26894_ = ~new_n25399_ & ~new_n26058_;
  assign new_n26895_ = ~new_n26893_ & ~new_n26894_;
  assign new_n26896_ = new_n13708_ & ~new_n26895_;
  assign new_n26897_ = ~new_n26885_ & ~new_n26896_;
  assign new_n26898_ = ~ys__n1598 & ~new_n26897_;
  assign new_n26899_ = ys__n24816 & ys__n1598;
  assign ys__n24817 = new_n26898_ | new_n26899_;
  assign new_n26901_ = ys__n368 & ~new_n26625_;
  assign new_n26902_ = ~ys__n366 & ys__n384;
  assign new_n26903_ = ~ys__n366 & ~new_n26902_;
  assign new_n26904_ = ~ys__n366 & ~ys__n384;
  assign new_n26905_ = ~new_n26849_ & new_n26904_;
  assign new_n26906_ = new_n26903_ & ~new_n26905_;
  assign new_n26907_ = ys__n368 & ~new_n26906_;
  assign new_n26908_ = ~ys__n368 & new_n26906_;
  assign new_n26909_ = ~new_n26907_ & ~new_n26908_;
  assign new_n26910_ = new_n26625_ & ~new_n26909_;
  assign new_n26911_ = ~new_n26901_ & ~new_n26910_;
  assign new_n26912_ = new_n25371_ & ~new_n26911_;
  assign new_n26913_ = ys__n2535 & ~new_n26161_;
  assign new_n26914_ = ~new_n26912_ & ~new_n26913_;
  assign new_n26915_ = ~new_n13708_ & ~new_n26914_;
  assign new_n26916_ = ys__n47100 & new_n25384_;
  assign new_n26917_ = ys__n47036 & new_n25386_;
  assign new_n26918_ = ~new_n26916_ & ~new_n26917_;
  assign new_n26919_ = ~new_n25389_ & ~new_n26918_;
  assign new_n26920_ = new_n25383_ & new_n26919_;
  assign new_n26921_ = ~new_n25383_ & ~new_n26130_;
  assign new_n26922_ = ~new_n26920_ & ~new_n26921_;
  assign new_n26923_ = new_n25399_ & ~new_n26922_;
  assign new_n26924_ = ~new_n25399_ & ~new_n26138_;
  assign new_n26925_ = ~new_n26923_ & ~new_n26924_;
  assign new_n26926_ = new_n13708_ & ~new_n26925_;
  assign new_n26927_ = ~new_n26915_ & ~new_n26926_;
  assign new_n26928_ = ~ys__n1598 & ~new_n26927_;
  assign new_n26929_ = ys__n24819 & ys__n1598;
  assign ys__n24820 = new_n26928_ | new_n26929_;
  assign new_n26931_ = ys__n364 & ~new_n26625_;
  assign new_n26932_ = ~ys__n368 & ~new_n26906_;
  assign new_n26933_ = ~ys__n368 & ~new_n26932_;
  assign new_n26934_ = ys__n364 & ~new_n26933_;
  assign new_n26935_ = ~ys__n364 & new_n26933_;
  assign new_n26936_ = ~new_n26934_ & ~new_n26935_;
  assign new_n26937_ = new_n26625_ & ~new_n26936_;
  assign new_n26938_ = ~new_n26931_ & ~new_n26937_;
  assign new_n26939_ = new_n25371_ & ~new_n26938_;
  assign new_n26940_ = ys__n2535 & ~new_n26237_;
  assign new_n26941_ = ~new_n26939_ & ~new_n26940_;
  assign new_n26942_ = ~new_n13708_ & ~new_n26941_;
  assign new_n26943_ = ys__n47101 & new_n25384_;
  assign new_n26944_ = ys__n47037 & new_n25386_;
  assign new_n26945_ = ~new_n26943_ & ~new_n26944_;
  assign new_n26946_ = ~new_n25389_ & ~new_n26945_;
  assign new_n26947_ = new_n25383_ & new_n26946_;
  assign new_n26948_ = ~new_n25383_ & ~new_n26206_;
  assign new_n26949_ = ~new_n26947_ & ~new_n26948_;
  assign new_n26950_ = new_n25399_ & ~new_n26949_;
  assign new_n26951_ = ~new_n25399_ & ~new_n26214_;
  assign new_n26952_ = ~new_n26950_ & ~new_n26951_;
  assign new_n26953_ = new_n13708_ & ~new_n26952_;
  assign new_n26954_ = ~new_n26942_ & ~new_n26953_;
  assign new_n26955_ = ~ys__n1598 & ~new_n26954_;
  assign new_n26956_ = ys__n24822 & ys__n1598;
  assign ys__n24823 = new_n26955_ | new_n26956_;
  assign new_n26958_ = ys__n370 & ~new_n26625_;
  assign new_n26959_ = ~ys__n364 & ~ys__n368;
  assign new_n26960_ = ~new_n26903_ & new_n26959_;
  assign new_n26961_ = ~ys__n364 & ys__n368;
  assign new_n26962_ = ~ys__n364 & ~new_n26961_;
  assign new_n26963_ = ~new_n26960_ & new_n26962_;
  assign new_n26964_ = new_n26904_ & new_n26959_;
  assign new_n26965_ = ~new_n26849_ & new_n26964_;
  assign new_n26966_ = new_n26963_ & ~new_n26965_;
  assign new_n26967_ = ys__n370 & ~new_n26966_;
  assign new_n26968_ = ~ys__n370 & new_n26966_;
  assign new_n26969_ = ~new_n26967_ & ~new_n26968_;
  assign new_n26970_ = new_n26625_ & ~new_n26969_;
  assign new_n26971_ = ~new_n26958_ & ~new_n26970_;
  assign new_n26972_ = new_n25371_ & ~new_n26971_;
  assign new_n26973_ = ys__n2535 & ~new_n26321_;
  assign new_n26974_ = ~new_n26972_ & ~new_n26973_;
  assign new_n26975_ = ~new_n13708_ & ~new_n26974_;
  assign new_n26976_ = ys__n47102 & new_n25384_;
  assign new_n26977_ = ys__n47038 & new_n25386_;
  assign new_n26978_ = ~new_n26976_ & ~new_n26977_;
  assign new_n26979_ = ~new_n25389_ & ~new_n26978_;
  assign new_n26980_ = new_n25383_ & new_n26979_;
  assign new_n26981_ = ~new_n25383_ & ~new_n26290_;
  assign new_n26982_ = ~new_n26980_ & ~new_n26981_;
  assign new_n26983_ = new_n25399_ & ~new_n26982_;
  assign new_n26984_ = ~new_n25399_ & ~new_n26298_;
  assign new_n26985_ = ~new_n26983_ & ~new_n26984_;
  assign new_n26986_ = new_n13708_ & ~new_n26985_;
  assign new_n26987_ = ~new_n26975_ & ~new_n26986_;
  assign new_n26988_ = ~ys__n1598 & ~new_n26987_;
  assign new_n26989_ = ys__n24825 & ys__n1598;
  assign ys__n24826 = new_n26988_ | new_n26989_;
  assign new_n26991_ = ys__n360 & ~new_n26625_;
  assign new_n26992_ = ~ys__n370 & ~new_n26966_;
  assign new_n26993_ = ~ys__n370 & ~new_n26992_;
  assign new_n26994_ = ys__n360 & ~new_n26993_;
  assign new_n26995_ = ~ys__n360 & new_n26993_;
  assign new_n26996_ = ~new_n26994_ & ~new_n26995_;
  assign new_n26997_ = new_n26625_ & ~new_n26996_;
  assign new_n26998_ = ~new_n26991_ & ~new_n26997_;
  assign new_n26999_ = new_n25371_ & ~new_n26998_;
  assign new_n27000_ = ys__n2535 & ~new_n26397_;
  assign new_n27001_ = ~new_n26999_ & ~new_n27000_;
  assign new_n27002_ = ~new_n13708_ & ~new_n27001_;
  assign new_n27003_ = ys__n47103 & new_n25384_;
  assign new_n27004_ = ys__n47039 & new_n25386_;
  assign new_n27005_ = ~new_n27003_ & ~new_n27004_;
  assign new_n27006_ = ~new_n25389_ & ~new_n27005_;
  assign new_n27007_ = new_n25383_ & new_n27006_;
  assign new_n27008_ = ~new_n25383_ & ~new_n26366_;
  assign new_n27009_ = ~new_n27007_ & ~new_n27008_;
  assign new_n27010_ = new_n25399_ & ~new_n27009_;
  assign new_n27011_ = ~new_n25399_ & ~new_n26374_;
  assign new_n27012_ = ~new_n27010_ & ~new_n27011_;
  assign new_n27013_ = new_n13708_ & ~new_n27012_;
  assign new_n27014_ = ~new_n27002_ & ~new_n27013_;
  assign new_n27015_ = ~ys__n1598 & ~new_n27014_;
  assign new_n27016_ = ys__n24828 & ys__n1598;
  assign ys__n24829 = new_n27015_ | new_n27016_;
  assign new_n27018_ = ys__n362 & ~new_n26625_;
  assign new_n27019_ = ~ys__n360 & ys__n370;
  assign new_n27020_ = ~ys__n360 & ~new_n27019_;
  assign new_n27021_ = ~ys__n360 & ~ys__n370;
  assign new_n27022_ = ~new_n26966_ & new_n27021_;
  assign new_n27023_ = new_n27020_ & ~new_n27022_;
  assign new_n27024_ = ys__n362 & ~new_n27023_;
  assign new_n27025_ = ~ys__n362 & new_n27023_;
  assign new_n27026_ = ~new_n27024_ & ~new_n27025_;
  assign new_n27027_ = new_n26625_ & ~new_n27026_;
  assign new_n27028_ = ~new_n27018_ & ~new_n27027_;
  assign new_n27029_ = new_n25371_ & ~new_n27028_;
  assign new_n27030_ = ys__n2535 & ~new_n26477_;
  assign new_n27031_ = ~new_n27029_ & ~new_n27030_;
  assign new_n27032_ = ~new_n13708_ & ~new_n27031_;
  assign new_n27033_ = ys__n47104 & new_n25384_;
  assign new_n27034_ = ys__n47040 & new_n25386_;
  assign new_n27035_ = ~new_n27033_ & ~new_n27034_;
  assign new_n27036_ = ~new_n25389_ & ~new_n27035_;
  assign new_n27037_ = new_n25383_ & new_n27036_;
  assign new_n27038_ = ~new_n25383_ & ~new_n26446_;
  assign new_n27039_ = ~new_n27037_ & ~new_n27038_;
  assign new_n27040_ = new_n25399_ & ~new_n27039_;
  assign new_n27041_ = ~new_n25399_ & ~new_n26454_;
  assign new_n27042_ = ~new_n27040_ & ~new_n27041_;
  assign new_n27043_ = new_n13708_ & ~new_n27042_;
  assign new_n27044_ = ~new_n27032_ & ~new_n27043_;
  assign new_n27045_ = ~ys__n1598 & ~new_n27044_;
  assign new_n27046_ = ys__n24831 & ys__n1598;
  assign ys__n24832 = new_n27045_ | new_n27046_;
  assign new_n27048_ = ys__n358 & ~new_n26625_;
  assign new_n27049_ = ~ys__n362 & ~new_n27023_;
  assign new_n27050_ = ~ys__n362 & ~new_n27049_;
  assign new_n27051_ = ys__n358 & ~new_n27050_;
  assign new_n27052_ = ~ys__n358 & new_n27050_;
  assign new_n27053_ = ~new_n27051_ & ~new_n27052_;
  assign new_n27054_ = new_n26625_ & ~new_n27053_;
  assign new_n27055_ = ~new_n27048_ & ~new_n27054_;
  assign new_n27056_ = new_n25371_ & ~new_n27055_;
  assign new_n27057_ = ys__n2535 & ~new_n26551_;
  assign new_n27058_ = ~new_n27056_ & ~new_n27057_;
  assign new_n27059_ = ~new_n13708_ & ~new_n27058_;
  assign new_n27060_ = ys__n47105 & new_n25384_;
  assign new_n27061_ = ys__n47041 & new_n25386_;
  assign new_n27062_ = ~new_n27060_ & ~new_n27061_;
  assign new_n27063_ = ~new_n25389_ & ~new_n27062_;
  assign new_n27064_ = new_n25383_ & new_n27063_;
  assign new_n27065_ = ~new_n25383_ & ~new_n26520_;
  assign new_n27066_ = ~new_n27064_ & ~new_n27065_;
  assign new_n27067_ = new_n25399_ & ~new_n27066_;
  assign new_n27068_ = ~new_n25399_ & ~new_n26528_;
  assign new_n27069_ = ~new_n27067_ & ~new_n27068_;
  assign new_n27070_ = new_n13708_ & ~new_n27069_;
  assign new_n27071_ = ~new_n27059_ & ~new_n27070_;
  assign new_n27072_ = ~ys__n1598 & ~new_n27071_;
  assign new_n27073_ = ys__n24834 & ys__n1598;
  assign ys__n24835 = new_n27072_ | new_n27073_;
  assign new_n27075_ = ys__n386 & ~new_n26625_;
  assign new_n27076_ = ~ys__n358 & ~ys__n362;
  assign new_n27077_ = new_n27021_ & new_n27076_;
  assign new_n27078_ = new_n26964_ & new_n27077_;
  assign new_n27079_ = ~new_n26849_ & new_n27078_;
  assign new_n27080_ = ~new_n26963_ & new_n27077_;
  assign new_n27081_ = ~new_n27020_ & new_n27076_;
  assign new_n27082_ = ~ys__n358 & ys__n362;
  assign new_n27083_ = ~ys__n358 & ~new_n27082_;
  assign new_n27084_ = ~new_n27081_ & new_n27083_;
  assign new_n27085_ = ~new_n27080_ & new_n27084_;
  assign new_n27086_ = ~new_n27079_ & new_n27085_;
  assign new_n27087_ = ys__n386 & ~new_n27086_;
  assign new_n27088_ = ~ys__n386 & new_n27086_;
  assign new_n27089_ = ~new_n27087_ & ~new_n27088_;
  assign new_n27090_ = new_n26625_ & ~new_n27089_;
  assign new_n27091_ = ~new_n27075_ & ~new_n27090_;
  assign new_n27092_ = ~new_n13708_ & new_n25371_;
  assign new_n27093_ = ~new_n27091_ & new_n27092_;
  assign new_n27094_ = ~new_n25383_ & new_n25399_;
  assign new_n27095_ = ~new_n26585_ & new_n27094_;
  assign new_n27096_ = new_n13708_ & new_n27095_;
  assign new_n27097_ = ~new_n27093_ & ~new_n27096_;
  assign new_n27098_ = ~ys__n1598 & ~new_n27097_;
  assign ys__n24837 = new_n27073_ | new_n27098_;
  assign new_n27100_ = ys__n356 & ~new_n26625_;
  assign new_n27101_ = ~ys__n386 & ~new_n27086_;
  assign new_n27102_ = ~ys__n386 & ~new_n27101_;
  assign new_n27103_ = ys__n356 & ~new_n27102_;
  assign new_n27104_ = ~ys__n356 & new_n27102_;
  assign new_n27105_ = ~new_n27103_ & ~new_n27104_;
  assign new_n27106_ = new_n26625_ & ~new_n27105_;
  assign new_n27107_ = ~new_n27100_ & ~new_n27106_;
  assign new_n27108_ = new_n27092_ & ~new_n27107_;
  assign ys__n24907 = ~new_n26624_ & new_n27094_;
  assign new_n27110_ = new_n13708_ & ys__n24907;
  assign new_n27111_ = ~new_n27108_ & ~new_n27110_;
  assign new_n27112_ = ~ys__n1598 & ~new_n27111_;
  assign ys__n24839 = new_n27073_ | new_n27112_;
  assign new_n27114_ = ys__n31031 & ys__n47010;
  assign new_n27115_ = new_n24614_ & new_n27114_;
  assign new_n27116_ = ~new_n24614_ & ~new_n25394_;
  assign new_n27117_ = ~new_n27115_ & ~new_n27116_;
  assign new_n27118_ = ~new_n25364_ & ~new_n27117_;
  assign new_n27119_ = ys__n314 & new_n25364_;
  assign new_n27120_ = ~new_n27118_ & ~new_n27119_;
  assign new_n27121_ = new_n25371_ & ~new_n27120_;
  assign new_n27122_ = ys__n2535 & ~new_n27120_;
  assign ys__n24910 = new_n27121_ | new_n27122_;
  assign new_n27124_ = ys__n31031 & ys__n47011;
  assign new_n27125_ = new_n24614_ & new_n27124_;
  assign new_n27126_ = ~new_n24614_ & ~new_n25463_;
  assign new_n27127_ = ~new_n27125_ & ~new_n27126_;
  assign new_n27128_ = ~new_n25364_ & ~new_n27127_;
  assign new_n27129_ = ys__n170 & new_n25364_;
  assign new_n27130_ = ~new_n27128_ & ~new_n27129_;
  assign new_n27131_ = new_n25371_ & ~new_n27130_;
  assign new_n27132_ = ys__n2535 & ~new_n27130_;
  assign ys__n24913 = new_n27131_ | new_n27132_;
  assign new_n27134_ = ys__n31031 & ys__n47012;
  assign new_n27135_ = new_n24614_ & new_n27134_;
  assign new_n27136_ = ~new_n24614_ & ~new_n25535_;
  assign new_n27137_ = ~new_n27135_ & ~new_n27136_;
  assign new_n27138_ = ~new_n25364_ & ~new_n27137_;
  assign new_n27139_ = ys__n380 & new_n25364_;
  assign new_n27140_ = ~new_n27138_ & ~new_n27139_;
  assign new_n27141_ = new_n25371_ & ~new_n27140_;
  assign new_n27142_ = ys__n2535 & ~new_n27140_;
  assign ys__n24916 = new_n27141_ | new_n27142_;
  assign new_n27144_ = ys__n31031 & ys__n47013;
  assign new_n27145_ = new_n24614_ & new_n27144_;
  assign new_n27146_ = ~new_n24614_ & ~new_n25610_;
  assign new_n27147_ = ~new_n27145_ & ~new_n27146_;
  assign new_n27148_ = ~new_n25364_ & ~new_n27147_;
  assign new_n27149_ = ys__n378 & new_n25364_;
  assign new_n27150_ = ~new_n27148_ & ~new_n27149_;
  assign new_n27151_ = new_n25371_ & ~new_n27150_;
  assign new_n27152_ = ys__n2535 & ~new_n27150_;
  assign ys__n24919 = new_n27151_ | new_n27152_;
  assign new_n27154_ = ys__n31031 & ys__n47014;
  assign new_n27155_ = new_n24614_ & new_n27154_;
  assign new_n27156_ = ~new_n24614_ & ~new_n25687_;
  assign new_n27157_ = ~new_n27155_ & ~new_n27156_;
  assign new_n27158_ = ~new_n25364_ & ~new_n27157_;
  assign new_n27159_ = ys__n382 & new_n25364_;
  assign new_n27160_ = ~new_n27158_ & ~new_n27159_;
  assign new_n27161_ = new_n25371_ & ~new_n27160_;
  assign new_n27162_ = ys__n2535 & ~new_n27160_;
  assign ys__n24922 = new_n27161_ | new_n27162_;
  assign new_n27164_ = ys__n31031 & ys__n47015;
  assign new_n27165_ = new_n24614_ & new_n27164_;
  assign new_n27166_ = ~new_n24614_ & ~new_n25763_;
  assign new_n27167_ = ~new_n27165_ & ~new_n27166_;
  assign new_n27168_ = ~new_n25364_ & ~new_n27167_;
  assign new_n27169_ = ys__n374 & new_n25364_;
  assign new_n27170_ = ~new_n27168_ & ~new_n27169_;
  assign new_n27171_ = new_n25371_ & ~new_n27170_;
  assign new_n27172_ = ys__n2535 & ~new_n27170_;
  assign ys__n24925 = new_n27171_ | new_n27172_;
  assign new_n27174_ = ys__n31031 & ys__n47016;
  assign new_n27175_ = new_n24614_ & new_n27174_;
  assign new_n27176_ = ~new_n24614_ & ~new_n25843_;
  assign new_n27177_ = ~new_n27175_ & ~new_n27176_;
  assign new_n27178_ = ~new_n25364_ & ~new_n27177_;
  assign new_n27179_ = ys__n376 & new_n25364_;
  assign new_n27180_ = ~new_n27178_ & ~new_n27179_;
  assign new_n27181_ = new_n25371_ & ~new_n27180_;
  assign new_n27182_ = ys__n2535 & ~new_n27180_;
  assign ys__n24928 = new_n27181_ | new_n27182_;
  assign new_n27184_ = ys__n31031 & ys__n47017;
  assign new_n27185_ = new_n24614_ & new_n27184_;
  assign new_n27186_ = ~new_n24614_ & ~new_n25919_;
  assign new_n27187_ = ~new_n27185_ & ~new_n27186_;
  assign new_n27188_ = ~new_n25364_ & ~new_n27187_;
  assign new_n27189_ = ys__n372 & new_n25364_;
  assign new_n27190_ = ~new_n27188_ & ~new_n27189_;
  assign new_n27191_ = new_n25371_ & ~new_n27190_;
  assign new_n27192_ = ys__n2535 & ~new_n27190_;
  assign ys__n24931 = new_n27191_ | new_n27192_;
  assign new_n27194_ = ys__n31031 & ys__n47018;
  assign new_n27195_ = new_n24614_ & new_n27194_;
  assign new_n27196_ = ~new_n24614_ & ~new_n26000_;
  assign new_n27197_ = ~new_n27195_ & ~new_n27196_;
  assign new_n27198_ = ~new_n25364_ & ~new_n27197_;
  assign new_n27199_ = ys__n384 & new_n25364_;
  assign new_n27200_ = ~new_n27198_ & ~new_n27199_;
  assign new_n27201_ = new_n25371_ & ~new_n27200_;
  assign new_n27202_ = ys__n2535 & ~new_n27200_;
  assign ys__n24934 = new_n27201_ | new_n27202_;
  assign new_n27204_ = ys__n31031 & ys__n47019;
  assign new_n27205_ = new_n24614_ & new_n27204_;
  assign new_n27206_ = ~new_n24614_ & ~new_n26076_;
  assign new_n27207_ = ~new_n27205_ & ~new_n27206_;
  assign new_n27208_ = ~new_n25364_ & ~new_n27207_;
  assign new_n27209_ = ys__n366 & new_n25364_;
  assign new_n27210_ = ~new_n27208_ & ~new_n27209_;
  assign new_n27211_ = new_n25371_ & ~new_n27210_;
  assign new_n27212_ = ys__n2535 & ~new_n27210_;
  assign ys__n24937 = new_n27211_ | new_n27212_;
  assign new_n27214_ = ys__n31031 & ys__n47020;
  assign new_n27215_ = new_n24614_ & new_n27214_;
  assign new_n27216_ = ~new_n24614_ & ~new_n26156_;
  assign new_n27217_ = ~new_n27215_ & ~new_n27216_;
  assign new_n27218_ = ~new_n25364_ & ~new_n27217_;
  assign new_n27219_ = ys__n368 & new_n25364_;
  assign new_n27220_ = ~new_n27218_ & ~new_n27219_;
  assign new_n27221_ = new_n25371_ & ~new_n27220_;
  assign new_n27222_ = ys__n2535 & ~new_n27220_;
  assign ys__n24940 = new_n27221_ | new_n27222_;
  assign new_n27224_ = ys__n31031 & ys__n47021;
  assign new_n27225_ = new_n24614_ & new_n27224_;
  assign new_n27226_ = ~new_n24614_ & ~new_n26232_;
  assign new_n27227_ = ~new_n27225_ & ~new_n27226_;
  assign new_n27228_ = ~new_n25364_ & ~new_n27227_;
  assign new_n27229_ = ys__n364 & new_n25364_;
  assign new_n27230_ = ~new_n27228_ & ~new_n27229_;
  assign new_n27231_ = new_n25371_ & ~new_n27230_;
  assign new_n27232_ = ys__n2535 & ~new_n27230_;
  assign ys__n24943 = new_n27231_ | new_n27232_;
  assign new_n27234_ = ys__n31031 & ys__n47022;
  assign new_n27235_ = new_n24614_ & new_n27234_;
  assign new_n27236_ = ~new_n24614_ & ~new_n26316_;
  assign new_n27237_ = ~new_n27235_ & ~new_n27236_;
  assign new_n27238_ = ~new_n25364_ & ~new_n27237_;
  assign new_n27239_ = ys__n370 & new_n25364_;
  assign new_n27240_ = ~new_n27238_ & ~new_n27239_;
  assign new_n27241_ = new_n25371_ & ~new_n27240_;
  assign new_n27242_ = ys__n2535 & ~new_n27240_;
  assign ys__n24946 = new_n27241_ | new_n27242_;
  assign new_n27244_ = ys__n31031 & ys__n47023;
  assign new_n27245_ = new_n24614_ & new_n27244_;
  assign new_n27246_ = ~new_n24614_ & ~new_n26392_;
  assign new_n27247_ = ~new_n27245_ & ~new_n27246_;
  assign new_n27248_ = ~new_n25364_ & ~new_n27247_;
  assign new_n27249_ = ys__n360 & new_n25364_;
  assign new_n27250_ = ~new_n27248_ & ~new_n27249_;
  assign new_n27251_ = new_n25371_ & ~new_n27250_;
  assign new_n27252_ = ys__n2535 & ~new_n27250_;
  assign ys__n24949 = new_n27251_ | new_n27252_;
  assign new_n27254_ = ys__n31031 & ys__n47024;
  assign new_n27255_ = new_n24614_ & new_n27254_;
  assign new_n27256_ = ~new_n24614_ & ~new_n26472_;
  assign new_n27257_ = ~new_n27255_ & ~new_n27256_;
  assign new_n27258_ = ~new_n25364_ & ~new_n27257_;
  assign new_n27259_ = ys__n362 & new_n25364_;
  assign new_n27260_ = ~new_n27258_ & ~new_n27259_;
  assign new_n27261_ = new_n25371_ & ~new_n27260_;
  assign new_n27262_ = ys__n2535 & ~new_n27260_;
  assign ys__n24952 = new_n27261_ | new_n27262_;
  assign new_n27264_ = ys__n31031 & ys__n47025;
  assign new_n27265_ = new_n24614_ & new_n27264_;
  assign new_n27266_ = ~new_n24614_ & ~new_n26546_;
  assign new_n27267_ = ~new_n27265_ & ~new_n27266_;
  assign new_n27268_ = ~new_n25364_ & ~new_n27267_;
  assign new_n27269_ = ys__n358 & new_n25364_;
  assign new_n27270_ = ~new_n27268_ & ~new_n27269_;
  assign new_n27271_ = new_n25371_ & ~new_n27270_;
  assign new_n27272_ = ys__n2535 & ~new_n27270_;
  assign ys__n24955 = new_n27271_ | new_n27272_;
  assign new_n27274_ = ys__n698 & ys__n25300;
  assign new_n27275_ = new_n17034_ & new_n27274_;
  assign new_n27276_ = new_n15064_ & new_n17035_;
  assign ys__n25294 = new_n27275_ & new_n27276_;
  assign new_n27278_ = new_n15068_ & new_n17037_;
  assign new_n27279_ = new_n15067_ & new_n27278_;
  assign new_n27280_ = ~ys__n780 & ys__n2644;
  assign new_n27281_ = ys__n25292 & new_n27280_;
  assign new_n27282_ = ~ys__n772 & ~ys__n782;
  assign new_n27283_ = new_n17034_ & new_n27282_;
  assign new_n27284_ = new_n27276_ & new_n27283_;
  assign new_n27285_ = new_n27281_ & new_n27284_;
  assign new_n27286_ = new_n27279_ & new_n27285_;
  assign ys__n25302 = ys__n4168 | new_n27286_;
  assign new_n27288_ = ys__n25381 & new_n27280_;
  assign new_n27289_ = new_n27284_ & new_n27288_;
  assign ys__n25304 = new_n27279_ & new_n27289_;
  assign new_n27291_ = ys__n25382 & new_n27280_;
  assign new_n27292_ = new_n27284_ & new_n27291_;
  assign ys__n25306 = new_n27279_ & new_n27292_;
  assign new_n27294_ = ys__n25383 & new_n27280_;
  assign new_n27295_ = new_n27284_ & new_n27294_;
  assign ys__n25308 = new_n27279_ & new_n27295_;
  assign new_n27297_ = ys__n25384 & new_n27280_;
  assign new_n27298_ = new_n27284_ & new_n27297_;
  assign ys__n25310 = new_n27279_ & new_n27298_;
  assign new_n27300_ = ys__n29883 & ~new_n11737_;
  assign new_n27301_ = ~new_n11735_ & new_n27300_;
  assign new_n27302_ = ~ys__n23764 & new_n27301_;
  assign new_n27303_ = ys__n29899 & ~new_n11737_;
  assign new_n27304_ = ~new_n11735_ & new_n27303_;
  assign new_n27305_ = ~ys__n22466 & new_n27304_;
  assign new_n27306_ = ys__n22466 & new_n27301_;
  assign new_n27307_ = ~new_n27305_ & ~new_n27306_;
  assign new_n27308_ = ys__n23764 & ~new_n27307_;
  assign new_n27309_ = ~new_n27302_ & ~new_n27308_;
  assign ys__n25385 = new_n12000_ & ~new_n27309_;
  assign new_n27311_ = ys__n29884 & ~new_n11737_;
  assign new_n27312_ = ~new_n11735_ & new_n27311_;
  assign new_n27313_ = ~ys__n23764 & new_n27312_;
  assign new_n27314_ = ys__n29900 & ~new_n11737_;
  assign new_n27315_ = ~new_n11735_ & new_n27314_;
  assign new_n27316_ = ~ys__n22466 & new_n27315_;
  assign new_n27317_ = ys__n22466 & new_n27312_;
  assign new_n27318_ = ~new_n27316_ & ~new_n27317_;
  assign new_n27319_ = ys__n23764 & ~new_n27318_;
  assign new_n27320_ = ~new_n27313_ & ~new_n27319_;
  assign ys__n25386 = new_n12000_ & ~new_n27320_;
  assign new_n27322_ = ys__n29885 & ~new_n11737_;
  assign new_n27323_ = ~new_n11735_ & new_n27322_;
  assign new_n27324_ = ~ys__n23764 & new_n27323_;
  assign new_n27325_ = ys__n29901 & ~new_n11737_;
  assign new_n27326_ = ~new_n11735_ & new_n27325_;
  assign new_n27327_ = ~ys__n22466 & new_n27326_;
  assign new_n27328_ = ys__n22466 & new_n27323_;
  assign new_n27329_ = ~new_n27327_ & ~new_n27328_;
  assign new_n27330_ = ys__n23764 & ~new_n27329_;
  assign new_n27331_ = ~new_n27324_ & ~new_n27330_;
  assign ys__n25387 = new_n12000_ & ~new_n27331_;
  assign new_n27333_ = ~ys__n782 & ys__n2644;
  assign new_n27334_ = ys__n25300 & new_n27333_;
  assign new_n27335_ = new_n17040_ & new_n17050_;
  assign new_n27336_ = new_n27334_ & new_n27335_;
  assign new_n27337_ = ys__n598 & ys__n25300;
  assign new_n27338_ = ~new_n27336_ & ~new_n27337_;
  assign new_n27339_ = ~ys__n778 & new_n15061_;
  assign new_n27340_ = new_n15066_ & new_n27339_;
  assign new_n27341_ = ~new_n27338_ & new_n27340_;
  assign new_n27342_ = ys__n776 & ys__n25300;
  assign new_n27343_ = ~new_n27341_ & ~new_n27342_;
  assign ys__n25390 = ~ys__n4168 & ~new_n27343_;
  assign new_n27345_ = new_n15064_ & new_n15067_;
  assign new_n27346_ = new_n27278_ & new_n27345_;
  assign new_n27347_ = ys__n25300 & new_n17054_;
  assign new_n27348_ = new_n17036_ & new_n27347_;
  assign ys__n25406 = new_n27346_ & new_n27348_;
  assign new_n27350_ = ys__n25300 & new_n17034_;
  assign new_n27351_ = new_n17037_ & new_n17043_;
  assign new_n27352_ = new_n27276_ & new_n27351_;
  assign new_n27353_ = new_n27350_ & new_n27352_;
  assign new_n27354_ = ys__n4168 & ys__n25300;
  assign ys__n25421 = new_n27353_ | new_n27354_;
  assign new_n27356_ = new_n13277_ & ~ys__n18360;
  assign new_n27357_ = new_n13204_ & new_n27356_;
  assign ys__n25430 = new_n13261_ & new_n27357_;
  assign new_n27359_ = ~ys__n19256 & ys__n25386;
  assign new_n27360_ = ys__n524 & ys__n19256;
  assign new_n27361_ = ~new_n27359_ & ~new_n27360_;
  assign new_n27362_ = ys__n874 & ~new_n27361_;
  assign new_n27363_ = ~ys__n19256 & ys__n25385;
  assign new_n27364_ = ys__n526 & ys__n19256;
  assign new_n27365_ = ~new_n27363_ & ~new_n27364_;
  assign new_n27366_ = ys__n874 & ~new_n27365_;
  assign new_n27367_ = ~ys__n19256 & ys__n25387;
  assign new_n27368_ = ys__n522 & ys__n19256;
  assign new_n27369_ = ~new_n27367_ & ~new_n27368_;
  assign new_n27370_ = ys__n874 & ~new_n27369_;
  assign new_n27371_ = ~new_n27366_ & new_n27370_;
  assign ys__n25431 = ~new_n27362_ & new_n27371_;
  assign new_n27373_ = ys__n604 & ~ys__n776;
  assign new_n27374_ = ~ys__n4168 & ~ys__n25300;
  assign ys__n25438 = new_n27373_ & new_n27374_;
  assign new_n27376_ = ~ys__n25300 & new_n17071_;
  assign new_n27377_ = new_n15064_ & new_n27376_;
  assign new_n27378_ = ys__n602 & ~ys__n25300;
  assign new_n27379_ = ~new_n27377_ & ~new_n27378_;
  assign new_n27380_ = ~ys__n778 & ~new_n27379_;
  assign new_n27381_ = ys__n778 & ~ys__n25300;
  assign new_n27382_ = ~new_n27380_ & ~new_n27381_;
  assign new_n27383_ = ~ys__n604 & ~ys__n776;
  assign new_n27384_ = ~ys__n4168 & new_n27383_;
  assign ys__n25441 = ~new_n27382_ & new_n27384_;
  assign new_n27386_ = ~ys__n600 & ys__n698;
  assign new_n27387_ = ~ys__n25300 & new_n27386_;
  assign new_n27388_ = ys__n600 & ~ys__n25300;
  assign new_n27389_ = ~new_n27387_ & ~new_n27388_;
  assign new_n27390_ = ~ys__n602 & ~ys__n604;
  assign new_n27391_ = ~ys__n778 & new_n17034_;
  assign new_n27392_ = new_n27390_ & new_n27391_;
  assign ys__n25449 = ~new_n27389_ & new_n27392_;
  assign new_n27394_ = ys__n602 & ~ys__n778;
  assign new_n27395_ = ys__n25300 & new_n27394_;
  assign new_n27396_ = ys__n778 & ys__n25300;
  assign new_n27397_ = ~new_n27395_ & ~new_n27396_;
  assign ys__n25456 = new_n27384_ & ~new_n27397_;
  assign new_n27399_ = ys__n25381 & new_n17045_;
  assign ys__n25461 = ys__n784 | new_n27399_;
  assign ys__n25463 = ys__n25382 & new_n17045_;
  assign ys__n25465 = ys__n25383 & new_n17045_;
  assign ys__n25467 = ys__n25384 & new_n17045_;
  assign ys__n25469 = ys__n25470 & new_n17045_;
  assign new_n27405_ = ~ys__n25300 & new_n17054_;
  assign new_n27406_ = ys__n772 & ~ys__n25300;
  assign new_n27407_ = ~new_n27405_ & ~new_n27406_;
  assign new_n27408_ = ~ys__n600 & ~ys__n778;
  assign new_n27409_ = new_n17034_ & new_n27408_;
  assign new_n27410_ = new_n15067_ & new_n27390_;
  assign new_n27411_ = new_n27278_ & new_n27410_;
  assign new_n27412_ = new_n27409_ & new_n27411_;
  assign ys__n25472 = ~new_n27407_ & new_n27412_;
  assign new_n27414_ = ~ys__n25300 & new_n17034_;
  assign new_n27415_ = new_n17037_ & new_n27408_;
  assign new_n27416_ = new_n17043_ & new_n27390_;
  assign new_n27417_ = new_n27415_ & new_n27416_;
  assign ys__n25486 = new_n27414_ & new_n27417_;
  assign new_n27419_ = ~ys__n600 & ~ys__n698;
  assign new_n27420_ = ys__n768 & ys__n25300;
  assign new_n27421_ = new_n27419_ & new_n27420_;
  assign new_n27422_ = ys__n600 & ys__n25300;
  assign new_n27423_ = ~new_n27421_ & ~new_n27422_;
  assign ys__n25496 = new_n27392_ & ~new_n27423_;
  assign new_n27425_ = ~ys__n770 & ~ys__n772;
  assign new_n27426_ = ~ys__n780 & ys__n782;
  assign new_n27427_ = ~ys__n25300 & new_n27426_;
  assign new_n27428_ = new_n27425_ & new_n27427_;
  assign new_n27429_ = ys__n770 & ~ys__n25300;
  assign new_n27430_ = ~new_n27428_ & ~new_n27429_;
  assign new_n27431_ = ~ys__n784 & ~new_n27430_;
  assign new_n27432_ = ys__n784 & ~ys__n25300;
  assign new_n27433_ = ~new_n27431_ & ~new_n27432_;
  assign new_n27434_ = new_n17037_ & new_n27390_;
  assign new_n27435_ = new_n15067_ & new_n27434_;
  assign new_n27436_ = new_n27409_ & new_n27435_;
  assign ys__n25504 = ~new_n27433_ & new_n27436_;
  assign new_n27438_ = ~ys__n4168 & ys__n25300;
  assign ys__n25519 = new_n27373_ & new_n27438_;
  assign new_n27440_ = ys__n25300 & new_n17045_;
  assign new_n27441_ = ys__n784 & ys__n25300;
  assign new_n27442_ = ~new_n27440_ & ~new_n27441_;
  assign ys__n25522 = new_n27436_ & ~new_n27442_;
  assign new_n27444_ = ~ys__n782 & ~ys__n784;
  assign new_n27445_ = ~ys__n25300 & new_n27444_;
  assign new_n27446_ = new_n27280_ & new_n27425_;
  assign new_n27447_ = new_n15067_ & new_n27446_;
  assign new_n27448_ = new_n27445_ & new_n27447_;
  assign new_n27449_ = ys__n598 & ~ys__n25300;
  assign new_n27450_ = ~new_n27448_ & ~new_n27449_;
  assign new_n27451_ = new_n27340_ & ~new_n27450_;
  assign new_n27452_ = ys__n776 & ~ys__n25300;
  assign new_n27453_ = ~new_n27451_ & ~new_n27452_;
  assign new_n27454_ = ~ys__n4168 & ~new_n27453_;
  assign new_n27455_ = ys__n4168 & ~ys__n25300;
  assign ys__n25534 = new_n27454_ | new_n27455_;
  assign new_n27457_ = ys__n782 & ys__n25300;
  assign new_n27458_ = new_n17050_ & new_n27457_;
  assign new_n27459_ = ys__n772 & ys__n25300;
  assign new_n27460_ = ~new_n27458_ & ~new_n27459_;
  assign ys__n25550 = new_n27412_ & ~new_n27460_;
  assign new_n27462_ = ~ys__n778 & ys__n25564;
  assign new_n27463_ = ~ys__n326 & ~ys__n332;
  assign new_n27464_ = ~ys__n336 & new_n13450_;
  assign new_n27465_ = new_n27463_ & new_n27464_;
  assign new_n27466_ = ys__n25564 & ~new_n27465_;
  assign new_n27467_ = ~new_n27465_ & ~new_n27466_;
  assign new_n27468_ = ys__n778 & ~new_n27467_;
  assign new_n27469_ = ~new_n27462_ & ~new_n27468_;
  assign new_n27470_ = ~ys__n602 & ~new_n27469_;
  assign new_n27471_ = ys__n25567 & new_n27465_;
  assign new_n27472_ = ~new_n27465_ & ~new_n27469_;
  assign new_n27473_ = ~new_n27471_ & ~new_n27472_;
  assign new_n27474_ = ys__n602 & ~new_n27473_;
  assign ys__n25661 = new_n27470_ | new_n27474_;
  assign new_n27476_ = ~ys__n778 & ys__n25567;
  assign new_n27477_ = ys__n778 & ys__n25567;
  assign new_n27478_ = ~new_n27465_ & new_n27477_;
  assign new_n27479_ = ~new_n27476_ & ~new_n27478_;
  assign new_n27480_ = ~ys__n602 & ~new_n27479_;
  assign new_n27481_ = ys__n25570 & new_n27465_;
  assign new_n27482_ = ~new_n27465_ & ~new_n27479_;
  assign new_n27483_ = ~new_n27481_ & ~new_n27482_;
  assign new_n27484_ = ys__n602 & ~new_n27483_;
  assign ys__n25663 = new_n27480_ | new_n27484_;
  assign new_n27486_ = ~ys__n778 & ys__n25570;
  assign new_n27487_ = ys__n25570 & ~new_n27465_;
  assign new_n27488_ = ~new_n27465_ & ~new_n27487_;
  assign new_n27489_ = ys__n778 & ~new_n27488_;
  assign new_n27490_ = ~new_n27486_ & ~new_n27489_;
  assign new_n27491_ = ~ys__n602 & ~new_n27490_;
  assign new_n27492_ = ys__n25573 & new_n27465_;
  assign new_n27493_ = ~new_n27465_ & ~new_n27490_;
  assign new_n27494_ = ~new_n27492_ & ~new_n27493_;
  assign new_n27495_ = ys__n602 & ~new_n27494_;
  assign ys__n25665 = new_n27491_ | new_n27495_;
  assign new_n27497_ = ~ys__n778 & ys__n25573;
  assign new_n27498_ = ys__n25573 & ~new_n27465_;
  assign new_n27499_ = ~new_n27465_ & ~new_n27498_;
  assign new_n27500_ = ys__n778 & ~new_n27499_;
  assign new_n27501_ = ~new_n27497_ & ~new_n27500_;
  assign new_n27502_ = ~ys__n602 & ~new_n27501_;
  assign new_n27503_ = ys__n25576 & new_n27465_;
  assign new_n27504_ = ~new_n27465_ & ~new_n27501_;
  assign new_n27505_ = ~new_n27503_ & ~new_n27504_;
  assign new_n27506_ = ys__n602 & ~new_n27505_;
  assign ys__n25667 = new_n27502_ | new_n27506_;
  assign new_n27508_ = ~ys__n778 & ys__n25576;
  assign new_n27509_ = ys__n778 & ys__n25576;
  assign new_n27510_ = ~new_n27465_ & new_n27509_;
  assign new_n27511_ = ~new_n27508_ & ~new_n27510_;
  assign new_n27512_ = ~ys__n602 & ~new_n27511_;
  assign new_n27513_ = ys__n25579 & new_n27465_;
  assign new_n27514_ = ~new_n27465_ & ~new_n27511_;
  assign new_n27515_ = ~new_n27513_ & ~new_n27514_;
  assign new_n27516_ = ys__n602 & ~new_n27515_;
  assign ys__n25669 = new_n27512_ | new_n27516_;
  assign new_n27518_ = ~ys__n778 & ys__n25579;
  assign new_n27519_ = ys__n778 & ys__n25579;
  assign new_n27520_ = ~new_n27465_ & new_n27519_;
  assign new_n27521_ = ~new_n27518_ & ~new_n27520_;
  assign new_n27522_ = ~ys__n602 & ~new_n27521_;
  assign new_n27523_ = ys__n25582 & new_n27465_;
  assign new_n27524_ = ~new_n27465_ & ~new_n27521_;
  assign new_n27525_ = ~new_n27523_ & ~new_n27524_;
  assign new_n27526_ = ys__n602 & ~new_n27525_;
  assign ys__n25671 = new_n27522_ | new_n27526_;
  assign new_n27528_ = ~ys__n778 & ys__n25582;
  assign new_n27529_ = ys__n778 & ys__n25582;
  assign new_n27530_ = ~new_n27465_ & new_n27529_;
  assign new_n27531_ = ~new_n27528_ & ~new_n27530_;
  assign new_n27532_ = ~ys__n602 & ~new_n27531_;
  assign new_n27533_ = ys__n25585 & new_n27465_;
  assign new_n27534_ = ~new_n27465_ & ~new_n27531_;
  assign new_n27535_ = ~new_n27533_ & ~new_n27534_;
  assign new_n27536_ = ys__n602 & ~new_n27535_;
  assign ys__n25673 = new_n27532_ | new_n27536_;
  assign new_n27538_ = ~ys__n778 & ys__n25585;
  assign new_n27539_ = ys__n778 & ys__n25585;
  assign new_n27540_ = ~new_n27465_ & new_n27539_;
  assign new_n27541_ = ~new_n27538_ & ~new_n27540_;
  assign new_n27542_ = ~ys__n602 & ~new_n27541_;
  assign new_n27543_ = ys__n25588 & new_n27465_;
  assign new_n27544_ = ~new_n27465_ & ~new_n27541_;
  assign new_n27545_ = ~new_n27543_ & ~new_n27544_;
  assign new_n27546_ = ys__n602 & ~new_n27545_;
  assign ys__n25675 = new_n27542_ | new_n27546_;
  assign new_n27548_ = ~ys__n778 & ys__n25588;
  assign new_n27549_ = ys__n778 & ys__n25588;
  assign new_n27550_ = ~new_n27465_ & new_n27549_;
  assign new_n27551_ = ~new_n27548_ & ~new_n27550_;
  assign new_n27552_ = ~ys__n602 & ~new_n27551_;
  assign new_n27553_ = ys__n25591 & new_n27465_;
  assign new_n27554_ = ~new_n27465_ & ~new_n27551_;
  assign new_n27555_ = ~new_n27553_ & ~new_n27554_;
  assign new_n27556_ = ys__n602 & ~new_n27555_;
  assign ys__n25677 = new_n27552_ | new_n27556_;
  assign new_n27558_ = ~ys__n778 & ys__n25591;
  assign new_n27559_ = ys__n778 & ys__n25591;
  assign new_n27560_ = ~new_n27465_ & new_n27559_;
  assign new_n27561_ = ~new_n27558_ & ~new_n27560_;
  assign new_n27562_ = ~ys__n602 & ~new_n27561_;
  assign new_n27563_ = ys__n25594 & new_n27465_;
  assign new_n27564_ = ~new_n27465_ & ~new_n27561_;
  assign new_n27565_ = ~new_n27563_ & ~new_n27564_;
  assign new_n27566_ = ys__n602 & ~new_n27565_;
  assign ys__n25679 = new_n27562_ | new_n27566_;
  assign new_n27568_ = ~ys__n778 & ys__n25594;
  assign new_n27569_ = ys__n778 & ys__n25594;
  assign new_n27570_ = ~new_n27465_ & new_n27569_;
  assign new_n27571_ = ~new_n27568_ & ~new_n27570_;
  assign new_n27572_ = ~ys__n602 & ~new_n27571_;
  assign new_n27573_ = ys__n25597 & new_n27465_;
  assign new_n27574_ = ~new_n27465_ & ~new_n27571_;
  assign new_n27575_ = ~new_n27573_ & ~new_n27574_;
  assign new_n27576_ = ys__n602 & ~new_n27575_;
  assign ys__n25681 = new_n27572_ | new_n27576_;
  assign new_n27578_ = ~ys__n778 & ys__n25597;
  assign new_n27579_ = ys__n778 & ys__n25597;
  assign new_n27580_ = ~new_n27465_ & new_n27579_;
  assign new_n27581_ = ~new_n27578_ & ~new_n27580_;
  assign new_n27582_ = ~ys__n602 & ~new_n27581_;
  assign new_n27583_ = ys__n25600 & new_n27465_;
  assign new_n27584_ = ~new_n27465_ & ~new_n27581_;
  assign new_n27585_ = ~new_n27583_ & ~new_n27584_;
  assign new_n27586_ = ys__n602 & ~new_n27585_;
  assign ys__n25683 = new_n27582_ | new_n27586_;
  assign new_n27588_ = ~ys__n778 & ys__n25600;
  assign new_n27589_ = ys__n778 & ys__n25600;
  assign new_n27590_ = ~new_n27465_ & new_n27589_;
  assign new_n27591_ = ~new_n27588_ & ~new_n27590_;
  assign new_n27592_ = ~ys__n602 & ~new_n27591_;
  assign new_n27593_ = ys__n25603 & new_n27465_;
  assign new_n27594_ = ~new_n27465_ & ~new_n27591_;
  assign new_n27595_ = ~new_n27593_ & ~new_n27594_;
  assign new_n27596_ = ys__n602 & ~new_n27595_;
  assign ys__n25685 = new_n27592_ | new_n27596_;
  assign new_n27598_ = ~ys__n778 & ys__n25603;
  assign new_n27599_ = ys__n778 & ys__n25603;
  assign new_n27600_ = ~new_n27465_ & new_n27599_;
  assign new_n27601_ = ~new_n27598_ & ~new_n27600_;
  assign new_n27602_ = ~ys__n602 & ~new_n27601_;
  assign new_n27603_ = ys__n25606 & new_n27465_;
  assign new_n27604_ = ~new_n27465_ & ~new_n27601_;
  assign new_n27605_ = ~new_n27603_ & ~new_n27604_;
  assign new_n27606_ = ys__n602 & ~new_n27605_;
  assign ys__n25687 = new_n27602_ | new_n27606_;
  assign new_n27608_ = ~ys__n778 & ys__n25606;
  assign new_n27609_ = ys__n778 & ys__n25606;
  assign new_n27610_ = ~new_n27465_ & new_n27609_;
  assign new_n27611_ = ~new_n27608_ & ~new_n27610_;
  assign new_n27612_ = ~ys__n602 & ~new_n27611_;
  assign new_n27613_ = ys__n25609 & new_n27465_;
  assign new_n27614_ = ~new_n27465_ & ~new_n27611_;
  assign new_n27615_ = ~new_n27613_ & ~new_n27614_;
  assign new_n27616_ = ys__n602 & ~new_n27615_;
  assign ys__n25689 = new_n27612_ | new_n27616_;
  assign new_n27618_ = ~ys__n778 & ys__n25609;
  assign new_n27619_ = ys__n778 & ys__n25609;
  assign new_n27620_ = ~new_n27465_ & new_n27619_;
  assign new_n27621_ = ~new_n27618_ & ~new_n27620_;
  assign new_n27622_ = ~ys__n602 & ~new_n27621_;
  assign new_n27623_ = ys__n25612 & new_n27465_;
  assign new_n27624_ = ~new_n27465_ & ~new_n27621_;
  assign new_n27625_ = ~new_n27623_ & ~new_n27624_;
  assign new_n27626_ = ys__n602 & ~new_n27625_;
  assign ys__n25691 = new_n27622_ | new_n27626_;
  assign new_n27628_ = ~ys__n778 & ys__n25612;
  assign new_n27629_ = ys__n778 & ys__n25612;
  assign new_n27630_ = ~new_n27465_ & new_n27629_;
  assign new_n27631_ = ~new_n27628_ & ~new_n27630_;
  assign new_n27632_ = ~ys__n602 & ~new_n27631_;
  assign new_n27633_ = ys__n25615 & new_n27465_;
  assign new_n27634_ = ~new_n27465_ & ~new_n27631_;
  assign new_n27635_ = ~new_n27633_ & ~new_n27634_;
  assign new_n27636_ = ys__n602 & ~new_n27635_;
  assign ys__n25693 = new_n27632_ | new_n27636_;
  assign new_n27638_ = ~ys__n778 & ys__n25615;
  assign new_n27639_ = ys__n778 & ys__n25615;
  assign new_n27640_ = ~new_n27465_ & new_n27639_;
  assign new_n27641_ = ~new_n27638_ & ~new_n27640_;
  assign new_n27642_ = ~ys__n602 & ~new_n27641_;
  assign new_n27643_ = ys__n25618 & new_n27465_;
  assign new_n27644_ = ~new_n27465_ & ~new_n27641_;
  assign new_n27645_ = ~new_n27643_ & ~new_n27644_;
  assign new_n27646_ = ys__n602 & ~new_n27645_;
  assign ys__n25695 = new_n27642_ | new_n27646_;
  assign new_n27648_ = ~ys__n778 & ys__n25618;
  assign new_n27649_ = ys__n778 & ys__n25618;
  assign new_n27650_ = ~new_n27465_ & new_n27649_;
  assign new_n27651_ = ~new_n27648_ & ~new_n27650_;
  assign new_n27652_ = ~ys__n602 & ~new_n27651_;
  assign new_n27653_ = ys__n25621 & new_n27465_;
  assign new_n27654_ = ~new_n27465_ & ~new_n27651_;
  assign new_n27655_ = ~new_n27653_ & ~new_n27654_;
  assign new_n27656_ = ys__n602 & ~new_n27655_;
  assign ys__n25697 = new_n27652_ | new_n27656_;
  assign new_n27658_ = ~ys__n778 & ys__n25621;
  assign new_n27659_ = ys__n25621 & ~new_n27465_;
  assign new_n27660_ = ~new_n27465_ & ~new_n27659_;
  assign new_n27661_ = ys__n778 & ~new_n27660_;
  assign new_n27662_ = ~new_n27658_ & ~new_n27661_;
  assign new_n27663_ = ~ys__n602 & ~new_n27662_;
  assign new_n27664_ = ys__n25624 & new_n27465_;
  assign new_n27665_ = ~new_n27465_ & ~new_n27662_;
  assign new_n27666_ = ~new_n27664_ & ~new_n27665_;
  assign new_n27667_ = ys__n602 & ~new_n27666_;
  assign ys__n25699 = new_n27663_ | new_n27667_;
  assign new_n27669_ = ~ys__n778 & ys__n25624;
  assign new_n27670_ = ys__n25624 & ~new_n27465_;
  assign new_n27671_ = ~new_n27465_ & ~new_n27670_;
  assign new_n27672_ = ys__n778 & ~new_n27671_;
  assign new_n27673_ = ~new_n27669_ & ~new_n27672_;
  assign new_n27674_ = ~ys__n602 & ~new_n27673_;
  assign new_n27675_ = ys__n25627 & new_n27465_;
  assign new_n27676_ = ~new_n27465_ & ~new_n27673_;
  assign new_n27677_ = ~new_n27675_ & ~new_n27676_;
  assign new_n27678_ = ys__n602 & ~new_n27677_;
  assign ys__n25701 = new_n27674_ | new_n27678_;
  assign new_n27680_ = ~ys__n778 & ys__n25627;
  assign new_n27681_ = ys__n778 & ys__n25627;
  assign new_n27682_ = ~new_n27465_ & new_n27681_;
  assign new_n27683_ = ~new_n27680_ & ~new_n27682_;
  assign new_n27684_ = ~ys__n602 & ~new_n27683_;
  assign new_n27685_ = ys__n25630 & new_n27465_;
  assign new_n27686_ = ~new_n27465_ & ~new_n27683_;
  assign new_n27687_ = ~new_n27685_ & ~new_n27686_;
  assign new_n27688_ = ys__n602 & ~new_n27687_;
  assign ys__n25703 = new_n27684_ | new_n27688_;
  assign new_n27690_ = ~ys__n778 & ys__n25630;
  assign new_n27691_ = ys__n778 & ys__n25630;
  assign new_n27692_ = ~new_n27465_ & new_n27691_;
  assign new_n27693_ = ~new_n27690_ & ~new_n27692_;
  assign new_n27694_ = ~ys__n602 & ~new_n27693_;
  assign new_n27695_ = ys__n25633 & new_n27465_;
  assign new_n27696_ = ~new_n27465_ & ~new_n27693_;
  assign new_n27697_ = ~new_n27695_ & ~new_n27696_;
  assign new_n27698_ = ys__n602 & ~new_n27697_;
  assign ys__n25705 = new_n27694_ | new_n27698_;
  assign new_n27700_ = ~ys__n778 & ys__n25633;
  assign new_n27701_ = ys__n778 & ys__n25633;
  assign new_n27702_ = ~new_n27465_ & new_n27701_;
  assign new_n27703_ = ~new_n27700_ & ~new_n27702_;
  assign new_n27704_ = ~ys__n602 & ~new_n27703_;
  assign new_n27705_ = ys__n25636 & new_n27465_;
  assign new_n27706_ = ~new_n27465_ & ~new_n27703_;
  assign new_n27707_ = ~new_n27705_ & ~new_n27706_;
  assign new_n27708_ = ys__n602 & ~new_n27707_;
  assign ys__n25707 = new_n27704_ | new_n27708_;
  assign new_n27710_ = ~ys__n778 & ys__n25636;
  assign new_n27711_ = ys__n778 & ys__n25636;
  assign new_n27712_ = ~new_n27465_ & new_n27711_;
  assign new_n27713_ = ~new_n27710_ & ~new_n27712_;
  assign new_n27714_ = ~ys__n602 & ~new_n27713_;
  assign new_n27715_ = ys__n25639 & new_n27465_;
  assign new_n27716_ = ~new_n27465_ & ~new_n27713_;
  assign new_n27717_ = ~new_n27715_ & ~new_n27716_;
  assign new_n27718_ = ys__n602 & ~new_n27717_;
  assign ys__n25709 = new_n27714_ | new_n27718_;
  assign new_n27720_ = ~ys__n778 & ys__n25639;
  assign new_n27721_ = ys__n778 & ys__n25639;
  assign new_n27722_ = ~new_n27465_ & new_n27721_;
  assign new_n27723_ = ~new_n27720_ & ~new_n27722_;
  assign new_n27724_ = ~ys__n602 & ~new_n27723_;
  assign new_n27725_ = ys__n25642 & new_n27465_;
  assign new_n27726_ = ~new_n27465_ & ~new_n27723_;
  assign new_n27727_ = ~new_n27725_ & ~new_n27726_;
  assign new_n27728_ = ys__n602 & ~new_n27727_;
  assign ys__n25711 = new_n27724_ | new_n27728_;
  assign new_n27730_ = ~ys__n778 & ys__n25642;
  assign new_n27731_ = ys__n25642 & ~new_n27465_;
  assign new_n27732_ = ~new_n27465_ & ~new_n27731_;
  assign new_n27733_ = ys__n778 & ~new_n27732_;
  assign new_n27734_ = ~new_n27730_ & ~new_n27733_;
  assign new_n27735_ = ~ys__n602 & ~new_n27734_;
  assign new_n27736_ = ys__n25645 & new_n27465_;
  assign new_n27737_ = ~new_n27465_ & ~new_n27734_;
  assign new_n27738_ = ~new_n27736_ & ~new_n27737_;
  assign new_n27739_ = ys__n602 & ~new_n27738_;
  assign ys__n25713 = new_n27735_ | new_n27739_;
  assign new_n27741_ = ~ys__n778 & ys__n25645;
  assign new_n27742_ = ys__n778 & ys__n25645;
  assign new_n27743_ = ~new_n27465_ & new_n27742_;
  assign new_n27744_ = ~new_n27741_ & ~new_n27743_;
  assign new_n27745_ = ~ys__n602 & ~new_n27744_;
  assign new_n27746_ = ys__n25648 & new_n27465_;
  assign new_n27747_ = ~new_n27465_ & ~new_n27744_;
  assign new_n27748_ = ~new_n27746_ & ~new_n27747_;
  assign new_n27749_ = ys__n602 & ~new_n27748_;
  assign ys__n25715 = new_n27745_ | new_n27749_;
  assign new_n27751_ = ~ys__n778 & ys__n25648;
  assign new_n27752_ = ys__n778 & ys__n25648;
  assign new_n27753_ = ~new_n27465_ & new_n27752_;
  assign new_n27754_ = ~new_n27751_ & ~new_n27753_;
  assign new_n27755_ = ~ys__n602 & ~new_n27754_;
  assign new_n27756_ = ys__n25651 & new_n27465_;
  assign new_n27757_ = ~new_n27465_ & ~new_n27754_;
  assign new_n27758_ = ~new_n27756_ & ~new_n27757_;
  assign new_n27759_ = ys__n602 & ~new_n27758_;
  assign ys__n25717 = new_n27755_ | new_n27759_;
  assign new_n27761_ = ~ys__n778 & ys__n25651;
  assign new_n27762_ = ys__n25651 & ~new_n27465_;
  assign new_n27763_ = ~new_n27465_ & ~new_n27762_;
  assign new_n27764_ = ys__n778 & ~new_n27763_;
  assign new_n27765_ = ~new_n27761_ & ~new_n27764_;
  assign new_n27766_ = ~ys__n602 & ~new_n27765_;
  assign new_n27767_ = ys__n25654 & new_n27465_;
  assign new_n27768_ = ~new_n27465_ & ~new_n27765_;
  assign new_n27769_ = ~new_n27767_ & ~new_n27768_;
  assign new_n27770_ = ys__n602 & ~new_n27769_;
  assign ys__n25719 = new_n27766_ | new_n27770_;
  assign new_n27772_ = ~ys__n778 & ys__n25654;
  assign new_n27773_ = ys__n778 & ys__n25654;
  assign new_n27774_ = ~new_n27465_ & new_n27773_;
  assign new_n27775_ = ~new_n27772_ & ~new_n27774_;
  assign new_n27776_ = ~ys__n602 & ~new_n27775_;
  assign new_n27777_ = ys__n25657 & new_n27465_;
  assign new_n27778_ = ~new_n27465_ & ~new_n27775_;
  assign new_n27779_ = ~new_n27777_ & ~new_n27778_;
  assign new_n27780_ = ys__n602 & ~new_n27779_;
  assign ys__n25721 = new_n27776_ | new_n27780_;
  assign new_n27782_ = ~ys__n778 & ys__n25657;
  assign new_n27783_ = ys__n778 & ys__n25657;
  assign new_n27784_ = ~new_n27465_ & new_n27783_;
  assign new_n27785_ = ~new_n27782_ & ~new_n27784_;
  assign new_n27786_ = ~ys__n602 & ~new_n27785_;
  assign new_n27787_ = ys__n25470 & new_n27465_;
  assign new_n27788_ = ~new_n27465_ & ~new_n27785_;
  assign new_n27789_ = ~new_n27787_ & ~new_n27788_;
  assign new_n27790_ = ys__n602 & ~new_n27789_;
  assign ys__n25723 = new_n27786_ | new_n27790_;
  assign new_n27792_ = ys__n25292 & new_n27408_;
  assign new_n27793_ = new_n17034_ & new_n17045_;
  assign new_n27794_ = new_n27792_ & new_n27793_;
  assign new_n27795_ = new_n27435_ & new_n27794_;
  assign new_n27796_ = ~ys__n336 & new_n13454_;
  assign new_n27797_ = new_n27463_ & new_n27796_;
  assign new_n27798_ = ys__n336 & new_n17847_;
  assign new_n27799_ = ys__n336 & new_n17845_;
  assign new_n27800_ = ~new_n27798_ & ~new_n27799_;
  assign new_n27801_ = ~new_n27797_ & new_n27800_;
  assign new_n27802_ = new_n13447_ & new_n27463_;
  assign new_n27803_ = ~ys__n336 & new_n27802_;
  assign new_n27804_ = ~new_n27465_ & ~new_n27803_;
  assign new_n27805_ = ys__n336 & new_n17855_;
  assign new_n27806_ = ys__n336 & new_n17860_;
  assign new_n27807_ = ~new_n27805_ & ~new_n27806_;
  assign new_n27808_ = new_n27804_ & new_n27807_;
  assign new_n27809_ = new_n27801_ & new_n27808_;
  assign new_n27810_ = new_n13463_ & new_n27809_;
  assign new_n27811_ = ~ys__n336 & new_n13456_;
  assign new_n27812_ = new_n27463_ & new_n27811_;
  assign new_n27813_ = ~new_n17861_ & ~new_n27812_;
  assign new_n27814_ = ys__n25980 & ~new_n27813_;
  assign new_n27815_ = ys__n26425 & ~new_n17849_;
  assign new_n27816_ = ys__n26359 & new_n17856_;
  assign new_n27817_ = ~new_n27815_ & ~new_n27816_;
  assign new_n27818_ = ~new_n27814_ & new_n27817_;
  assign new_n27819_ = new_n17849_ & ~new_n17856_;
  assign new_n27820_ = new_n27813_ & new_n27819_;
  assign new_n27821_ = ~new_n27818_ & ~new_n27820_;
  assign new_n27822_ = new_n27810_ & new_n27821_;
  assign new_n27823_ = ys__n25564 & new_n27465_;
  assign new_n27824_ = ys__n46955 & ~new_n13463_;
  assign new_n27825_ = ~new_n27823_ & ~new_n27824_;
  assign new_n27826_ = ~new_n27810_ & ~new_n27825_;
  assign new_n27827_ = ~new_n27822_ & ~new_n27826_;
  assign new_n27828_ = ys__n602 & ~new_n27827_;
  assign ys__n25725 = new_n27795_ | new_n27828_;
  assign new_n27830_ = ~ys__n25727 & ~ys__n44988;
  assign new_n27831_ = ys__n18317 & new_n13376_;
  assign new_n27832_ = new_n15151_ & new_n27831_;
  assign new_n27833_ = new_n15150_ & new_n27832_;
  assign new_n27834_ = new_n15148_ & new_n27833_;
  assign new_n27835_ = new_n13419_ & new_n27834_;
  assign new_n27836_ = ~new_n27830_ & ~new_n27835_;
  assign new_n27837_ = ~ys__n18208 & ys__n18210;
  assign new_n27838_ = ~new_n27830_ & ~new_n27837_;
  assign new_n27839_ = ys__n18448 & new_n27837_;
  assign new_n27840_ = ~new_n27838_ & ~new_n27839_;
  assign new_n27841_ = new_n27835_ & ~new_n27840_;
  assign ys__n25830 = new_n27836_ | new_n27841_;
  assign new_n27843_ = ~ys__n25730 & ~ys__n44989;
  assign new_n27844_ = ~new_n27835_ & ~new_n27843_;
  assign new_n27845_ = ~new_n27837_ & ~new_n27843_;
  assign new_n27846_ = ys__n18451 & new_n27837_;
  assign new_n27847_ = ~new_n27845_ & ~new_n27846_;
  assign new_n27848_ = new_n27835_ & ~new_n27847_;
  assign ys__n25833 = new_n27844_ | new_n27848_;
  assign new_n27850_ = ~ys__n25733 & ~ys__n44990;
  assign new_n27851_ = ~new_n27835_ & ~new_n27850_;
  assign new_n27852_ = ~new_n27837_ & ~new_n27850_;
  assign new_n27853_ = ys__n18454 & new_n27837_;
  assign new_n27854_ = ~new_n27852_ & ~new_n27853_;
  assign new_n27855_ = new_n27835_ & ~new_n27854_;
  assign ys__n25836 = new_n27851_ | new_n27855_;
  assign new_n27857_ = ~ys__n25736 & ~ys__n44991;
  assign new_n27858_ = ~new_n27835_ & ~new_n27857_;
  assign new_n27859_ = ~new_n27837_ & ~new_n27857_;
  assign new_n27860_ = ys__n18457 & new_n27837_;
  assign new_n27861_ = ~new_n27859_ & ~new_n27860_;
  assign new_n27862_ = new_n27835_ & ~new_n27861_;
  assign ys__n25839 = new_n27858_ | new_n27862_;
  assign ys__n25842 = new_n15010_ & ~new_n15017_;
  assign ys__n25844 = new_n14700_ & ~new_n15017_;
  assign ys__n25846 = new_n14389_ & ~new_n15017_;
  assign ys__n25852 = new_n14079_ & ~new_n15017_;
  assign new_n27868_ = ~ys__n25853 & ~ys__n45707;
  assign new_n27869_ = ys__n18317 & new_n13384_;
  assign new_n27870_ = new_n15151_ & new_n27869_;
  assign new_n27871_ = new_n15150_ & new_n27870_;
  assign new_n27872_ = new_n15148_ & new_n27871_;
  assign new_n27873_ = new_n13419_ & new_n27872_;
  assign new_n27874_ = ~new_n27868_ & ~new_n27873_;
  assign new_n27875_ = ~new_n27837_ & ~new_n27868_;
  assign new_n27876_ = ~new_n27839_ & ~new_n27875_;
  assign new_n27877_ = new_n27873_ & ~new_n27876_;
  assign ys__n25957 = new_n27874_ | new_n27877_;
  assign new_n27879_ = ~ys__n25856 & ~ys__n45708;
  assign new_n27880_ = ~new_n27873_ & ~new_n27879_;
  assign new_n27881_ = ~new_n27837_ & ~new_n27879_;
  assign new_n27882_ = ~new_n27846_ & ~new_n27881_;
  assign new_n27883_ = new_n27873_ & ~new_n27882_;
  assign ys__n25960 = new_n27880_ | new_n27883_;
  assign new_n27885_ = ~ys__n25859 & ~ys__n45709;
  assign new_n27886_ = ~new_n27873_ & ~new_n27885_;
  assign new_n27887_ = ~new_n27837_ & ~new_n27885_;
  assign new_n27888_ = ~new_n27853_ & ~new_n27887_;
  assign new_n27889_ = new_n27873_ & ~new_n27888_;
  assign ys__n25963 = new_n27886_ | new_n27889_;
  assign new_n27891_ = ~ys__n25862 & ~ys__n45710;
  assign new_n27892_ = ~new_n27873_ & ~new_n27891_;
  assign new_n27893_ = ~new_n27837_ & ~new_n27891_;
  assign new_n27894_ = ~new_n27860_ & ~new_n27893_;
  assign new_n27895_ = new_n27873_ & ~new_n27894_;
  assign ys__n25966 = new_n27892_ | new_n27895_;
  assign new_n27897_ = ys__n18317 & new_n13374_;
  assign new_n27898_ = new_n15151_ & new_n27897_;
  assign new_n27899_ = new_n15150_ & new_n27898_;
  assign new_n27900_ = new_n15148_ & new_n27899_;
  assign new_n27901_ = new_n13419_ & new_n27900_;
  assign new_n27902_ = ~new_n13499_ & ~new_n27901_;
  assign new_n27903_ = ys__n26002 & new_n27902_;
  assign new_n27904_ = ys__n18041 & new_n13490_;
  assign new_n27905_ = ys__n18047 & new_n13382_;
  assign new_n27906_ = ~new_n27904_ & ~new_n27905_;
  assign new_n27907_ = ys__n18053 & new_n13379_;
  assign new_n27908_ = ys__n18061 & new_n13380_;
  assign new_n27909_ = ~new_n27907_ & ~new_n27908_;
  assign new_n27910_ = new_n27906_ & new_n27909_;
  assign new_n27911_ = ~new_n13382_ & ~new_n13490_;
  assign new_n27912_ = new_n13381_ & new_n27911_;
  assign new_n27913_ = new_n13374_ & ~new_n27912_;
  assign new_n27914_ = ~new_n27910_ & new_n27913_;
  assign new_n27915_ = ys__n46266 & new_n13490_;
  assign new_n27916_ = ys__n46442 & new_n13382_;
  assign new_n27917_ = ~new_n27915_ & ~new_n27916_;
  assign new_n27918_ = ys__n46618 & new_n13379_;
  assign new_n27919_ = ys__n46794 & new_n13380_;
  assign new_n27920_ = ~new_n27918_ & ~new_n27919_;
  assign new_n27921_ = new_n27917_ & new_n27920_;
  assign new_n27922_ = new_n13376_ & ~new_n27912_;
  assign new_n27923_ = ~new_n27921_ & new_n27922_;
  assign new_n27924_ = ~new_n27914_ & ~new_n27923_;
  assign new_n27925_ = ys__n46322 & new_n13490_;
  assign new_n27926_ = ys__n46498 & new_n13382_;
  assign new_n27927_ = ~new_n27925_ & ~new_n27926_;
  assign new_n27928_ = ys__n46674 & new_n13379_;
  assign new_n27929_ = ys__n46850 & new_n13380_;
  assign new_n27930_ = ~new_n27928_ & ~new_n27929_;
  assign new_n27931_ = new_n27927_ & new_n27930_;
  assign new_n27932_ = new_n13384_ & ~new_n27912_;
  assign new_n27933_ = ~new_n27931_ & new_n27932_;
  assign new_n27934_ = ys__n46399 & new_n13490_;
  assign new_n27935_ = ys__n46575 & new_n13382_;
  assign new_n27936_ = ~new_n27934_ & ~new_n27935_;
  assign new_n27937_ = ys__n46751 & new_n13379_;
  assign new_n27938_ = ys__n46927 & new_n13380_;
  assign new_n27939_ = ~new_n27937_ & ~new_n27938_;
  assign new_n27940_ = new_n27936_ & new_n27939_;
  assign new_n27941_ = new_n13375_ & ~new_n27912_;
  assign new_n27942_ = ~new_n27940_ & new_n27941_;
  assign new_n27943_ = ~new_n27933_ & ~new_n27942_;
  assign new_n27944_ = new_n27924_ & new_n27943_;
  assign new_n27945_ = ~new_n13374_ & ~new_n13376_;
  assign new_n27946_ = new_n13488_ & new_n27945_;
  assign new_n27947_ = new_n13380_ & new_n13393_;
  assign new_n27948_ = ~new_n13394_ & ~new_n27947_;
  assign new_n27949_ = ~new_n27947_ & ~new_n27948_;
  assign new_n27950_ = ~new_n27946_ & new_n27949_;
  assign new_n27951_ = new_n13499_ & new_n27950_;
  assign new_n27952_ = ~new_n27902_ & new_n27951_;
  assign new_n27953_ = ~new_n27944_ & new_n27952_;
  assign new_n27954_ = ~new_n27903_ & ~new_n27953_;
  assign new_n27955_ = ~new_n13420_ & ~new_n27835_;
  assign new_n27956_ = ~new_n27954_ & new_n27955_;
  assign new_n27957_ = ys__n45648 & new_n13490_;
  assign new_n27958_ = ys__n45484 & new_n13382_;
  assign new_n27959_ = ~new_n27957_ & ~new_n27958_;
  assign new_n27960_ = ys__n45320 & new_n13379_;
  assign new_n27961_ = ys__n45134 & new_n13380_;
  assign new_n27962_ = ~new_n27960_ & ~new_n27961_;
  assign new_n27963_ = new_n27959_ & new_n27962_;
  assign new_n27964_ = new_n27913_ & ~new_n27963_;
  assign new_n27965_ = ys__n45609 & new_n13490_;
  assign new_n27966_ = ys__n45445 & new_n13382_;
  assign new_n27967_ = ~new_n27965_ & ~new_n27966_;
  assign new_n27968_ = ys__n45281 & new_n13379_;
  assign new_n27969_ = ys__n45087 & new_n13380_;
  assign new_n27970_ = ~new_n27968_ & ~new_n27969_;
  assign new_n27971_ = new_n27967_ & new_n27970_;
  assign new_n27972_ = new_n27922_ & ~new_n27971_;
  assign new_n27973_ = ~new_n27964_ & ~new_n27972_;
  assign new_n27974_ = ys__n45701 & new_n13490_;
  assign new_n27975_ = ys__n45537 & new_n13382_;
  assign new_n27976_ = ~new_n27974_ & ~new_n27975_;
  assign new_n27977_ = ys__n45373 & new_n13379_;
  assign new_n27978_ = ys__n45211 & new_n13380_;
  assign new_n27979_ = ~new_n27977_ & ~new_n27978_;
  assign new_n27980_ = new_n27976_ & new_n27979_;
  assign new_n27981_ = new_n27932_ & ~new_n27980_;
  assign new_n27982_ = ys__n45554 & new_n13490_;
  assign new_n27983_ = ys__n45390 & new_n13382_;
  assign new_n27984_ = ~new_n27982_ & ~new_n27983_;
  assign new_n27985_ = ys__n45226 & new_n13379_;
  assign new_n27986_ = ys__n45008 & new_n13380_;
  assign new_n27987_ = ~new_n27985_ & ~new_n27986_;
  assign new_n27988_ = new_n27984_ & new_n27987_;
  assign new_n27989_ = new_n27941_ & ~new_n27988_;
  assign new_n27990_ = ~new_n27981_ & ~new_n27989_;
  assign new_n27991_ = new_n27973_ & new_n27990_;
  assign new_n27992_ = new_n13420_ & new_n27950_;
  assign new_n27993_ = ~new_n27955_ & new_n27992_;
  assign new_n27994_ = ~new_n27991_ & new_n27993_;
  assign new_n27995_ = ~new_n27956_ & ~new_n27994_;
  assign new_n27996_ = ~new_n13529_ & ~new_n27873_;
  assign new_n27997_ = ~new_n27995_ & new_n27996_;
  assign new_n27998_ = ys__n46102 & new_n13490_;
  assign new_n27999_ = ys__n46004 & new_n13382_;
  assign new_n28000_ = ~new_n27998_ & ~new_n27999_;
  assign new_n28001_ = ys__n45906 & new_n13379_;
  assign new_n28002_ = ys__n45810 & new_n13380_;
  assign new_n28003_ = ~new_n28001_ & ~new_n28002_;
  assign new_n28004_ = new_n28000_ & new_n28003_;
  assign new_n28005_ = new_n27922_ & ~new_n28004_;
  assign new_n28006_ = ys__n46046 & new_n13490_;
  assign new_n28007_ = ys__n45948 & new_n13382_;
  assign new_n28008_ = ~new_n28006_ & ~new_n28007_;
  assign new_n28009_ = ys__n45850 & new_n13379_;
  assign new_n28010_ = ys__n45730 & new_n13380_;
  assign new_n28011_ = ~new_n28009_ & ~new_n28010_;
  assign new_n28012_ = new_n28008_ & new_n28011_;
  assign new_n28013_ = new_n27941_ & ~new_n28012_;
  assign new_n28014_ = ~new_n28005_ & ~new_n28013_;
  assign new_n28015_ = ~new_n13377_ & new_n27949_;
  assign new_n28016_ = new_n13529_ & new_n28015_;
  assign new_n28017_ = ~new_n28014_ & new_n28016_;
  assign new_n28018_ = ~new_n27996_ & new_n28017_;
  assign ys__n26118 = new_n27997_ | new_n28018_;
  assign new_n28020_ = ys__n26005 & new_n27902_;
  assign new_n28021_ = ys__n47110 & new_n13490_;
  assign new_n28022_ = ys__n47113 & new_n13382_;
  assign new_n28023_ = ~new_n28021_ & ~new_n28022_;
  assign new_n28024_ = ys__n47116 & new_n13379_;
  assign new_n28025_ = ys__n47119 & new_n13380_;
  assign new_n28026_ = ~new_n28024_ & ~new_n28025_;
  assign new_n28027_ = new_n28023_ & new_n28026_;
  assign new_n28028_ = new_n27913_ & ~new_n28027_;
  assign new_n28029_ = ys__n46268 & new_n13490_;
  assign new_n28030_ = ys__n46444 & new_n13382_;
  assign new_n28031_ = ~new_n28029_ & ~new_n28030_;
  assign new_n28032_ = ys__n46620 & new_n13379_;
  assign new_n28033_ = ys__n46796 & new_n13380_;
  assign new_n28034_ = ~new_n28032_ & ~new_n28033_;
  assign new_n28035_ = new_n28031_ & new_n28034_;
  assign new_n28036_ = new_n27922_ & ~new_n28035_;
  assign new_n28037_ = ~new_n28028_ & ~new_n28036_;
  assign new_n28038_ = ys__n46323 & new_n13490_;
  assign new_n28039_ = ys__n46499 & new_n13382_;
  assign new_n28040_ = ~new_n28038_ & ~new_n28039_;
  assign new_n28041_ = ys__n46675 & new_n13379_;
  assign new_n28042_ = ys__n46851 & new_n13380_;
  assign new_n28043_ = ~new_n28041_ & ~new_n28042_;
  assign new_n28044_ = new_n28040_ & new_n28043_;
  assign new_n28045_ = new_n27932_ & ~new_n28044_;
  assign new_n28046_ = ys__n46400 & new_n13490_;
  assign new_n28047_ = ys__n46576 & new_n13382_;
  assign new_n28048_ = ~new_n28046_ & ~new_n28047_;
  assign new_n28049_ = ys__n46752 & new_n13379_;
  assign new_n28050_ = ys__n46928 & new_n13380_;
  assign new_n28051_ = ~new_n28049_ & ~new_n28050_;
  assign new_n28052_ = new_n28048_ & new_n28051_;
  assign new_n28053_ = new_n27941_ & ~new_n28052_;
  assign new_n28054_ = ~new_n28045_ & ~new_n28053_;
  assign new_n28055_ = new_n28037_ & new_n28054_;
  assign new_n28056_ = new_n27952_ & ~new_n28055_;
  assign new_n28057_ = ~new_n28020_ & ~new_n28056_;
  assign new_n28058_ = new_n27955_ & ~new_n28057_;
  assign new_n28059_ = ys__n45556 & new_n13490_;
  assign new_n28060_ = ys__n45392 & new_n13382_;
  assign new_n28061_ = ~new_n28059_ & ~new_n28060_;
  assign new_n28062_ = ys__n45228 & new_n13379_;
  assign new_n28063_ = ys__n45011 & new_n13380_;
  assign new_n28064_ = ~new_n28062_ & ~new_n28063_;
  assign new_n28065_ = new_n28061_ & new_n28064_;
  assign new_n28066_ = new_n27941_ & ~new_n28065_;
  assign new_n28067_ = ys__n45650 & new_n13490_;
  assign new_n28068_ = ys__n45486 & new_n13382_;
  assign new_n28069_ = ~new_n28067_ & ~new_n28068_;
  assign new_n28070_ = ys__n45322 & new_n13379_;
  assign new_n28071_ = ys__n45137 & new_n13380_;
  assign new_n28072_ = ~new_n28070_ & ~new_n28071_;
  assign new_n28073_ = new_n28069_ & new_n28072_;
  assign new_n28074_ = new_n27913_ & ~new_n28073_;
  assign new_n28075_ = ys__n45610 & new_n13490_;
  assign new_n28076_ = ys__n45446 & new_n13382_;
  assign new_n28077_ = ~new_n28075_ & ~new_n28076_;
  assign new_n28078_ = ys__n45282 & new_n13379_;
  assign new_n28079_ = ys__n45088 & new_n13380_;
  assign new_n28080_ = ~new_n28078_ & ~new_n28079_;
  assign new_n28081_ = new_n28077_ & new_n28080_;
  assign new_n28082_ = new_n27922_ & ~new_n28081_;
  assign new_n28083_ = ~new_n28074_ & ~new_n28082_;
  assign new_n28084_ = ~new_n28066_ & new_n28083_;
  assign new_n28085_ = new_n27993_ & ~new_n28084_;
  assign new_n28086_ = ~new_n28058_ & ~new_n28085_;
  assign new_n28087_ = new_n27996_ & ~new_n28086_;
  assign new_n28088_ = ys__n46103 & new_n13490_;
  assign new_n28089_ = ys__n46005 & new_n13382_;
  assign new_n28090_ = ~new_n28088_ & ~new_n28089_;
  assign new_n28091_ = ys__n45907 & new_n13379_;
  assign new_n28092_ = ys__n45811 & new_n13380_;
  assign new_n28093_ = ~new_n28091_ & ~new_n28092_;
  assign new_n28094_ = new_n28090_ & new_n28093_;
  assign new_n28095_ = new_n27922_ & ~new_n28094_;
  assign new_n28096_ = ys__n46048 & new_n13490_;
  assign new_n28097_ = ys__n45950 & new_n13382_;
  assign new_n28098_ = ~new_n28096_ & ~new_n28097_;
  assign new_n28099_ = ys__n45852 & new_n13379_;
  assign new_n28100_ = ys__n45733 & new_n13380_;
  assign new_n28101_ = ~new_n28099_ & ~new_n28100_;
  assign new_n28102_ = new_n28098_ & new_n28101_;
  assign new_n28103_ = new_n27941_ & ~new_n28102_;
  assign new_n28104_ = ~new_n28095_ & ~new_n28103_;
  assign new_n28105_ = new_n28016_ & ~new_n28104_;
  assign new_n28106_ = ~new_n27996_ & new_n28105_;
  assign ys__n26119 = new_n28087_ | new_n28106_;
  assign new_n28108_ = ys__n26008 & new_n27902_;
  assign new_n28109_ = ys__n46348 & new_n13490_;
  assign new_n28110_ = ys__n46524 & new_n13382_;
  assign new_n28111_ = ~new_n28109_ & ~new_n28110_;
  assign new_n28112_ = ys__n46700 & new_n13379_;
  assign new_n28113_ = ys__n46876 & new_n13380_;
  assign new_n28114_ = ~new_n28112_ & ~new_n28113_;
  assign new_n28115_ = new_n28111_ & new_n28114_;
  assign new_n28116_ = new_n27913_ & ~new_n28115_;
  assign new_n28117_ = ys__n46270 & new_n13490_;
  assign new_n28118_ = ys__n46446 & new_n13382_;
  assign new_n28119_ = ~new_n28117_ & ~new_n28118_;
  assign new_n28120_ = ys__n46622 & new_n13379_;
  assign new_n28121_ = ys__n46798 & new_n13380_;
  assign new_n28122_ = ~new_n28120_ & ~new_n28121_;
  assign new_n28123_ = new_n28119_ & new_n28122_;
  assign new_n28124_ = new_n27922_ & ~new_n28123_;
  assign new_n28125_ = ~new_n28116_ & ~new_n28124_;
  assign new_n28126_ = ys__n46324 & new_n13490_;
  assign new_n28127_ = ys__n46500 & new_n13382_;
  assign new_n28128_ = ~new_n28126_ & ~new_n28127_;
  assign new_n28129_ = ys__n46676 & new_n13379_;
  assign new_n28130_ = ys__n46852 & new_n13380_;
  assign new_n28131_ = ~new_n28129_ & ~new_n28130_;
  assign new_n28132_ = new_n28128_ & new_n28131_;
  assign new_n28133_ = new_n27932_ & ~new_n28132_;
  assign new_n28134_ = ys__n46401 & new_n13490_;
  assign new_n28135_ = ys__n46577 & new_n13382_;
  assign new_n28136_ = ~new_n28134_ & ~new_n28135_;
  assign new_n28137_ = ys__n46753 & new_n13379_;
  assign new_n28138_ = ys__n46929 & new_n13380_;
  assign new_n28139_ = ~new_n28137_ & ~new_n28138_;
  assign new_n28140_ = new_n28136_ & new_n28139_;
  assign new_n28141_ = new_n27941_ & ~new_n28140_;
  assign new_n28142_ = ~new_n28133_ & ~new_n28141_;
  assign new_n28143_ = new_n28125_ & new_n28142_;
  assign new_n28144_ = new_n27952_ & ~new_n28143_;
  assign new_n28145_ = ~new_n28108_ & ~new_n28144_;
  assign new_n28146_ = new_n27955_ & ~new_n28145_;
  assign new_n28147_ = ys__n45558 & new_n13490_;
  assign new_n28148_ = ys__n45394 & new_n13382_;
  assign new_n28149_ = ~new_n28147_ & ~new_n28148_;
  assign new_n28150_ = ys__n45230 & new_n13379_;
  assign new_n28151_ = ys__n45014 & new_n13380_;
  assign new_n28152_ = ~new_n28150_ & ~new_n28151_;
  assign new_n28153_ = new_n28149_ & new_n28152_;
  assign new_n28154_ = new_n27941_ & ~new_n28153_;
  assign new_n28155_ = ys__n45652 & new_n13490_;
  assign new_n28156_ = ys__n45488 & new_n13382_;
  assign new_n28157_ = ~new_n28155_ & ~new_n28156_;
  assign new_n28158_ = ys__n45324 & new_n13379_;
  assign new_n28159_ = ys__n45140 & new_n13380_;
  assign new_n28160_ = ~new_n28158_ & ~new_n28159_;
  assign new_n28161_ = new_n28157_ & new_n28160_;
  assign new_n28162_ = new_n27913_ & ~new_n28161_;
  assign new_n28163_ = ys__n45611 & new_n13490_;
  assign new_n28164_ = ys__n45447 & new_n13382_;
  assign new_n28165_ = ~new_n28163_ & ~new_n28164_;
  assign new_n28166_ = ys__n45283 & new_n13379_;
  assign new_n28167_ = ys__n45089 & new_n13380_;
  assign new_n28168_ = ~new_n28166_ & ~new_n28167_;
  assign new_n28169_ = new_n28165_ & new_n28168_;
  assign new_n28170_ = new_n27922_ & ~new_n28169_;
  assign new_n28171_ = ~new_n28162_ & ~new_n28170_;
  assign new_n28172_ = ~new_n28154_ & new_n28171_;
  assign new_n28173_ = new_n27993_ & ~new_n28172_;
  assign new_n28174_ = ~new_n28146_ & ~new_n28173_;
  assign new_n28175_ = new_n27996_ & ~new_n28174_;
  assign new_n28176_ = ys__n46104 & new_n13490_;
  assign new_n28177_ = ys__n46006 & new_n13382_;
  assign new_n28178_ = ~new_n28176_ & ~new_n28177_;
  assign new_n28179_ = ys__n45908 & new_n13379_;
  assign new_n28180_ = ys__n45812 & new_n13380_;
  assign new_n28181_ = ~new_n28179_ & ~new_n28180_;
  assign new_n28182_ = new_n28178_ & new_n28181_;
  assign new_n28183_ = new_n27922_ & ~new_n28182_;
  assign new_n28184_ = ys__n46050 & new_n13490_;
  assign new_n28185_ = ys__n45952 & new_n13382_;
  assign new_n28186_ = ~new_n28184_ & ~new_n28185_;
  assign new_n28187_ = ys__n45854 & new_n13379_;
  assign new_n28188_ = ys__n45736 & new_n13380_;
  assign new_n28189_ = ~new_n28187_ & ~new_n28188_;
  assign new_n28190_ = new_n28186_ & new_n28189_;
  assign new_n28191_ = new_n27941_ & ~new_n28190_;
  assign new_n28192_ = ~new_n28183_ & ~new_n28191_;
  assign new_n28193_ = new_n28016_ & ~new_n28192_;
  assign new_n28194_ = ~new_n27996_ & new_n28193_;
  assign ys__n26120 = new_n28175_ | new_n28194_;
  assign new_n28196_ = ys__n26011 & new_n27902_;
  assign new_n28197_ = ys__n46350 & new_n13490_;
  assign new_n28198_ = ys__n46526 & new_n13382_;
  assign new_n28199_ = ~new_n28197_ & ~new_n28198_;
  assign new_n28200_ = ys__n46702 & new_n13379_;
  assign new_n28201_ = ys__n46878 & new_n13380_;
  assign new_n28202_ = ~new_n28200_ & ~new_n28201_;
  assign new_n28203_ = new_n28199_ & new_n28202_;
  assign new_n28204_ = new_n27913_ & ~new_n28203_;
  assign new_n28205_ = ys__n46272 & new_n13490_;
  assign new_n28206_ = ys__n46448 & new_n13382_;
  assign new_n28207_ = ~new_n28205_ & ~new_n28206_;
  assign new_n28208_ = ys__n46624 & new_n13379_;
  assign new_n28209_ = ys__n46800 & new_n13380_;
  assign new_n28210_ = ~new_n28208_ & ~new_n28209_;
  assign new_n28211_ = new_n28207_ & new_n28210_;
  assign new_n28212_ = new_n27922_ & ~new_n28211_;
  assign new_n28213_ = ~new_n28204_ & ~new_n28212_;
  assign new_n28214_ = ys__n46325 & new_n13490_;
  assign new_n28215_ = ys__n46501 & new_n13382_;
  assign new_n28216_ = ~new_n28214_ & ~new_n28215_;
  assign new_n28217_ = ys__n46677 & new_n13379_;
  assign new_n28218_ = ys__n46853 & new_n13380_;
  assign new_n28219_ = ~new_n28217_ & ~new_n28218_;
  assign new_n28220_ = new_n28216_ & new_n28219_;
  assign new_n28221_ = new_n27932_ & ~new_n28220_;
  assign new_n28222_ = ys__n46402 & new_n13490_;
  assign new_n28223_ = ys__n46578 & new_n13382_;
  assign new_n28224_ = ~new_n28222_ & ~new_n28223_;
  assign new_n28225_ = ys__n46754 & new_n13379_;
  assign new_n28226_ = ys__n46930 & new_n13380_;
  assign new_n28227_ = ~new_n28225_ & ~new_n28226_;
  assign new_n28228_ = new_n28224_ & new_n28227_;
  assign new_n28229_ = new_n27941_ & ~new_n28228_;
  assign new_n28230_ = ~new_n28221_ & ~new_n28229_;
  assign new_n28231_ = new_n28213_ & new_n28230_;
  assign new_n28232_ = new_n27952_ & ~new_n28231_;
  assign new_n28233_ = ~new_n28196_ & ~new_n28232_;
  assign new_n28234_ = new_n27955_ & ~new_n28233_;
  assign new_n28235_ = ys__n45560 & new_n13490_;
  assign new_n28236_ = ys__n45396 & new_n13382_;
  assign new_n28237_ = ~new_n28235_ & ~new_n28236_;
  assign new_n28238_ = ys__n45232 & new_n13379_;
  assign new_n28239_ = ys__n45017 & new_n13380_;
  assign new_n28240_ = ~new_n28238_ & ~new_n28239_;
  assign new_n28241_ = new_n28237_ & new_n28240_;
  assign new_n28242_ = new_n27941_ & ~new_n28241_;
  assign new_n28243_ = ys__n45654 & new_n13490_;
  assign new_n28244_ = ys__n45490 & new_n13382_;
  assign new_n28245_ = ~new_n28243_ & ~new_n28244_;
  assign new_n28246_ = ys__n45326 & new_n13379_;
  assign new_n28247_ = ys__n45143 & new_n13380_;
  assign new_n28248_ = ~new_n28246_ & ~new_n28247_;
  assign new_n28249_ = new_n28245_ & new_n28248_;
  assign new_n28250_ = new_n27913_ & ~new_n28249_;
  assign new_n28251_ = ys__n45612 & new_n13490_;
  assign new_n28252_ = ys__n45448 & new_n13382_;
  assign new_n28253_ = ~new_n28251_ & ~new_n28252_;
  assign new_n28254_ = ys__n45284 & new_n13379_;
  assign new_n28255_ = ys__n45090 & new_n13380_;
  assign new_n28256_ = ~new_n28254_ & ~new_n28255_;
  assign new_n28257_ = new_n28253_ & new_n28256_;
  assign new_n28258_ = new_n27922_ & ~new_n28257_;
  assign new_n28259_ = ~new_n28250_ & ~new_n28258_;
  assign new_n28260_ = ~new_n28242_ & new_n28259_;
  assign new_n28261_ = new_n27993_ & ~new_n28260_;
  assign new_n28262_ = ~new_n28234_ & ~new_n28261_;
  assign new_n28263_ = new_n27996_ & ~new_n28262_;
  assign new_n28264_ = ys__n46105 & new_n13490_;
  assign new_n28265_ = ys__n46007 & new_n13382_;
  assign new_n28266_ = ~new_n28264_ & ~new_n28265_;
  assign new_n28267_ = ys__n45909 & new_n13379_;
  assign new_n28268_ = ys__n45813 & new_n13380_;
  assign new_n28269_ = ~new_n28267_ & ~new_n28268_;
  assign new_n28270_ = new_n28266_ & new_n28269_;
  assign new_n28271_ = new_n27922_ & ~new_n28270_;
  assign new_n28272_ = ys__n46052 & new_n13490_;
  assign new_n28273_ = ys__n45954 & new_n13382_;
  assign new_n28274_ = ~new_n28272_ & ~new_n28273_;
  assign new_n28275_ = ys__n45856 & new_n13379_;
  assign new_n28276_ = ys__n45739 & new_n13380_;
  assign new_n28277_ = ~new_n28275_ & ~new_n28276_;
  assign new_n28278_ = new_n28274_ & new_n28277_;
  assign new_n28279_ = new_n27941_ & ~new_n28278_;
  assign new_n28280_ = ~new_n28271_ & ~new_n28279_;
  assign new_n28281_ = new_n28016_ & ~new_n28280_;
  assign new_n28282_ = ~new_n27996_ & new_n28281_;
  assign ys__n26121 = new_n28263_ | new_n28282_;
  assign new_n28284_ = ys__n26014 & new_n27902_;
  assign new_n28285_ = ys__n46352 & new_n13490_;
  assign new_n28286_ = ys__n46528 & new_n13382_;
  assign new_n28287_ = ~new_n28285_ & ~new_n28286_;
  assign new_n28288_ = ys__n46704 & new_n13379_;
  assign new_n28289_ = ys__n46880 & new_n13380_;
  assign new_n28290_ = ~new_n28288_ & ~new_n28289_;
  assign new_n28291_ = new_n28287_ & new_n28290_;
  assign new_n28292_ = new_n27913_ & ~new_n28291_;
  assign new_n28293_ = ys__n46274 & new_n13490_;
  assign new_n28294_ = ys__n46450 & new_n13382_;
  assign new_n28295_ = ~new_n28293_ & ~new_n28294_;
  assign new_n28296_ = ys__n46626 & new_n13379_;
  assign new_n28297_ = ys__n46802 & new_n13380_;
  assign new_n28298_ = ~new_n28296_ & ~new_n28297_;
  assign new_n28299_ = new_n28295_ & new_n28298_;
  assign new_n28300_ = new_n27922_ & ~new_n28299_;
  assign new_n28301_ = ~new_n28292_ & ~new_n28300_;
  assign new_n28302_ = ys__n46326 & new_n13490_;
  assign new_n28303_ = ys__n46502 & new_n13382_;
  assign new_n28304_ = ~new_n28302_ & ~new_n28303_;
  assign new_n28305_ = ys__n46678 & new_n13379_;
  assign new_n28306_ = ys__n46854 & new_n13380_;
  assign new_n28307_ = ~new_n28305_ & ~new_n28306_;
  assign new_n28308_ = new_n28304_ & new_n28307_;
  assign new_n28309_ = new_n27932_ & ~new_n28308_;
  assign new_n28310_ = ys__n46403 & new_n13490_;
  assign new_n28311_ = ys__n46579 & new_n13382_;
  assign new_n28312_ = ~new_n28310_ & ~new_n28311_;
  assign new_n28313_ = ys__n46755 & new_n13379_;
  assign new_n28314_ = ys__n46931 & new_n13380_;
  assign new_n28315_ = ~new_n28313_ & ~new_n28314_;
  assign new_n28316_ = new_n28312_ & new_n28315_;
  assign new_n28317_ = new_n27941_ & ~new_n28316_;
  assign new_n28318_ = ~new_n28309_ & ~new_n28317_;
  assign new_n28319_ = new_n28301_ & new_n28318_;
  assign new_n28320_ = new_n27952_ & ~new_n28319_;
  assign new_n28321_ = ~new_n28284_ & ~new_n28320_;
  assign new_n28322_ = new_n27955_ & ~new_n28321_;
  assign new_n28323_ = ys__n45562 & new_n13490_;
  assign new_n28324_ = ys__n45398 & new_n13382_;
  assign new_n28325_ = ~new_n28323_ & ~new_n28324_;
  assign new_n28326_ = ys__n45234 & new_n13379_;
  assign new_n28327_ = ys__n45020 & new_n13380_;
  assign new_n28328_ = ~new_n28326_ & ~new_n28327_;
  assign new_n28329_ = new_n28325_ & new_n28328_;
  assign new_n28330_ = new_n27941_ & ~new_n28329_;
  assign new_n28331_ = ys__n45656 & new_n13490_;
  assign new_n28332_ = ys__n45492 & new_n13382_;
  assign new_n28333_ = ~new_n28331_ & ~new_n28332_;
  assign new_n28334_ = ys__n45328 & new_n13379_;
  assign new_n28335_ = ys__n45146 & new_n13380_;
  assign new_n28336_ = ~new_n28334_ & ~new_n28335_;
  assign new_n28337_ = new_n28333_ & new_n28336_;
  assign new_n28338_ = new_n27913_ & ~new_n28337_;
  assign new_n28339_ = ys__n45613 & new_n13490_;
  assign new_n28340_ = ys__n45449 & new_n13382_;
  assign new_n28341_ = ~new_n28339_ & ~new_n28340_;
  assign new_n28342_ = ys__n45285 & new_n13379_;
  assign new_n28343_ = ys__n45091 & new_n13380_;
  assign new_n28344_ = ~new_n28342_ & ~new_n28343_;
  assign new_n28345_ = new_n28341_ & new_n28344_;
  assign new_n28346_ = new_n27922_ & ~new_n28345_;
  assign new_n28347_ = ~new_n28338_ & ~new_n28346_;
  assign new_n28348_ = ~new_n28330_ & new_n28347_;
  assign new_n28349_ = new_n27993_ & ~new_n28348_;
  assign new_n28350_ = ~new_n28322_ & ~new_n28349_;
  assign new_n28351_ = new_n27996_ & ~new_n28350_;
  assign new_n28352_ = ys__n46106 & new_n13490_;
  assign new_n28353_ = ys__n46008 & new_n13382_;
  assign new_n28354_ = ~new_n28352_ & ~new_n28353_;
  assign new_n28355_ = ys__n45910 & new_n13379_;
  assign new_n28356_ = ys__n45814 & new_n13380_;
  assign new_n28357_ = ~new_n28355_ & ~new_n28356_;
  assign new_n28358_ = new_n28354_ & new_n28357_;
  assign new_n28359_ = new_n27922_ & ~new_n28358_;
  assign new_n28360_ = ys__n46054 & new_n13490_;
  assign new_n28361_ = ys__n45956 & new_n13382_;
  assign new_n28362_ = ~new_n28360_ & ~new_n28361_;
  assign new_n28363_ = ys__n45858 & new_n13379_;
  assign new_n28364_ = ys__n45742 & new_n13380_;
  assign new_n28365_ = ~new_n28363_ & ~new_n28364_;
  assign new_n28366_ = new_n28362_ & new_n28365_;
  assign new_n28367_ = new_n27941_ & ~new_n28366_;
  assign new_n28368_ = ~new_n28359_ & ~new_n28367_;
  assign new_n28369_ = new_n28016_ & ~new_n28368_;
  assign new_n28370_ = ~new_n27996_ & new_n28369_;
  assign ys__n26122 = new_n28351_ | new_n28370_;
  assign new_n28372_ = ys__n26017 & new_n27902_;
  assign new_n28373_ = ys__n46354 & new_n13490_;
  assign new_n28374_ = ys__n46530 & new_n13382_;
  assign new_n28375_ = ~new_n28373_ & ~new_n28374_;
  assign new_n28376_ = ys__n46706 & new_n13379_;
  assign new_n28377_ = ys__n46882 & new_n13380_;
  assign new_n28378_ = ~new_n28376_ & ~new_n28377_;
  assign new_n28379_ = new_n28375_ & new_n28378_;
  assign new_n28380_ = new_n27913_ & ~new_n28379_;
  assign new_n28381_ = ys__n46276 & new_n13490_;
  assign new_n28382_ = ys__n46452 & new_n13382_;
  assign new_n28383_ = ~new_n28381_ & ~new_n28382_;
  assign new_n28384_ = ys__n46628 & new_n13379_;
  assign new_n28385_ = ys__n46804 & new_n13380_;
  assign new_n28386_ = ~new_n28384_ & ~new_n28385_;
  assign new_n28387_ = new_n28383_ & new_n28386_;
  assign new_n28388_ = new_n27922_ & ~new_n28387_;
  assign new_n28389_ = ~new_n28380_ & ~new_n28388_;
  assign new_n28390_ = ys__n46327 & new_n13490_;
  assign new_n28391_ = ys__n46503 & new_n13382_;
  assign new_n28392_ = ~new_n28390_ & ~new_n28391_;
  assign new_n28393_ = ys__n46679 & new_n13379_;
  assign new_n28394_ = ys__n46855 & new_n13380_;
  assign new_n28395_ = ~new_n28393_ & ~new_n28394_;
  assign new_n28396_ = new_n28392_ & new_n28395_;
  assign new_n28397_ = new_n27932_ & ~new_n28396_;
  assign new_n28398_ = ys__n46404 & new_n13490_;
  assign new_n28399_ = ys__n46580 & new_n13382_;
  assign new_n28400_ = ~new_n28398_ & ~new_n28399_;
  assign new_n28401_ = ys__n46756 & new_n13379_;
  assign new_n28402_ = ys__n46932 & new_n13380_;
  assign new_n28403_ = ~new_n28401_ & ~new_n28402_;
  assign new_n28404_ = new_n28400_ & new_n28403_;
  assign new_n28405_ = new_n27941_ & ~new_n28404_;
  assign new_n28406_ = ~new_n28397_ & ~new_n28405_;
  assign new_n28407_ = new_n28389_ & new_n28406_;
  assign new_n28408_ = new_n27952_ & ~new_n28407_;
  assign new_n28409_ = ~new_n28372_ & ~new_n28408_;
  assign new_n28410_ = new_n27955_ & ~new_n28409_;
  assign new_n28411_ = ys__n45564 & new_n13490_;
  assign new_n28412_ = ys__n45400 & new_n13382_;
  assign new_n28413_ = ~new_n28411_ & ~new_n28412_;
  assign new_n28414_ = ys__n45236 & new_n13379_;
  assign new_n28415_ = ys__n45023 & new_n13380_;
  assign new_n28416_ = ~new_n28414_ & ~new_n28415_;
  assign new_n28417_ = new_n28413_ & new_n28416_;
  assign new_n28418_ = new_n27941_ & ~new_n28417_;
  assign new_n28419_ = ys__n45658 & new_n13490_;
  assign new_n28420_ = ys__n45494 & new_n13382_;
  assign new_n28421_ = ~new_n28419_ & ~new_n28420_;
  assign new_n28422_ = ys__n45330 & new_n13379_;
  assign new_n28423_ = ys__n45149 & new_n13380_;
  assign new_n28424_ = ~new_n28422_ & ~new_n28423_;
  assign new_n28425_ = new_n28421_ & new_n28424_;
  assign new_n28426_ = new_n27913_ & ~new_n28425_;
  assign new_n28427_ = ys__n45614 & new_n13490_;
  assign new_n28428_ = ys__n45450 & new_n13382_;
  assign new_n28429_ = ~new_n28427_ & ~new_n28428_;
  assign new_n28430_ = ys__n45286 & new_n13379_;
  assign new_n28431_ = ys__n45092 & new_n13380_;
  assign new_n28432_ = ~new_n28430_ & ~new_n28431_;
  assign new_n28433_ = new_n28429_ & new_n28432_;
  assign new_n28434_ = new_n27922_ & ~new_n28433_;
  assign new_n28435_ = ~new_n28426_ & ~new_n28434_;
  assign new_n28436_ = ~new_n28418_ & new_n28435_;
  assign new_n28437_ = new_n27993_ & ~new_n28436_;
  assign new_n28438_ = ~new_n28410_ & ~new_n28437_;
  assign new_n28439_ = new_n27996_ & ~new_n28438_;
  assign new_n28440_ = ys__n46107 & new_n13490_;
  assign new_n28441_ = ys__n46009 & new_n13382_;
  assign new_n28442_ = ~new_n28440_ & ~new_n28441_;
  assign new_n28443_ = ys__n45911 & new_n13379_;
  assign new_n28444_ = ys__n45815 & new_n13380_;
  assign new_n28445_ = ~new_n28443_ & ~new_n28444_;
  assign new_n28446_ = new_n28442_ & new_n28445_;
  assign new_n28447_ = new_n27922_ & ~new_n28446_;
  assign new_n28448_ = ys__n46056 & new_n13490_;
  assign new_n28449_ = ys__n45958 & new_n13382_;
  assign new_n28450_ = ~new_n28448_ & ~new_n28449_;
  assign new_n28451_ = ys__n45860 & new_n13379_;
  assign new_n28452_ = ys__n45745 & new_n13380_;
  assign new_n28453_ = ~new_n28451_ & ~new_n28452_;
  assign new_n28454_ = new_n28450_ & new_n28453_;
  assign new_n28455_ = new_n27941_ & ~new_n28454_;
  assign new_n28456_ = ~new_n28447_ & ~new_n28455_;
  assign new_n28457_ = new_n28016_ & ~new_n28456_;
  assign new_n28458_ = ~new_n27996_ & new_n28457_;
  assign ys__n26123 = new_n28439_ | new_n28458_;
  assign new_n28460_ = ys__n26020 & new_n27902_;
  assign new_n28461_ = ys__n46356 & new_n13490_;
  assign new_n28462_ = ys__n46532 & new_n13382_;
  assign new_n28463_ = ~new_n28461_ & ~new_n28462_;
  assign new_n28464_ = ys__n46708 & new_n13379_;
  assign new_n28465_ = ys__n46884 & new_n13380_;
  assign new_n28466_ = ~new_n28464_ & ~new_n28465_;
  assign new_n28467_ = new_n28463_ & new_n28466_;
  assign new_n28468_ = new_n27913_ & ~new_n28467_;
  assign new_n28469_ = ys__n46278 & new_n13490_;
  assign new_n28470_ = ys__n46454 & new_n13382_;
  assign new_n28471_ = ~new_n28469_ & ~new_n28470_;
  assign new_n28472_ = ys__n46630 & new_n13379_;
  assign new_n28473_ = ys__n46806 & new_n13380_;
  assign new_n28474_ = ~new_n28472_ & ~new_n28473_;
  assign new_n28475_ = new_n28471_ & new_n28474_;
  assign new_n28476_ = new_n27922_ & ~new_n28475_;
  assign new_n28477_ = ~new_n28468_ & ~new_n28476_;
  assign new_n28478_ = ys__n46328 & new_n13490_;
  assign new_n28479_ = ys__n46504 & new_n13382_;
  assign new_n28480_ = ~new_n28478_ & ~new_n28479_;
  assign new_n28481_ = ys__n46680 & new_n13379_;
  assign new_n28482_ = ys__n46856 & new_n13380_;
  assign new_n28483_ = ~new_n28481_ & ~new_n28482_;
  assign new_n28484_ = new_n28480_ & new_n28483_;
  assign new_n28485_ = new_n27932_ & ~new_n28484_;
  assign new_n28486_ = ys__n46405 & new_n13490_;
  assign new_n28487_ = ys__n46581 & new_n13382_;
  assign new_n28488_ = ~new_n28486_ & ~new_n28487_;
  assign new_n28489_ = ys__n46757 & new_n13379_;
  assign new_n28490_ = ys__n46933 & new_n13380_;
  assign new_n28491_ = ~new_n28489_ & ~new_n28490_;
  assign new_n28492_ = new_n28488_ & new_n28491_;
  assign new_n28493_ = new_n27941_ & ~new_n28492_;
  assign new_n28494_ = ~new_n28485_ & ~new_n28493_;
  assign new_n28495_ = new_n28477_ & new_n28494_;
  assign new_n28496_ = new_n27952_ & ~new_n28495_;
  assign new_n28497_ = ~new_n28460_ & ~new_n28496_;
  assign new_n28498_ = new_n27955_ & ~new_n28497_;
  assign new_n28499_ = ys__n45566 & new_n13490_;
  assign new_n28500_ = ys__n45402 & new_n13382_;
  assign new_n28501_ = ~new_n28499_ & ~new_n28500_;
  assign new_n28502_ = ys__n45238 & new_n13379_;
  assign new_n28503_ = ys__n45026 & new_n13380_;
  assign new_n28504_ = ~new_n28502_ & ~new_n28503_;
  assign new_n28505_ = new_n28501_ & new_n28504_;
  assign new_n28506_ = new_n27941_ & ~new_n28505_;
  assign new_n28507_ = ys__n45660 & new_n13490_;
  assign new_n28508_ = ys__n45496 & new_n13382_;
  assign new_n28509_ = ~new_n28507_ & ~new_n28508_;
  assign new_n28510_ = ys__n45332 & new_n13379_;
  assign new_n28511_ = ys__n45152 & new_n13380_;
  assign new_n28512_ = ~new_n28510_ & ~new_n28511_;
  assign new_n28513_ = new_n28509_ & new_n28512_;
  assign new_n28514_ = new_n27913_ & ~new_n28513_;
  assign new_n28515_ = ys__n45615 & new_n13490_;
  assign new_n28516_ = ys__n45451 & new_n13382_;
  assign new_n28517_ = ~new_n28515_ & ~new_n28516_;
  assign new_n28518_ = ys__n45287 & new_n13379_;
  assign new_n28519_ = ys__n45093 & new_n13380_;
  assign new_n28520_ = ~new_n28518_ & ~new_n28519_;
  assign new_n28521_ = new_n28517_ & new_n28520_;
  assign new_n28522_ = new_n27922_ & ~new_n28521_;
  assign new_n28523_ = ~new_n28514_ & ~new_n28522_;
  assign new_n28524_ = ~new_n28506_ & new_n28523_;
  assign new_n28525_ = new_n27993_ & ~new_n28524_;
  assign new_n28526_ = ~new_n28498_ & ~new_n28525_;
  assign new_n28527_ = new_n27996_ & ~new_n28526_;
  assign new_n28528_ = ys__n46108 & new_n13490_;
  assign new_n28529_ = ys__n46010 & new_n13382_;
  assign new_n28530_ = ~new_n28528_ & ~new_n28529_;
  assign new_n28531_ = ys__n45912 & new_n13379_;
  assign new_n28532_ = ys__n45816 & new_n13380_;
  assign new_n28533_ = ~new_n28531_ & ~new_n28532_;
  assign new_n28534_ = new_n28530_ & new_n28533_;
  assign new_n28535_ = new_n27922_ & ~new_n28534_;
  assign new_n28536_ = ys__n46058 & new_n13490_;
  assign new_n28537_ = ys__n45960 & new_n13382_;
  assign new_n28538_ = ~new_n28536_ & ~new_n28537_;
  assign new_n28539_ = ys__n45862 & new_n13379_;
  assign new_n28540_ = ys__n45748 & new_n13380_;
  assign new_n28541_ = ~new_n28539_ & ~new_n28540_;
  assign new_n28542_ = new_n28538_ & new_n28541_;
  assign new_n28543_ = new_n27941_ & ~new_n28542_;
  assign new_n28544_ = ~new_n28535_ & ~new_n28543_;
  assign new_n28545_ = new_n28016_ & ~new_n28544_;
  assign new_n28546_ = ~new_n27996_ & new_n28545_;
  assign ys__n26124 = new_n28527_ | new_n28546_;
  assign new_n28548_ = ys__n26023 & new_n27902_;
  assign new_n28549_ = ys__n46358 & new_n13490_;
  assign new_n28550_ = ys__n46534 & new_n13382_;
  assign new_n28551_ = ~new_n28549_ & ~new_n28550_;
  assign new_n28552_ = ys__n46710 & new_n13379_;
  assign new_n28553_ = ys__n46886 & new_n13380_;
  assign new_n28554_ = ~new_n28552_ & ~new_n28553_;
  assign new_n28555_ = new_n28551_ & new_n28554_;
  assign new_n28556_ = new_n27913_ & ~new_n28555_;
  assign new_n28557_ = ys__n46280 & new_n13490_;
  assign new_n28558_ = ys__n46456 & new_n13382_;
  assign new_n28559_ = ~new_n28557_ & ~new_n28558_;
  assign new_n28560_ = ys__n46632 & new_n13379_;
  assign new_n28561_ = ys__n46808 & new_n13380_;
  assign new_n28562_ = ~new_n28560_ & ~new_n28561_;
  assign new_n28563_ = new_n28559_ & new_n28562_;
  assign new_n28564_ = new_n27922_ & ~new_n28563_;
  assign new_n28565_ = ~new_n28556_ & ~new_n28564_;
  assign new_n28566_ = ys__n46329 & new_n13490_;
  assign new_n28567_ = ys__n46505 & new_n13382_;
  assign new_n28568_ = ~new_n28566_ & ~new_n28567_;
  assign new_n28569_ = ys__n46681 & new_n13379_;
  assign new_n28570_ = ys__n46857 & new_n13380_;
  assign new_n28571_ = ~new_n28569_ & ~new_n28570_;
  assign new_n28572_ = new_n28568_ & new_n28571_;
  assign new_n28573_ = new_n27932_ & ~new_n28572_;
  assign new_n28574_ = ys__n46406 & new_n13490_;
  assign new_n28575_ = ys__n46582 & new_n13382_;
  assign new_n28576_ = ~new_n28574_ & ~new_n28575_;
  assign new_n28577_ = ys__n46758 & new_n13379_;
  assign new_n28578_ = ys__n46934 & new_n13380_;
  assign new_n28579_ = ~new_n28577_ & ~new_n28578_;
  assign new_n28580_ = new_n28576_ & new_n28579_;
  assign new_n28581_ = new_n27941_ & ~new_n28580_;
  assign new_n28582_ = ~new_n28573_ & ~new_n28581_;
  assign new_n28583_ = new_n28565_ & new_n28582_;
  assign new_n28584_ = new_n27952_ & ~new_n28583_;
  assign new_n28585_ = ~new_n28548_ & ~new_n28584_;
  assign new_n28586_ = new_n27955_ & ~new_n28585_;
  assign new_n28587_ = ys__n45568 & new_n13490_;
  assign new_n28588_ = ys__n45404 & new_n13382_;
  assign new_n28589_ = ~new_n28587_ & ~new_n28588_;
  assign new_n28590_ = ys__n45240 & new_n13379_;
  assign new_n28591_ = ys__n45029 & new_n13380_;
  assign new_n28592_ = ~new_n28590_ & ~new_n28591_;
  assign new_n28593_ = new_n28589_ & new_n28592_;
  assign new_n28594_ = new_n27941_ & ~new_n28593_;
  assign new_n28595_ = ys__n45662 & new_n13490_;
  assign new_n28596_ = ys__n45498 & new_n13382_;
  assign new_n28597_ = ~new_n28595_ & ~new_n28596_;
  assign new_n28598_ = ys__n45334 & new_n13379_;
  assign new_n28599_ = ys__n45155 & new_n13380_;
  assign new_n28600_ = ~new_n28598_ & ~new_n28599_;
  assign new_n28601_ = new_n28597_ & new_n28600_;
  assign new_n28602_ = new_n27913_ & ~new_n28601_;
  assign new_n28603_ = ys__n45616 & new_n13490_;
  assign new_n28604_ = ys__n45452 & new_n13382_;
  assign new_n28605_ = ~new_n28603_ & ~new_n28604_;
  assign new_n28606_ = ys__n45288 & new_n13379_;
  assign new_n28607_ = ys__n45094 & new_n13380_;
  assign new_n28608_ = ~new_n28606_ & ~new_n28607_;
  assign new_n28609_ = new_n28605_ & new_n28608_;
  assign new_n28610_ = new_n27922_ & ~new_n28609_;
  assign new_n28611_ = ~new_n28602_ & ~new_n28610_;
  assign new_n28612_ = ~new_n28594_ & new_n28611_;
  assign new_n28613_ = new_n27993_ & ~new_n28612_;
  assign new_n28614_ = ~new_n28586_ & ~new_n28613_;
  assign new_n28615_ = new_n27996_ & ~new_n28614_;
  assign new_n28616_ = ys__n46109 & new_n13490_;
  assign new_n28617_ = ys__n46011 & new_n13382_;
  assign new_n28618_ = ~new_n28616_ & ~new_n28617_;
  assign new_n28619_ = ys__n45913 & new_n13379_;
  assign new_n28620_ = ys__n45817 & new_n13380_;
  assign new_n28621_ = ~new_n28619_ & ~new_n28620_;
  assign new_n28622_ = new_n28618_ & new_n28621_;
  assign new_n28623_ = new_n27922_ & ~new_n28622_;
  assign new_n28624_ = ys__n46060 & new_n13490_;
  assign new_n28625_ = ys__n45962 & new_n13382_;
  assign new_n28626_ = ~new_n28624_ & ~new_n28625_;
  assign new_n28627_ = ys__n45864 & new_n13379_;
  assign new_n28628_ = ys__n45751 & new_n13380_;
  assign new_n28629_ = ~new_n28627_ & ~new_n28628_;
  assign new_n28630_ = new_n28626_ & new_n28629_;
  assign new_n28631_ = new_n27941_ & ~new_n28630_;
  assign new_n28632_ = ~new_n28623_ & ~new_n28631_;
  assign new_n28633_ = new_n28016_ & ~new_n28632_;
  assign new_n28634_ = ~new_n27996_ & new_n28633_;
  assign ys__n26125 = new_n28615_ | new_n28634_;
  assign new_n28636_ = ys__n26026 & new_n27902_;
  assign new_n28637_ = ys__n46360 & new_n13490_;
  assign new_n28638_ = ys__n46536 & new_n13382_;
  assign new_n28639_ = ~new_n28637_ & ~new_n28638_;
  assign new_n28640_ = ys__n46712 & new_n13379_;
  assign new_n28641_ = ys__n46888 & new_n13380_;
  assign new_n28642_ = ~new_n28640_ & ~new_n28641_;
  assign new_n28643_ = new_n28639_ & new_n28642_;
  assign new_n28644_ = new_n27913_ & ~new_n28643_;
  assign new_n28645_ = ys__n46282 & new_n13490_;
  assign new_n28646_ = ys__n46458 & new_n13382_;
  assign new_n28647_ = ~new_n28645_ & ~new_n28646_;
  assign new_n28648_ = ys__n46634 & new_n13379_;
  assign new_n28649_ = ys__n46810 & new_n13380_;
  assign new_n28650_ = ~new_n28648_ & ~new_n28649_;
  assign new_n28651_ = new_n28647_ & new_n28650_;
  assign new_n28652_ = new_n27922_ & ~new_n28651_;
  assign new_n28653_ = ~new_n28644_ & ~new_n28652_;
  assign new_n28654_ = ys__n46330 & new_n13490_;
  assign new_n28655_ = ys__n46506 & new_n13382_;
  assign new_n28656_ = ~new_n28654_ & ~new_n28655_;
  assign new_n28657_ = ys__n46682 & new_n13379_;
  assign new_n28658_ = ys__n46858 & new_n13380_;
  assign new_n28659_ = ~new_n28657_ & ~new_n28658_;
  assign new_n28660_ = new_n28656_ & new_n28659_;
  assign new_n28661_ = new_n27932_ & ~new_n28660_;
  assign new_n28662_ = ys__n46407 & new_n13490_;
  assign new_n28663_ = ys__n46583 & new_n13382_;
  assign new_n28664_ = ~new_n28662_ & ~new_n28663_;
  assign new_n28665_ = ys__n46759 & new_n13379_;
  assign new_n28666_ = ys__n46935 & new_n13380_;
  assign new_n28667_ = ~new_n28665_ & ~new_n28666_;
  assign new_n28668_ = new_n28664_ & new_n28667_;
  assign new_n28669_ = new_n27941_ & ~new_n28668_;
  assign new_n28670_ = ~new_n28661_ & ~new_n28669_;
  assign new_n28671_ = new_n28653_ & new_n28670_;
  assign new_n28672_ = new_n27952_ & ~new_n28671_;
  assign new_n28673_ = ~new_n28636_ & ~new_n28672_;
  assign new_n28674_ = new_n27955_ & ~new_n28673_;
  assign new_n28675_ = ys__n45570 & new_n13490_;
  assign new_n28676_ = ys__n45406 & new_n13382_;
  assign new_n28677_ = ~new_n28675_ & ~new_n28676_;
  assign new_n28678_ = ys__n45242 & new_n13379_;
  assign new_n28679_ = ys__n45032 & new_n13380_;
  assign new_n28680_ = ~new_n28678_ & ~new_n28679_;
  assign new_n28681_ = new_n28677_ & new_n28680_;
  assign new_n28682_ = new_n27941_ & ~new_n28681_;
  assign new_n28683_ = ys__n45664 & new_n13490_;
  assign new_n28684_ = ys__n45500 & new_n13382_;
  assign new_n28685_ = ~new_n28683_ & ~new_n28684_;
  assign new_n28686_ = ys__n45336 & new_n13379_;
  assign new_n28687_ = ys__n45158 & new_n13380_;
  assign new_n28688_ = ~new_n28686_ & ~new_n28687_;
  assign new_n28689_ = new_n28685_ & new_n28688_;
  assign new_n28690_ = new_n27913_ & ~new_n28689_;
  assign new_n28691_ = ys__n45617 & new_n13490_;
  assign new_n28692_ = ys__n45453 & new_n13382_;
  assign new_n28693_ = ~new_n28691_ & ~new_n28692_;
  assign new_n28694_ = ys__n45289 & new_n13379_;
  assign new_n28695_ = ys__n45095 & new_n13380_;
  assign new_n28696_ = ~new_n28694_ & ~new_n28695_;
  assign new_n28697_ = new_n28693_ & new_n28696_;
  assign new_n28698_ = new_n27922_ & ~new_n28697_;
  assign new_n28699_ = ~new_n28690_ & ~new_n28698_;
  assign new_n28700_ = ~new_n28682_ & new_n28699_;
  assign new_n28701_ = new_n27993_ & ~new_n28700_;
  assign new_n28702_ = ~new_n28674_ & ~new_n28701_;
  assign new_n28703_ = new_n27996_ & ~new_n28702_;
  assign new_n28704_ = ys__n46110 & new_n13490_;
  assign new_n28705_ = ys__n46012 & new_n13382_;
  assign new_n28706_ = ~new_n28704_ & ~new_n28705_;
  assign new_n28707_ = ys__n45914 & new_n13379_;
  assign new_n28708_ = ys__n45818 & new_n13380_;
  assign new_n28709_ = ~new_n28707_ & ~new_n28708_;
  assign new_n28710_ = new_n28706_ & new_n28709_;
  assign new_n28711_ = new_n27922_ & ~new_n28710_;
  assign new_n28712_ = ys__n46062 & new_n13490_;
  assign new_n28713_ = ys__n45964 & new_n13382_;
  assign new_n28714_ = ~new_n28712_ & ~new_n28713_;
  assign new_n28715_ = ys__n45866 & new_n13379_;
  assign new_n28716_ = ys__n45754 & new_n13380_;
  assign new_n28717_ = ~new_n28715_ & ~new_n28716_;
  assign new_n28718_ = new_n28714_ & new_n28717_;
  assign new_n28719_ = new_n27941_ & ~new_n28718_;
  assign new_n28720_ = ~new_n28711_ & ~new_n28719_;
  assign new_n28721_ = new_n28016_ & ~new_n28720_;
  assign new_n28722_ = ~new_n27996_ & new_n28721_;
  assign ys__n26126 = new_n28703_ | new_n28722_;
  assign new_n28724_ = ys__n26029 & new_n27902_;
  assign new_n28725_ = ys__n46362 & new_n13490_;
  assign new_n28726_ = ys__n46538 & new_n13382_;
  assign new_n28727_ = ~new_n28725_ & ~new_n28726_;
  assign new_n28728_ = ys__n46714 & new_n13379_;
  assign new_n28729_ = ys__n46890 & new_n13380_;
  assign new_n28730_ = ~new_n28728_ & ~new_n28729_;
  assign new_n28731_ = new_n28727_ & new_n28730_;
  assign new_n28732_ = new_n27913_ & ~new_n28731_;
  assign new_n28733_ = ys__n46284 & new_n13490_;
  assign new_n28734_ = ys__n46460 & new_n13382_;
  assign new_n28735_ = ~new_n28733_ & ~new_n28734_;
  assign new_n28736_ = ys__n46636 & new_n13379_;
  assign new_n28737_ = ys__n46812 & new_n13380_;
  assign new_n28738_ = ~new_n28736_ & ~new_n28737_;
  assign new_n28739_ = new_n28735_ & new_n28738_;
  assign new_n28740_ = new_n27922_ & ~new_n28739_;
  assign new_n28741_ = ~new_n28732_ & ~new_n28740_;
  assign new_n28742_ = ys__n46331 & new_n13490_;
  assign new_n28743_ = ys__n46507 & new_n13382_;
  assign new_n28744_ = ~new_n28742_ & ~new_n28743_;
  assign new_n28745_ = ys__n46683 & new_n13379_;
  assign new_n28746_ = ys__n46859 & new_n13380_;
  assign new_n28747_ = ~new_n28745_ & ~new_n28746_;
  assign new_n28748_ = new_n28744_ & new_n28747_;
  assign new_n28749_ = new_n27932_ & ~new_n28748_;
  assign new_n28750_ = ys__n46408 & new_n13490_;
  assign new_n28751_ = ys__n46584 & new_n13382_;
  assign new_n28752_ = ~new_n28750_ & ~new_n28751_;
  assign new_n28753_ = ys__n46760 & new_n13379_;
  assign new_n28754_ = ys__n46936 & new_n13380_;
  assign new_n28755_ = ~new_n28753_ & ~new_n28754_;
  assign new_n28756_ = new_n28752_ & new_n28755_;
  assign new_n28757_ = new_n27941_ & ~new_n28756_;
  assign new_n28758_ = ~new_n28749_ & ~new_n28757_;
  assign new_n28759_ = new_n28741_ & new_n28758_;
  assign new_n28760_ = new_n27952_ & ~new_n28759_;
  assign new_n28761_ = ~new_n28724_ & ~new_n28760_;
  assign new_n28762_ = new_n27955_ & ~new_n28761_;
  assign new_n28763_ = ys__n45572 & new_n13490_;
  assign new_n28764_ = ys__n45408 & new_n13382_;
  assign new_n28765_ = ~new_n28763_ & ~new_n28764_;
  assign new_n28766_ = ys__n45244 & new_n13379_;
  assign new_n28767_ = ys__n45035 & new_n13380_;
  assign new_n28768_ = ~new_n28766_ & ~new_n28767_;
  assign new_n28769_ = new_n28765_ & new_n28768_;
  assign new_n28770_ = new_n27941_ & ~new_n28769_;
  assign new_n28771_ = ys__n45666 & new_n13490_;
  assign new_n28772_ = ys__n45502 & new_n13382_;
  assign new_n28773_ = ~new_n28771_ & ~new_n28772_;
  assign new_n28774_ = ys__n45338 & new_n13379_;
  assign new_n28775_ = ys__n45161 & new_n13380_;
  assign new_n28776_ = ~new_n28774_ & ~new_n28775_;
  assign new_n28777_ = new_n28773_ & new_n28776_;
  assign new_n28778_ = new_n27913_ & ~new_n28777_;
  assign new_n28779_ = ys__n45618 & new_n13490_;
  assign new_n28780_ = ys__n45454 & new_n13382_;
  assign new_n28781_ = ~new_n28779_ & ~new_n28780_;
  assign new_n28782_ = ys__n45290 & new_n13379_;
  assign new_n28783_ = ys__n45096 & new_n13380_;
  assign new_n28784_ = ~new_n28782_ & ~new_n28783_;
  assign new_n28785_ = new_n28781_ & new_n28784_;
  assign new_n28786_ = new_n27922_ & ~new_n28785_;
  assign new_n28787_ = ~new_n28778_ & ~new_n28786_;
  assign new_n28788_ = ~new_n28770_ & new_n28787_;
  assign new_n28789_ = new_n27993_ & ~new_n28788_;
  assign new_n28790_ = ~new_n28762_ & ~new_n28789_;
  assign new_n28791_ = new_n27996_ & ~new_n28790_;
  assign new_n28792_ = ys__n46111 & new_n13490_;
  assign new_n28793_ = ys__n46013 & new_n13382_;
  assign new_n28794_ = ~new_n28792_ & ~new_n28793_;
  assign new_n28795_ = ys__n45915 & new_n13379_;
  assign new_n28796_ = ys__n45819 & new_n13380_;
  assign new_n28797_ = ~new_n28795_ & ~new_n28796_;
  assign new_n28798_ = new_n28794_ & new_n28797_;
  assign new_n28799_ = new_n27922_ & ~new_n28798_;
  assign new_n28800_ = ys__n46064 & new_n13490_;
  assign new_n28801_ = ys__n45966 & new_n13382_;
  assign new_n28802_ = ~new_n28800_ & ~new_n28801_;
  assign new_n28803_ = ys__n45868 & new_n13379_;
  assign new_n28804_ = ys__n45757 & new_n13380_;
  assign new_n28805_ = ~new_n28803_ & ~new_n28804_;
  assign new_n28806_ = new_n28802_ & new_n28805_;
  assign new_n28807_ = new_n27941_ & ~new_n28806_;
  assign new_n28808_ = ~new_n28799_ & ~new_n28807_;
  assign new_n28809_ = new_n28016_ & ~new_n28808_;
  assign new_n28810_ = ~new_n27996_ & new_n28809_;
  assign ys__n26127 = new_n28791_ | new_n28810_;
  assign new_n28812_ = ys__n26032 & new_n27902_;
  assign new_n28813_ = ys__n46364 & new_n13490_;
  assign new_n28814_ = ys__n46540 & new_n13382_;
  assign new_n28815_ = ~new_n28813_ & ~new_n28814_;
  assign new_n28816_ = ys__n46716 & new_n13379_;
  assign new_n28817_ = ys__n46892 & new_n13380_;
  assign new_n28818_ = ~new_n28816_ & ~new_n28817_;
  assign new_n28819_ = new_n28815_ & new_n28818_;
  assign new_n28820_ = new_n27913_ & ~new_n28819_;
  assign new_n28821_ = ys__n46286 & new_n13490_;
  assign new_n28822_ = ys__n46462 & new_n13382_;
  assign new_n28823_ = ~new_n28821_ & ~new_n28822_;
  assign new_n28824_ = ys__n46638 & new_n13379_;
  assign new_n28825_ = ys__n46814 & new_n13380_;
  assign new_n28826_ = ~new_n28824_ & ~new_n28825_;
  assign new_n28827_ = new_n28823_ & new_n28826_;
  assign new_n28828_ = new_n27922_ & ~new_n28827_;
  assign new_n28829_ = ~new_n28820_ & ~new_n28828_;
  assign new_n28830_ = ys__n46332 & new_n13490_;
  assign new_n28831_ = ys__n46508 & new_n13382_;
  assign new_n28832_ = ~new_n28830_ & ~new_n28831_;
  assign new_n28833_ = ys__n46684 & new_n13379_;
  assign new_n28834_ = ys__n46860 & new_n13380_;
  assign new_n28835_ = ~new_n28833_ & ~new_n28834_;
  assign new_n28836_ = new_n28832_ & new_n28835_;
  assign new_n28837_ = new_n27932_ & ~new_n28836_;
  assign new_n28838_ = ys__n46409 & new_n13490_;
  assign new_n28839_ = ys__n46585 & new_n13382_;
  assign new_n28840_ = ~new_n28838_ & ~new_n28839_;
  assign new_n28841_ = ys__n46761 & new_n13379_;
  assign new_n28842_ = ys__n46937 & new_n13380_;
  assign new_n28843_ = ~new_n28841_ & ~new_n28842_;
  assign new_n28844_ = new_n28840_ & new_n28843_;
  assign new_n28845_ = new_n27941_ & ~new_n28844_;
  assign new_n28846_ = ~new_n28837_ & ~new_n28845_;
  assign new_n28847_ = new_n28829_ & new_n28846_;
  assign new_n28848_ = new_n27952_ & ~new_n28847_;
  assign new_n28849_ = ~new_n28812_ & ~new_n28848_;
  assign new_n28850_ = new_n27955_ & ~new_n28849_;
  assign new_n28851_ = ys__n45574 & new_n13490_;
  assign new_n28852_ = ys__n45410 & new_n13382_;
  assign new_n28853_ = ~new_n28851_ & ~new_n28852_;
  assign new_n28854_ = ys__n45246 & new_n13379_;
  assign new_n28855_ = ys__n45038 & new_n13380_;
  assign new_n28856_ = ~new_n28854_ & ~new_n28855_;
  assign new_n28857_ = new_n28853_ & new_n28856_;
  assign new_n28858_ = new_n27941_ & ~new_n28857_;
  assign new_n28859_ = ys__n45668 & new_n13490_;
  assign new_n28860_ = ys__n45504 & new_n13382_;
  assign new_n28861_ = ~new_n28859_ & ~new_n28860_;
  assign new_n28862_ = ys__n45340 & new_n13379_;
  assign new_n28863_ = ys__n45164 & new_n13380_;
  assign new_n28864_ = ~new_n28862_ & ~new_n28863_;
  assign new_n28865_ = new_n28861_ & new_n28864_;
  assign new_n28866_ = new_n27913_ & ~new_n28865_;
  assign new_n28867_ = ys__n45619 & new_n13490_;
  assign new_n28868_ = ys__n45455 & new_n13382_;
  assign new_n28869_ = ~new_n28867_ & ~new_n28868_;
  assign new_n28870_ = ys__n45291 & new_n13379_;
  assign new_n28871_ = ys__n45097 & new_n13380_;
  assign new_n28872_ = ~new_n28870_ & ~new_n28871_;
  assign new_n28873_ = new_n28869_ & new_n28872_;
  assign new_n28874_ = new_n27922_ & ~new_n28873_;
  assign new_n28875_ = ~new_n28866_ & ~new_n28874_;
  assign new_n28876_ = ~new_n28858_ & new_n28875_;
  assign new_n28877_ = new_n27993_ & ~new_n28876_;
  assign new_n28878_ = ~new_n28850_ & ~new_n28877_;
  assign new_n28879_ = new_n27996_ & ~new_n28878_;
  assign new_n28880_ = ys__n46112 & new_n13490_;
  assign new_n28881_ = ys__n46014 & new_n13382_;
  assign new_n28882_ = ~new_n28880_ & ~new_n28881_;
  assign new_n28883_ = ys__n45916 & new_n13379_;
  assign new_n28884_ = ys__n45820 & new_n13380_;
  assign new_n28885_ = ~new_n28883_ & ~new_n28884_;
  assign new_n28886_ = new_n28882_ & new_n28885_;
  assign new_n28887_ = new_n27922_ & ~new_n28886_;
  assign new_n28888_ = ys__n46066 & new_n13490_;
  assign new_n28889_ = ys__n45968 & new_n13382_;
  assign new_n28890_ = ~new_n28888_ & ~new_n28889_;
  assign new_n28891_ = ys__n45870 & new_n13379_;
  assign new_n28892_ = ys__n45760 & new_n13380_;
  assign new_n28893_ = ~new_n28891_ & ~new_n28892_;
  assign new_n28894_ = new_n28890_ & new_n28893_;
  assign new_n28895_ = new_n27941_ & ~new_n28894_;
  assign new_n28896_ = ~new_n28887_ & ~new_n28895_;
  assign new_n28897_ = new_n28016_ & ~new_n28896_;
  assign new_n28898_ = ~new_n27996_ & new_n28897_;
  assign ys__n26128 = new_n28879_ | new_n28898_;
  assign new_n28900_ = ys__n26035 & new_n27902_;
  assign new_n28901_ = ys__n46366 & new_n13490_;
  assign new_n28902_ = ys__n46542 & new_n13382_;
  assign new_n28903_ = ~new_n28901_ & ~new_n28902_;
  assign new_n28904_ = ys__n46718 & new_n13379_;
  assign new_n28905_ = ys__n46894 & new_n13380_;
  assign new_n28906_ = ~new_n28904_ & ~new_n28905_;
  assign new_n28907_ = new_n28903_ & new_n28906_;
  assign new_n28908_ = new_n27913_ & ~new_n28907_;
  assign new_n28909_ = ys__n46288 & new_n13490_;
  assign new_n28910_ = ys__n46464 & new_n13382_;
  assign new_n28911_ = ~new_n28909_ & ~new_n28910_;
  assign new_n28912_ = ys__n46640 & new_n13379_;
  assign new_n28913_ = ys__n46816 & new_n13380_;
  assign new_n28914_ = ~new_n28912_ & ~new_n28913_;
  assign new_n28915_ = new_n28911_ & new_n28914_;
  assign new_n28916_ = new_n27922_ & ~new_n28915_;
  assign new_n28917_ = ~new_n28908_ & ~new_n28916_;
  assign new_n28918_ = ys__n46333 & new_n13490_;
  assign new_n28919_ = ys__n46509 & new_n13382_;
  assign new_n28920_ = ~new_n28918_ & ~new_n28919_;
  assign new_n28921_ = ys__n46685 & new_n13379_;
  assign new_n28922_ = ys__n46861 & new_n13380_;
  assign new_n28923_ = ~new_n28921_ & ~new_n28922_;
  assign new_n28924_ = new_n28920_ & new_n28923_;
  assign new_n28925_ = new_n27932_ & ~new_n28924_;
  assign new_n28926_ = ys__n46410 & new_n13490_;
  assign new_n28927_ = ys__n46586 & new_n13382_;
  assign new_n28928_ = ~new_n28926_ & ~new_n28927_;
  assign new_n28929_ = ys__n46762 & new_n13379_;
  assign new_n28930_ = ys__n46938 & new_n13380_;
  assign new_n28931_ = ~new_n28929_ & ~new_n28930_;
  assign new_n28932_ = new_n28928_ & new_n28931_;
  assign new_n28933_ = new_n27941_ & ~new_n28932_;
  assign new_n28934_ = ~new_n28925_ & ~new_n28933_;
  assign new_n28935_ = new_n28917_ & new_n28934_;
  assign new_n28936_ = new_n27952_ & ~new_n28935_;
  assign new_n28937_ = ~new_n28900_ & ~new_n28936_;
  assign new_n28938_ = new_n27955_ & ~new_n28937_;
  assign new_n28939_ = ys__n45576 & new_n13490_;
  assign new_n28940_ = ys__n45412 & new_n13382_;
  assign new_n28941_ = ~new_n28939_ & ~new_n28940_;
  assign new_n28942_ = ys__n45248 & new_n13379_;
  assign new_n28943_ = ys__n45041 & new_n13380_;
  assign new_n28944_ = ~new_n28942_ & ~new_n28943_;
  assign new_n28945_ = new_n28941_ & new_n28944_;
  assign new_n28946_ = new_n27941_ & ~new_n28945_;
  assign new_n28947_ = ys__n45670 & new_n13490_;
  assign new_n28948_ = ys__n45506 & new_n13382_;
  assign new_n28949_ = ~new_n28947_ & ~new_n28948_;
  assign new_n28950_ = ys__n45342 & new_n13379_;
  assign new_n28951_ = ys__n45167 & new_n13380_;
  assign new_n28952_ = ~new_n28950_ & ~new_n28951_;
  assign new_n28953_ = new_n28949_ & new_n28952_;
  assign new_n28954_ = new_n27913_ & ~new_n28953_;
  assign new_n28955_ = ys__n45620 & new_n13490_;
  assign new_n28956_ = ys__n45456 & new_n13382_;
  assign new_n28957_ = ~new_n28955_ & ~new_n28956_;
  assign new_n28958_ = ys__n45292 & new_n13379_;
  assign new_n28959_ = ys__n45098 & new_n13380_;
  assign new_n28960_ = ~new_n28958_ & ~new_n28959_;
  assign new_n28961_ = new_n28957_ & new_n28960_;
  assign new_n28962_ = new_n27922_ & ~new_n28961_;
  assign new_n28963_ = ~new_n28954_ & ~new_n28962_;
  assign new_n28964_ = ~new_n28946_ & new_n28963_;
  assign new_n28965_ = new_n27993_ & ~new_n28964_;
  assign new_n28966_ = ~new_n28938_ & ~new_n28965_;
  assign new_n28967_ = new_n27996_ & ~new_n28966_;
  assign new_n28968_ = ys__n46113 & new_n13490_;
  assign new_n28969_ = ys__n46015 & new_n13382_;
  assign new_n28970_ = ~new_n28968_ & ~new_n28969_;
  assign new_n28971_ = ys__n45917 & new_n13379_;
  assign new_n28972_ = ys__n45821 & new_n13380_;
  assign new_n28973_ = ~new_n28971_ & ~new_n28972_;
  assign new_n28974_ = new_n28970_ & new_n28973_;
  assign new_n28975_ = new_n27922_ & ~new_n28974_;
  assign new_n28976_ = ys__n46068 & new_n13490_;
  assign new_n28977_ = ys__n45970 & new_n13382_;
  assign new_n28978_ = ~new_n28976_ & ~new_n28977_;
  assign new_n28979_ = ys__n45872 & new_n13379_;
  assign new_n28980_ = ys__n45763 & new_n13380_;
  assign new_n28981_ = ~new_n28979_ & ~new_n28980_;
  assign new_n28982_ = new_n28978_ & new_n28981_;
  assign new_n28983_ = new_n27941_ & ~new_n28982_;
  assign new_n28984_ = ~new_n28975_ & ~new_n28983_;
  assign new_n28985_ = new_n28016_ & ~new_n28984_;
  assign new_n28986_ = ~new_n27996_ & new_n28985_;
  assign ys__n26129 = new_n28967_ | new_n28986_;
  assign new_n28988_ = ys__n26038 & new_n27902_;
  assign new_n28989_ = ys__n46368 & new_n13490_;
  assign new_n28990_ = ys__n46544 & new_n13382_;
  assign new_n28991_ = ~new_n28989_ & ~new_n28990_;
  assign new_n28992_ = ys__n46720 & new_n13379_;
  assign new_n28993_ = ys__n46896 & new_n13380_;
  assign new_n28994_ = ~new_n28992_ & ~new_n28993_;
  assign new_n28995_ = new_n28991_ & new_n28994_;
  assign new_n28996_ = new_n27913_ & ~new_n28995_;
  assign new_n28997_ = ys__n46290 & new_n13490_;
  assign new_n28998_ = ys__n46466 & new_n13382_;
  assign new_n28999_ = ~new_n28997_ & ~new_n28998_;
  assign new_n29000_ = ys__n46642 & new_n13379_;
  assign new_n29001_ = ys__n46818 & new_n13380_;
  assign new_n29002_ = ~new_n29000_ & ~new_n29001_;
  assign new_n29003_ = new_n28999_ & new_n29002_;
  assign new_n29004_ = new_n27922_ & ~new_n29003_;
  assign new_n29005_ = ~new_n28996_ & ~new_n29004_;
  assign new_n29006_ = ys__n46334 & new_n13490_;
  assign new_n29007_ = ys__n46510 & new_n13382_;
  assign new_n29008_ = ~new_n29006_ & ~new_n29007_;
  assign new_n29009_ = ys__n46686 & new_n13379_;
  assign new_n29010_ = ys__n46862 & new_n13380_;
  assign new_n29011_ = ~new_n29009_ & ~new_n29010_;
  assign new_n29012_ = new_n29008_ & new_n29011_;
  assign new_n29013_ = new_n27932_ & ~new_n29012_;
  assign new_n29014_ = ys__n46411 & new_n13490_;
  assign new_n29015_ = ys__n46587 & new_n13382_;
  assign new_n29016_ = ~new_n29014_ & ~new_n29015_;
  assign new_n29017_ = ys__n46763 & new_n13379_;
  assign new_n29018_ = ys__n46939 & new_n13380_;
  assign new_n29019_ = ~new_n29017_ & ~new_n29018_;
  assign new_n29020_ = new_n29016_ & new_n29019_;
  assign new_n29021_ = new_n27941_ & ~new_n29020_;
  assign new_n29022_ = ~new_n29013_ & ~new_n29021_;
  assign new_n29023_ = new_n29005_ & new_n29022_;
  assign new_n29024_ = new_n27952_ & ~new_n29023_;
  assign new_n29025_ = ~new_n28988_ & ~new_n29024_;
  assign new_n29026_ = new_n27955_ & ~new_n29025_;
  assign new_n29027_ = ys__n45578 & new_n13490_;
  assign new_n29028_ = ys__n45414 & new_n13382_;
  assign new_n29029_ = ~new_n29027_ & ~new_n29028_;
  assign new_n29030_ = ys__n45250 & new_n13379_;
  assign new_n29031_ = ys__n45044 & new_n13380_;
  assign new_n29032_ = ~new_n29030_ & ~new_n29031_;
  assign new_n29033_ = new_n29029_ & new_n29032_;
  assign new_n29034_ = new_n27941_ & ~new_n29033_;
  assign new_n29035_ = ys__n45672 & new_n13490_;
  assign new_n29036_ = ys__n45508 & new_n13382_;
  assign new_n29037_ = ~new_n29035_ & ~new_n29036_;
  assign new_n29038_ = ys__n45344 & new_n13379_;
  assign new_n29039_ = ys__n45170 & new_n13380_;
  assign new_n29040_ = ~new_n29038_ & ~new_n29039_;
  assign new_n29041_ = new_n29037_ & new_n29040_;
  assign new_n29042_ = new_n27913_ & ~new_n29041_;
  assign new_n29043_ = ys__n45621 & new_n13490_;
  assign new_n29044_ = ys__n45457 & new_n13382_;
  assign new_n29045_ = ~new_n29043_ & ~new_n29044_;
  assign new_n29046_ = ys__n45293 & new_n13379_;
  assign new_n29047_ = ys__n45099 & new_n13380_;
  assign new_n29048_ = ~new_n29046_ & ~new_n29047_;
  assign new_n29049_ = new_n29045_ & new_n29048_;
  assign new_n29050_ = new_n27922_ & ~new_n29049_;
  assign new_n29051_ = ~new_n29042_ & ~new_n29050_;
  assign new_n29052_ = ~new_n29034_ & new_n29051_;
  assign new_n29053_ = new_n27993_ & ~new_n29052_;
  assign new_n29054_ = ~new_n29026_ & ~new_n29053_;
  assign new_n29055_ = new_n27996_ & ~new_n29054_;
  assign new_n29056_ = ys__n46114 & new_n13490_;
  assign new_n29057_ = ys__n46016 & new_n13382_;
  assign new_n29058_ = ~new_n29056_ & ~new_n29057_;
  assign new_n29059_ = ys__n45918 & new_n13379_;
  assign new_n29060_ = ys__n45822 & new_n13380_;
  assign new_n29061_ = ~new_n29059_ & ~new_n29060_;
  assign new_n29062_ = new_n29058_ & new_n29061_;
  assign new_n29063_ = new_n27922_ & ~new_n29062_;
  assign new_n29064_ = ys__n46070 & new_n13490_;
  assign new_n29065_ = ys__n45972 & new_n13382_;
  assign new_n29066_ = ~new_n29064_ & ~new_n29065_;
  assign new_n29067_ = ys__n45874 & new_n13379_;
  assign new_n29068_ = ys__n45766 & new_n13380_;
  assign new_n29069_ = ~new_n29067_ & ~new_n29068_;
  assign new_n29070_ = new_n29066_ & new_n29069_;
  assign new_n29071_ = new_n27941_ & ~new_n29070_;
  assign new_n29072_ = ~new_n29063_ & ~new_n29071_;
  assign new_n29073_ = new_n28016_ & ~new_n29072_;
  assign new_n29074_ = ~new_n27996_ & new_n29073_;
  assign ys__n26130 = new_n29055_ | new_n29074_;
  assign new_n29076_ = ys__n26041 & new_n27902_;
  assign new_n29077_ = ys__n46370 & new_n13490_;
  assign new_n29078_ = ys__n46546 & new_n13382_;
  assign new_n29079_ = ~new_n29077_ & ~new_n29078_;
  assign new_n29080_ = ys__n46722 & new_n13379_;
  assign new_n29081_ = ys__n46898 & new_n13380_;
  assign new_n29082_ = ~new_n29080_ & ~new_n29081_;
  assign new_n29083_ = new_n29079_ & new_n29082_;
  assign new_n29084_ = new_n27913_ & ~new_n29083_;
  assign new_n29085_ = ys__n46292 & new_n13490_;
  assign new_n29086_ = ys__n46468 & new_n13382_;
  assign new_n29087_ = ~new_n29085_ & ~new_n29086_;
  assign new_n29088_ = ys__n46644 & new_n13379_;
  assign new_n29089_ = ys__n46820 & new_n13380_;
  assign new_n29090_ = ~new_n29088_ & ~new_n29089_;
  assign new_n29091_ = new_n29087_ & new_n29090_;
  assign new_n29092_ = new_n27922_ & ~new_n29091_;
  assign new_n29093_ = ~new_n29084_ & ~new_n29092_;
  assign new_n29094_ = ys__n46335 & new_n13490_;
  assign new_n29095_ = ys__n46511 & new_n13382_;
  assign new_n29096_ = ~new_n29094_ & ~new_n29095_;
  assign new_n29097_ = ys__n46687 & new_n13379_;
  assign new_n29098_ = ys__n46863 & new_n13380_;
  assign new_n29099_ = ~new_n29097_ & ~new_n29098_;
  assign new_n29100_ = new_n29096_ & new_n29099_;
  assign new_n29101_ = new_n27932_ & ~new_n29100_;
  assign new_n29102_ = ys__n46412 & new_n13490_;
  assign new_n29103_ = ys__n46588 & new_n13382_;
  assign new_n29104_ = ~new_n29102_ & ~new_n29103_;
  assign new_n29105_ = ys__n46764 & new_n13379_;
  assign new_n29106_ = ys__n46940 & new_n13380_;
  assign new_n29107_ = ~new_n29105_ & ~new_n29106_;
  assign new_n29108_ = new_n29104_ & new_n29107_;
  assign new_n29109_ = new_n27941_ & ~new_n29108_;
  assign new_n29110_ = ~new_n29101_ & ~new_n29109_;
  assign new_n29111_ = new_n29093_ & new_n29110_;
  assign new_n29112_ = new_n27952_ & ~new_n29111_;
  assign new_n29113_ = ~new_n29076_ & ~new_n29112_;
  assign new_n29114_ = new_n27955_ & ~new_n29113_;
  assign new_n29115_ = ys__n45580 & new_n13490_;
  assign new_n29116_ = ys__n45416 & new_n13382_;
  assign new_n29117_ = ~new_n29115_ & ~new_n29116_;
  assign new_n29118_ = ys__n45252 & new_n13379_;
  assign new_n29119_ = ys__n45047 & new_n13380_;
  assign new_n29120_ = ~new_n29118_ & ~new_n29119_;
  assign new_n29121_ = new_n29117_ & new_n29120_;
  assign new_n29122_ = new_n27941_ & ~new_n29121_;
  assign new_n29123_ = ys__n45674 & new_n13490_;
  assign new_n29124_ = ys__n45510 & new_n13382_;
  assign new_n29125_ = ~new_n29123_ & ~new_n29124_;
  assign new_n29126_ = ys__n45346 & new_n13379_;
  assign new_n29127_ = ys__n45173 & new_n13380_;
  assign new_n29128_ = ~new_n29126_ & ~new_n29127_;
  assign new_n29129_ = new_n29125_ & new_n29128_;
  assign new_n29130_ = new_n27913_ & ~new_n29129_;
  assign new_n29131_ = ys__n45622 & new_n13490_;
  assign new_n29132_ = ys__n45458 & new_n13382_;
  assign new_n29133_ = ~new_n29131_ & ~new_n29132_;
  assign new_n29134_ = ys__n45294 & new_n13379_;
  assign new_n29135_ = ys__n45100 & new_n13380_;
  assign new_n29136_ = ~new_n29134_ & ~new_n29135_;
  assign new_n29137_ = new_n29133_ & new_n29136_;
  assign new_n29138_ = new_n27922_ & ~new_n29137_;
  assign new_n29139_ = ~new_n29130_ & ~new_n29138_;
  assign new_n29140_ = ~new_n29122_ & new_n29139_;
  assign new_n29141_ = new_n27993_ & ~new_n29140_;
  assign new_n29142_ = ~new_n29114_ & ~new_n29141_;
  assign new_n29143_ = new_n27996_ & ~new_n29142_;
  assign new_n29144_ = ys__n46115 & new_n13490_;
  assign new_n29145_ = ys__n46017 & new_n13382_;
  assign new_n29146_ = ~new_n29144_ & ~new_n29145_;
  assign new_n29147_ = ys__n45919 & new_n13379_;
  assign new_n29148_ = ys__n45823 & new_n13380_;
  assign new_n29149_ = ~new_n29147_ & ~new_n29148_;
  assign new_n29150_ = new_n29146_ & new_n29149_;
  assign new_n29151_ = new_n27922_ & ~new_n29150_;
  assign new_n29152_ = ys__n46072 & new_n13490_;
  assign new_n29153_ = ys__n45974 & new_n13382_;
  assign new_n29154_ = ~new_n29152_ & ~new_n29153_;
  assign new_n29155_ = ys__n45876 & new_n13379_;
  assign new_n29156_ = ys__n45769 & new_n13380_;
  assign new_n29157_ = ~new_n29155_ & ~new_n29156_;
  assign new_n29158_ = new_n29154_ & new_n29157_;
  assign new_n29159_ = new_n27941_ & ~new_n29158_;
  assign new_n29160_ = ~new_n29151_ & ~new_n29159_;
  assign new_n29161_ = new_n28016_ & ~new_n29160_;
  assign new_n29162_ = ~new_n27996_ & new_n29161_;
  assign ys__n26131 = new_n29143_ | new_n29162_;
  assign new_n29164_ = ys__n26044 & new_n27902_;
  assign new_n29165_ = ys__n46372 & new_n13490_;
  assign new_n29166_ = ys__n46548 & new_n13382_;
  assign new_n29167_ = ~new_n29165_ & ~new_n29166_;
  assign new_n29168_ = ys__n46724 & new_n13379_;
  assign new_n29169_ = ys__n46900 & new_n13380_;
  assign new_n29170_ = ~new_n29168_ & ~new_n29169_;
  assign new_n29171_ = new_n29167_ & new_n29170_;
  assign new_n29172_ = new_n27913_ & ~new_n29171_;
  assign new_n29173_ = ys__n46294 & new_n13490_;
  assign new_n29174_ = ys__n46470 & new_n13382_;
  assign new_n29175_ = ~new_n29173_ & ~new_n29174_;
  assign new_n29176_ = ys__n46646 & new_n13379_;
  assign new_n29177_ = ys__n46822 & new_n13380_;
  assign new_n29178_ = ~new_n29176_ & ~new_n29177_;
  assign new_n29179_ = new_n29175_ & new_n29178_;
  assign new_n29180_ = new_n27922_ & ~new_n29179_;
  assign new_n29181_ = ~new_n29172_ & ~new_n29180_;
  assign new_n29182_ = ys__n46336 & new_n13490_;
  assign new_n29183_ = ys__n46512 & new_n13382_;
  assign new_n29184_ = ~new_n29182_ & ~new_n29183_;
  assign new_n29185_ = ys__n46688 & new_n13379_;
  assign new_n29186_ = ys__n46864 & new_n13380_;
  assign new_n29187_ = ~new_n29185_ & ~new_n29186_;
  assign new_n29188_ = new_n29184_ & new_n29187_;
  assign new_n29189_ = new_n27932_ & ~new_n29188_;
  assign new_n29190_ = ys__n46413 & new_n13490_;
  assign new_n29191_ = ys__n46589 & new_n13382_;
  assign new_n29192_ = ~new_n29190_ & ~new_n29191_;
  assign new_n29193_ = ys__n46765 & new_n13379_;
  assign new_n29194_ = ys__n46941 & new_n13380_;
  assign new_n29195_ = ~new_n29193_ & ~new_n29194_;
  assign new_n29196_ = new_n29192_ & new_n29195_;
  assign new_n29197_ = new_n27941_ & ~new_n29196_;
  assign new_n29198_ = ~new_n29189_ & ~new_n29197_;
  assign new_n29199_ = new_n29181_ & new_n29198_;
  assign new_n29200_ = new_n27952_ & ~new_n29199_;
  assign new_n29201_ = ~new_n29164_ & ~new_n29200_;
  assign new_n29202_ = new_n27955_ & ~new_n29201_;
  assign new_n29203_ = ys__n45582 & new_n13490_;
  assign new_n29204_ = ys__n45418 & new_n13382_;
  assign new_n29205_ = ~new_n29203_ & ~new_n29204_;
  assign new_n29206_ = ys__n45254 & new_n13379_;
  assign new_n29207_ = ys__n45050 & new_n13380_;
  assign new_n29208_ = ~new_n29206_ & ~new_n29207_;
  assign new_n29209_ = new_n29205_ & new_n29208_;
  assign new_n29210_ = new_n27941_ & ~new_n29209_;
  assign new_n29211_ = ys__n45676 & new_n13490_;
  assign new_n29212_ = ys__n45512 & new_n13382_;
  assign new_n29213_ = ~new_n29211_ & ~new_n29212_;
  assign new_n29214_ = ys__n45348 & new_n13379_;
  assign new_n29215_ = ys__n45176 & new_n13380_;
  assign new_n29216_ = ~new_n29214_ & ~new_n29215_;
  assign new_n29217_ = new_n29213_ & new_n29216_;
  assign new_n29218_ = new_n27913_ & ~new_n29217_;
  assign new_n29219_ = ys__n45623 & new_n13490_;
  assign new_n29220_ = ys__n45459 & new_n13382_;
  assign new_n29221_ = ~new_n29219_ & ~new_n29220_;
  assign new_n29222_ = ys__n45295 & new_n13379_;
  assign new_n29223_ = ys__n45101 & new_n13380_;
  assign new_n29224_ = ~new_n29222_ & ~new_n29223_;
  assign new_n29225_ = new_n29221_ & new_n29224_;
  assign new_n29226_ = new_n27922_ & ~new_n29225_;
  assign new_n29227_ = ~new_n29218_ & ~new_n29226_;
  assign new_n29228_ = ~new_n29210_ & new_n29227_;
  assign new_n29229_ = new_n27993_ & ~new_n29228_;
  assign new_n29230_ = ~new_n29202_ & ~new_n29229_;
  assign new_n29231_ = new_n27996_ & ~new_n29230_;
  assign new_n29232_ = ys__n46116 & new_n13490_;
  assign new_n29233_ = ys__n46018 & new_n13382_;
  assign new_n29234_ = ~new_n29232_ & ~new_n29233_;
  assign new_n29235_ = ys__n45920 & new_n13379_;
  assign new_n29236_ = ys__n45824 & new_n13380_;
  assign new_n29237_ = ~new_n29235_ & ~new_n29236_;
  assign new_n29238_ = new_n29234_ & new_n29237_;
  assign new_n29239_ = new_n27922_ & ~new_n29238_;
  assign new_n29240_ = ys__n46074 & new_n13490_;
  assign new_n29241_ = ys__n45976 & new_n13382_;
  assign new_n29242_ = ~new_n29240_ & ~new_n29241_;
  assign new_n29243_ = ys__n45878 & new_n13379_;
  assign new_n29244_ = ys__n45772 & new_n13380_;
  assign new_n29245_ = ~new_n29243_ & ~new_n29244_;
  assign new_n29246_ = new_n29242_ & new_n29245_;
  assign new_n29247_ = new_n27941_ & ~new_n29246_;
  assign new_n29248_ = ~new_n29239_ & ~new_n29247_;
  assign new_n29249_ = new_n28016_ & ~new_n29248_;
  assign new_n29250_ = ~new_n27996_ & new_n29249_;
  assign ys__n26132 = new_n29231_ | new_n29250_;
  assign new_n29252_ = ys__n26047 & new_n27902_;
  assign new_n29253_ = ys__n46374 & new_n13490_;
  assign new_n29254_ = ys__n46550 & new_n13382_;
  assign new_n29255_ = ~new_n29253_ & ~new_n29254_;
  assign new_n29256_ = ys__n46726 & new_n13379_;
  assign new_n29257_ = ys__n46902 & new_n13380_;
  assign new_n29258_ = ~new_n29256_ & ~new_n29257_;
  assign new_n29259_ = new_n29255_ & new_n29258_;
  assign new_n29260_ = new_n27913_ & ~new_n29259_;
  assign new_n29261_ = ys__n46296 & new_n13490_;
  assign new_n29262_ = ys__n46472 & new_n13382_;
  assign new_n29263_ = ~new_n29261_ & ~new_n29262_;
  assign new_n29264_ = ys__n46648 & new_n13379_;
  assign new_n29265_ = ys__n46824 & new_n13380_;
  assign new_n29266_ = ~new_n29264_ & ~new_n29265_;
  assign new_n29267_ = new_n29263_ & new_n29266_;
  assign new_n29268_ = new_n27922_ & ~new_n29267_;
  assign new_n29269_ = ~new_n29260_ & ~new_n29268_;
  assign new_n29270_ = ys__n46337 & new_n13490_;
  assign new_n29271_ = ys__n46513 & new_n13382_;
  assign new_n29272_ = ~new_n29270_ & ~new_n29271_;
  assign new_n29273_ = ys__n46689 & new_n13379_;
  assign new_n29274_ = ys__n46865 & new_n13380_;
  assign new_n29275_ = ~new_n29273_ & ~new_n29274_;
  assign new_n29276_ = new_n29272_ & new_n29275_;
  assign new_n29277_ = new_n27932_ & ~new_n29276_;
  assign new_n29278_ = ys__n46414 & new_n13490_;
  assign new_n29279_ = ys__n46590 & new_n13382_;
  assign new_n29280_ = ~new_n29278_ & ~new_n29279_;
  assign new_n29281_ = ys__n46766 & new_n13379_;
  assign new_n29282_ = ys__n46942 & new_n13380_;
  assign new_n29283_ = ~new_n29281_ & ~new_n29282_;
  assign new_n29284_ = new_n29280_ & new_n29283_;
  assign new_n29285_ = new_n27941_ & ~new_n29284_;
  assign new_n29286_ = ~new_n29277_ & ~new_n29285_;
  assign new_n29287_ = new_n29269_ & new_n29286_;
  assign new_n29288_ = new_n27952_ & ~new_n29287_;
  assign new_n29289_ = ~new_n29252_ & ~new_n29288_;
  assign new_n29290_ = new_n27955_ & ~new_n29289_;
  assign new_n29291_ = ys__n45584 & new_n13490_;
  assign new_n29292_ = ys__n45420 & new_n13382_;
  assign new_n29293_ = ~new_n29291_ & ~new_n29292_;
  assign new_n29294_ = ys__n45256 & new_n13379_;
  assign new_n29295_ = ys__n45053 & new_n13380_;
  assign new_n29296_ = ~new_n29294_ & ~new_n29295_;
  assign new_n29297_ = new_n29293_ & new_n29296_;
  assign new_n29298_ = new_n27941_ & ~new_n29297_;
  assign new_n29299_ = ys__n45678 & new_n13490_;
  assign new_n29300_ = ys__n45514 & new_n13382_;
  assign new_n29301_ = ~new_n29299_ & ~new_n29300_;
  assign new_n29302_ = ys__n45350 & new_n13379_;
  assign new_n29303_ = ys__n45179 & new_n13380_;
  assign new_n29304_ = ~new_n29302_ & ~new_n29303_;
  assign new_n29305_ = new_n29301_ & new_n29304_;
  assign new_n29306_ = new_n27913_ & ~new_n29305_;
  assign new_n29307_ = ys__n45624 & new_n13490_;
  assign new_n29308_ = ys__n45460 & new_n13382_;
  assign new_n29309_ = ~new_n29307_ & ~new_n29308_;
  assign new_n29310_ = ys__n45296 & new_n13379_;
  assign new_n29311_ = ys__n45102 & new_n13380_;
  assign new_n29312_ = ~new_n29310_ & ~new_n29311_;
  assign new_n29313_ = new_n29309_ & new_n29312_;
  assign new_n29314_ = new_n27922_ & ~new_n29313_;
  assign new_n29315_ = ~new_n29306_ & ~new_n29314_;
  assign new_n29316_ = ~new_n29298_ & new_n29315_;
  assign new_n29317_ = new_n27993_ & ~new_n29316_;
  assign new_n29318_ = ~new_n29290_ & ~new_n29317_;
  assign new_n29319_ = new_n27996_ & ~new_n29318_;
  assign new_n29320_ = ys__n46117 & new_n13490_;
  assign new_n29321_ = ys__n46019 & new_n13382_;
  assign new_n29322_ = ~new_n29320_ & ~new_n29321_;
  assign new_n29323_ = ys__n45921 & new_n13379_;
  assign new_n29324_ = ys__n45825 & new_n13380_;
  assign new_n29325_ = ~new_n29323_ & ~new_n29324_;
  assign new_n29326_ = new_n29322_ & new_n29325_;
  assign new_n29327_ = new_n27922_ & ~new_n29326_;
  assign new_n29328_ = ys__n46076 & new_n13490_;
  assign new_n29329_ = ys__n45978 & new_n13382_;
  assign new_n29330_ = ~new_n29328_ & ~new_n29329_;
  assign new_n29331_ = ys__n45880 & new_n13379_;
  assign new_n29332_ = ys__n45775 & new_n13380_;
  assign new_n29333_ = ~new_n29331_ & ~new_n29332_;
  assign new_n29334_ = new_n29330_ & new_n29333_;
  assign new_n29335_ = new_n27941_ & ~new_n29334_;
  assign new_n29336_ = ~new_n29327_ & ~new_n29335_;
  assign new_n29337_ = new_n28016_ & ~new_n29336_;
  assign new_n29338_ = ~new_n27996_ & new_n29337_;
  assign ys__n26133 = new_n29319_ | new_n29338_;
  assign new_n29340_ = ys__n26050 & new_n27902_;
  assign new_n29341_ = ys__n46376 & new_n13490_;
  assign new_n29342_ = ys__n46552 & new_n13382_;
  assign new_n29343_ = ~new_n29341_ & ~new_n29342_;
  assign new_n29344_ = ys__n46728 & new_n13379_;
  assign new_n29345_ = ys__n46904 & new_n13380_;
  assign new_n29346_ = ~new_n29344_ & ~new_n29345_;
  assign new_n29347_ = new_n29343_ & new_n29346_;
  assign new_n29348_ = new_n27913_ & ~new_n29347_;
  assign new_n29349_ = ys__n46298 & new_n13490_;
  assign new_n29350_ = ys__n46474 & new_n13382_;
  assign new_n29351_ = ~new_n29349_ & ~new_n29350_;
  assign new_n29352_ = ys__n46650 & new_n13379_;
  assign new_n29353_ = ys__n46826 & new_n13380_;
  assign new_n29354_ = ~new_n29352_ & ~new_n29353_;
  assign new_n29355_ = new_n29351_ & new_n29354_;
  assign new_n29356_ = new_n27922_ & ~new_n29355_;
  assign new_n29357_ = ~new_n29348_ & ~new_n29356_;
  assign new_n29358_ = ys__n46338 & new_n13490_;
  assign new_n29359_ = ys__n46514 & new_n13382_;
  assign new_n29360_ = ~new_n29358_ & ~new_n29359_;
  assign new_n29361_ = ys__n46690 & new_n13379_;
  assign new_n29362_ = ys__n46866 & new_n13380_;
  assign new_n29363_ = ~new_n29361_ & ~new_n29362_;
  assign new_n29364_ = new_n29360_ & new_n29363_;
  assign new_n29365_ = new_n27932_ & ~new_n29364_;
  assign new_n29366_ = ys__n46415 & new_n13490_;
  assign new_n29367_ = ys__n46591 & new_n13382_;
  assign new_n29368_ = ~new_n29366_ & ~new_n29367_;
  assign new_n29369_ = ys__n46767 & new_n13379_;
  assign new_n29370_ = ys__n46943 & new_n13380_;
  assign new_n29371_ = ~new_n29369_ & ~new_n29370_;
  assign new_n29372_ = new_n29368_ & new_n29371_;
  assign new_n29373_ = new_n27941_ & ~new_n29372_;
  assign new_n29374_ = ~new_n29365_ & ~new_n29373_;
  assign new_n29375_ = new_n29357_ & new_n29374_;
  assign new_n29376_ = new_n27952_ & ~new_n29375_;
  assign new_n29377_ = ~new_n29340_ & ~new_n29376_;
  assign new_n29378_ = new_n27955_ & ~new_n29377_;
  assign new_n29379_ = ys__n45586 & new_n13490_;
  assign new_n29380_ = ys__n45422 & new_n13382_;
  assign new_n29381_ = ~new_n29379_ & ~new_n29380_;
  assign new_n29382_ = ys__n45258 & new_n13379_;
  assign new_n29383_ = ys__n45056 & new_n13380_;
  assign new_n29384_ = ~new_n29382_ & ~new_n29383_;
  assign new_n29385_ = new_n29381_ & new_n29384_;
  assign new_n29386_ = new_n27941_ & ~new_n29385_;
  assign new_n29387_ = ys__n45680 & new_n13490_;
  assign new_n29388_ = ys__n45516 & new_n13382_;
  assign new_n29389_ = ~new_n29387_ & ~new_n29388_;
  assign new_n29390_ = ys__n45352 & new_n13379_;
  assign new_n29391_ = ys__n45182 & new_n13380_;
  assign new_n29392_ = ~new_n29390_ & ~new_n29391_;
  assign new_n29393_ = new_n29389_ & new_n29392_;
  assign new_n29394_ = new_n27913_ & ~new_n29393_;
  assign new_n29395_ = ys__n45625 & new_n13490_;
  assign new_n29396_ = ys__n45461 & new_n13382_;
  assign new_n29397_ = ~new_n29395_ & ~new_n29396_;
  assign new_n29398_ = ys__n45297 & new_n13379_;
  assign new_n29399_ = ys__n45103 & new_n13380_;
  assign new_n29400_ = ~new_n29398_ & ~new_n29399_;
  assign new_n29401_ = new_n29397_ & new_n29400_;
  assign new_n29402_ = new_n27922_ & ~new_n29401_;
  assign new_n29403_ = ~new_n29394_ & ~new_n29402_;
  assign new_n29404_ = ~new_n29386_ & new_n29403_;
  assign new_n29405_ = new_n27993_ & ~new_n29404_;
  assign new_n29406_ = ~new_n29378_ & ~new_n29405_;
  assign new_n29407_ = new_n27996_ & ~new_n29406_;
  assign new_n29408_ = ys__n46118 & new_n13490_;
  assign new_n29409_ = ys__n46020 & new_n13382_;
  assign new_n29410_ = ~new_n29408_ & ~new_n29409_;
  assign new_n29411_ = ys__n45922 & new_n13379_;
  assign new_n29412_ = ys__n45826 & new_n13380_;
  assign new_n29413_ = ~new_n29411_ & ~new_n29412_;
  assign new_n29414_ = new_n29410_ & new_n29413_;
  assign new_n29415_ = new_n27922_ & ~new_n29414_;
  assign new_n29416_ = ys__n46078 & new_n13490_;
  assign new_n29417_ = ys__n45980 & new_n13382_;
  assign new_n29418_ = ~new_n29416_ & ~new_n29417_;
  assign new_n29419_ = ys__n45882 & new_n13379_;
  assign new_n29420_ = ys__n45778 & new_n13380_;
  assign new_n29421_ = ~new_n29419_ & ~new_n29420_;
  assign new_n29422_ = new_n29418_ & new_n29421_;
  assign new_n29423_ = new_n27941_ & ~new_n29422_;
  assign new_n29424_ = ~new_n29415_ & ~new_n29423_;
  assign new_n29425_ = new_n28016_ & ~new_n29424_;
  assign new_n29426_ = ~new_n27996_ & new_n29425_;
  assign ys__n26134 = new_n29407_ | new_n29426_;
  assign new_n29428_ = ys__n26053 & new_n27902_;
  assign new_n29429_ = ys__n46378 & new_n13490_;
  assign new_n29430_ = ys__n46554 & new_n13382_;
  assign new_n29431_ = ~new_n29429_ & ~new_n29430_;
  assign new_n29432_ = ys__n46730 & new_n13379_;
  assign new_n29433_ = ys__n46906 & new_n13380_;
  assign new_n29434_ = ~new_n29432_ & ~new_n29433_;
  assign new_n29435_ = new_n29431_ & new_n29434_;
  assign new_n29436_ = new_n27913_ & ~new_n29435_;
  assign new_n29437_ = ys__n46300 & new_n13490_;
  assign new_n29438_ = ys__n46476 & new_n13382_;
  assign new_n29439_ = ~new_n29437_ & ~new_n29438_;
  assign new_n29440_ = ys__n46652 & new_n13379_;
  assign new_n29441_ = ys__n46828 & new_n13380_;
  assign new_n29442_ = ~new_n29440_ & ~new_n29441_;
  assign new_n29443_ = new_n29439_ & new_n29442_;
  assign new_n29444_ = new_n27922_ & ~new_n29443_;
  assign new_n29445_ = ~new_n29436_ & ~new_n29444_;
  assign new_n29446_ = ys__n46339 & new_n13490_;
  assign new_n29447_ = ys__n46515 & new_n13382_;
  assign new_n29448_ = ~new_n29446_ & ~new_n29447_;
  assign new_n29449_ = ys__n46691 & new_n13379_;
  assign new_n29450_ = ys__n46867 & new_n13380_;
  assign new_n29451_ = ~new_n29449_ & ~new_n29450_;
  assign new_n29452_ = new_n29448_ & new_n29451_;
  assign new_n29453_ = new_n27932_ & ~new_n29452_;
  assign new_n29454_ = ys__n46416 & new_n13490_;
  assign new_n29455_ = ys__n46592 & new_n13382_;
  assign new_n29456_ = ~new_n29454_ & ~new_n29455_;
  assign new_n29457_ = ys__n46768 & new_n13379_;
  assign new_n29458_ = ys__n46944 & new_n13380_;
  assign new_n29459_ = ~new_n29457_ & ~new_n29458_;
  assign new_n29460_ = new_n29456_ & new_n29459_;
  assign new_n29461_ = new_n27941_ & ~new_n29460_;
  assign new_n29462_ = ~new_n29453_ & ~new_n29461_;
  assign new_n29463_ = new_n29445_ & new_n29462_;
  assign new_n29464_ = new_n27952_ & ~new_n29463_;
  assign new_n29465_ = ~new_n29428_ & ~new_n29464_;
  assign new_n29466_ = new_n27955_ & ~new_n29465_;
  assign new_n29467_ = ys__n45588 & new_n13490_;
  assign new_n29468_ = ys__n45424 & new_n13382_;
  assign new_n29469_ = ~new_n29467_ & ~new_n29468_;
  assign new_n29470_ = ys__n45260 & new_n13379_;
  assign new_n29471_ = ys__n45059 & new_n13380_;
  assign new_n29472_ = ~new_n29470_ & ~new_n29471_;
  assign new_n29473_ = new_n29469_ & new_n29472_;
  assign new_n29474_ = new_n27941_ & ~new_n29473_;
  assign new_n29475_ = ys__n45682 & new_n13490_;
  assign new_n29476_ = ys__n45518 & new_n13382_;
  assign new_n29477_ = ~new_n29475_ & ~new_n29476_;
  assign new_n29478_ = ys__n45354 & new_n13379_;
  assign new_n29479_ = ys__n45185 & new_n13380_;
  assign new_n29480_ = ~new_n29478_ & ~new_n29479_;
  assign new_n29481_ = new_n29477_ & new_n29480_;
  assign new_n29482_ = new_n27913_ & ~new_n29481_;
  assign new_n29483_ = ys__n45626 & new_n13490_;
  assign new_n29484_ = ys__n45462 & new_n13382_;
  assign new_n29485_ = ~new_n29483_ & ~new_n29484_;
  assign new_n29486_ = ys__n45298 & new_n13379_;
  assign new_n29487_ = ys__n45104 & new_n13380_;
  assign new_n29488_ = ~new_n29486_ & ~new_n29487_;
  assign new_n29489_ = new_n29485_ & new_n29488_;
  assign new_n29490_ = new_n27922_ & ~new_n29489_;
  assign new_n29491_ = ~new_n29482_ & ~new_n29490_;
  assign new_n29492_ = ~new_n29474_ & new_n29491_;
  assign new_n29493_ = new_n27993_ & ~new_n29492_;
  assign new_n29494_ = ~new_n29466_ & ~new_n29493_;
  assign new_n29495_ = new_n27996_ & ~new_n29494_;
  assign new_n29496_ = ys__n46119 & new_n13490_;
  assign new_n29497_ = ys__n46021 & new_n13382_;
  assign new_n29498_ = ~new_n29496_ & ~new_n29497_;
  assign new_n29499_ = ys__n45923 & new_n13379_;
  assign new_n29500_ = ys__n45827 & new_n13380_;
  assign new_n29501_ = ~new_n29499_ & ~new_n29500_;
  assign new_n29502_ = new_n29498_ & new_n29501_;
  assign new_n29503_ = new_n27922_ & ~new_n29502_;
  assign new_n29504_ = ys__n46080 & new_n13490_;
  assign new_n29505_ = ys__n45982 & new_n13382_;
  assign new_n29506_ = ~new_n29504_ & ~new_n29505_;
  assign new_n29507_ = ys__n45884 & new_n13379_;
  assign new_n29508_ = ys__n45781 & new_n13380_;
  assign new_n29509_ = ~new_n29507_ & ~new_n29508_;
  assign new_n29510_ = new_n29506_ & new_n29509_;
  assign new_n29511_ = new_n27941_ & ~new_n29510_;
  assign new_n29512_ = ~new_n29503_ & ~new_n29511_;
  assign new_n29513_ = new_n28016_ & ~new_n29512_;
  assign new_n29514_ = ~new_n27996_ & new_n29513_;
  assign ys__n26135 = new_n29495_ | new_n29514_;
  assign new_n29516_ = ys__n26056 & new_n27902_;
  assign new_n29517_ = ys__n46380 & new_n13490_;
  assign new_n29518_ = ys__n46556 & new_n13382_;
  assign new_n29519_ = ~new_n29517_ & ~new_n29518_;
  assign new_n29520_ = ys__n46732 & new_n13379_;
  assign new_n29521_ = ys__n46908 & new_n13380_;
  assign new_n29522_ = ~new_n29520_ & ~new_n29521_;
  assign new_n29523_ = new_n29519_ & new_n29522_;
  assign new_n29524_ = new_n27913_ & ~new_n29523_;
  assign new_n29525_ = ys__n46302 & new_n13490_;
  assign new_n29526_ = ys__n46478 & new_n13382_;
  assign new_n29527_ = ~new_n29525_ & ~new_n29526_;
  assign new_n29528_ = ys__n46654 & new_n13379_;
  assign new_n29529_ = ys__n46830 & new_n13380_;
  assign new_n29530_ = ~new_n29528_ & ~new_n29529_;
  assign new_n29531_ = new_n29527_ & new_n29530_;
  assign new_n29532_ = new_n27922_ & ~new_n29531_;
  assign new_n29533_ = ~new_n29524_ & ~new_n29532_;
  assign new_n29534_ = ys__n46340 & new_n13490_;
  assign new_n29535_ = ys__n46516 & new_n13382_;
  assign new_n29536_ = ~new_n29534_ & ~new_n29535_;
  assign new_n29537_ = ys__n46692 & new_n13379_;
  assign new_n29538_ = ys__n46868 & new_n13380_;
  assign new_n29539_ = ~new_n29537_ & ~new_n29538_;
  assign new_n29540_ = new_n29536_ & new_n29539_;
  assign new_n29541_ = new_n27932_ & ~new_n29540_;
  assign new_n29542_ = ys__n46417 & new_n13490_;
  assign new_n29543_ = ys__n46593 & new_n13382_;
  assign new_n29544_ = ~new_n29542_ & ~new_n29543_;
  assign new_n29545_ = ys__n46769 & new_n13379_;
  assign new_n29546_ = ys__n46945 & new_n13380_;
  assign new_n29547_ = ~new_n29545_ & ~new_n29546_;
  assign new_n29548_ = new_n29544_ & new_n29547_;
  assign new_n29549_ = new_n27941_ & ~new_n29548_;
  assign new_n29550_ = ~new_n29541_ & ~new_n29549_;
  assign new_n29551_ = new_n29533_ & new_n29550_;
  assign new_n29552_ = new_n27952_ & ~new_n29551_;
  assign new_n29553_ = ~new_n29516_ & ~new_n29552_;
  assign new_n29554_ = new_n27955_ & ~new_n29553_;
  assign new_n29555_ = ys__n45590 & new_n13490_;
  assign new_n29556_ = ys__n45426 & new_n13382_;
  assign new_n29557_ = ~new_n29555_ & ~new_n29556_;
  assign new_n29558_ = ys__n45262 & new_n13379_;
  assign new_n29559_ = ys__n45062 & new_n13380_;
  assign new_n29560_ = ~new_n29558_ & ~new_n29559_;
  assign new_n29561_ = new_n29557_ & new_n29560_;
  assign new_n29562_ = new_n27941_ & ~new_n29561_;
  assign new_n29563_ = ys__n45684 & new_n13490_;
  assign new_n29564_ = ys__n45520 & new_n13382_;
  assign new_n29565_ = ~new_n29563_ & ~new_n29564_;
  assign new_n29566_ = ys__n45356 & new_n13379_;
  assign new_n29567_ = ys__n45188 & new_n13380_;
  assign new_n29568_ = ~new_n29566_ & ~new_n29567_;
  assign new_n29569_ = new_n29565_ & new_n29568_;
  assign new_n29570_ = new_n27913_ & ~new_n29569_;
  assign new_n29571_ = ys__n45627 & new_n13490_;
  assign new_n29572_ = ys__n45463 & new_n13382_;
  assign new_n29573_ = ~new_n29571_ & ~new_n29572_;
  assign new_n29574_ = ys__n45299 & new_n13379_;
  assign new_n29575_ = ys__n45105 & new_n13380_;
  assign new_n29576_ = ~new_n29574_ & ~new_n29575_;
  assign new_n29577_ = new_n29573_ & new_n29576_;
  assign new_n29578_ = new_n27922_ & ~new_n29577_;
  assign new_n29579_ = ~new_n29570_ & ~new_n29578_;
  assign new_n29580_ = ~new_n29562_ & new_n29579_;
  assign new_n29581_ = new_n27993_ & ~new_n29580_;
  assign new_n29582_ = ~new_n29554_ & ~new_n29581_;
  assign new_n29583_ = new_n27996_ & ~new_n29582_;
  assign new_n29584_ = ys__n46120 & new_n13490_;
  assign new_n29585_ = ys__n46022 & new_n13382_;
  assign new_n29586_ = ~new_n29584_ & ~new_n29585_;
  assign new_n29587_ = ys__n45924 & new_n13379_;
  assign new_n29588_ = ys__n45828 & new_n13380_;
  assign new_n29589_ = ~new_n29587_ & ~new_n29588_;
  assign new_n29590_ = new_n29586_ & new_n29589_;
  assign new_n29591_ = new_n27922_ & ~new_n29590_;
  assign new_n29592_ = ys__n46082 & new_n13490_;
  assign new_n29593_ = ys__n45984 & new_n13382_;
  assign new_n29594_ = ~new_n29592_ & ~new_n29593_;
  assign new_n29595_ = ys__n45886 & new_n13379_;
  assign new_n29596_ = ys__n45784 & new_n13380_;
  assign new_n29597_ = ~new_n29595_ & ~new_n29596_;
  assign new_n29598_ = new_n29594_ & new_n29597_;
  assign new_n29599_ = new_n27941_ & ~new_n29598_;
  assign new_n29600_ = ~new_n29591_ & ~new_n29599_;
  assign new_n29601_ = new_n28016_ & ~new_n29600_;
  assign new_n29602_ = ~new_n27996_ & new_n29601_;
  assign ys__n26136 = new_n29583_ | new_n29602_;
  assign new_n29604_ = ys__n26059 & new_n27902_;
  assign new_n29605_ = ys__n46382 & new_n13490_;
  assign new_n29606_ = ys__n46558 & new_n13382_;
  assign new_n29607_ = ~new_n29605_ & ~new_n29606_;
  assign new_n29608_ = ys__n46734 & new_n13379_;
  assign new_n29609_ = ys__n46910 & new_n13380_;
  assign new_n29610_ = ~new_n29608_ & ~new_n29609_;
  assign new_n29611_ = new_n29607_ & new_n29610_;
  assign new_n29612_ = new_n27913_ & ~new_n29611_;
  assign new_n29613_ = ys__n46304 & new_n13490_;
  assign new_n29614_ = ys__n46480 & new_n13382_;
  assign new_n29615_ = ~new_n29613_ & ~new_n29614_;
  assign new_n29616_ = ys__n46656 & new_n13379_;
  assign new_n29617_ = ys__n46832 & new_n13380_;
  assign new_n29618_ = ~new_n29616_ & ~new_n29617_;
  assign new_n29619_ = new_n29615_ & new_n29618_;
  assign new_n29620_ = new_n27922_ & ~new_n29619_;
  assign new_n29621_ = ~new_n29612_ & ~new_n29620_;
  assign new_n29622_ = ys__n46341 & new_n13490_;
  assign new_n29623_ = ys__n46517 & new_n13382_;
  assign new_n29624_ = ~new_n29622_ & ~new_n29623_;
  assign new_n29625_ = ys__n46693 & new_n13379_;
  assign new_n29626_ = ys__n46869 & new_n13380_;
  assign new_n29627_ = ~new_n29625_ & ~new_n29626_;
  assign new_n29628_ = new_n29624_ & new_n29627_;
  assign new_n29629_ = new_n27932_ & ~new_n29628_;
  assign new_n29630_ = ys__n46418 & new_n13490_;
  assign new_n29631_ = ys__n46594 & new_n13382_;
  assign new_n29632_ = ~new_n29630_ & ~new_n29631_;
  assign new_n29633_ = ys__n46770 & new_n13379_;
  assign new_n29634_ = ys__n46946 & new_n13380_;
  assign new_n29635_ = ~new_n29633_ & ~new_n29634_;
  assign new_n29636_ = new_n29632_ & new_n29635_;
  assign new_n29637_ = new_n27941_ & ~new_n29636_;
  assign new_n29638_ = ~new_n29629_ & ~new_n29637_;
  assign new_n29639_ = new_n29621_ & new_n29638_;
  assign new_n29640_ = new_n27951_ & ~new_n29639_;
  assign new_n29641_ = new_n13499_ & ~new_n29640_;
  assign new_n29642_ = ~new_n27902_ & ~new_n29641_;
  assign new_n29643_ = ~new_n29604_ & ~new_n29642_;
  assign new_n29644_ = new_n27955_ & ~new_n29643_;
  assign new_n29645_ = ys__n45592 & new_n13490_;
  assign new_n29646_ = ys__n45428 & new_n13382_;
  assign new_n29647_ = ~new_n29645_ & ~new_n29646_;
  assign new_n29648_ = ys__n45264 & new_n13379_;
  assign new_n29649_ = ys__n45065 & new_n13380_;
  assign new_n29650_ = ~new_n29648_ & ~new_n29649_;
  assign new_n29651_ = new_n29647_ & new_n29650_;
  assign new_n29652_ = new_n27941_ & ~new_n29651_;
  assign new_n29653_ = ys__n45686 & new_n13490_;
  assign new_n29654_ = ys__n45522 & new_n13382_;
  assign new_n29655_ = ~new_n29653_ & ~new_n29654_;
  assign new_n29656_ = ys__n45358 & new_n13379_;
  assign new_n29657_ = ys__n45191 & new_n13380_;
  assign new_n29658_ = ~new_n29656_ & ~new_n29657_;
  assign new_n29659_ = new_n29655_ & new_n29658_;
  assign new_n29660_ = new_n27913_ & ~new_n29659_;
  assign new_n29661_ = ys__n45628 & new_n13490_;
  assign new_n29662_ = ys__n45464 & new_n13382_;
  assign new_n29663_ = ~new_n29661_ & ~new_n29662_;
  assign new_n29664_ = ys__n45300 & new_n13379_;
  assign new_n29665_ = ys__n45106 & new_n13380_;
  assign new_n29666_ = ~new_n29664_ & ~new_n29665_;
  assign new_n29667_ = new_n29663_ & new_n29666_;
  assign new_n29668_ = new_n27922_ & ~new_n29667_;
  assign new_n29669_ = ~new_n29660_ & ~new_n29668_;
  assign new_n29670_ = ~new_n29652_ & new_n29669_;
  assign new_n29671_ = new_n27992_ & ~new_n29670_;
  assign new_n29672_ = new_n13420_ & ~new_n29671_;
  assign new_n29673_ = ~new_n27955_ & ~new_n29672_;
  assign new_n29674_ = ~new_n29644_ & ~new_n29673_;
  assign new_n29675_ = new_n27996_ & ~new_n29674_;
  assign new_n29676_ = ys__n46121 & new_n13490_;
  assign new_n29677_ = ys__n46023 & new_n13382_;
  assign new_n29678_ = ~new_n29676_ & ~new_n29677_;
  assign new_n29679_ = ys__n45925 & new_n13379_;
  assign new_n29680_ = ys__n45829 & new_n13380_;
  assign new_n29681_ = ~new_n29679_ & ~new_n29680_;
  assign new_n29682_ = new_n29678_ & new_n29681_;
  assign new_n29683_ = new_n27922_ & ~new_n29682_;
  assign new_n29684_ = ys__n46084 & new_n13490_;
  assign new_n29685_ = ys__n45986 & new_n13382_;
  assign new_n29686_ = ~new_n29684_ & ~new_n29685_;
  assign new_n29687_ = ys__n45888 & new_n13379_;
  assign new_n29688_ = ys__n45787 & new_n13380_;
  assign new_n29689_ = ~new_n29687_ & ~new_n29688_;
  assign new_n29690_ = new_n29686_ & new_n29689_;
  assign new_n29691_ = new_n27941_ & ~new_n29690_;
  assign new_n29692_ = ~new_n29683_ & ~new_n29691_;
  assign new_n29693_ = new_n28016_ & ~new_n29692_;
  assign new_n29694_ = new_n13529_ & ~new_n29693_;
  assign new_n29695_ = ~new_n27996_ & ~new_n29694_;
  assign ys__n26137 = new_n29675_ | new_n29695_;
  assign new_n29697_ = ys__n26062 & new_n27902_;
  assign new_n29698_ = ys__n46384 & new_n13490_;
  assign new_n29699_ = ys__n46560 & new_n13382_;
  assign new_n29700_ = ~new_n29698_ & ~new_n29699_;
  assign new_n29701_ = ys__n46736 & new_n13379_;
  assign new_n29702_ = ys__n46912 & new_n13380_;
  assign new_n29703_ = ~new_n29701_ & ~new_n29702_;
  assign new_n29704_ = new_n29700_ & new_n29703_;
  assign new_n29705_ = new_n27913_ & ~new_n29704_;
  assign new_n29706_ = ys__n46306 & new_n13490_;
  assign new_n29707_ = ys__n46482 & new_n13382_;
  assign new_n29708_ = ~new_n29706_ & ~new_n29707_;
  assign new_n29709_ = ys__n46658 & new_n13379_;
  assign new_n29710_ = ys__n46834 & new_n13380_;
  assign new_n29711_ = ~new_n29709_ & ~new_n29710_;
  assign new_n29712_ = new_n29708_ & new_n29711_;
  assign new_n29713_ = new_n27922_ & ~new_n29712_;
  assign new_n29714_ = ~new_n29705_ & ~new_n29713_;
  assign new_n29715_ = ys__n46342 & new_n13490_;
  assign new_n29716_ = ys__n46518 & new_n13382_;
  assign new_n29717_ = ~new_n29715_ & ~new_n29716_;
  assign new_n29718_ = ys__n46694 & new_n13379_;
  assign new_n29719_ = ys__n46870 & new_n13380_;
  assign new_n29720_ = ~new_n29718_ & ~new_n29719_;
  assign new_n29721_ = new_n29717_ & new_n29720_;
  assign new_n29722_ = new_n27932_ & ~new_n29721_;
  assign new_n29723_ = ys__n46419 & new_n13490_;
  assign new_n29724_ = ys__n46595 & new_n13382_;
  assign new_n29725_ = ~new_n29723_ & ~new_n29724_;
  assign new_n29726_ = ys__n46771 & new_n13379_;
  assign new_n29727_ = ys__n46947 & new_n13380_;
  assign new_n29728_ = ~new_n29726_ & ~new_n29727_;
  assign new_n29729_ = new_n29725_ & new_n29728_;
  assign new_n29730_ = new_n27941_ & ~new_n29729_;
  assign new_n29731_ = ~new_n29722_ & ~new_n29730_;
  assign new_n29732_ = new_n29714_ & new_n29731_;
  assign new_n29733_ = new_n27952_ & ~new_n29732_;
  assign new_n29734_ = ~new_n29697_ & ~new_n29733_;
  assign new_n29735_ = new_n27955_ & ~new_n29734_;
  assign new_n29736_ = ys__n45594 & new_n13490_;
  assign new_n29737_ = ys__n45430 & new_n13382_;
  assign new_n29738_ = ~new_n29736_ & ~new_n29737_;
  assign new_n29739_ = ys__n45266 & new_n13379_;
  assign new_n29740_ = ys__n45068 & new_n13380_;
  assign new_n29741_ = ~new_n29739_ & ~new_n29740_;
  assign new_n29742_ = new_n29738_ & new_n29741_;
  assign new_n29743_ = new_n27941_ & ~new_n29742_;
  assign new_n29744_ = ys__n45688 & new_n13490_;
  assign new_n29745_ = ys__n45524 & new_n13382_;
  assign new_n29746_ = ~new_n29744_ & ~new_n29745_;
  assign new_n29747_ = ys__n45360 & new_n13379_;
  assign new_n29748_ = ys__n45194 & new_n13380_;
  assign new_n29749_ = ~new_n29747_ & ~new_n29748_;
  assign new_n29750_ = new_n29746_ & new_n29749_;
  assign new_n29751_ = new_n27913_ & ~new_n29750_;
  assign new_n29752_ = ys__n45629 & new_n13490_;
  assign new_n29753_ = ys__n45465 & new_n13382_;
  assign new_n29754_ = ~new_n29752_ & ~new_n29753_;
  assign new_n29755_ = ys__n45301 & new_n13379_;
  assign new_n29756_ = ys__n45107 & new_n13380_;
  assign new_n29757_ = ~new_n29755_ & ~new_n29756_;
  assign new_n29758_ = new_n29754_ & new_n29757_;
  assign new_n29759_ = new_n27922_ & ~new_n29758_;
  assign new_n29760_ = ~new_n29751_ & ~new_n29759_;
  assign new_n29761_ = ~new_n29743_ & new_n29760_;
  assign new_n29762_ = new_n27993_ & ~new_n29761_;
  assign new_n29763_ = ~new_n29735_ & ~new_n29762_;
  assign new_n29764_ = new_n27996_ & ~new_n29763_;
  assign new_n29765_ = ys__n46122 & new_n13490_;
  assign new_n29766_ = ys__n46024 & new_n13382_;
  assign new_n29767_ = ~new_n29765_ & ~new_n29766_;
  assign new_n29768_ = ys__n45926 & new_n13379_;
  assign new_n29769_ = ys__n45830 & new_n13380_;
  assign new_n29770_ = ~new_n29768_ & ~new_n29769_;
  assign new_n29771_ = new_n29767_ & new_n29770_;
  assign new_n29772_ = new_n27922_ & ~new_n29771_;
  assign new_n29773_ = ys__n46086 & new_n13490_;
  assign new_n29774_ = ys__n45988 & new_n13382_;
  assign new_n29775_ = ~new_n29773_ & ~new_n29774_;
  assign new_n29776_ = ys__n45890 & new_n13379_;
  assign new_n29777_ = ys__n45790 & new_n13380_;
  assign new_n29778_ = ~new_n29776_ & ~new_n29777_;
  assign new_n29779_ = new_n29775_ & new_n29778_;
  assign new_n29780_ = new_n27941_ & ~new_n29779_;
  assign new_n29781_ = ~new_n29772_ & ~new_n29780_;
  assign new_n29782_ = new_n28016_ & ~new_n29781_;
  assign new_n29783_ = ~new_n27996_ & new_n29782_;
  assign ys__n26138 = new_n29764_ | new_n29783_;
  assign new_n29785_ = ys__n26065 & new_n27902_;
  assign new_n29786_ = ys__n46386 & new_n13490_;
  assign new_n29787_ = ys__n46562 & new_n13382_;
  assign new_n29788_ = ~new_n29786_ & ~new_n29787_;
  assign new_n29789_ = ys__n46738 & new_n13379_;
  assign new_n29790_ = ys__n46914 & new_n13380_;
  assign new_n29791_ = ~new_n29789_ & ~new_n29790_;
  assign new_n29792_ = new_n29788_ & new_n29791_;
  assign new_n29793_ = new_n27913_ & ~new_n29792_;
  assign new_n29794_ = ys__n46308 & new_n13490_;
  assign new_n29795_ = ys__n46484 & new_n13382_;
  assign new_n29796_ = ~new_n29794_ & ~new_n29795_;
  assign new_n29797_ = ys__n46660 & new_n13379_;
  assign new_n29798_ = ys__n46836 & new_n13380_;
  assign new_n29799_ = ~new_n29797_ & ~new_n29798_;
  assign new_n29800_ = new_n29796_ & new_n29799_;
  assign new_n29801_ = new_n27922_ & ~new_n29800_;
  assign new_n29802_ = ~new_n29793_ & ~new_n29801_;
  assign new_n29803_ = ys__n46343 & new_n13490_;
  assign new_n29804_ = ys__n46519 & new_n13382_;
  assign new_n29805_ = ~new_n29803_ & ~new_n29804_;
  assign new_n29806_ = ys__n46695 & new_n13379_;
  assign new_n29807_ = ys__n46871 & new_n13380_;
  assign new_n29808_ = ~new_n29806_ & ~new_n29807_;
  assign new_n29809_ = new_n29805_ & new_n29808_;
  assign new_n29810_ = new_n27932_ & ~new_n29809_;
  assign new_n29811_ = ys__n46420 & new_n13490_;
  assign new_n29812_ = ys__n46596 & new_n13382_;
  assign new_n29813_ = ~new_n29811_ & ~new_n29812_;
  assign new_n29814_ = ys__n46772 & new_n13379_;
  assign new_n29815_ = ys__n46948 & new_n13380_;
  assign new_n29816_ = ~new_n29814_ & ~new_n29815_;
  assign new_n29817_ = new_n29813_ & new_n29816_;
  assign new_n29818_ = new_n27941_ & ~new_n29817_;
  assign new_n29819_ = ~new_n29810_ & ~new_n29818_;
  assign new_n29820_ = new_n29802_ & new_n29819_;
  assign new_n29821_ = new_n27952_ & ~new_n29820_;
  assign new_n29822_ = ~new_n29785_ & ~new_n29821_;
  assign new_n29823_ = new_n27955_ & ~new_n29822_;
  assign new_n29824_ = ys__n45596 & new_n13490_;
  assign new_n29825_ = ys__n45432 & new_n13382_;
  assign new_n29826_ = ~new_n29824_ & ~new_n29825_;
  assign new_n29827_ = ys__n45268 & new_n13379_;
  assign new_n29828_ = ys__n45071 & new_n13380_;
  assign new_n29829_ = ~new_n29827_ & ~new_n29828_;
  assign new_n29830_ = new_n29826_ & new_n29829_;
  assign new_n29831_ = new_n27941_ & ~new_n29830_;
  assign new_n29832_ = ys__n45690 & new_n13490_;
  assign new_n29833_ = ys__n45526 & new_n13382_;
  assign new_n29834_ = ~new_n29832_ & ~new_n29833_;
  assign new_n29835_ = ys__n45362 & new_n13379_;
  assign new_n29836_ = ys__n45197 & new_n13380_;
  assign new_n29837_ = ~new_n29835_ & ~new_n29836_;
  assign new_n29838_ = new_n29834_ & new_n29837_;
  assign new_n29839_ = new_n27913_ & ~new_n29838_;
  assign new_n29840_ = ys__n45630 & new_n13490_;
  assign new_n29841_ = ys__n45466 & new_n13382_;
  assign new_n29842_ = ~new_n29840_ & ~new_n29841_;
  assign new_n29843_ = ys__n45302 & new_n13379_;
  assign new_n29844_ = ys__n45108 & new_n13380_;
  assign new_n29845_ = ~new_n29843_ & ~new_n29844_;
  assign new_n29846_ = new_n29842_ & new_n29845_;
  assign new_n29847_ = new_n27922_ & ~new_n29846_;
  assign new_n29848_ = ~new_n29839_ & ~new_n29847_;
  assign new_n29849_ = ~new_n29831_ & new_n29848_;
  assign new_n29850_ = new_n27993_ & ~new_n29849_;
  assign new_n29851_ = ~new_n29823_ & ~new_n29850_;
  assign new_n29852_ = new_n27996_ & ~new_n29851_;
  assign new_n29853_ = ys__n46123 & new_n13490_;
  assign new_n29854_ = ys__n46025 & new_n13382_;
  assign new_n29855_ = ~new_n29853_ & ~new_n29854_;
  assign new_n29856_ = ys__n45927 & new_n13379_;
  assign new_n29857_ = ys__n45831 & new_n13380_;
  assign new_n29858_ = ~new_n29856_ & ~new_n29857_;
  assign new_n29859_ = new_n29855_ & new_n29858_;
  assign new_n29860_ = new_n27922_ & ~new_n29859_;
  assign new_n29861_ = ys__n46088 & new_n13490_;
  assign new_n29862_ = ys__n45990 & new_n13382_;
  assign new_n29863_ = ~new_n29861_ & ~new_n29862_;
  assign new_n29864_ = ys__n45892 & new_n13379_;
  assign new_n29865_ = ys__n45793 & new_n13380_;
  assign new_n29866_ = ~new_n29864_ & ~new_n29865_;
  assign new_n29867_ = new_n29863_ & new_n29866_;
  assign new_n29868_ = new_n27941_ & ~new_n29867_;
  assign new_n29869_ = ~new_n29860_ & ~new_n29868_;
  assign new_n29870_ = new_n28016_ & ~new_n29869_;
  assign new_n29871_ = ~new_n27996_ & new_n29870_;
  assign ys__n26139 = new_n29852_ | new_n29871_;
  assign new_n29873_ = ys__n26071 & new_n27902_;
  assign new_n29874_ = ys__n46390 & new_n13490_;
  assign new_n29875_ = ys__n46566 & new_n13382_;
  assign new_n29876_ = ~new_n29874_ & ~new_n29875_;
  assign new_n29877_ = ys__n46742 & new_n13379_;
  assign new_n29878_ = ys__n46918 & new_n13380_;
  assign new_n29879_ = ~new_n29877_ & ~new_n29878_;
  assign new_n29880_ = new_n29876_ & new_n29879_;
  assign new_n29881_ = new_n27913_ & ~new_n29880_;
  assign new_n29882_ = ys__n46312 & new_n13490_;
  assign new_n29883_ = ys__n46488 & new_n13382_;
  assign new_n29884_ = ~new_n29882_ & ~new_n29883_;
  assign new_n29885_ = ys__n46664 & new_n13379_;
  assign new_n29886_ = ys__n46840 & new_n13380_;
  assign new_n29887_ = ~new_n29885_ & ~new_n29886_;
  assign new_n29888_ = new_n29884_ & new_n29887_;
  assign new_n29889_ = new_n27922_ & ~new_n29888_;
  assign new_n29890_ = ~new_n29881_ & ~new_n29889_;
  assign new_n29891_ = ys__n46345 & new_n13490_;
  assign new_n29892_ = ys__n46521 & new_n13382_;
  assign new_n29893_ = ~new_n29891_ & ~new_n29892_;
  assign new_n29894_ = ys__n46697 & new_n13379_;
  assign new_n29895_ = ys__n46873 & new_n13380_;
  assign new_n29896_ = ~new_n29894_ & ~new_n29895_;
  assign new_n29897_ = new_n29893_ & new_n29896_;
  assign new_n29898_ = new_n27932_ & ~new_n29897_;
  assign new_n29899_ = ys__n46422 & new_n13490_;
  assign new_n29900_ = ys__n46598 & new_n13382_;
  assign new_n29901_ = ~new_n29899_ & ~new_n29900_;
  assign new_n29902_ = ys__n46774 & new_n13379_;
  assign new_n29903_ = ys__n46950 & new_n13380_;
  assign new_n29904_ = ~new_n29902_ & ~new_n29903_;
  assign new_n29905_ = new_n29901_ & new_n29904_;
  assign new_n29906_ = new_n27941_ & ~new_n29905_;
  assign new_n29907_ = ~new_n29898_ & ~new_n29906_;
  assign new_n29908_ = new_n29890_ & new_n29907_;
  assign new_n29909_ = new_n27952_ & ~new_n29908_;
  assign new_n29910_ = ~new_n29873_ & ~new_n29909_;
  assign new_n29911_ = new_n27955_ & ~new_n29910_;
  assign new_n29912_ = ys__n45600 & new_n13490_;
  assign new_n29913_ = ys__n45436 & new_n13382_;
  assign new_n29914_ = ~new_n29912_ & ~new_n29913_;
  assign new_n29915_ = ys__n45272 & new_n13379_;
  assign new_n29916_ = ys__n45077 & new_n13380_;
  assign new_n29917_ = ~new_n29915_ & ~new_n29916_;
  assign new_n29918_ = new_n29914_ & new_n29917_;
  assign new_n29919_ = new_n27941_ & ~new_n29918_;
  assign new_n29920_ = ys__n45694 & new_n13490_;
  assign new_n29921_ = ys__n45530 & new_n13382_;
  assign new_n29922_ = ~new_n29920_ & ~new_n29921_;
  assign new_n29923_ = ys__n45366 & new_n13379_;
  assign new_n29924_ = ys__n45203 & new_n13380_;
  assign new_n29925_ = ~new_n29923_ & ~new_n29924_;
  assign new_n29926_ = new_n29922_ & new_n29925_;
  assign new_n29927_ = new_n27913_ & ~new_n29926_;
  assign new_n29928_ = ys__n45632 & new_n13490_;
  assign new_n29929_ = ys__n45468 & new_n13382_;
  assign new_n29930_ = ~new_n29928_ & ~new_n29929_;
  assign new_n29931_ = ys__n45304 & new_n13379_;
  assign new_n29932_ = ys__n45110 & new_n13380_;
  assign new_n29933_ = ~new_n29931_ & ~new_n29932_;
  assign new_n29934_ = new_n29930_ & new_n29933_;
  assign new_n29935_ = new_n27922_ & ~new_n29934_;
  assign new_n29936_ = ~new_n29927_ & ~new_n29935_;
  assign new_n29937_ = ~new_n29919_ & new_n29936_;
  assign new_n29938_ = new_n27993_ & ~new_n29937_;
  assign new_n29939_ = ~new_n29911_ & ~new_n29938_;
  assign new_n29940_ = new_n27996_ & ~new_n29939_;
  assign new_n29941_ = ys__n46125 & new_n13490_;
  assign new_n29942_ = ys__n46027 & new_n13382_;
  assign new_n29943_ = ~new_n29941_ & ~new_n29942_;
  assign new_n29944_ = ys__n45929 & new_n13379_;
  assign new_n29945_ = ys__n45833 & new_n13380_;
  assign new_n29946_ = ~new_n29944_ & ~new_n29945_;
  assign new_n29947_ = new_n29943_ & new_n29946_;
  assign new_n29948_ = new_n27922_ & ~new_n29947_;
  assign new_n29949_ = ys__n46092 & new_n13490_;
  assign new_n29950_ = ys__n45994 & new_n13382_;
  assign new_n29951_ = ~new_n29949_ & ~new_n29950_;
  assign new_n29952_ = ys__n45896 & new_n13379_;
  assign new_n29953_ = ys__n45799 & new_n13380_;
  assign new_n29954_ = ~new_n29952_ & ~new_n29953_;
  assign new_n29955_ = new_n29951_ & new_n29954_;
  assign new_n29956_ = new_n27941_ & ~new_n29955_;
  assign new_n29957_ = ~new_n29948_ & ~new_n29956_;
  assign new_n29958_ = new_n28016_ & ~new_n29957_;
  assign new_n29959_ = ~new_n27996_ & new_n29958_;
  assign ys__n26141 = new_n29940_ | new_n29959_;
  assign new_n29961_ = ys__n25980 & new_n27902_;
  assign new_n29962_ = ys__n26766 & ~new_n13499_;
  assign new_n29963_ = ys__n46315 & new_n13490_;
  assign new_n29964_ = ys__n46491 & new_n13382_;
  assign new_n29965_ = ~new_n29963_ & ~new_n29964_;
  assign new_n29966_ = ys__n46667 & new_n13379_;
  assign new_n29967_ = ys__n46843 & new_n13380_;
  assign new_n29968_ = ~new_n29966_ & ~new_n29967_;
  assign new_n29969_ = new_n29965_ & new_n29968_;
  assign new_n29970_ = new_n27932_ & ~new_n29969_;
  assign new_n29971_ = ys__n27518 & new_n13490_;
  assign new_n29972_ = ys__n27507 & new_n13382_;
  assign new_n29973_ = ~new_n29971_ & ~new_n29972_;
  assign new_n29974_ = ys__n27496 & new_n13379_;
  assign new_n29975_ = ys__n27481 & new_n13380_;
  assign new_n29976_ = ~new_n29974_ & ~new_n29975_;
  assign new_n29977_ = new_n29973_ & new_n29976_;
  assign new_n29978_ = new_n27913_ & ~new_n29977_;
  assign new_n29979_ = ys__n46252 & new_n13490_;
  assign new_n29980_ = ys__n46428 & new_n13382_;
  assign new_n29981_ = ~new_n29979_ & ~new_n29980_;
  assign new_n29982_ = ys__n46604 & new_n13379_;
  assign new_n29983_ = ys__n46780 & new_n13380_;
  assign new_n29984_ = ~new_n29982_ & ~new_n29983_;
  assign new_n29985_ = new_n29981_ & new_n29984_;
  assign new_n29986_ = new_n27922_ & ~new_n29985_;
  assign new_n29987_ = ~new_n29978_ & ~new_n29986_;
  assign new_n29988_ = ~new_n29970_ & new_n29987_;
  assign new_n29989_ = new_n27951_ & ~new_n29988_;
  assign new_n29990_ = ~new_n29962_ & ~new_n29989_;
  assign new_n29991_ = ~new_n27902_ & ~new_n29990_;
  assign new_n29992_ = ~new_n29961_ & ~new_n29991_;
  assign new_n29993_ = new_n27955_ & ~new_n29992_;
  assign new_n29994_ = ys__n25727 & ~new_n13420_;
  assign new_n29995_ = ys__n45634 & new_n13490_;
  assign new_n29996_ = ys__n45470 & new_n13382_;
  assign new_n29997_ = ~new_n29995_ & ~new_n29996_;
  assign new_n29998_ = ys__n45306 & new_n13379_;
  assign new_n29999_ = ys__n45113 & new_n13380_;
  assign new_n30000_ = ~new_n29998_ & ~new_n29999_;
  assign new_n30001_ = new_n29997_ & new_n30000_;
  assign new_n30002_ = new_n27913_ & ~new_n30001_;
  assign new_n30003_ = ys__n45702 & new_n13490_;
  assign new_n30004_ = ys__n45538 & new_n13382_;
  assign new_n30005_ = ~new_n30003_ & ~new_n30004_;
  assign new_n30006_ = ys__n45374 & new_n13379_;
  assign new_n30007_ = ys__n45212 & new_n13380_;
  assign new_n30008_ = ~new_n30006_ & ~new_n30007_;
  assign new_n30009_ = new_n30005_ & new_n30008_;
  assign new_n30010_ = new_n27932_ & ~new_n30009_;
  assign new_n30011_ = ~new_n30002_ & ~new_n30010_;
  assign new_n30012_ = new_n13378_ & ~new_n13384_;
  assign new_n30013_ = new_n27949_ & ~new_n30012_;
  assign new_n30014_ = new_n13420_ & new_n30013_;
  assign new_n30015_ = ~new_n30011_ & new_n30014_;
  assign new_n30016_ = ~new_n29994_ & ~new_n30015_;
  assign new_n30017_ = ~new_n27955_ & ~new_n30016_;
  assign new_n30018_ = ~new_n29993_ & ~new_n30017_;
  assign new_n30019_ = new_n27996_ & ~new_n30018_;
  assign new_n30020_ = ys__n25853 & ~new_n13529_;
  assign new_n30021_ = ys__n46127 & new_n13490_;
  assign new_n30022_ = ys__n46029 & new_n13382_;
  assign new_n30023_ = ~new_n30021_ & ~new_n30022_;
  assign new_n30024_ = ys__n45931 & new_n13379_;
  assign new_n30025_ = ys__n45835 & new_n13380_;
  assign new_n30026_ = ~new_n30024_ & ~new_n30025_;
  assign new_n30027_ = new_n30023_ & new_n30026_;
  assign new_n30028_ = new_n27932_ & new_n27949_;
  assign new_n30029_ = ~new_n30027_ & new_n30028_;
  assign new_n30030_ = new_n13529_ & new_n30029_;
  assign new_n30031_ = ~new_n30020_ & ~new_n30030_;
  assign new_n30032_ = ~new_n27996_ & ~new_n30031_;
  assign new_n30033_ = ~new_n30019_ & ~new_n30032_;
  assign new_n30034_ = ~new_n15156_ & ~new_n30033_;
  assign new_n30035_ = ys__n26143 & new_n15156_;
  assign ys__n26144 = new_n30034_ | new_n30035_;
  assign new_n30037_ = ys__n25984 & new_n27902_;
  assign new_n30038_ = ys__n26768 & ~new_n13499_;
  assign new_n30039_ = ys__n47108 & new_n13490_;
  assign new_n30040_ = ys__n47111 & new_n13382_;
  assign new_n30041_ = ~new_n30039_ & ~new_n30040_;
  assign new_n30042_ = ys__n47114 & new_n13379_;
  assign new_n30043_ = ys__n47117 & new_n13380_;
  assign new_n30044_ = ~new_n30042_ & ~new_n30043_;
  assign new_n30045_ = new_n30041_ & new_n30044_;
  assign new_n30046_ = new_n27913_ & ~new_n30045_;
  assign new_n30047_ = ys__n46254 & new_n13490_;
  assign new_n30048_ = ys__n46430 & new_n13382_;
  assign new_n30049_ = ~new_n30047_ & ~new_n30048_;
  assign new_n30050_ = ys__n46606 & new_n13379_;
  assign new_n30051_ = ys__n46782 & new_n13380_;
  assign new_n30052_ = ~new_n30050_ & ~new_n30051_;
  assign new_n30053_ = new_n30049_ & new_n30052_;
  assign new_n30054_ = new_n27922_ & ~new_n30053_;
  assign new_n30055_ = ~new_n30046_ & ~new_n30054_;
  assign new_n30056_ = ys__n46316 & new_n13490_;
  assign new_n30057_ = ys__n46492 & new_n13382_;
  assign new_n30058_ = ~new_n30056_ & ~new_n30057_;
  assign new_n30059_ = ys__n46668 & new_n13379_;
  assign new_n30060_ = ys__n46844 & new_n13380_;
  assign new_n30061_ = ~new_n30059_ & ~new_n30060_;
  assign new_n30062_ = new_n30058_ & new_n30061_;
  assign new_n30063_ = new_n27932_ & ~new_n30062_;
  assign new_n30064_ = ys__n46393 & new_n13490_;
  assign new_n30065_ = ys__n46569 & new_n13382_;
  assign new_n30066_ = ~new_n30064_ & ~new_n30065_;
  assign new_n30067_ = ys__n46745 & new_n13379_;
  assign new_n30068_ = ys__n46921 & new_n13380_;
  assign new_n30069_ = ~new_n30067_ & ~new_n30068_;
  assign new_n30070_ = new_n30066_ & new_n30069_;
  assign new_n30071_ = new_n27941_ & ~new_n30070_;
  assign new_n30072_ = ~new_n30063_ & ~new_n30071_;
  assign new_n30073_ = new_n30055_ & new_n30072_;
  assign new_n30074_ = new_n27951_ & ~new_n30073_;
  assign new_n30075_ = ~new_n30038_ & ~new_n30074_;
  assign new_n30076_ = ~new_n27902_ & ~new_n30075_;
  assign new_n30077_ = ~new_n30037_ & ~new_n30076_;
  assign new_n30078_ = new_n27955_ & ~new_n30077_;
  assign new_n30079_ = ys__n25730 & ~new_n13420_;
  assign new_n30080_ = new_n27913_ & new_n27949_;
  assign new_n30081_ = ys__n45636 & new_n13490_;
  assign new_n30082_ = ys__n45472 & new_n13382_;
  assign new_n30083_ = ~new_n30081_ & ~new_n30082_;
  assign new_n30084_ = ys__n45308 & new_n13379_;
  assign new_n30085_ = ys__n45116 & new_n13380_;
  assign new_n30086_ = ~new_n30084_ & ~new_n30085_;
  assign new_n30087_ = new_n30083_ & new_n30086_;
  assign new_n30088_ = ~new_n13374_ & new_n13489_;
  assign new_n30089_ = ~new_n30087_ & ~new_n30088_;
  assign new_n30090_ = new_n30080_ & new_n30089_;
  assign new_n30091_ = new_n13420_ & new_n30090_;
  assign new_n30092_ = ~new_n30079_ & ~new_n30091_;
  assign new_n30093_ = ~new_n27955_ & ~new_n30092_;
  assign new_n30094_ = ~new_n30078_ & ~new_n30093_;
  assign new_n30095_ = new_n27996_ & ~new_n30094_;
  assign new_n30096_ = ys__n25856 & ~new_n13529_;
  assign new_n30097_ = ys__n46096 & new_n13490_;
  assign new_n30098_ = ys__n45998 & new_n13382_;
  assign new_n30099_ = ~new_n30097_ & ~new_n30098_;
  assign new_n30100_ = ys__n45900 & new_n13379_;
  assign new_n30101_ = ys__n45804 & new_n13380_;
  assign new_n30102_ = ~new_n30100_ & ~new_n30101_;
  assign new_n30103_ = new_n30099_ & new_n30102_;
  assign new_n30104_ = new_n27922_ & ~new_n30103_;
  assign new_n30105_ = ys__n46034 & new_n13490_;
  assign new_n30106_ = ys__n45936 & new_n13382_;
  assign new_n30107_ = ~new_n30105_ & ~new_n30106_;
  assign new_n30108_ = ys__n45838 & new_n13379_;
  assign new_n30109_ = ys__n45712 & new_n13380_;
  assign new_n30110_ = ~new_n30108_ & ~new_n30109_;
  assign new_n30111_ = new_n30107_ & new_n30110_;
  assign new_n30112_ = new_n27941_ & ~new_n30111_;
  assign new_n30113_ = ~new_n30104_ & ~new_n30112_;
  assign new_n30114_ = new_n28016_ & ~new_n30113_;
  assign new_n30115_ = ~new_n30096_ & ~new_n30114_;
  assign new_n30116_ = ~new_n27996_ & ~new_n30115_;
  assign new_n30117_ = ~new_n30095_ & ~new_n30116_;
  assign new_n30118_ = ~new_n15156_ & ~new_n30117_;
  assign new_n30119_ = ys__n26145 & new_n15156_;
  assign ys__n26146 = new_n30118_ | new_n30119_;
  assign new_n30121_ = ys__n25987 & new_n27902_;
  assign new_n30122_ = ys__n26770 & ~new_n13499_;
  assign new_n30123_ = ys__n27520 & new_n13490_;
  assign new_n30124_ = ys__n27509 & new_n13382_;
  assign new_n30125_ = ~new_n30123_ & ~new_n30124_;
  assign new_n30126_ = ys__n27498 & new_n13379_;
  assign new_n30127_ = ys__n27485 & new_n13380_;
  assign new_n30128_ = ~new_n30126_ & ~new_n30127_;
  assign new_n30129_ = new_n30125_ & new_n30128_;
  assign new_n30130_ = new_n27913_ & ~new_n30129_;
  assign new_n30131_ = ys__n46256 & new_n13490_;
  assign new_n30132_ = ys__n46432 & new_n13382_;
  assign new_n30133_ = ~new_n30131_ & ~new_n30132_;
  assign new_n30134_ = ys__n46608 & new_n13379_;
  assign new_n30135_ = ys__n46784 & new_n13380_;
  assign new_n30136_ = ~new_n30134_ & ~new_n30135_;
  assign new_n30137_ = new_n30133_ & new_n30136_;
  assign new_n30138_ = new_n27922_ & ~new_n30137_;
  assign new_n30139_ = ~new_n30130_ & ~new_n30138_;
  assign new_n30140_ = ys__n46317 & new_n13490_;
  assign new_n30141_ = ys__n46493 & new_n13382_;
  assign new_n30142_ = ~new_n30140_ & ~new_n30141_;
  assign new_n30143_ = ys__n46669 & new_n13379_;
  assign new_n30144_ = ys__n46845 & new_n13380_;
  assign new_n30145_ = ~new_n30143_ & ~new_n30144_;
  assign new_n30146_ = new_n30142_ & new_n30145_;
  assign new_n30147_ = new_n27932_ & ~new_n30146_;
  assign new_n30148_ = ys__n46394 & new_n13490_;
  assign new_n30149_ = ys__n46570 & new_n13382_;
  assign new_n30150_ = ~new_n30148_ & ~new_n30149_;
  assign new_n30151_ = ys__n46746 & new_n13379_;
  assign new_n30152_ = ys__n46922 & new_n13380_;
  assign new_n30153_ = ~new_n30151_ & ~new_n30152_;
  assign new_n30154_ = new_n30150_ & new_n30153_;
  assign new_n30155_ = new_n27941_ & ~new_n30154_;
  assign new_n30156_ = ~new_n30147_ & ~new_n30155_;
  assign new_n30157_ = new_n30139_ & new_n30156_;
  assign new_n30158_ = new_n27951_ & ~new_n30157_;
  assign new_n30159_ = ~new_n30122_ & ~new_n30158_;
  assign new_n30160_ = ~new_n27902_ & ~new_n30159_;
  assign new_n30161_ = ~new_n30121_ & ~new_n30160_;
  assign new_n30162_ = new_n27955_ & ~new_n30161_;
  assign new_n30163_ = ys__n25733 & ~new_n13420_;
  assign new_n30164_ = ys__n45638 & new_n13490_;
  assign new_n30165_ = ys__n45474 & new_n13382_;
  assign new_n30166_ = ~new_n30164_ & ~new_n30165_;
  assign new_n30167_ = ys__n45310 & new_n13379_;
  assign new_n30168_ = ys__n45119 & new_n13380_;
  assign new_n30169_ = ~new_n30167_ & ~new_n30168_;
  assign new_n30170_ = new_n30166_ & new_n30169_;
  assign new_n30171_ = new_n27913_ & ~new_n30170_;
  assign new_n30172_ = ys__n45604 & new_n13490_;
  assign new_n30173_ = ys__n45440 & new_n13382_;
  assign new_n30174_ = ~new_n30172_ & ~new_n30173_;
  assign new_n30175_ = ys__n45276 & new_n13379_;
  assign new_n30176_ = ys__n45082 & new_n13380_;
  assign new_n30177_ = ~new_n30175_ & ~new_n30176_;
  assign new_n30178_ = new_n30174_ & new_n30177_;
  assign new_n30179_ = new_n27922_ & ~new_n30178_;
  assign new_n30180_ = ~new_n30171_ & ~new_n30179_;
  assign new_n30181_ = ys__n45704 & new_n13490_;
  assign new_n30182_ = ys__n45541 & new_n13382_;
  assign new_n30183_ = ~new_n30181_ & ~new_n30182_;
  assign new_n30184_ = ys__n45377 & new_n13379_;
  assign new_n30185_ = ys__n45214 & new_n13380_;
  assign new_n30186_ = ~new_n30184_ & ~new_n30185_;
  assign new_n30187_ = new_n30183_ & new_n30186_;
  assign new_n30188_ = new_n27932_ & ~new_n30187_;
  assign new_n30189_ = ys__n45544 & new_n13490_;
  assign new_n30190_ = ys__n45380 & new_n13382_;
  assign new_n30191_ = ~new_n30189_ & ~new_n30190_;
  assign new_n30192_ = ys__n45216 & new_n13379_;
  assign new_n30193_ = ys__n44993 & new_n13380_;
  assign new_n30194_ = ~new_n30192_ & ~new_n30193_;
  assign new_n30195_ = new_n30191_ & new_n30194_;
  assign new_n30196_ = new_n27941_ & ~new_n30195_;
  assign new_n30197_ = ~new_n30188_ & ~new_n30196_;
  assign new_n30198_ = new_n30180_ & new_n30197_;
  assign new_n30199_ = new_n27992_ & ~new_n30198_;
  assign new_n30200_ = ~new_n30163_ & ~new_n30199_;
  assign new_n30201_ = ~new_n27955_ & ~new_n30200_;
  assign new_n30202_ = ~new_n30162_ & ~new_n30201_;
  assign new_n30203_ = new_n27996_ & ~new_n30202_;
  assign new_n30204_ = ys__n25859 & ~new_n13529_;
  assign new_n30205_ = ys__n46036 & new_n13490_;
  assign new_n30206_ = ys__n45938 & new_n13382_;
  assign new_n30207_ = ~new_n30205_ & ~new_n30206_;
  assign new_n30208_ = ys__n45840 & new_n13379_;
  assign new_n30209_ = ys__n45715 & new_n13380_;
  assign new_n30210_ = ~new_n30208_ & ~new_n30209_;
  assign new_n30211_ = new_n30207_ & new_n30210_;
  assign new_n30212_ = new_n27941_ & ~new_n30211_;
  assign new_n30213_ = ys__n46097 & new_n13490_;
  assign new_n30214_ = ys__n45999 & new_n13382_;
  assign new_n30215_ = ~new_n30213_ & ~new_n30214_;
  assign new_n30216_ = ys__n45901 & new_n13379_;
  assign new_n30217_ = ys__n45805 & new_n13380_;
  assign new_n30218_ = ~new_n30216_ & ~new_n30217_;
  assign new_n30219_ = new_n30215_ & new_n30218_;
  assign new_n30220_ = new_n27922_ & ~new_n30219_;
  assign new_n30221_ = ys__n46128 & new_n13490_;
  assign new_n30222_ = ys__n46031 & new_n13382_;
  assign new_n30223_ = ~new_n30221_ & ~new_n30222_;
  assign new_n30224_ = ys__n45933 & new_n13379_;
  assign new_n30225_ = ys__n45836 & new_n13380_;
  assign new_n30226_ = ~new_n30224_ & ~new_n30225_;
  assign new_n30227_ = new_n30223_ & new_n30226_;
  assign new_n30228_ = new_n27932_ & ~new_n30227_;
  assign new_n30229_ = ~new_n30220_ & ~new_n30228_;
  assign new_n30230_ = ~new_n30212_ & new_n30229_;
  assign new_n30231_ = ~new_n13375_ & new_n13511_;
  assign new_n30232_ = new_n27949_ & ~new_n30231_;
  assign new_n30233_ = new_n13529_ & new_n30232_;
  assign new_n30234_ = ~new_n30230_ & new_n30233_;
  assign new_n30235_ = ~new_n30204_ & ~new_n30234_;
  assign new_n30236_ = ~new_n27996_ & ~new_n30235_;
  assign new_n30237_ = ~new_n30203_ & ~new_n30236_;
  assign new_n30238_ = ~new_n15156_ & ~new_n30237_;
  assign new_n30239_ = ys__n26147 & new_n15156_;
  assign ys__n26148 = new_n30238_ | new_n30239_;
  assign new_n30241_ = ys__n25990 & new_n27902_;
  assign new_n30242_ = ys__n26772 & ~new_n13499_;
  assign new_n30243_ = ys__n47109 & new_n13490_;
  assign new_n30244_ = ys__n47112 & new_n13382_;
  assign new_n30245_ = ~new_n30243_ & ~new_n30244_;
  assign new_n30246_ = ys__n47115 & new_n13379_;
  assign new_n30247_ = ys__n47118 & new_n13380_;
  assign new_n30248_ = ~new_n30246_ & ~new_n30247_;
  assign new_n30249_ = new_n30245_ & new_n30248_;
  assign new_n30250_ = new_n27913_ & ~new_n30249_;
  assign new_n30251_ = ys__n46258 & new_n13490_;
  assign new_n30252_ = ys__n46434 & new_n13382_;
  assign new_n30253_ = ~new_n30251_ & ~new_n30252_;
  assign new_n30254_ = ys__n46610 & new_n13379_;
  assign new_n30255_ = ys__n46786 & new_n13380_;
  assign new_n30256_ = ~new_n30254_ & ~new_n30255_;
  assign new_n30257_ = new_n30253_ & new_n30256_;
  assign new_n30258_ = new_n27922_ & ~new_n30257_;
  assign new_n30259_ = ~new_n30250_ & ~new_n30258_;
  assign new_n30260_ = ys__n46318 & new_n13490_;
  assign new_n30261_ = ys__n46494 & new_n13382_;
  assign new_n30262_ = ~new_n30260_ & ~new_n30261_;
  assign new_n30263_ = ys__n46670 & new_n13379_;
  assign new_n30264_ = ys__n46846 & new_n13380_;
  assign new_n30265_ = ~new_n30263_ & ~new_n30264_;
  assign new_n30266_ = new_n30262_ & new_n30265_;
  assign new_n30267_ = new_n27932_ & ~new_n30266_;
  assign new_n30268_ = ys__n46395 & new_n13490_;
  assign new_n30269_ = ys__n46571 & new_n13382_;
  assign new_n30270_ = ~new_n30268_ & ~new_n30269_;
  assign new_n30271_ = ys__n46747 & new_n13379_;
  assign new_n30272_ = ys__n46923 & new_n13380_;
  assign new_n30273_ = ~new_n30271_ & ~new_n30272_;
  assign new_n30274_ = new_n30270_ & new_n30273_;
  assign new_n30275_ = new_n27941_ & ~new_n30274_;
  assign new_n30276_ = ~new_n30267_ & ~new_n30275_;
  assign new_n30277_ = new_n30259_ & new_n30276_;
  assign new_n30278_ = new_n27951_ & ~new_n30277_;
  assign new_n30279_ = ~new_n30242_ & ~new_n30278_;
  assign new_n30280_ = ~new_n27902_ & ~new_n30279_;
  assign new_n30281_ = ~new_n30241_ & ~new_n30280_;
  assign new_n30282_ = new_n27955_ & ~new_n30281_;
  assign new_n30283_ = ys__n25736 & ~new_n13420_;
  assign new_n30284_ = ys__n45546 & new_n13490_;
  assign new_n30285_ = ys__n45382 & new_n13382_;
  assign new_n30286_ = ~new_n30284_ & ~new_n30285_;
  assign new_n30287_ = ys__n45218 & new_n13379_;
  assign new_n30288_ = ys__n44996 & new_n13380_;
  assign new_n30289_ = ~new_n30287_ & ~new_n30288_;
  assign new_n30290_ = new_n30286_ & new_n30289_;
  assign new_n30291_ = new_n27941_ & ~new_n30290_;
  assign new_n30292_ = ys__n45640 & new_n13490_;
  assign new_n30293_ = ys__n45476 & new_n13382_;
  assign new_n30294_ = ~new_n30292_ & ~new_n30293_;
  assign new_n30295_ = ys__n45312 & new_n13379_;
  assign new_n30296_ = ys__n45122 & new_n13380_;
  assign new_n30297_ = ~new_n30295_ & ~new_n30296_;
  assign new_n30298_ = new_n30294_ & new_n30297_;
  assign new_n30299_ = new_n27913_ & ~new_n30298_;
  assign new_n30300_ = ys__n45605 & new_n13490_;
  assign new_n30301_ = ys__n45441 & new_n13382_;
  assign new_n30302_ = ~new_n30300_ & ~new_n30301_;
  assign new_n30303_ = ys__n45277 & new_n13379_;
  assign new_n30304_ = ys__n45083 & new_n13380_;
  assign new_n30305_ = ~new_n30303_ & ~new_n30304_;
  assign new_n30306_ = new_n30302_ & new_n30305_;
  assign new_n30307_ = new_n27922_ & ~new_n30306_;
  assign new_n30308_ = ~new_n30299_ & ~new_n30307_;
  assign new_n30309_ = ~new_n30291_ & new_n30308_;
  assign new_n30310_ = new_n27992_ & ~new_n30309_;
  assign new_n30311_ = ~new_n30283_ & ~new_n30310_;
  assign new_n30312_ = ~new_n27955_ & ~new_n30311_;
  assign new_n30313_ = ~new_n30282_ & ~new_n30312_;
  assign new_n30314_ = new_n27996_ & ~new_n30313_;
  assign new_n30315_ = ys__n25862 & ~new_n13529_;
  assign new_n30316_ = ys__n46098 & new_n13490_;
  assign new_n30317_ = ys__n46000 & new_n13382_;
  assign new_n30318_ = ~new_n30316_ & ~new_n30317_;
  assign new_n30319_ = ys__n45902 & new_n13379_;
  assign new_n30320_ = ys__n45806 & new_n13380_;
  assign new_n30321_ = ~new_n30319_ & ~new_n30320_;
  assign new_n30322_ = new_n30318_ & new_n30321_;
  assign new_n30323_ = new_n27922_ & ~new_n30322_;
  assign new_n30324_ = ys__n46038 & new_n13490_;
  assign new_n30325_ = ys__n45940 & new_n13382_;
  assign new_n30326_ = ~new_n30324_ & ~new_n30325_;
  assign new_n30327_ = ys__n45842 & new_n13379_;
  assign new_n30328_ = ys__n45718 & new_n13380_;
  assign new_n30329_ = ~new_n30327_ & ~new_n30328_;
  assign new_n30330_ = new_n30326_ & new_n30329_;
  assign new_n30331_ = new_n27941_ & ~new_n30330_;
  assign new_n30332_ = ~new_n30323_ & ~new_n30331_;
  assign new_n30333_ = new_n28016_ & ~new_n30332_;
  assign new_n30334_ = ~new_n30315_ & ~new_n30333_;
  assign new_n30335_ = ~new_n27996_ & ~new_n30334_;
  assign new_n30336_ = ~new_n30314_ & ~new_n30335_;
  assign new_n30337_ = ~new_n15156_ & ~new_n30336_;
  assign new_n30338_ = ys__n26149 & new_n15156_;
  assign ys__n26150 = new_n30337_ | new_n30338_;
  assign new_n30340_ = ys__n25993 & new_n27902_;
  assign new_n30341_ = ys__n27510 & new_n13490_;
  assign new_n30342_ = ys__n27499 & new_n13382_;
  assign new_n30343_ = ~new_n30341_ & ~new_n30342_;
  assign new_n30344_ = ys__n27488 & new_n13379_;
  assign new_n30345_ = ys__n27479 & new_n13380_;
  assign new_n30346_ = ~new_n30344_ & ~new_n30345_;
  assign new_n30347_ = new_n30343_ & new_n30346_;
  assign new_n30348_ = new_n27913_ & ~new_n30347_;
  assign new_n30349_ = ys__n46260 & new_n13490_;
  assign new_n30350_ = ys__n46436 & new_n13382_;
  assign new_n30351_ = ~new_n30349_ & ~new_n30350_;
  assign new_n30352_ = ys__n46612 & new_n13379_;
  assign new_n30353_ = ys__n46788 & new_n13380_;
  assign new_n30354_ = ~new_n30352_ & ~new_n30353_;
  assign new_n30355_ = new_n30351_ & new_n30354_;
  assign new_n30356_ = new_n27922_ & ~new_n30355_;
  assign new_n30357_ = ~new_n30348_ & ~new_n30356_;
  assign new_n30358_ = ys__n46319 & new_n13490_;
  assign new_n30359_ = ys__n46495 & new_n13382_;
  assign new_n30360_ = ~new_n30358_ & ~new_n30359_;
  assign new_n30361_ = ys__n46671 & new_n13379_;
  assign new_n30362_ = ys__n46847 & new_n13380_;
  assign new_n30363_ = ~new_n30361_ & ~new_n30362_;
  assign new_n30364_ = new_n30360_ & new_n30363_;
  assign new_n30365_ = new_n27932_ & ~new_n30364_;
  assign new_n30366_ = ys__n46396 & new_n13490_;
  assign new_n30367_ = ys__n46572 & new_n13382_;
  assign new_n30368_ = ~new_n30366_ & ~new_n30367_;
  assign new_n30369_ = ys__n46748 & new_n13379_;
  assign new_n30370_ = ys__n46924 & new_n13380_;
  assign new_n30371_ = ~new_n30369_ & ~new_n30370_;
  assign new_n30372_ = new_n30368_ & new_n30371_;
  assign new_n30373_ = new_n27941_ & ~new_n30372_;
  assign new_n30374_ = ~new_n30365_ & ~new_n30373_;
  assign new_n30375_ = new_n30357_ & new_n30374_;
  assign new_n30376_ = new_n27952_ & ~new_n30375_;
  assign new_n30377_ = ~new_n30340_ & ~new_n30376_;
  assign new_n30378_ = new_n27955_ & ~new_n30377_;
  assign new_n30379_ = ys__n45642 & new_n13490_;
  assign new_n30380_ = ys__n45478 & new_n13382_;
  assign new_n30381_ = ~new_n30379_ & ~new_n30380_;
  assign new_n30382_ = ys__n45314 & new_n13379_;
  assign new_n30383_ = ys__n45125 & new_n13380_;
  assign new_n30384_ = ~new_n30382_ & ~new_n30383_;
  assign new_n30385_ = new_n30381_ & new_n30384_;
  assign new_n30386_ = new_n27913_ & ~new_n30385_;
  assign new_n30387_ = ys__n45606 & new_n13490_;
  assign new_n30388_ = ys__n45442 & new_n13382_;
  assign new_n30389_ = ~new_n30387_ & ~new_n30388_;
  assign new_n30390_ = ys__n45278 & new_n13379_;
  assign new_n30391_ = ys__n45084 & new_n13380_;
  assign new_n30392_ = ~new_n30390_ & ~new_n30391_;
  assign new_n30393_ = new_n30389_ & new_n30392_;
  assign new_n30394_ = new_n27922_ & ~new_n30393_;
  assign new_n30395_ = ~new_n30386_ & ~new_n30394_;
  assign new_n30396_ = ys__n45698 & new_n13490_;
  assign new_n30397_ = ys__n45534 & new_n13382_;
  assign new_n30398_ = ~new_n30396_ & ~new_n30397_;
  assign new_n30399_ = ys__n45370 & new_n13379_;
  assign new_n30400_ = ys__n45208 & new_n13380_;
  assign new_n30401_ = ~new_n30399_ & ~new_n30400_;
  assign new_n30402_ = new_n30398_ & new_n30401_;
  assign new_n30403_ = new_n27932_ & ~new_n30402_;
  assign new_n30404_ = ys__n45548 & new_n13490_;
  assign new_n30405_ = ys__n45384 & new_n13382_;
  assign new_n30406_ = ~new_n30404_ & ~new_n30405_;
  assign new_n30407_ = ys__n45220 & new_n13379_;
  assign new_n30408_ = ys__n44999 & new_n13380_;
  assign new_n30409_ = ~new_n30407_ & ~new_n30408_;
  assign new_n30410_ = new_n30406_ & new_n30409_;
  assign new_n30411_ = new_n27941_ & ~new_n30410_;
  assign new_n30412_ = ~new_n30403_ & ~new_n30411_;
  assign new_n30413_ = new_n30395_ & new_n30412_;
  assign new_n30414_ = new_n27993_ & ~new_n30413_;
  assign new_n30415_ = ~new_n30378_ & ~new_n30414_;
  assign new_n30416_ = new_n27996_ & ~new_n30415_;
  assign new_n30417_ = ys__n46099 & new_n13490_;
  assign new_n30418_ = ys__n46001 & new_n13382_;
  assign new_n30419_ = ~new_n30417_ & ~new_n30418_;
  assign new_n30420_ = ys__n45903 & new_n13379_;
  assign new_n30421_ = ys__n45807 & new_n13380_;
  assign new_n30422_ = ~new_n30420_ & ~new_n30421_;
  assign new_n30423_ = new_n30419_ & new_n30422_;
  assign new_n30424_ = new_n27922_ & ~new_n30423_;
  assign new_n30425_ = ys__n46040 & new_n13490_;
  assign new_n30426_ = ys__n45942 & new_n13382_;
  assign new_n30427_ = ~new_n30425_ & ~new_n30426_;
  assign new_n30428_ = ys__n45844 & new_n13379_;
  assign new_n30429_ = ys__n45721 & new_n13380_;
  assign new_n30430_ = ~new_n30428_ & ~new_n30429_;
  assign new_n30431_ = new_n30427_ & new_n30430_;
  assign new_n30432_ = new_n27941_ & ~new_n30431_;
  assign new_n30433_ = ~new_n30424_ & ~new_n30432_;
  assign new_n30434_ = new_n28016_ & ~new_n30433_;
  assign new_n30435_ = ~new_n27996_ & new_n30434_;
  assign new_n30436_ = ~new_n30416_ & ~new_n30435_;
  assign new_n30437_ = ~new_n15156_ & ~new_n30436_;
  assign new_n30438_ = ys__n26151 & new_n15156_;
  assign ys__n26152 = new_n30437_ | new_n30438_;
  assign new_n30440_ = ys__n25996 & new_n27902_;
  assign new_n30441_ = ys__n18045 & new_n13490_;
  assign new_n30442_ = ys__n18051 & new_n13382_;
  assign new_n30443_ = ~new_n30441_ & ~new_n30442_;
  assign new_n30444_ = ys__n18057 & new_n13379_;
  assign new_n30445_ = ys__n18067 & new_n13380_;
  assign new_n30446_ = ~new_n30444_ & ~new_n30445_;
  assign new_n30447_ = new_n30443_ & new_n30446_;
  assign new_n30448_ = new_n27913_ & ~new_n30447_;
  assign new_n30449_ = ys__n46262 & new_n13490_;
  assign new_n30450_ = ys__n46438 & new_n13382_;
  assign new_n30451_ = ~new_n30449_ & ~new_n30450_;
  assign new_n30452_ = ys__n46614 & new_n13379_;
  assign new_n30453_ = ys__n46790 & new_n13380_;
  assign new_n30454_ = ~new_n30452_ & ~new_n30453_;
  assign new_n30455_ = new_n30451_ & new_n30454_;
  assign new_n30456_ = new_n27922_ & ~new_n30455_;
  assign new_n30457_ = ~new_n30448_ & ~new_n30456_;
  assign new_n30458_ = ys__n46320 & new_n13490_;
  assign new_n30459_ = ys__n46496 & new_n13382_;
  assign new_n30460_ = ~new_n30458_ & ~new_n30459_;
  assign new_n30461_ = ys__n46672 & new_n13379_;
  assign new_n30462_ = ys__n46848 & new_n13380_;
  assign new_n30463_ = ~new_n30461_ & ~new_n30462_;
  assign new_n30464_ = new_n30460_ & new_n30463_;
  assign new_n30465_ = new_n27932_ & ~new_n30464_;
  assign new_n30466_ = ys__n46397 & new_n13490_;
  assign new_n30467_ = ys__n46573 & new_n13382_;
  assign new_n30468_ = ~new_n30466_ & ~new_n30467_;
  assign new_n30469_ = ys__n46749 & new_n13379_;
  assign new_n30470_ = ys__n46925 & new_n13380_;
  assign new_n30471_ = ~new_n30469_ & ~new_n30470_;
  assign new_n30472_ = new_n30468_ & new_n30471_;
  assign new_n30473_ = new_n27941_ & ~new_n30472_;
  assign new_n30474_ = ~new_n30465_ & ~new_n30473_;
  assign new_n30475_ = new_n30457_ & new_n30474_;
  assign new_n30476_ = new_n27952_ & ~new_n30475_;
  assign new_n30477_ = ~new_n30440_ & ~new_n30476_;
  assign new_n30478_ = new_n27955_ & ~new_n30477_;
  assign new_n30479_ = ys__n45644 & new_n13490_;
  assign new_n30480_ = ys__n45480 & new_n13382_;
  assign new_n30481_ = ~new_n30479_ & ~new_n30480_;
  assign new_n30482_ = ys__n45316 & new_n13379_;
  assign new_n30483_ = ys__n45128 & new_n13380_;
  assign new_n30484_ = ~new_n30482_ & ~new_n30483_;
  assign new_n30485_ = new_n30481_ & new_n30484_;
  assign new_n30486_ = new_n27913_ & ~new_n30485_;
  assign new_n30487_ = ys__n45607 & new_n13490_;
  assign new_n30488_ = ys__n45443 & new_n13382_;
  assign new_n30489_ = ~new_n30487_ & ~new_n30488_;
  assign new_n30490_ = ys__n45279 & new_n13379_;
  assign new_n30491_ = ys__n45085 & new_n13380_;
  assign new_n30492_ = ~new_n30490_ & ~new_n30491_;
  assign new_n30493_ = new_n30489_ & new_n30492_;
  assign new_n30494_ = new_n27922_ & ~new_n30493_;
  assign new_n30495_ = ~new_n30486_ & ~new_n30494_;
  assign new_n30496_ = ys__n45699 & new_n13490_;
  assign new_n30497_ = ys__n45535 & new_n13382_;
  assign new_n30498_ = ~new_n30496_ & ~new_n30497_;
  assign new_n30499_ = ys__n45371 & new_n13379_;
  assign new_n30500_ = ys__n45209 & new_n13380_;
  assign new_n30501_ = ~new_n30499_ & ~new_n30500_;
  assign new_n30502_ = new_n30498_ & new_n30501_;
  assign new_n30503_ = new_n27932_ & ~new_n30502_;
  assign new_n30504_ = ys__n45550 & new_n13490_;
  assign new_n30505_ = ys__n45386 & new_n13382_;
  assign new_n30506_ = ~new_n30504_ & ~new_n30505_;
  assign new_n30507_ = ys__n45222 & new_n13379_;
  assign new_n30508_ = ys__n45002 & new_n13380_;
  assign new_n30509_ = ~new_n30507_ & ~new_n30508_;
  assign new_n30510_ = new_n30506_ & new_n30509_;
  assign new_n30511_ = new_n27941_ & ~new_n30510_;
  assign new_n30512_ = ~new_n30503_ & ~new_n30511_;
  assign new_n30513_ = new_n30495_ & new_n30512_;
  assign new_n30514_ = new_n27993_ & ~new_n30513_;
  assign new_n30515_ = ~new_n30478_ & ~new_n30514_;
  assign new_n30516_ = new_n27996_ & ~new_n30515_;
  assign new_n30517_ = ys__n46100 & new_n13490_;
  assign new_n30518_ = ys__n46002 & new_n13382_;
  assign new_n30519_ = ~new_n30517_ & ~new_n30518_;
  assign new_n30520_ = ys__n45904 & new_n13379_;
  assign new_n30521_ = ys__n45808 & new_n13380_;
  assign new_n30522_ = ~new_n30520_ & ~new_n30521_;
  assign new_n30523_ = new_n30519_ & new_n30522_;
  assign new_n30524_ = new_n27922_ & ~new_n30523_;
  assign new_n30525_ = ys__n46042 & new_n13490_;
  assign new_n30526_ = ys__n45944 & new_n13382_;
  assign new_n30527_ = ~new_n30525_ & ~new_n30526_;
  assign new_n30528_ = ys__n45846 & new_n13379_;
  assign new_n30529_ = ys__n45724 & new_n13380_;
  assign new_n30530_ = ~new_n30528_ & ~new_n30529_;
  assign new_n30531_ = new_n30527_ & new_n30530_;
  assign new_n30532_ = new_n27941_ & ~new_n30531_;
  assign new_n30533_ = ~new_n30524_ & ~new_n30532_;
  assign new_n30534_ = new_n28016_ & ~new_n30533_;
  assign new_n30535_ = ~new_n27996_ & new_n30534_;
  assign new_n30536_ = ~new_n30516_ & ~new_n30535_;
  assign new_n30537_ = ~new_n15156_ & ~new_n30536_;
  assign new_n30538_ = ys__n26153 & new_n15156_;
  assign ys__n26154 = new_n30537_ | new_n30538_;
  assign new_n30540_ = ys__n25999 & new_n27902_;
  assign new_n30541_ = ys__n18043 & new_n13490_;
  assign new_n30542_ = ys__n18049 & new_n13382_;
  assign new_n30543_ = ~new_n30541_ & ~new_n30542_;
  assign new_n30544_ = ys__n18055 & new_n13379_;
  assign new_n30545_ = ys__n18063 & new_n13380_;
  assign new_n30546_ = ~new_n30544_ & ~new_n30545_;
  assign new_n30547_ = new_n30543_ & new_n30546_;
  assign new_n30548_ = new_n27913_ & ~new_n30547_;
  assign new_n30549_ = ys__n46264 & new_n13490_;
  assign new_n30550_ = ys__n46440 & new_n13382_;
  assign new_n30551_ = ~new_n30549_ & ~new_n30550_;
  assign new_n30552_ = ys__n46616 & new_n13379_;
  assign new_n30553_ = ys__n46792 & new_n13380_;
  assign new_n30554_ = ~new_n30552_ & ~new_n30553_;
  assign new_n30555_ = new_n30551_ & new_n30554_;
  assign new_n30556_ = new_n27922_ & ~new_n30555_;
  assign new_n30557_ = ~new_n30548_ & ~new_n30556_;
  assign new_n30558_ = ys__n46321 & new_n13490_;
  assign new_n30559_ = ys__n46497 & new_n13382_;
  assign new_n30560_ = ~new_n30558_ & ~new_n30559_;
  assign new_n30561_ = ys__n46673 & new_n13379_;
  assign new_n30562_ = ys__n46849 & new_n13380_;
  assign new_n30563_ = ~new_n30561_ & ~new_n30562_;
  assign new_n30564_ = new_n30560_ & new_n30563_;
  assign new_n30565_ = new_n27932_ & ~new_n30564_;
  assign new_n30566_ = ys__n46398 & new_n13490_;
  assign new_n30567_ = ys__n46574 & new_n13382_;
  assign new_n30568_ = ~new_n30566_ & ~new_n30567_;
  assign new_n30569_ = ys__n46750 & new_n13379_;
  assign new_n30570_ = ys__n46926 & new_n13380_;
  assign new_n30571_ = ~new_n30569_ & ~new_n30570_;
  assign new_n30572_ = new_n30568_ & new_n30571_;
  assign new_n30573_ = new_n27941_ & ~new_n30572_;
  assign new_n30574_ = ~new_n30565_ & ~new_n30573_;
  assign new_n30575_ = new_n30557_ & new_n30574_;
  assign new_n30576_ = new_n27952_ & ~new_n30575_;
  assign new_n30577_ = ~new_n30540_ & ~new_n30576_;
  assign new_n30578_ = new_n27955_ & ~new_n30577_;
  assign new_n30579_ = ys__n45646 & new_n13490_;
  assign new_n30580_ = ys__n45482 & new_n13382_;
  assign new_n30581_ = ~new_n30579_ & ~new_n30580_;
  assign new_n30582_ = ys__n45318 & new_n13379_;
  assign new_n30583_ = ys__n45131 & new_n13380_;
  assign new_n30584_ = ~new_n30582_ & ~new_n30583_;
  assign new_n30585_ = new_n30581_ & new_n30584_;
  assign new_n30586_ = new_n27913_ & ~new_n30585_;
  assign new_n30587_ = ys__n45608 & new_n13490_;
  assign new_n30588_ = ys__n45444 & new_n13382_;
  assign new_n30589_ = ~new_n30587_ & ~new_n30588_;
  assign new_n30590_ = ys__n45280 & new_n13379_;
  assign new_n30591_ = ys__n45086 & new_n13380_;
  assign new_n30592_ = ~new_n30590_ & ~new_n30591_;
  assign new_n30593_ = new_n30589_ & new_n30592_;
  assign new_n30594_ = new_n27922_ & ~new_n30593_;
  assign new_n30595_ = ~new_n30586_ & ~new_n30594_;
  assign new_n30596_ = ys__n45700 & new_n13490_;
  assign new_n30597_ = ys__n45536 & new_n13382_;
  assign new_n30598_ = ~new_n30596_ & ~new_n30597_;
  assign new_n30599_ = ys__n45372 & new_n13379_;
  assign new_n30600_ = ys__n45210 & new_n13380_;
  assign new_n30601_ = ~new_n30599_ & ~new_n30600_;
  assign new_n30602_ = new_n30598_ & new_n30601_;
  assign new_n30603_ = new_n27932_ & ~new_n30602_;
  assign new_n30604_ = ys__n45552 & new_n13490_;
  assign new_n30605_ = ys__n45388 & new_n13382_;
  assign new_n30606_ = ~new_n30604_ & ~new_n30605_;
  assign new_n30607_ = ys__n45224 & new_n13379_;
  assign new_n30608_ = ys__n45005 & new_n13380_;
  assign new_n30609_ = ~new_n30607_ & ~new_n30608_;
  assign new_n30610_ = new_n30606_ & new_n30609_;
  assign new_n30611_ = new_n27941_ & ~new_n30610_;
  assign new_n30612_ = ~new_n30603_ & ~new_n30611_;
  assign new_n30613_ = new_n30595_ & new_n30612_;
  assign new_n30614_ = new_n27993_ & ~new_n30613_;
  assign new_n30615_ = ~new_n30578_ & ~new_n30614_;
  assign new_n30616_ = new_n27996_ & ~new_n30615_;
  assign new_n30617_ = ys__n46101 & new_n13490_;
  assign new_n30618_ = ys__n46003 & new_n13382_;
  assign new_n30619_ = ~new_n30617_ & ~new_n30618_;
  assign new_n30620_ = ys__n45905 & new_n13379_;
  assign new_n30621_ = ys__n45809 & new_n13380_;
  assign new_n30622_ = ~new_n30620_ & ~new_n30621_;
  assign new_n30623_ = new_n30619_ & new_n30622_;
  assign new_n30624_ = new_n27922_ & ~new_n30623_;
  assign new_n30625_ = ys__n46044 & new_n13490_;
  assign new_n30626_ = ys__n45946 & new_n13382_;
  assign new_n30627_ = ~new_n30625_ & ~new_n30626_;
  assign new_n30628_ = ys__n45848 & new_n13379_;
  assign new_n30629_ = ys__n45727 & new_n13380_;
  assign new_n30630_ = ~new_n30628_ & ~new_n30629_;
  assign new_n30631_ = new_n30627_ & new_n30630_;
  assign new_n30632_ = new_n27941_ & ~new_n30631_;
  assign new_n30633_ = ~new_n30624_ & ~new_n30632_;
  assign new_n30634_ = new_n28016_ & ~new_n30633_;
  assign new_n30635_ = ~new_n27996_ & new_n30634_;
  assign new_n30636_ = ~new_n30616_ & ~new_n30635_;
  assign new_n30637_ = ~new_n15156_ & ~new_n30636_;
  assign new_n30638_ = ys__n26155 & new_n15156_;
  assign ys__n26156 = new_n30637_ | new_n30638_;
  assign new_n30640_ = ys__n26068 & new_n27902_;
  assign new_n30641_ = ys__n46388 & new_n13490_;
  assign new_n30642_ = ys__n46564 & new_n13382_;
  assign new_n30643_ = ~new_n30641_ & ~new_n30642_;
  assign new_n30644_ = ys__n46740 & new_n13379_;
  assign new_n30645_ = ys__n46916 & new_n13380_;
  assign new_n30646_ = ~new_n30644_ & ~new_n30645_;
  assign new_n30647_ = new_n30643_ & new_n30646_;
  assign new_n30648_ = new_n27913_ & ~new_n30647_;
  assign new_n30649_ = ys__n46310 & new_n13490_;
  assign new_n30650_ = ys__n46486 & new_n13382_;
  assign new_n30651_ = ~new_n30649_ & ~new_n30650_;
  assign new_n30652_ = ys__n46662 & new_n13379_;
  assign new_n30653_ = ys__n46838 & new_n13380_;
  assign new_n30654_ = ~new_n30652_ & ~new_n30653_;
  assign new_n30655_ = new_n30651_ & new_n30654_;
  assign new_n30656_ = new_n27922_ & ~new_n30655_;
  assign new_n30657_ = ~new_n30648_ & ~new_n30656_;
  assign new_n30658_ = ys__n46344 & new_n13490_;
  assign new_n30659_ = ys__n46520 & new_n13382_;
  assign new_n30660_ = ~new_n30658_ & ~new_n30659_;
  assign new_n30661_ = ys__n46696 & new_n13379_;
  assign new_n30662_ = ys__n46872 & new_n13380_;
  assign new_n30663_ = ~new_n30661_ & ~new_n30662_;
  assign new_n30664_ = new_n30660_ & new_n30663_;
  assign new_n30665_ = new_n27932_ & ~new_n30664_;
  assign new_n30666_ = ys__n46421 & new_n13490_;
  assign new_n30667_ = ys__n46597 & new_n13382_;
  assign new_n30668_ = ~new_n30666_ & ~new_n30667_;
  assign new_n30669_ = ys__n46773 & new_n13379_;
  assign new_n30670_ = ys__n46949 & new_n13380_;
  assign new_n30671_ = ~new_n30669_ & ~new_n30670_;
  assign new_n30672_ = new_n30668_ & new_n30671_;
  assign new_n30673_ = new_n27941_ & ~new_n30672_;
  assign new_n30674_ = ~new_n30665_ & ~new_n30673_;
  assign new_n30675_ = new_n30657_ & new_n30674_;
  assign new_n30676_ = new_n27952_ & ~new_n30675_;
  assign new_n30677_ = ~new_n30640_ & ~new_n30676_;
  assign new_n30678_ = new_n27955_ & ~new_n30677_;
  assign new_n30679_ = ys__n45598 & new_n13490_;
  assign new_n30680_ = ys__n45434 & new_n13382_;
  assign new_n30681_ = ~new_n30679_ & ~new_n30680_;
  assign new_n30682_ = ys__n45270 & new_n13379_;
  assign new_n30683_ = ys__n45074 & new_n13380_;
  assign new_n30684_ = ~new_n30682_ & ~new_n30683_;
  assign new_n30685_ = new_n30681_ & new_n30684_;
  assign new_n30686_ = new_n27941_ & ~new_n30685_;
  assign new_n30687_ = ys__n45692 & new_n13490_;
  assign new_n30688_ = ys__n45528 & new_n13382_;
  assign new_n30689_ = ~new_n30687_ & ~new_n30688_;
  assign new_n30690_ = ys__n45364 & new_n13379_;
  assign new_n30691_ = ys__n45200 & new_n13380_;
  assign new_n30692_ = ~new_n30690_ & ~new_n30691_;
  assign new_n30693_ = new_n30689_ & new_n30692_;
  assign new_n30694_ = new_n27913_ & ~new_n30693_;
  assign new_n30695_ = ys__n45631 & new_n13490_;
  assign new_n30696_ = ys__n45467 & new_n13382_;
  assign new_n30697_ = ~new_n30695_ & ~new_n30696_;
  assign new_n30698_ = ys__n45303 & new_n13379_;
  assign new_n30699_ = ys__n45109 & new_n13380_;
  assign new_n30700_ = ~new_n30698_ & ~new_n30699_;
  assign new_n30701_ = new_n30697_ & new_n30700_;
  assign new_n30702_ = new_n27922_ & ~new_n30701_;
  assign new_n30703_ = ~new_n30694_ & ~new_n30702_;
  assign new_n30704_ = ~new_n30686_ & new_n30703_;
  assign new_n30705_ = new_n27993_ & ~new_n30704_;
  assign new_n30706_ = ~new_n30678_ & ~new_n30705_;
  assign new_n30707_ = new_n27996_ & ~new_n30706_;
  assign new_n30708_ = ys__n46124 & new_n13490_;
  assign new_n30709_ = ys__n46026 & new_n13382_;
  assign new_n30710_ = ~new_n30708_ & ~new_n30709_;
  assign new_n30711_ = ys__n45928 & new_n13379_;
  assign new_n30712_ = ys__n45832 & new_n13380_;
  assign new_n30713_ = ~new_n30711_ & ~new_n30712_;
  assign new_n30714_ = new_n30710_ & new_n30713_;
  assign new_n30715_ = new_n27922_ & ~new_n30714_;
  assign new_n30716_ = ys__n46090 & new_n13490_;
  assign new_n30717_ = ys__n45992 & new_n13382_;
  assign new_n30718_ = ~new_n30716_ & ~new_n30717_;
  assign new_n30719_ = ys__n45894 & new_n13379_;
  assign new_n30720_ = ys__n45796 & new_n13380_;
  assign new_n30721_ = ~new_n30719_ & ~new_n30720_;
  assign new_n30722_ = new_n30718_ & new_n30721_;
  assign new_n30723_ = new_n27941_ & ~new_n30722_;
  assign new_n30724_ = ~new_n30715_ & ~new_n30723_;
  assign new_n30725_ = new_n28016_ & ~new_n30724_;
  assign new_n30726_ = ~new_n27996_ & new_n30725_;
  assign new_n30727_ = ~new_n30707_ & ~new_n30726_;
  assign new_n30728_ = ~new_n15156_ & ~new_n30727_;
  assign new_n30729_ = ys__n26157 & new_n15156_;
  assign ys__n26158 = new_n30728_ | new_n30729_;
  assign new_n30731_ = ys__n26074 & new_n27902_;
  assign new_n30732_ = ys__n46392 & new_n13490_;
  assign new_n30733_ = ys__n46568 & new_n13382_;
  assign new_n30734_ = ~new_n30732_ & ~new_n30733_;
  assign new_n30735_ = ys__n46744 & new_n13379_;
  assign new_n30736_ = ys__n46920 & new_n13380_;
  assign new_n30737_ = ~new_n30735_ & ~new_n30736_;
  assign new_n30738_ = new_n30734_ & new_n30737_;
  assign new_n30739_ = new_n27913_ & ~new_n30738_;
  assign new_n30740_ = ys__n46314 & new_n13490_;
  assign new_n30741_ = ys__n46490 & new_n13382_;
  assign new_n30742_ = ~new_n30740_ & ~new_n30741_;
  assign new_n30743_ = ys__n46666 & new_n13379_;
  assign new_n30744_ = ys__n46842 & new_n13380_;
  assign new_n30745_ = ~new_n30743_ & ~new_n30744_;
  assign new_n30746_ = new_n30742_ & new_n30745_;
  assign new_n30747_ = new_n27922_ & ~new_n30746_;
  assign new_n30748_ = ~new_n30739_ & ~new_n30747_;
  assign new_n30749_ = ys__n46346 & new_n13490_;
  assign new_n30750_ = ys__n46522 & new_n13382_;
  assign new_n30751_ = ~new_n30749_ & ~new_n30750_;
  assign new_n30752_ = ys__n46698 & new_n13379_;
  assign new_n30753_ = ys__n46874 & new_n13380_;
  assign new_n30754_ = ~new_n30752_ & ~new_n30753_;
  assign new_n30755_ = new_n30751_ & new_n30754_;
  assign new_n30756_ = new_n27932_ & ~new_n30755_;
  assign new_n30757_ = ys__n46423 & new_n13490_;
  assign new_n30758_ = ys__n46599 & new_n13382_;
  assign new_n30759_ = ~new_n30757_ & ~new_n30758_;
  assign new_n30760_ = ys__n46775 & new_n13379_;
  assign new_n30761_ = ys__n46951 & new_n13380_;
  assign new_n30762_ = ~new_n30760_ & ~new_n30761_;
  assign new_n30763_ = new_n30759_ & new_n30762_;
  assign new_n30764_ = new_n27941_ & ~new_n30763_;
  assign new_n30765_ = ~new_n30756_ & ~new_n30764_;
  assign new_n30766_ = new_n30748_ & new_n30765_;
  assign new_n30767_ = new_n27952_ & ~new_n30766_;
  assign new_n30768_ = ~new_n30731_ & ~new_n30767_;
  assign new_n30769_ = new_n27955_ & ~new_n30768_;
  assign new_n30770_ = ys__n45602 & new_n13490_;
  assign new_n30771_ = ys__n45438 & new_n13382_;
  assign new_n30772_ = ~new_n30770_ & ~new_n30771_;
  assign new_n30773_ = ys__n45274 & new_n13379_;
  assign new_n30774_ = ys__n45080 & new_n13380_;
  assign new_n30775_ = ~new_n30773_ & ~new_n30774_;
  assign new_n30776_ = new_n30772_ & new_n30775_;
  assign new_n30777_ = new_n27941_ & ~new_n30776_;
  assign new_n30778_ = ys__n45696 & new_n13490_;
  assign new_n30779_ = ys__n45532 & new_n13382_;
  assign new_n30780_ = ~new_n30778_ & ~new_n30779_;
  assign new_n30781_ = ys__n45368 & new_n13379_;
  assign new_n30782_ = ys__n45206 & new_n13380_;
  assign new_n30783_ = ~new_n30781_ & ~new_n30782_;
  assign new_n30784_ = new_n30780_ & new_n30783_;
  assign new_n30785_ = new_n27913_ & ~new_n30784_;
  assign new_n30786_ = ys__n45633 & new_n13490_;
  assign new_n30787_ = ys__n45469 & new_n13382_;
  assign new_n30788_ = ~new_n30786_ & ~new_n30787_;
  assign new_n30789_ = ys__n45305 & new_n13379_;
  assign new_n30790_ = ys__n45111 & new_n13380_;
  assign new_n30791_ = ~new_n30789_ & ~new_n30790_;
  assign new_n30792_ = new_n30788_ & new_n30791_;
  assign new_n30793_ = new_n27922_ & ~new_n30792_;
  assign new_n30794_ = ~new_n30785_ & ~new_n30793_;
  assign new_n30795_ = ~new_n30777_ & new_n30794_;
  assign new_n30796_ = new_n27993_ & ~new_n30795_;
  assign new_n30797_ = ~new_n30769_ & ~new_n30796_;
  assign new_n30798_ = new_n27996_ & ~new_n30797_;
  assign new_n30799_ = ys__n46126 & new_n13490_;
  assign new_n30800_ = ys__n46028 & new_n13382_;
  assign new_n30801_ = ~new_n30799_ & ~new_n30800_;
  assign new_n30802_ = ys__n45930 & new_n13379_;
  assign new_n30803_ = ys__n45834 & new_n13380_;
  assign new_n30804_ = ~new_n30802_ & ~new_n30803_;
  assign new_n30805_ = new_n30801_ & new_n30804_;
  assign new_n30806_ = new_n27922_ & ~new_n30805_;
  assign new_n30807_ = ys__n46094 & new_n13490_;
  assign new_n30808_ = ys__n45996 & new_n13382_;
  assign new_n30809_ = ~new_n30807_ & ~new_n30808_;
  assign new_n30810_ = ys__n45898 & new_n13379_;
  assign new_n30811_ = ys__n45802 & new_n13380_;
  assign new_n30812_ = ~new_n30810_ & ~new_n30811_;
  assign new_n30813_ = new_n30809_ & new_n30812_;
  assign new_n30814_ = new_n27941_ & ~new_n30813_;
  assign new_n30815_ = ~new_n30806_ & ~new_n30814_;
  assign new_n30816_ = new_n28016_ & ~new_n30815_;
  assign new_n30817_ = ~new_n27996_ & new_n30816_;
  assign new_n30818_ = ~new_n30798_ & ~new_n30817_;
  assign new_n30819_ = ~new_n15156_ & ~new_n30818_;
  assign new_n30820_ = ys__n26159 & new_n15156_;
  assign ys__n26160 = new_n30819_ | new_n30820_;
  assign new_n30822_ = ys__n18833 & ~ys__n18174;
  assign new_n30823_ = ys__n26161 & ys__n18174;
  assign new_n30824_ = ~new_n30822_ & ~new_n30823_;
  assign new_n30825_ = ys__n18169 & ys__n18170;
  assign new_n30826_ = ~new_n30824_ & ~new_n30825_;
  assign new_n30827_ = new_n30824_ & new_n30825_;
  assign ys__n26220 = new_n30826_ | new_n30827_;
  assign new_n30829_ = ys__n18835 & ~ys__n18174;
  assign new_n30830_ = ys__n26162 & ys__n18174;
  assign new_n30831_ = ~new_n30829_ & ~new_n30830_;
  assign new_n30832_ = ~new_n30825_ & ~new_n30831_;
  assign new_n30833_ = ~new_n30824_ & new_n30831_;
  assign new_n30834_ = new_n30824_ & ~new_n30831_;
  assign new_n30835_ = ~new_n30833_ & ~new_n30834_;
  assign new_n30836_ = new_n30825_ & ~new_n30835_;
  assign ys__n26222 = new_n30832_ | new_n30836_;
  assign new_n30838_ = ys__n18837 & ~ys__n18174;
  assign new_n30839_ = ys__n26164 & ys__n18174;
  assign new_n30840_ = ~new_n30838_ & ~new_n30839_;
  assign new_n30841_ = ~new_n30825_ & ~new_n30840_;
  assign new_n30842_ = ~new_n30824_ & ~new_n30831_;
  assign new_n30843_ = new_n30840_ & new_n30842_;
  assign new_n30844_ = ~new_n30840_ & ~new_n30842_;
  assign new_n30845_ = ~new_n30843_ & ~new_n30844_;
  assign new_n30846_ = new_n30825_ & ~new_n30845_;
  assign ys__n26224 = new_n30841_ | new_n30846_;
  assign new_n30848_ = ys__n18839 & ~ys__n18174;
  assign new_n30849_ = ys__n26166 & ys__n18174;
  assign new_n30850_ = ~new_n30848_ & ~new_n30849_;
  assign new_n30851_ = ~new_n30825_ & ~new_n30850_;
  assign new_n30852_ = ~new_n30840_ & new_n30842_;
  assign new_n30853_ = new_n30850_ & new_n30852_;
  assign new_n30854_ = ~new_n30850_ & ~new_n30852_;
  assign new_n30855_ = ~new_n30853_ & ~new_n30854_;
  assign new_n30856_ = new_n30825_ & ~new_n30855_;
  assign ys__n26226 = new_n30851_ | new_n30856_;
  assign new_n30858_ = ys__n18841 & ~ys__n18174;
  assign new_n30859_ = ys__n26168 & ys__n18174;
  assign new_n30860_ = ~new_n30858_ & ~new_n30859_;
  assign new_n30861_ = ~new_n30825_ & ~new_n30860_;
  assign new_n30862_ = ~new_n30840_ & ~new_n30850_;
  assign new_n30863_ = new_n30842_ & new_n30862_;
  assign new_n30864_ = new_n30860_ & new_n30863_;
  assign new_n30865_ = ~new_n30860_ & ~new_n30863_;
  assign new_n30866_ = ~new_n30864_ & ~new_n30865_;
  assign new_n30867_ = new_n30825_ & ~new_n30866_;
  assign ys__n26228 = new_n30861_ | new_n30867_;
  assign new_n30869_ = ys__n18843 & ~ys__n18174;
  assign new_n30870_ = ys__n26170 & ys__n18174;
  assign new_n30871_ = ~new_n30869_ & ~new_n30870_;
  assign new_n30872_ = ~new_n30825_ & ~new_n30871_;
  assign new_n30873_ = ~new_n30860_ & new_n30863_;
  assign new_n30874_ = new_n30871_ & new_n30873_;
  assign new_n30875_ = ~new_n30871_ & ~new_n30873_;
  assign new_n30876_ = ~new_n30874_ & ~new_n30875_;
  assign new_n30877_ = new_n30825_ & ~new_n30876_;
  assign ys__n26230 = new_n30872_ | new_n30877_;
  assign new_n30879_ = ys__n18845 & ~ys__n18174;
  assign new_n30880_ = ys__n26172 & ys__n18174;
  assign new_n30881_ = ~new_n30879_ & ~new_n30880_;
  assign new_n30882_ = ~new_n30825_ & ~new_n30881_;
  assign new_n30883_ = ~new_n30860_ & ~new_n30871_;
  assign new_n30884_ = new_n30842_ & new_n30883_;
  assign new_n30885_ = new_n30862_ & new_n30884_;
  assign new_n30886_ = new_n30881_ & new_n30885_;
  assign new_n30887_ = ~new_n30881_ & ~new_n30885_;
  assign new_n30888_ = ~new_n30886_ & ~new_n30887_;
  assign new_n30889_ = new_n30825_ & ~new_n30888_;
  assign ys__n26232 = new_n30882_ | new_n30889_;
  assign new_n30891_ = ys__n18847 & ~ys__n18174;
  assign new_n30892_ = ys__n26174 & ys__n18174;
  assign new_n30893_ = ~new_n30891_ & ~new_n30892_;
  assign new_n30894_ = ~new_n30825_ & ~new_n30893_;
  assign new_n30895_ = ~new_n30881_ & new_n30885_;
  assign new_n30896_ = new_n30893_ & new_n30895_;
  assign new_n30897_ = ~new_n30893_ & ~new_n30895_;
  assign new_n30898_ = ~new_n30896_ & ~new_n30897_;
  assign new_n30899_ = new_n30825_ & ~new_n30898_;
  assign ys__n26234 = new_n30894_ | new_n30899_;
  assign new_n30901_ = ys__n18849 & ~ys__n18174;
  assign new_n30902_ = ys__n26176 & ys__n18174;
  assign new_n30903_ = ~new_n30901_ & ~new_n30902_;
  assign new_n30904_ = ~new_n30825_ & ~new_n30903_;
  assign new_n30905_ = ~new_n30881_ & ~new_n30893_;
  assign new_n30906_ = new_n30885_ & new_n30905_;
  assign new_n30907_ = new_n30903_ & new_n30906_;
  assign new_n30908_ = ~new_n30903_ & ~new_n30906_;
  assign new_n30909_ = ~new_n30907_ & ~new_n30908_;
  assign new_n30910_ = new_n30825_ & ~new_n30909_;
  assign ys__n26236 = new_n30904_ | new_n30910_;
  assign new_n30912_ = ys__n18851 & ~ys__n18174;
  assign new_n30913_ = ys__n26178 & ys__n18174;
  assign new_n30914_ = ~new_n30912_ & ~new_n30913_;
  assign new_n30915_ = ~new_n30825_ & ~new_n30914_;
  assign new_n30916_ = ~new_n30903_ & new_n30906_;
  assign new_n30917_ = new_n30914_ & new_n30916_;
  assign new_n30918_ = ~new_n30914_ & ~new_n30916_;
  assign new_n30919_ = ~new_n30917_ & ~new_n30918_;
  assign new_n30920_ = new_n30825_ & ~new_n30919_;
  assign ys__n26238 = new_n30915_ | new_n30920_;
  assign new_n30922_ = ys__n18853 & ~ys__n18174;
  assign new_n30923_ = ys__n26180 & ys__n18174;
  assign new_n30924_ = ~new_n30922_ & ~new_n30923_;
  assign new_n30925_ = ~new_n30825_ & ~new_n30924_;
  assign new_n30926_ = ~new_n30903_ & ~new_n30914_;
  assign new_n30927_ = new_n30905_ & new_n30926_;
  assign new_n30928_ = new_n30885_ & new_n30927_;
  assign new_n30929_ = new_n30924_ & new_n30928_;
  assign new_n30930_ = ~new_n30924_ & ~new_n30928_;
  assign new_n30931_ = ~new_n30929_ & ~new_n30930_;
  assign new_n30932_ = new_n30825_ & ~new_n30931_;
  assign ys__n26240 = new_n30925_ | new_n30932_;
  assign new_n30934_ = ys__n18855 & ~ys__n18174;
  assign new_n30935_ = ys__n26182 & ys__n18174;
  assign new_n30936_ = ~new_n30934_ & ~new_n30935_;
  assign new_n30937_ = ~new_n30825_ & ~new_n30936_;
  assign new_n30938_ = ~new_n30924_ & new_n30928_;
  assign new_n30939_ = new_n30936_ & new_n30938_;
  assign new_n30940_ = ~new_n30936_ & ~new_n30938_;
  assign new_n30941_ = ~new_n30939_ & ~new_n30940_;
  assign new_n30942_ = new_n30825_ & ~new_n30941_;
  assign ys__n26242 = new_n30937_ | new_n30942_;
  assign new_n30944_ = ys__n18857 & ~ys__n18174;
  assign new_n30945_ = ys__n26184 & ys__n18174;
  assign new_n30946_ = ~new_n30944_ & ~new_n30945_;
  assign new_n30947_ = ~new_n30825_ & ~new_n30946_;
  assign new_n30948_ = ~new_n30924_ & ~new_n30936_;
  assign new_n30949_ = new_n30928_ & new_n30948_;
  assign new_n30950_ = new_n30946_ & new_n30949_;
  assign new_n30951_ = ~new_n30946_ & ~new_n30949_;
  assign new_n30952_ = ~new_n30950_ & ~new_n30951_;
  assign new_n30953_ = new_n30825_ & ~new_n30952_;
  assign ys__n26244 = new_n30947_ | new_n30953_;
  assign new_n30955_ = ys__n18859 & ~ys__n18174;
  assign new_n30956_ = ys__n26186 & ys__n18174;
  assign new_n30957_ = ~new_n30955_ & ~new_n30956_;
  assign new_n30958_ = ~new_n30825_ & ~new_n30957_;
  assign new_n30959_ = ~new_n30946_ & new_n30949_;
  assign new_n30960_ = new_n30957_ & new_n30959_;
  assign new_n30961_ = ~new_n30957_ & ~new_n30959_;
  assign new_n30962_ = ~new_n30960_ & ~new_n30961_;
  assign new_n30963_ = new_n30825_ & ~new_n30962_;
  assign ys__n26246 = new_n30958_ | new_n30963_;
  assign new_n30965_ = ys__n18861 & ~ys__n18174;
  assign new_n30966_ = ys__n26188 & ys__n18174;
  assign new_n30967_ = ~new_n30965_ & ~new_n30966_;
  assign new_n30968_ = ~new_n30825_ & ~new_n30967_;
  assign new_n30969_ = ~new_n30946_ & ~new_n30957_;
  assign new_n30970_ = new_n30948_ & new_n30969_;
  assign new_n30971_ = new_n30927_ & new_n30970_;
  assign new_n30972_ = new_n30885_ & new_n30971_;
  assign new_n30973_ = new_n30967_ & new_n30972_;
  assign new_n30974_ = ~new_n30967_ & ~new_n30972_;
  assign new_n30975_ = ~new_n30973_ & ~new_n30974_;
  assign new_n30976_ = new_n30825_ & ~new_n30975_;
  assign ys__n26248 = new_n30968_ | new_n30976_;
  assign new_n30978_ = ys__n18863 & ~ys__n18174;
  assign new_n30979_ = ys__n26190 & ys__n18174;
  assign new_n30980_ = ~new_n30978_ & ~new_n30979_;
  assign new_n30981_ = ~new_n30825_ & ~new_n30980_;
  assign new_n30982_ = ~new_n30967_ & new_n30972_;
  assign new_n30983_ = new_n30980_ & new_n30982_;
  assign new_n30984_ = ~new_n30980_ & ~new_n30982_;
  assign new_n30985_ = ~new_n30983_ & ~new_n30984_;
  assign new_n30986_ = new_n30825_ & ~new_n30985_;
  assign ys__n26250 = new_n30981_ | new_n30986_;
  assign new_n30988_ = ys__n18865 & ~ys__n18174;
  assign new_n30989_ = ys__n26192 & ys__n18174;
  assign new_n30990_ = ~new_n30988_ & ~new_n30989_;
  assign new_n30991_ = ~new_n30825_ & ~new_n30990_;
  assign new_n30992_ = ~new_n30967_ & ~new_n30980_;
  assign new_n30993_ = new_n30972_ & new_n30992_;
  assign new_n30994_ = new_n30990_ & new_n30993_;
  assign new_n30995_ = ~new_n30990_ & ~new_n30993_;
  assign new_n30996_ = ~new_n30994_ & ~new_n30995_;
  assign new_n30997_ = new_n30825_ & ~new_n30996_;
  assign ys__n26252 = new_n30991_ | new_n30997_;
  assign new_n30999_ = ys__n18867 & ~ys__n18174;
  assign new_n31000_ = ys__n26194 & ys__n18174;
  assign new_n31001_ = ~new_n30999_ & ~new_n31000_;
  assign new_n31002_ = ~new_n30825_ & ~new_n31001_;
  assign new_n31003_ = ~new_n30990_ & new_n30993_;
  assign new_n31004_ = new_n31001_ & new_n31003_;
  assign new_n31005_ = ~new_n31001_ & ~new_n31003_;
  assign new_n31006_ = ~new_n31004_ & ~new_n31005_;
  assign new_n31007_ = new_n30825_ & ~new_n31006_;
  assign ys__n26254 = new_n31002_ | new_n31007_;
  assign new_n31009_ = ys__n18869 & ~ys__n18174;
  assign new_n31010_ = ys__n26196 & ys__n18174;
  assign new_n31011_ = ~new_n31009_ & ~new_n31010_;
  assign new_n31012_ = ~new_n30825_ & ~new_n31011_;
  assign new_n31013_ = ~new_n30990_ & ~new_n31001_;
  assign new_n31014_ = new_n30992_ & new_n31013_;
  assign new_n31015_ = new_n30972_ & new_n31014_;
  assign new_n31016_ = new_n31011_ & new_n31015_;
  assign new_n31017_ = ~new_n31011_ & ~new_n31015_;
  assign new_n31018_ = ~new_n31016_ & ~new_n31017_;
  assign new_n31019_ = new_n30825_ & ~new_n31018_;
  assign ys__n26256 = new_n31012_ | new_n31019_;
  assign new_n31021_ = ys__n18871 & ~ys__n18174;
  assign new_n31022_ = ys__n26198 & ys__n18174;
  assign new_n31023_ = ~new_n31021_ & ~new_n31022_;
  assign new_n31024_ = ~new_n30825_ & ~new_n31023_;
  assign new_n31025_ = ~new_n31011_ & new_n31015_;
  assign new_n31026_ = new_n31023_ & new_n31025_;
  assign new_n31027_ = ~new_n31023_ & ~new_n31025_;
  assign new_n31028_ = ~new_n31026_ & ~new_n31027_;
  assign new_n31029_ = new_n30825_ & ~new_n31028_;
  assign ys__n26258 = new_n31024_ | new_n31029_;
  assign new_n31031_ = ys__n18873 & ~ys__n18174;
  assign new_n31032_ = ys__n26200 & ys__n18174;
  assign new_n31033_ = ~new_n31031_ & ~new_n31032_;
  assign new_n31034_ = ~new_n30825_ & ~new_n31033_;
  assign new_n31035_ = ~new_n31011_ & ~new_n31023_;
  assign new_n31036_ = new_n31015_ & new_n31035_;
  assign new_n31037_ = new_n31033_ & new_n31036_;
  assign new_n31038_ = ~new_n31033_ & ~new_n31036_;
  assign new_n31039_ = ~new_n31037_ & ~new_n31038_;
  assign new_n31040_ = new_n30825_ & ~new_n31039_;
  assign ys__n26260 = new_n31034_ | new_n31040_;
  assign new_n31042_ = ys__n18875 & ~ys__n18174;
  assign new_n31043_ = ys__n26202 & ys__n18174;
  assign new_n31044_ = ~new_n31042_ & ~new_n31043_;
  assign new_n31045_ = ~new_n30825_ & ~new_n31044_;
  assign new_n31046_ = ~new_n31033_ & new_n31036_;
  assign new_n31047_ = new_n31044_ & new_n31046_;
  assign new_n31048_ = ~new_n31044_ & ~new_n31046_;
  assign new_n31049_ = ~new_n31047_ & ~new_n31048_;
  assign new_n31050_ = new_n30825_ & ~new_n31049_;
  assign ys__n26262 = new_n31045_ | new_n31050_;
  assign new_n31052_ = ys__n18877 & ~ys__n18174;
  assign new_n31053_ = ys__n26204 & ys__n18174;
  assign new_n31054_ = ~new_n31052_ & ~new_n31053_;
  assign new_n31055_ = ~new_n30825_ & ~new_n31054_;
  assign new_n31056_ = ~new_n31033_ & ~new_n31044_;
  assign new_n31057_ = new_n31035_ & new_n31056_;
  assign new_n31058_ = new_n31014_ & new_n31057_;
  assign new_n31059_ = new_n30972_ & new_n31058_;
  assign new_n31060_ = new_n31054_ & new_n31059_;
  assign new_n31061_ = ~new_n31054_ & ~new_n31059_;
  assign new_n31062_ = ~new_n31060_ & ~new_n31061_;
  assign new_n31063_ = new_n30825_ & ~new_n31062_;
  assign ys__n26264 = new_n31055_ | new_n31063_;
  assign new_n31065_ = ys__n18879 & ~ys__n18174;
  assign new_n31066_ = ys__n26206 & ys__n18174;
  assign new_n31067_ = ~new_n31065_ & ~new_n31066_;
  assign new_n31068_ = ~new_n30825_ & ~new_n31067_;
  assign new_n31069_ = ~new_n31054_ & new_n31059_;
  assign new_n31070_ = new_n31067_ & new_n31069_;
  assign new_n31071_ = ~new_n31067_ & ~new_n31069_;
  assign new_n31072_ = ~new_n31070_ & ~new_n31071_;
  assign new_n31073_ = new_n30825_ & ~new_n31072_;
  assign ys__n26266 = new_n31068_ | new_n31073_;
  assign new_n31075_ = ys__n18881 & ~ys__n18174;
  assign new_n31076_ = ys__n26208 & ys__n18174;
  assign new_n31077_ = ~new_n31075_ & ~new_n31076_;
  assign new_n31078_ = ~new_n30825_ & ~new_n31077_;
  assign new_n31079_ = ~new_n31054_ & ~new_n31067_;
  assign new_n31080_ = new_n31059_ & new_n31079_;
  assign new_n31081_ = new_n31077_ & new_n31080_;
  assign new_n31082_ = ~new_n31077_ & ~new_n31080_;
  assign new_n31083_ = ~new_n31081_ & ~new_n31082_;
  assign new_n31084_ = new_n30825_ & ~new_n31083_;
  assign ys__n26268 = new_n31078_ | new_n31084_;
  assign new_n31086_ = ys__n18883 & ~ys__n18174;
  assign new_n31087_ = ys__n26210 & ys__n18174;
  assign new_n31088_ = ~new_n31086_ & ~new_n31087_;
  assign new_n31089_ = ~new_n30825_ & ~new_n31088_;
  assign new_n31090_ = ~new_n31077_ & new_n31080_;
  assign new_n31091_ = new_n31088_ & new_n31090_;
  assign new_n31092_ = ~new_n31088_ & ~new_n31090_;
  assign new_n31093_ = ~new_n31091_ & ~new_n31092_;
  assign new_n31094_ = new_n30825_ & ~new_n31093_;
  assign ys__n26270 = new_n31089_ | new_n31094_;
  assign new_n31096_ = ys__n18885 & ~ys__n18174;
  assign new_n31097_ = ys__n26212 & ys__n18174;
  assign new_n31098_ = ~new_n31096_ & ~new_n31097_;
  assign new_n31099_ = ~new_n30825_ & ~new_n31098_;
  assign new_n31100_ = ~new_n31077_ & ~new_n31088_;
  assign new_n31101_ = new_n31079_ & new_n31100_;
  assign new_n31102_ = new_n31059_ & new_n31101_;
  assign new_n31103_ = new_n31098_ & new_n31102_;
  assign new_n31104_ = ~new_n31098_ & ~new_n31102_;
  assign new_n31105_ = ~new_n31103_ & ~new_n31104_;
  assign new_n31106_ = new_n30825_ & ~new_n31105_;
  assign ys__n26272 = new_n31099_ | new_n31106_;
  assign new_n31108_ = ys__n18887 & ~ys__n18174;
  assign new_n31109_ = ys__n26214 & ys__n18174;
  assign new_n31110_ = ~new_n31108_ & ~new_n31109_;
  assign new_n31111_ = ~new_n30825_ & ~new_n31110_;
  assign new_n31112_ = ~new_n31098_ & new_n31102_;
  assign new_n31113_ = new_n31110_ & new_n31112_;
  assign new_n31114_ = ~new_n31110_ & ~new_n31112_;
  assign new_n31115_ = ~new_n31113_ & ~new_n31114_;
  assign new_n31116_ = new_n30825_ & ~new_n31115_;
  assign ys__n26274 = new_n31111_ | new_n31116_;
  assign new_n31118_ = ys__n18889 & ~ys__n18174;
  assign new_n31119_ = ys__n26216 & ys__n18174;
  assign new_n31120_ = ~new_n31118_ & ~new_n31119_;
  assign new_n31121_ = ~new_n30825_ & ~new_n31120_;
  assign new_n31122_ = ~new_n31098_ & ~new_n31110_;
  assign new_n31123_ = new_n31102_ & new_n31122_;
  assign new_n31124_ = new_n31120_ & new_n31123_;
  assign new_n31125_ = ~new_n31120_ & ~new_n31123_;
  assign new_n31126_ = ~new_n31124_ & ~new_n31125_;
  assign new_n31127_ = new_n30825_ & ~new_n31126_;
  assign ys__n26276 = new_n31121_ | new_n31127_;
  assign new_n31129_ = ys__n18891 & ~ys__n18174;
  assign new_n31130_ = ys__n26218 & ys__n18174;
  assign new_n31131_ = ~new_n31129_ & ~new_n31130_;
  assign new_n31132_ = ~new_n30825_ & ~new_n31131_;
  assign new_n31133_ = ~new_n31120_ & new_n31123_;
  assign new_n31134_ = new_n31131_ & new_n31133_;
  assign new_n31135_ = ~new_n31131_ & ~new_n31133_;
  assign new_n31136_ = ~new_n31134_ & ~new_n31135_;
  assign new_n31137_ = new_n30825_ & ~new_n31136_;
  assign ys__n26278 = new_n31132_ | new_n31137_;
  assign new_n31139_ = ~ys__n26428 & ~ys__n30941;
  assign ys__n26282 = ys__n18169 & new_n31139_;
  assign new_n31141_ = ys__n26431 & ~ys__n30941;
  assign ys__n26284 = ys__n18169 & new_n31141_;
  assign ys__n26286 = ys__n26285 & ys__n18169;
  assign new_n31144_ = ys__n26460 & ~ys__n30941;
  assign ys__n26288 = ys__n18169 & new_n31144_;
  assign new_n31146_ = ys__n336 & ys__n776;
  assign ys__n26573 = new_n27802_ & new_n31146_;
  assign new_n31148_ = ys__n26569 & ~ys__n26573;
  assign new_n31149_ = ~ys__n18169 & new_n31148_;
  assign new_n31150_ = ~ys__n26478 & ys__n26493;
  assign new_n31151_ = ys__n35031 & new_n31150_;
  assign new_n31152_ = ys__n18169 & new_n31151_;
  assign ys__n26291 = new_n31149_ | new_n31152_;
  assign ys__n26293 = ~ys__n18466 & ys__n18178;
  assign ys__n26294 = ys__n18463 & ys__n18178;
  assign new_n31156_ = ~ys__n18208 & ~ys__n26565;
  assign new_n31157_ = ys__n26565 & ys__n30962;
  assign ys__n26566 = new_n31156_ | new_n31157_;
  assign new_n31159_ = ~ys__n778 & ys__n25980;
  assign new_n31160_ = new_n17862_ & ~new_n27812_;
  assign new_n31161_ = ys__n25980 & new_n31160_;
  assign new_n31162_ = ~ys__n18173 & ys__n18448;
  assign new_n31163_ = ys__n18173 & ys__n30877;
  assign new_n31164_ = ~new_n31162_ & ~new_n31163_;
  assign new_n31165_ = ~new_n17862_ & ~new_n31164_;
  assign new_n31166_ = ~new_n31160_ & new_n31165_;
  assign new_n31167_ = ~new_n31161_ & ~new_n31166_;
  assign new_n31168_ = ys__n778 & ~new_n31167_;
  assign new_n31169_ = ~new_n31159_ & ~new_n31168_;
  assign new_n31170_ = ~ys__n602 & ~new_n31169_;
  assign new_n31171_ = ~new_n17846_ & new_n27813_;
  assign new_n31172_ = ~new_n31169_ & new_n31171_;
  assign new_n31173_ = ys__n25984 & new_n17846_;
  assign new_n31174_ = ys__n25984 & ~new_n27813_;
  assign new_n31175_ = ~new_n31173_ & ~new_n31174_;
  assign new_n31176_ = ~new_n31171_ & ~new_n31175_;
  assign new_n31177_ = ~new_n31172_ & ~new_n31176_;
  assign new_n31178_ = ys__n602 & ~new_n31177_;
  assign ys__n26607 = new_n31170_ | new_n31178_;
  assign new_n31180_ = ~ys__n778 & ys__n25984;
  assign new_n31181_ = ys__n25984 & new_n31160_;
  assign new_n31182_ = ~ys__n18173 & ys__n18451;
  assign new_n31183_ = ys__n18173 & ys__n30879;
  assign new_n31184_ = ~new_n31182_ & ~new_n31183_;
  assign new_n31185_ = ~new_n17862_ & ~new_n31184_;
  assign new_n31186_ = ~new_n31160_ & new_n31185_;
  assign new_n31187_ = ~new_n31181_ & ~new_n31186_;
  assign new_n31188_ = ys__n778 & ~new_n31187_;
  assign new_n31189_ = ~new_n31180_ & ~new_n31188_;
  assign new_n31190_ = ~ys__n602 & ~new_n31189_;
  assign new_n31191_ = new_n31171_ & ~new_n31189_;
  assign new_n31192_ = ys__n25987 & new_n17846_;
  assign new_n31193_ = ys__n25987 & ~new_n27813_;
  assign new_n31194_ = ~new_n31192_ & ~new_n31193_;
  assign new_n31195_ = ~new_n31171_ & ~new_n31194_;
  assign new_n31196_ = ~new_n31191_ & ~new_n31195_;
  assign new_n31197_ = ys__n602 & ~new_n31196_;
  assign ys__n26609 = new_n31190_ | new_n31197_;
  assign new_n31199_ = ~ys__n778 & ys__n25987;
  assign new_n31200_ = ys__n25987 & new_n31160_;
  assign new_n31201_ = ~ys__n18173 & ys__n18454;
  assign new_n31202_ = ys__n18173 & ys__n30881;
  assign new_n31203_ = ~new_n31201_ & ~new_n31202_;
  assign new_n31204_ = ~new_n17862_ & ~new_n31203_;
  assign new_n31205_ = ~new_n31160_ & new_n31204_;
  assign new_n31206_ = ~new_n31200_ & ~new_n31205_;
  assign new_n31207_ = ys__n778 & ~new_n31206_;
  assign new_n31208_ = ~new_n31199_ & ~new_n31207_;
  assign new_n31209_ = ~ys__n602 & ~new_n31208_;
  assign new_n31210_ = new_n31171_ & ~new_n31208_;
  assign new_n31211_ = ys__n25990 & new_n17846_;
  assign new_n31212_ = ys__n25990 & ~new_n27813_;
  assign new_n31213_ = ~new_n31211_ & ~new_n31212_;
  assign new_n31214_ = ~new_n31171_ & ~new_n31213_;
  assign new_n31215_ = ~new_n31210_ & ~new_n31214_;
  assign new_n31216_ = ys__n602 & ~new_n31215_;
  assign ys__n26611 = new_n31209_ | new_n31216_;
  assign new_n31218_ = ~ys__n778 & ys__n25990;
  assign new_n31219_ = ys__n25990 & new_n31160_;
  assign new_n31220_ = ~ys__n18173 & ys__n18457;
  assign new_n31221_ = ys__n18173 & ys__n30883;
  assign new_n31222_ = ~new_n31220_ & ~new_n31221_;
  assign new_n31223_ = ~new_n17862_ & ~new_n31222_;
  assign new_n31224_ = ~new_n31160_ & new_n31223_;
  assign new_n31225_ = ~new_n31219_ & ~new_n31224_;
  assign new_n31226_ = ys__n778 & ~new_n31225_;
  assign new_n31227_ = ~new_n31218_ & ~new_n31226_;
  assign new_n31228_ = ~ys__n602 & ~new_n31227_;
  assign new_n31229_ = new_n31171_ & ~new_n31227_;
  assign new_n31230_ = ys__n25993 & new_n17846_;
  assign new_n31231_ = ys__n25993 & ~new_n27813_;
  assign new_n31232_ = ~new_n31230_ & ~new_n31231_;
  assign new_n31233_ = ~new_n31171_ & ~new_n31232_;
  assign new_n31234_ = ~new_n31229_ & ~new_n31233_;
  assign new_n31235_ = ys__n602 & ~new_n31234_;
  assign ys__n26613 = new_n31228_ | new_n31235_;
  assign new_n31237_ = ~ys__n778 & ys__n25993;
  assign new_n31238_ = ys__n25993 & new_n31160_;
  assign new_n31239_ = ~ys__n18173 & ys__n18460;
  assign new_n31240_ = ys__n18173 & ys__n30885;
  assign new_n31241_ = ~new_n31239_ & ~new_n31240_;
  assign new_n31242_ = ~new_n17862_ & ~new_n31241_;
  assign new_n31243_ = ~new_n31160_ & new_n31242_;
  assign new_n31244_ = ~new_n31238_ & ~new_n31243_;
  assign new_n31245_ = ys__n778 & ~new_n31244_;
  assign new_n31246_ = ~new_n31237_ & ~new_n31245_;
  assign new_n31247_ = ~ys__n602 & ~new_n31246_;
  assign new_n31248_ = new_n31171_ & ~new_n31246_;
  assign new_n31249_ = ys__n25996 & new_n17846_;
  assign new_n31250_ = ys__n25996 & ~new_n27813_;
  assign new_n31251_ = ~new_n31249_ & ~new_n31250_;
  assign new_n31252_ = ~new_n31171_ & ~new_n31251_;
  assign new_n31253_ = ~new_n31248_ & ~new_n31252_;
  assign new_n31254_ = ys__n602 & ~new_n31253_;
  assign ys__n26615 = new_n31247_ | new_n31254_;
  assign new_n31256_ = ~ys__n778 & ys__n25996;
  assign new_n31257_ = ys__n25996 & new_n31160_;
  assign new_n31258_ = ~ys__n18173 & ys__n18463;
  assign new_n31259_ = ys__n18173 & ys__n30887;
  assign new_n31260_ = ~new_n31258_ & ~new_n31259_;
  assign new_n31261_ = ~new_n17862_ & ~new_n31260_;
  assign new_n31262_ = ~new_n31160_ & new_n31261_;
  assign new_n31263_ = ~new_n31257_ & ~new_n31262_;
  assign new_n31264_ = ys__n778 & ~new_n31263_;
  assign new_n31265_ = ~new_n31256_ & ~new_n31264_;
  assign new_n31266_ = ~ys__n602 & ~new_n31265_;
  assign new_n31267_ = new_n31171_ & ~new_n31265_;
  assign new_n31268_ = ys__n25999 & new_n17846_;
  assign new_n31269_ = ys__n25999 & ~new_n27813_;
  assign new_n31270_ = ~new_n31268_ & ~new_n31269_;
  assign new_n31271_ = ~new_n31171_ & ~new_n31270_;
  assign new_n31272_ = ~new_n31267_ & ~new_n31271_;
  assign new_n31273_ = ys__n602 & ~new_n31272_;
  assign ys__n26617 = new_n31266_ | new_n31273_;
  assign new_n31275_ = ~ys__n778 & ys__n25999;
  assign new_n31276_ = ys__n25999 & new_n31160_;
  assign new_n31277_ = ~ys__n18173 & ys__n18466;
  assign new_n31278_ = ys__n18173 & ys__n30889;
  assign new_n31279_ = ~new_n31277_ & ~new_n31278_;
  assign new_n31280_ = ~new_n17862_ & ~new_n31279_;
  assign new_n31281_ = ~new_n31160_ & new_n31280_;
  assign new_n31282_ = ~new_n31276_ & ~new_n31281_;
  assign new_n31283_ = ys__n778 & ~new_n31282_;
  assign new_n31284_ = ~new_n31275_ & ~new_n31283_;
  assign new_n31285_ = ~ys__n602 & ~new_n31284_;
  assign new_n31286_ = new_n31171_ & ~new_n31284_;
  assign new_n31287_ = ys__n26002 & new_n17846_;
  assign new_n31288_ = ys__n26002 & ~new_n27813_;
  assign new_n31289_ = ~new_n31287_ & ~new_n31288_;
  assign new_n31290_ = ~new_n31171_ & ~new_n31289_;
  assign new_n31291_ = ~new_n31286_ & ~new_n31290_;
  assign new_n31292_ = ys__n602 & ~new_n31291_;
  assign ys__n26619 = new_n31285_ | new_n31292_;
  assign new_n31294_ = ~ys__n778 & ys__n26002;
  assign new_n31295_ = ys__n26002 & new_n31160_;
  assign new_n31296_ = ~ys__n18173 & ys__n18469;
  assign new_n31297_ = ys__n18173 & ys__n30891;
  assign new_n31298_ = ~new_n31296_ & ~new_n31297_;
  assign new_n31299_ = ~new_n17862_ & ~new_n31298_;
  assign new_n31300_ = ~new_n31160_ & new_n31299_;
  assign new_n31301_ = ~new_n31295_ & ~new_n31300_;
  assign new_n31302_ = ys__n778 & ~new_n31301_;
  assign new_n31303_ = ~new_n31294_ & ~new_n31302_;
  assign new_n31304_ = ~ys__n602 & ~new_n31303_;
  assign new_n31305_ = new_n31171_ & ~new_n31303_;
  assign new_n31306_ = ys__n26005 & new_n17846_;
  assign new_n31307_ = ys__n26005 & ~new_n27813_;
  assign new_n31308_ = ~new_n31306_ & ~new_n31307_;
  assign new_n31309_ = ~new_n31171_ & ~new_n31308_;
  assign new_n31310_ = ~new_n31305_ & ~new_n31309_;
  assign new_n31311_ = ys__n602 & ~new_n31310_;
  assign ys__n26621 = new_n31304_ | new_n31311_;
  assign new_n31313_ = ~ys__n778 & ys__n26005;
  assign new_n31314_ = ys__n26005 & new_n31160_;
  assign new_n31315_ = ys__n35059 & new_n27812_;
  assign new_n31316_ = ~ys__n18173 & ys__n18472;
  assign new_n31317_ = ys__n18173 & ys__n30893;
  assign new_n31318_ = ~new_n31316_ & ~new_n31317_;
  assign new_n31319_ = ~new_n17862_ & ~new_n31318_;
  assign new_n31320_ = ~new_n31315_ & ~new_n31319_;
  assign new_n31321_ = ~new_n31160_ & ~new_n31320_;
  assign new_n31322_ = ~new_n31314_ & ~new_n31321_;
  assign new_n31323_ = ys__n778 & ~new_n31322_;
  assign new_n31324_ = ~new_n31313_ & ~new_n31323_;
  assign new_n31325_ = ~ys__n602 & ~new_n31324_;
  assign new_n31326_ = new_n31171_ & ~new_n31324_;
  assign new_n31327_ = ys__n26008 & new_n17846_;
  assign new_n31328_ = ys__n26008 & ~new_n27813_;
  assign new_n31329_ = ~new_n31327_ & ~new_n31328_;
  assign new_n31330_ = ~new_n31171_ & ~new_n31329_;
  assign new_n31331_ = ~new_n31326_ & ~new_n31330_;
  assign new_n31332_ = ys__n602 & ~new_n31331_;
  assign ys__n26623 = new_n31325_ | new_n31332_;
  assign new_n31334_ = ~ys__n778 & ys__n26008;
  assign new_n31335_ = ys__n26008 & new_n31160_;
  assign new_n31336_ = ys__n35057 & new_n27812_;
  assign new_n31337_ = ~ys__n18173 & ys__n18475;
  assign new_n31338_ = ys__n18173 & ys__n30895;
  assign new_n31339_ = ~new_n31337_ & ~new_n31338_;
  assign new_n31340_ = ~new_n17862_ & ~new_n31339_;
  assign new_n31341_ = ~new_n31336_ & ~new_n31340_;
  assign new_n31342_ = ~new_n31160_ & ~new_n31341_;
  assign new_n31343_ = ~new_n31335_ & ~new_n31342_;
  assign new_n31344_ = ys__n778 & ~new_n31343_;
  assign new_n31345_ = ~new_n31334_ & ~new_n31344_;
  assign new_n31346_ = ~ys__n602 & ~new_n31345_;
  assign new_n31347_ = new_n31171_ & ~new_n31345_;
  assign new_n31348_ = ys__n26011 & new_n17846_;
  assign new_n31349_ = ys__n26011 & ~new_n27813_;
  assign new_n31350_ = ~new_n31348_ & ~new_n31349_;
  assign new_n31351_ = ~new_n31171_ & ~new_n31350_;
  assign new_n31352_ = ~new_n31347_ & ~new_n31351_;
  assign new_n31353_ = ys__n602 & ~new_n31352_;
  assign ys__n26625 = new_n31346_ | new_n31353_;
  assign new_n31355_ = ~ys__n778 & ys__n26011;
  assign new_n31356_ = ys__n26011 & new_n31160_;
  assign new_n31357_ = ~ys__n18173 & ys__n18478;
  assign new_n31358_ = ys__n18173 & ys__n30897;
  assign new_n31359_ = ~new_n31357_ & ~new_n31358_;
  assign new_n31360_ = ~new_n17862_ & ~new_n31359_;
  assign new_n31361_ = ~new_n31160_ & new_n31360_;
  assign new_n31362_ = ~new_n31356_ & ~new_n31361_;
  assign new_n31363_ = ys__n778 & ~new_n31362_;
  assign new_n31364_ = ~new_n31355_ & ~new_n31363_;
  assign new_n31365_ = ~ys__n602 & ~new_n31364_;
  assign new_n31366_ = new_n31171_ & ~new_n31364_;
  assign new_n31367_ = ys__n26014 & new_n17846_;
  assign new_n31368_ = ys__n26014 & ~new_n27813_;
  assign new_n31369_ = ~new_n31367_ & ~new_n31368_;
  assign new_n31370_ = ~new_n31171_ & ~new_n31369_;
  assign new_n31371_ = ~new_n31366_ & ~new_n31370_;
  assign new_n31372_ = ys__n602 & ~new_n31371_;
  assign ys__n26627 = new_n31365_ | new_n31372_;
  assign new_n31374_ = ~ys__n778 & ys__n26014;
  assign new_n31375_ = ys__n26014 & new_n31160_;
  assign new_n31376_ = ys__n184 & new_n27812_;
  assign new_n31377_ = ~ys__n18173 & ys__n18481;
  assign new_n31378_ = ys__n18173 & ys__n30899;
  assign new_n31379_ = ~new_n31377_ & ~new_n31378_;
  assign new_n31380_ = ~new_n17862_ & ~new_n31379_;
  assign new_n31381_ = ~new_n31376_ & ~new_n31380_;
  assign new_n31382_ = ~new_n31160_ & ~new_n31381_;
  assign new_n31383_ = ~new_n31375_ & ~new_n31382_;
  assign new_n31384_ = ys__n778 & ~new_n31383_;
  assign new_n31385_ = ~new_n31374_ & ~new_n31384_;
  assign new_n31386_ = ~ys__n602 & ~new_n31385_;
  assign new_n31387_ = new_n31171_ & ~new_n31385_;
  assign new_n31388_ = ys__n26017 & new_n17846_;
  assign new_n31389_ = ys__n26017 & ~new_n27813_;
  assign new_n31390_ = ~new_n31388_ & ~new_n31389_;
  assign new_n31391_ = ~new_n31171_ & ~new_n31390_;
  assign new_n31392_ = ~new_n31387_ & ~new_n31391_;
  assign new_n31393_ = ys__n602 & ~new_n31392_;
  assign ys__n26629 = new_n31386_ | new_n31393_;
  assign new_n31395_ = ~ys__n778 & ys__n26017;
  assign new_n31396_ = ys__n26017 & new_n31160_;
  assign new_n31397_ = ys__n182 & new_n27812_;
  assign new_n31398_ = ~ys__n18173 & ys__n18484;
  assign new_n31399_ = ys__n18173 & ys__n30901;
  assign new_n31400_ = ~new_n31398_ & ~new_n31399_;
  assign new_n31401_ = ~new_n17862_ & ~new_n31400_;
  assign new_n31402_ = ~new_n31397_ & ~new_n31401_;
  assign new_n31403_ = ~new_n31160_ & ~new_n31402_;
  assign new_n31404_ = ~new_n31396_ & ~new_n31403_;
  assign new_n31405_ = ys__n778 & ~new_n31404_;
  assign new_n31406_ = ~new_n31395_ & ~new_n31405_;
  assign new_n31407_ = ~ys__n602 & ~new_n31406_;
  assign new_n31408_ = new_n31171_ & ~new_n31406_;
  assign new_n31409_ = ys__n26020 & new_n17846_;
  assign new_n31410_ = ys__n26020 & ~new_n27813_;
  assign new_n31411_ = ~new_n31409_ & ~new_n31410_;
  assign new_n31412_ = ~new_n31171_ & ~new_n31411_;
  assign new_n31413_ = ~new_n31408_ & ~new_n31412_;
  assign new_n31414_ = ys__n602 & ~new_n31413_;
  assign ys__n26631 = new_n31407_ | new_n31414_;
  assign new_n31416_ = ~ys__n778 & ys__n26020;
  assign new_n31417_ = ys__n26020 & new_n31160_;
  assign new_n31418_ = ~ys__n18173 & ys__n18487;
  assign new_n31419_ = ys__n18173 & ys__n30903;
  assign new_n31420_ = ~new_n31418_ & ~new_n31419_;
  assign new_n31421_ = ~new_n17862_ & ~new_n31420_;
  assign new_n31422_ = ~new_n31160_ & new_n31421_;
  assign new_n31423_ = ~new_n31417_ & ~new_n31422_;
  assign new_n31424_ = ys__n778 & ~new_n31423_;
  assign new_n31425_ = ~new_n31416_ & ~new_n31424_;
  assign new_n31426_ = ~ys__n602 & ~new_n31425_;
  assign new_n31427_ = new_n31171_ & ~new_n31425_;
  assign new_n31428_ = ys__n26023 & new_n17846_;
  assign new_n31429_ = ys__n26023 & ~new_n27813_;
  assign new_n31430_ = ~new_n31428_ & ~new_n31429_;
  assign new_n31431_ = ~new_n31171_ & ~new_n31430_;
  assign new_n31432_ = ~new_n31427_ & ~new_n31431_;
  assign new_n31433_ = ys__n602 & ~new_n31432_;
  assign ys__n26633 = new_n31426_ | new_n31433_;
  assign new_n31435_ = ~ys__n778 & ys__n26023;
  assign new_n31436_ = ys__n26023 & new_n31160_;
  assign new_n31437_ = ~ys__n18173 & ys__n18490;
  assign new_n31438_ = ys__n18173 & ys__n30905;
  assign new_n31439_ = ~new_n31437_ & ~new_n31438_;
  assign new_n31440_ = ~new_n17862_ & ~new_n31439_;
  assign new_n31441_ = ~new_n31160_ & new_n31440_;
  assign new_n31442_ = ~new_n31436_ & ~new_n31441_;
  assign new_n31443_ = ys__n778 & ~new_n31442_;
  assign new_n31444_ = ~new_n31435_ & ~new_n31443_;
  assign new_n31445_ = ~ys__n602 & ~new_n31444_;
  assign new_n31446_ = new_n31171_ & ~new_n31444_;
  assign new_n31447_ = ys__n26026 & new_n17846_;
  assign new_n31448_ = ys__n26026 & ~new_n27813_;
  assign new_n31449_ = ~new_n31447_ & ~new_n31448_;
  assign new_n31450_ = ~new_n31171_ & ~new_n31449_;
  assign new_n31451_ = ~new_n31446_ & ~new_n31450_;
  assign new_n31452_ = ys__n602 & ~new_n31451_;
  assign ys__n26635 = new_n31445_ | new_n31452_;
  assign new_n31454_ = ~ys__n778 & ys__n26026;
  assign new_n31455_ = ys__n26026 & new_n31160_;
  assign new_n31456_ = ~ys__n18173 & ys__n18493;
  assign new_n31457_ = ys__n18173 & ys__n30907;
  assign new_n31458_ = ~new_n31456_ & ~new_n31457_;
  assign new_n31459_ = ~new_n17862_ & ~new_n31458_;
  assign new_n31460_ = ~new_n31160_ & new_n31459_;
  assign new_n31461_ = ~new_n31455_ & ~new_n31460_;
  assign new_n31462_ = ys__n778 & ~new_n31461_;
  assign new_n31463_ = ~new_n31454_ & ~new_n31462_;
  assign new_n31464_ = ~ys__n602 & ~new_n31463_;
  assign new_n31465_ = new_n31171_ & ~new_n31463_;
  assign new_n31466_ = ys__n26029 & new_n17846_;
  assign new_n31467_ = ys__n26029 & ~new_n27813_;
  assign new_n31468_ = ~new_n31466_ & ~new_n31467_;
  assign new_n31469_ = ~new_n31171_ & ~new_n31468_;
  assign new_n31470_ = ~new_n31465_ & ~new_n31469_;
  assign new_n31471_ = ys__n602 & ~new_n31470_;
  assign ys__n26637 = new_n31464_ | new_n31471_;
  assign new_n31473_ = ~ys__n778 & ys__n26029;
  assign new_n31474_ = ys__n26029 & new_n31160_;
  assign new_n31475_ = ~ys__n18173 & ys__n18496;
  assign new_n31476_ = ys__n18173 & ys__n30909;
  assign new_n31477_ = ~new_n31475_ & ~new_n31476_;
  assign new_n31478_ = ~new_n17862_ & ~new_n31477_;
  assign new_n31479_ = ~new_n27812_ & ~new_n31478_;
  assign new_n31480_ = ~new_n31160_ & ~new_n31479_;
  assign new_n31481_ = ~new_n31474_ & ~new_n31480_;
  assign new_n31482_ = ys__n778 & ~new_n31481_;
  assign new_n31483_ = ~new_n31473_ & ~new_n31482_;
  assign new_n31484_ = ~ys__n602 & ~new_n31483_;
  assign new_n31485_ = new_n31171_ & ~new_n31483_;
  assign new_n31486_ = ys__n26032 & new_n17846_;
  assign new_n31487_ = ys__n26032 & ~new_n27813_;
  assign new_n31488_ = ~new_n31486_ & ~new_n31487_;
  assign new_n31489_ = ~new_n31171_ & ~new_n31488_;
  assign new_n31490_ = ~new_n31485_ & ~new_n31489_;
  assign new_n31491_ = ys__n602 & ~new_n31490_;
  assign ys__n26639 = new_n31484_ | new_n31491_;
  assign new_n31493_ = ~ys__n778 & ys__n26032;
  assign new_n31494_ = ys__n26032 & new_n31160_;
  assign new_n31495_ = ~ys__n18173 & ys__n18499;
  assign new_n31496_ = ys__n18173 & ys__n30911;
  assign new_n31497_ = ~new_n31495_ & ~new_n31496_;
  assign new_n31498_ = ~new_n17862_ & ~new_n31497_;
  assign new_n31499_ = ~new_n31160_ & new_n31498_;
  assign new_n31500_ = ~new_n31494_ & ~new_n31499_;
  assign new_n31501_ = ys__n778 & ~new_n31500_;
  assign new_n31502_ = ~new_n31493_ & ~new_n31501_;
  assign new_n31503_ = ~ys__n602 & ~new_n31502_;
  assign new_n31504_ = new_n31171_ & ~new_n31502_;
  assign new_n31505_ = ys__n26035 & new_n17846_;
  assign new_n31506_ = ys__n26035 & ~new_n27813_;
  assign new_n31507_ = ~new_n31505_ & ~new_n31506_;
  assign new_n31508_ = ~new_n31171_ & ~new_n31507_;
  assign new_n31509_ = ~new_n31504_ & ~new_n31508_;
  assign new_n31510_ = ys__n602 & ~new_n31509_;
  assign ys__n26641 = new_n31503_ | new_n31510_;
  assign new_n31512_ = ~ys__n778 & ys__n26035;
  assign new_n31513_ = ys__n26035 & new_n31160_;
  assign new_n31514_ = ~ys__n18173 & ys__n18502;
  assign new_n31515_ = ys__n18173 & ys__n30913;
  assign new_n31516_ = ~new_n31514_ & ~new_n31515_;
  assign new_n31517_ = ~new_n17862_ & ~new_n31516_;
  assign new_n31518_ = ~new_n31160_ & new_n31517_;
  assign new_n31519_ = ~new_n31513_ & ~new_n31518_;
  assign new_n31520_ = ys__n778 & ~new_n31519_;
  assign new_n31521_ = ~new_n31512_ & ~new_n31520_;
  assign new_n31522_ = ~ys__n602 & ~new_n31521_;
  assign new_n31523_ = new_n31171_ & ~new_n31521_;
  assign new_n31524_ = ys__n26038 & new_n17846_;
  assign new_n31525_ = ys__n26038 & ~new_n27813_;
  assign new_n31526_ = ~new_n31524_ & ~new_n31525_;
  assign new_n31527_ = ~new_n31171_ & ~new_n31526_;
  assign new_n31528_ = ~new_n31523_ & ~new_n31527_;
  assign new_n31529_ = ys__n602 & ~new_n31528_;
  assign ys__n26643 = new_n31522_ | new_n31529_;
  assign new_n31531_ = ~ys__n778 & ys__n26038;
  assign new_n31532_ = ys__n26038 & new_n31160_;
  assign new_n31533_ = ~ys__n18173 & ys__n18505;
  assign new_n31534_ = ys__n18173 & ys__n30915;
  assign new_n31535_ = ~new_n31533_ & ~new_n31534_;
  assign new_n31536_ = ~new_n17862_ & ~new_n31535_;
  assign new_n31537_ = ~new_n31160_ & new_n31536_;
  assign new_n31538_ = ~new_n31532_ & ~new_n31537_;
  assign new_n31539_ = ys__n778 & ~new_n31538_;
  assign new_n31540_ = ~new_n31531_ & ~new_n31539_;
  assign new_n31541_ = ~ys__n602 & ~new_n31540_;
  assign new_n31542_ = new_n31171_ & ~new_n31540_;
  assign new_n31543_ = ys__n26041 & new_n17846_;
  assign new_n31544_ = ys__n26041 & ~new_n27813_;
  assign new_n31545_ = ~new_n31543_ & ~new_n31544_;
  assign new_n31546_ = ~new_n31171_ & ~new_n31545_;
  assign new_n31547_ = ~new_n31542_ & ~new_n31546_;
  assign new_n31548_ = ys__n602 & ~new_n31547_;
  assign ys__n26645 = new_n31541_ | new_n31548_;
  assign new_n31550_ = ~ys__n778 & ys__n26041;
  assign new_n31551_ = ys__n26041 & new_n31160_;
  assign new_n31552_ = ~ys__n18173 & ys__n18508;
  assign new_n31553_ = ys__n18173 & ys__n30917;
  assign new_n31554_ = ~new_n31552_ & ~new_n31553_;
  assign new_n31555_ = ~new_n17862_ & ~new_n31554_;
  assign new_n31556_ = ~new_n31160_ & new_n31555_;
  assign new_n31557_ = ~new_n31551_ & ~new_n31556_;
  assign new_n31558_ = ys__n778 & ~new_n31557_;
  assign new_n31559_ = ~new_n31550_ & ~new_n31558_;
  assign new_n31560_ = ~ys__n602 & ~new_n31559_;
  assign new_n31561_ = new_n31171_ & ~new_n31559_;
  assign new_n31562_ = ys__n26044 & new_n17846_;
  assign new_n31563_ = ys__n26044 & ~new_n27813_;
  assign new_n31564_ = ~new_n31562_ & ~new_n31563_;
  assign new_n31565_ = ~new_n31171_ & ~new_n31564_;
  assign new_n31566_ = ~new_n31561_ & ~new_n31565_;
  assign new_n31567_ = ys__n602 & ~new_n31566_;
  assign ys__n26647 = new_n31560_ | new_n31567_;
  assign new_n31569_ = ~ys__n778 & ys__n26044;
  assign new_n31570_ = ys__n26044 & new_n31160_;
  assign new_n31571_ = ~ys__n18173 & ys__n18511;
  assign new_n31572_ = ys__n18173 & ys__n30919;
  assign new_n31573_ = ~new_n31571_ & ~new_n31572_;
  assign new_n31574_ = ~new_n17862_ & ~new_n31573_;
  assign new_n31575_ = ~new_n31160_ & new_n31574_;
  assign new_n31576_ = ~new_n31570_ & ~new_n31575_;
  assign new_n31577_ = ys__n778 & ~new_n31576_;
  assign new_n31578_ = ~new_n31569_ & ~new_n31577_;
  assign new_n31579_ = ~ys__n602 & ~new_n31578_;
  assign new_n31580_ = new_n31171_ & ~new_n31578_;
  assign new_n31581_ = ys__n26047 & new_n17846_;
  assign new_n31582_ = ys__n26047 & ~new_n27813_;
  assign new_n31583_ = ~new_n31581_ & ~new_n31582_;
  assign new_n31584_ = ~new_n31171_ & ~new_n31583_;
  assign new_n31585_ = ~new_n31580_ & ~new_n31584_;
  assign new_n31586_ = ys__n602 & ~new_n31585_;
  assign ys__n26649 = new_n31579_ | new_n31586_;
  assign new_n31588_ = ~ys__n778 & ys__n26047;
  assign new_n31589_ = ys__n26047 & new_n31160_;
  assign new_n31590_ = ~ys__n18173 & ys__n18514;
  assign new_n31591_ = ys__n18173 & ys__n30921;
  assign new_n31592_ = ~new_n31590_ & ~new_n31591_;
  assign new_n31593_ = ~new_n17862_ & ~new_n31592_;
  assign new_n31594_ = ~new_n31160_ & new_n31593_;
  assign new_n31595_ = ~new_n31589_ & ~new_n31594_;
  assign new_n31596_ = ys__n778 & ~new_n31595_;
  assign new_n31597_ = ~new_n31588_ & ~new_n31596_;
  assign new_n31598_ = ~ys__n602 & ~new_n31597_;
  assign new_n31599_ = new_n31171_ & ~new_n31597_;
  assign new_n31600_ = ys__n26050 & new_n17846_;
  assign new_n31601_ = ys__n26050 & ~new_n27813_;
  assign new_n31602_ = ~new_n31600_ & ~new_n31601_;
  assign new_n31603_ = ~new_n31171_ & ~new_n31602_;
  assign new_n31604_ = ~new_n31599_ & ~new_n31603_;
  assign new_n31605_ = ys__n602 & ~new_n31604_;
  assign ys__n26651 = new_n31598_ | new_n31605_;
  assign new_n31607_ = ~ys__n778 & ys__n26050;
  assign new_n31608_ = ys__n26050 & new_n31160_;
  assign new_n31609_ = ~ys__n18173 & ys__n18517;
  assign new_n31610_ = ys__n18173 & ys__n30923;
  assign new_n31611_ = ~new_n31609_ & ~new_n31610_;
  assign new_n31612_ = ~new_n17862_ & ~new_n31611_;
  assign new_n31613_ = ~new_n27812_ & ~new_n31612_;
  assign new_n31614_ = ~new_n31160_ & ~new_n31613_;
  assign new_n31615_ = ~new_n31608_ & ~new_n31614_;
  assign new_n31616_ = ys__n778 & ~new_n31615_;
  assign new_n31617_ = ~new_n31607_ & ~new_n31616_;
  assign new_n31618_ = ~ys__n602 & ~new_n31617_;
  assign new_n31619_ = new_n31171_ & ~new_n31617_;
  assign new_n31620_ = ys__n26053 & new_n17846_;
  assign new_n31621_ = ys__n26053 & ~new_n27813_;
  assign new_n31622_ = ~new_n31620_ & ~new_n31621_;
  assign new_n31623_ = ~new_n31171_ & ~new_n31622_;
  assign new_n31624_ = ~new_n31619_ & ~new_n31623_;
  assign new_n31625_ = ys__n602 & ~new_n31624_;
  assign ys__n26653 = new_n31618_ | new_n31625_;
  assign new_n31627_ = ~ys__n778 & ys__n26053;
  assign new_n31628_ = ys__n26053 & new_n31160_;
  assign new_n31629_ = ~ys__n18173 & ys__n18520;
  assign new_n31630_ = ys__n18173 & ys__n30925;
  assign new_n31631_ = ~new_n31629_ & ~new_n31630_;
  assign new_n31632_ = ~new_n17862_ & ~new_n31631_;
  assign new_n31633_ = ~new_n31160_ & new_n31632_;
  assign new_n31634_ = ~new_n31628_ & ~new_n31633_;
  assign new_n31635_ = ys__n778 & ~new_n31634_;
  assign new_n31636_ = ~new_n31627_ & ~new_n31635_;
  assign new_n31637_ = ~ys__n602 & ~new_n31636_;
  assign new_n31638_ = new_n31171_ & ~new_n31636_;
  assign new_n31639_ = ys__n26056 & new_n17846_;
  assign new_n31640_ = ys__n26056 & ~new_n27813_;
  assign new_n31641_ = ~new_n31639_ & ~new_n31640_;
  assign new_n31642_ = ~new_n31171_ & ~new_n31641_;
  assign new_n31643_ = ~new_n31638_ & ~new_n31642_;
  assign new_n31644_ = ys__n602 & ~new_n31643_;
  assign ys__n26655 = new_n31637_ | new_n31644_;
  assign new_n31646_ = ~ys__n778 & ys__n26056;
  assign new_n31647_ = ys__n26056 & new_n31160_;
  assign new_n31648_ = ~ys__n18173 & ys__n18523;
  assign new_n31649_ = ys__n18173 & ys__n30927;
  assign new_n31650_ = ~new_n31648_ & ~new_n31649_;
  assign new_n31651_ = ~new_n17862_ & ~new_n31650_;
  assign new_n31652_ = ~new_n31160_ & new_n31651_;
  assign new_n31653_ = ~new_n31647_ & ~new_n31652_;
  assign new_n31654_ = ys__n778 & ~new_n31653_;
  assign new_n31655_ = ~new_n31646_ & ~new_n31654_;
  assign new_n31656_ = ~ys__n602 & ~new_n31655_;
  assign new_n31657_ = new_n31171_ & ~new_n31655_;
  assign new_n31658_ = ys__n26059 & new_n17846_;
  assign new_n31659_ = ys__n26059 & ~new_n27813_;
  assign new_n31660_ = ~new_n31658_ & ~new_n31659_;
  assign new_n31661_ = ~new_n31171_ & ~new_n31660_;
  assign new_n31662_ = ~new_n31657_ & ~new_n31661_;
  assign new_n31663_ = ys__n602 & ~new_n31662_;
  assign ys__n26657 = new_n31656_ | new_n31663_;
  assign new_n31665_ = ~ys__n778 & ys__n26059;
  assign new_n31666_ = ys__n26059 & new_n31160_;
  assign new_n31667_ = ys__n30941 & new_n27812_;
  assign new_n31668_ = ~ys__n18173 & ys__n18526;
  assign new_n31669_ = ys__n18173 & ys__n30929;
  assign new_n31670_ = ~new_n31668_ & ~new_n31669_;
  assign new_n31671_ = ~new_n17862_ & ~new_n31670_;
  assign new_n31672_ = ~new_n31667_ & ~new_n31671_;
  assign new_n31673_ = ~new_n31160_ & ~new_n31672_;
  assign new_n31674_ = ~new_n31666_ & ~new_n31673_;
  assign new_n31675_ = ys__n778 & ~new_n31674_;
  assign new_n31676_ = ~new_n31665_ & ~new_n31675_;
  assign new_n31677_ = ~ys__n602 & ~new_n31676_;
  assign new_n31678_ = new_n31171_ & ~new_n31676_;
  assign new_n31679_ = ys__n26062 & new_n17846_;
  assign new_n31680_ = ys__n26062 & ~new_n27813_;
  assign new_n31681_ = ~new_n31679_ & ~new_n31680_;
  assign new_n31682_ = ~new_n31171_ & ~new_n31681_;
  assign new_n31683_ = ~new_n31678_ & ~new_n31682_;
  assign new_n31684_ = ys__n602 & ~new_n31683_;
  assign ys__n26659 = new_n31677_ | new_n31684_;
  assign new_n31686_ = ~ys__n778 & ys__n26062;
  assign new_n31687_ = ys__n26062 & new_n31160_;
  assign new_n31688_ = ys__n202 & new_n27812_;
  assign new_n31689_ = ~ys__n18173 & ys__n18529;
  assign new_n31690_ = ys__n18173 & ys__n30931;
  assign new_n31691_ = ~new_n31689_ & ~new_n31690_;
  assign new_n31692_ = ~new_n17862_ & ~new_n31691_;
  assign new_n31693_ = ~new_n31688_ & ~new_n31692_;
  assign new_n31694_ = ~new_n31160_ & ~new_n31693_;
  assign new_n31695_ = ~new_n31687_ & ~new_n31694_;
  assign new_n31696_ = ys__n778 & ~new_n31695_;
  assign new_n31697_ = ~new_n31686_ & ~new_n31696_;
  assign new_n31698_ = ~ys__n602 & ~new_n31697_;
  assign new_n31699_ = new_n31171_ & ~new_n31697_;
  assign new_n31700_ = ys__n26065 & new_n17846_;
  assign new_n31701_ = ys__n26065 & ~new_n27813_;
  assign new_n31702_ = ~new_n31700_ & ~new_n31701_;
  assign new_n31703_ = ~new_n31171_ & ~new_n31702_;
  assign new_n31704_ = ~new_n31699_ & ~new_n31703_;
  assign new_n31705_ = ys__n602 & ~new_n31704_;
  assign ys__n26661 = new_n31698_ | new_n31705_;
  assign new_n31707_ = ~ys__n778 & ys__n26065;
  assign new_n31708_ = ys__n26065 & new_n31160_;
  assign new_n31709_ = ~ys__n18173 & ys__n18532;
  assign new_n31710_ = ys__n18173 & ys__n30933;
  assign new_n31711_ = ~new_n31709_ & ~new_n31710_;
  assign new_n31712_ = ~new_n17862_ & ~new_n31711_;
  assign new_n31713_ = ~new_n31160_ & new_n31712_;
  assign new_n31714_ = ~new_n31708_ & ~new_n31713_;
  assign new_n31715_ = ys__n778 & ~new_n31714_;
  assign new_n31716_ = ~new_n31707_ & ~new_n31715_;
  assign new_n31717_ = ~ys__n602 & ~new_n31716_;
  assign new_n31718_ = new_n31171_ & ~new_n31716_;
  assign new_n31719_ = ys__n26068 & new_n17846_;
  assign new_n31720_ = ys__n26068 & ~new_n27813_;
  assign new_n31721_ = ~new_n31719_ & ~new_n31720_;
  assign new_n31722_ = ~new_n31171_ & ~new_n31721_;
  assign new_n31723_ = ~new_n31718_ & ~new_n31722_;
  assign new_n31724_ = ys__n602 & ~new_n31723_;
  assign ys__n26663 = new_n31717_ | new_n31724_;
  assign new_n31726_ = ~ys__n778 & ys__n26068;
  assign new_n31727_ = ys__n26068 & new_n31160_;
  assign new_n31728_ = ~ys__n18173 & ys__n18535;
  assign new_n31729_ = ys__n18173 & ys__n30935;
  assign new_n31730_ = ~new_n31728_ & ~new_n31729_;
  assign new_n31731_ = ~new_n17862_ & ~new_n31730_;
  assign new_n31732_ = ~new_n31160_ & new_n31731_;
  assign new_n31733_ = ~new_n31727_ & ~new_n31732_;
  assign new_n31734_ = ys__n778 & ~new_n31733_;
  assign new_n31735_ = ~new_n31726_ & ~new_n31734_;
  assign new_n31736_ = ~ys__n602 & ~new_n31735_;
  assign new_n31737_ = new_n31171_ & ~new_n31735_;
  assign new_n31738_ = ys__n26071 & new_n17846_;
  assign new_n31739_ = ys__n26071 & ~new_n27813_;
  assign new_n31740_ = ~new_n31738_ & ~new_n31739_;
  assign new_n31741_ = ~new_n31171_ & ~new_n31740_;
  assign new_n31742_ = ~new_n31737_ & ~new_n31741_;
  assign new_n31743_ = ys__n602 & ~new_n31742_;
  assign ys__n26665 = new_n31736_ | new_n31743_;
  assign new_n31745_ = ~ys__n778 & ys__n26071;
  assign new_n31746_ = ys__n26071 & new_n31160_;
  assign new_n31747_ = ~ys__n18173 & ys__n18538;
  assign new_n31748_ = ys__n18173 & ys__n30937;
  assign new_n31749_ = ~new_n31747_ & ~new_n31748_;
  assign new_n31750_ = ~new_n17862_ & ~new_n31749_;
  assign new_n31751_ = ~new_n31160_ & new_n31750_;
  assign new_n31752_ = ~new_n31746_ & ~new_n31751_;
  assign new_n31753_ = ys__n778 & ~new_n31752_;
  assign new_n31754_ = ~new_n31745_ & ~new_n31753_;
  assign new_n31755_ = ~ys__n602 & ~new_n31754_;
  assign new_n31756_ = new_n31171_ & ~new_n31754_;
  assign new_n31757_ = ys__n26074 & new_n17846_;
  assign new_n31758_ = ys__n26074 & ~new_n27813_;
  assign new_n31759_ = ~new_n31757_ & ~new_n31758_;
  assign new_n31760_ = ~new_n31171_ & ~new_n31759_;
  assign new_n31761_ = ~new_n31756_ & ~new_n31760_;
  assign new_n31762_ = ys__n602 & ~new_n31761_;
  assign ys__n26667 = new_n31755_ | new_n31762_;
  assign new_n31764_ = ~ys__n778 & ys__n26074;
  assign new_n31765_ = ys__n26074 & new_n31160_;
  assign new_n31766_ = ~ys__n18173 & ys__n18541;
  assign new_n31767_ = ys__n18173 & ys__n30939;
  assign new_n31768_ = ~new_n31766_ & ~new_n31767_;
  assign new_n31769_ = ~new_n17862_ & ~new_n31768_;
  assign new_n31770_ = ~new_n31160_ & new_n31769_;
  assign new_n31771_ = ~new_n31765_ & ~new_n31770_;
  assign new_n31772_ = ys__n778 & ~new_n31771_;
  assign new_n31773_ = ~new_n31764_ & ~new_n31772_;
  assign new_n31774_ = ~ys__n602 & ~new_n31773_;
  assign new_n31775_ = new_n31171_ & ~new_n31773_;
  assign new_n31776_ = ys__n26359 & new_n17846_;
  assign new_n31777_ = ys__n25470 & ~new_n13462_;
  assign new_n31778_ = new_n27808_ & new_n31777_;
  assign new_n31779_ = new_n13459_ & new_n27801_;
  assign new_n31780_ = new_n31778_ & new_n31779_;
  assign new_n31781_ = ~new_n27813_ & new_n31780_;
  assign new_n31782_ = ~new_n31776_ & ~new_n31781_;
  assign new_n31783_ = ~new_n31171_ & ~new_n31782_;
  assign new_n31784_ = ~new_n31775_ & ~new_n31783_;
  assign new_n31785_ = ys__n602 & ~new_n31784_;
  assign ys__n26669 = new_n31774_ | new_n31785_;
  assign new_n31787_ = ~ys__n778 & ys__n26425;
  assign new_n31788_ = ys__n26425 & new_n17849_;
  assign new_n31789_ = ys__n26552 & ~new_n17849_;
  assign new_n31790_ = ~new_n31788_ & ~new_n31789_;
  assign new_n31791_ = ys__n778 & ~new_n31790_;
  assign new_n31792_ = ~new_n31787_ & ~new_n31791_;
  assign new_n31793_ = ~ys__n602 & ~new_n31792_;
  assign new_n31794_ = new_n17849_ & ~new_n31792_;
  assign new_n31795_ = ys__n26428 & new_n17846_;
  assign new_n31796_ = ys__n26428 & new_n17848_;
  assign new_n31797_ = ~new_n31795_ & ~new_n31796_;
  assign new_n31798_ = ~new_n17849_ & ~new_n31797_;
  assign new_n31799_ = ~new_n31794_ & ~new_n31798_;
  assign new_n31800_ = ys__n602 & ~new_n31799_;
  assign ys__n26671 = new_n31793_ | new_n31800_;
  assign new_n31802_ = ~ys__n778 & ys__n26428;
  assign new_n31803_ = ys__n26428 & new_n17849_;
  assign new_n31804_ = ys__n26553 & ~new_n17849_;
  assign new_n31805_ = ~new_n31803_ & ~new_n31804_;
  assign new_n31806_ = ys__n778 & ~new_n31805_;
  assign new_n31807_ = ~new_n31802_ & ~new_n31806_;
  assign new_n31808_ = ~ys__n602 & ~new_n31807_;
  assign new_n31809_ = new_n17849_ & ~new_n31807_;
  assign new_n31810_ = ys__n26431 & new_n17846_;
  assign new_n31811_ = ys__n26431 & new_n17848_;
  assign new_n31812_ = ~new_n31810_ & ~new_n31811_;
  assign new_n31813_ = ~new_n17849_ & ~new_n31812_;
  assign new_n31814_ = ~new_n31809_ & ~new_n31813_;
  assign new_n31815_ = ys__n602 & ~new_n31814_;
  assign ys__n26673 = new_n31808_ | new_n31815_;
  assign new_n31817_ = ~ys__n778 & ys__n26431;
  assign new_n31818_ = ys__n26431 & new_n17849_;
  assign new_n31819_ = ys__n26554 & ~new_n17849_;
  assign new_n31820_ = ~new_n31818_ & ~new_n31819_;
  assign new_n31821_ = ys__n778 & ~new_n31820_;
  assign new_n31822_ = ~new_n31817_ & ~new_n31821_;
  assign new_n31823_ = ~ys__n602 & ~new_n31822_;
  assign new_n31824_ = new_n17849_ & ~new_n31822_;
  assign new_n31825_ = ys__n26434 & new_n17846_;
  assign new_n31826_ = ys__n26434 & new_n17848_;
  assign new_n31827_ = ~new_n31825_ & ~new_n31826_;
  assign new_n31828_ = ~new_n17849_ & ~new_n31827_;
  assign new_n31829_ = ~new_n31824_ & ~new_n31828_;
  assign new_n31830_ = ys__n602 & ~new_n31829_;
  assign ys__n26675 = new_n31823_ | new_n31830_;
  assign new_n31832_ = ~ys__n778 & ys__n26434;
  assign new_n31833_ = ys__n26434 & new_n17849_;
  assign new_n31834_ = ys__n26555 & ~new_n17849_;
  assign new_n31835_ = ~new_n31833_ & ~new_n31834_;
  assign new_n31836_ = ys__n778 & ~new_n31835_;
  assign new_n31837_ = ~new_n31832_ & ~new_n31836_;
  assign new_n31838_ = ~ys__n602 & ~new_n31837_;
  assign new_n31839_ = new_n17849_ & ~new_n31837_;
  assign new_n31840_ = ys__n26437 & new_n17846_;
  assign new_n31841_ = ys__n26437 & new_n17848_;
  assign new_n31842_ = ~new_n31840_ & ~new_n31841_;
  assign new_n31843_ = ~new_n17849_ & ~new_n31842_;
  assign new_n31844_ = ~new_n31839_ & ~new_n31843_;
  assign new_n31845_ = ys__n602 & ~new_n31844_;
  assign ys__n26677 = new_n31838_ | new_n31845_;
  assign new_n31847_ = ~ys__n778 & ys__n26437;
  assign new_n31848_ = ys__n26437 & new_n17849_;
  assign new_n31849_ = ys__n26279 & ~new_n17849_;
  assign new_n31850_ = ~new_n31848_ & ~new_n31849_;
  assign new_n31851_ = ys__n778 & ~new_n31850_;
  assign new_n31852_ = ~new_n31847_ & ~new_n31851_;
  assign new_n31853_ = ~ys__n602 & ~new_n31852_;
  assign new_n31854_ = new_n17849_ & ~new_n31852_;
  assign new_n31855_ = ys__n26440 & new_n17846_;
  assign new_n31856_ = ys__n26440 & new_n17848_;
  assign new_n31857_ = ~new_n31855_ & ~new_n31856_;
  assign new_n31858_ = ~new_n17849_ & ~new_n31857_;
  assign new_n31859_ = ~new_n31854_ & ~new_n31858_;
  assign new_n31860_ = ys__n602 & ~new_n31859_;
  assign ys__n26679 = new_n31853_ | new_n31860_;
  assign new_n31862_ = ~ys__n778 & ys__n26440;
  assign new_n31863_ = ys__n26440 & new_n17849_;
  assign new_n31864_ = ys__n26556 & ~new_n17849_;
  assign new_n31865_ = ~new_n31863_ & ~new_n31864_;
  assign new_n31866_ = ys__n778 & ~new_n31865_;
  assign new_n31867_ = ~new_n31862_ & ~new_n31866_;
  assign new_n31868_ = ~ys__n602 & ~new_n31867_;
  assign new_n31869_ = new_n17849_ & ~new_n31867_;
  assign new_n31870_ = ys__n26443 & new_n17846_;
  assign new_n31871_ = ys__n26443 & new_n17848_;
  assign new_n31872_ = ~new_n31870_ & ~new_n31871_;
  assign new_n31873_ = ~new_n17849_ & ~new_n31872_;
  assign new_n31874_ = ~new_n31869_ & ~new_n31873_;
  assign new_n31875_ = ys__n602 & ~new_n31874_;
  assign ys__n26681 = new_n31868_ | new_n31875_;
  assign new_n31877_ = ~ys__n778 & ys__n26443;
  assign new_n31878_ = ys__n778 & ys__n26443;
  assign new_n31879_ = new_n17849_ & new_n31878_;
  assign new_n31880_ = ~new_n31877_ & ~new_n31879_;
  assign new_n31881_ = ~ys__n602 & ~new_n31880_;
  assign new_n31882_ = new_n17849_ & ~new_n31880_;
  assign new_n31883_ = ys__n26446 & new_n17846_;
  assign new_n31884_ = ys__n26446 & new_n17848_;
  assign new_n31885_ = ~new_n31883_ & ~new_n31884_;
  assign new_n31886_ = ~new_n17849_ & ~new_n31885_;
  assign new_n31887_ = ~new_n31882_ & ~new_n31886_;
  assign new_n31888_ = ys__n602 & ~new_n31887_;
  assign ys__n26683 = new_n31881_ | new_n31888_;
  assign new_n31890_ = ~ys__n778 & ys__n26446;
  assign new_n31891_ = ys__n26446 & new_n17849_;
  assign new_n31892_ = ys__n26557 & ~new_n17849_;
  assign new_n31893_ = ~new_n31891_ & ~new_n31892_;
  assign new_n31894_ = ys__n778 & ~new_n31893_;
  assign new_n31895_ = ~new_n31890_ & ~new_n31894_;
  assign new_n31896_ = ~ys__n602 & ~new_n31895_;
  assign new_n31897_ = new_n17849_ & ~new_n31895_;
  assign new_n31898_ = ys__n26449 & new_n17846_;
  assign new_n31899_ = ys__n26449 & new_n17848_;
  assign new_n31900_ = ~new_n31898_ & ~new_n31899_;
  assign new_n31901_ = ~new_n17849_ & ~new_n31900_;
  assign new_n31902_ = ~new_n31897_ & ~new_n31901_;
  assign new_n31903_ = ys__n602 & ~new_n31902_;
  assign ys__n26685 = new_n31896_ | new_n31903_;
  assign new_n31905_ = ~ys__n778 & ys__n26449;
  assign new_n31906_ = ys__n26449 & new_n17849_;
  assign new_n31907_ = ys__n26558 & ~new_n17849_;
  assign new_n31908_ = ~new_n31906_ & ~new_n31907_;
  assign new_n31909_ = ys__n778 & ~new_n31908_;
  assign new_n31910_ = ~new_n31905_ & ~new_n31909_;
  assign new_n31911_ = ~ys__n602 & ~new_n31910_;
  assign new_n31912_ = new_n17849_ & ~new_n31910_;
  assign new_n31913_ = ys__n26452 & new_n17846_;
  assign new_n31914_ = ys__n26452 & new_n17848_;
  assign new_n31915_ = ~new_n31913_ & ~new_n31914_;
  assign new_n31916_ = ~new_n17849_ & ~new_n31915_;
  assign new_n31917_ = ~new_n31912_ & ~new_n31916_;
  assign new_n31918_ = ys__n602 & ~new_n31917_;
  assign ys__n26687 = new_n31911_ | new_n31918_;
  assign new_n31920_ = ~ys__n778 & ys__n26452;
  assign new_n31921_ = ys__n26452 & new_n17849_;
  assign new_n31922_ = ys__n26559 & ~new_n17849_;
  assign new_n31923_ = ~new_n31921_ & ~new_n31922_;
  assign new_n31924_ = ys__n778 & ~new_n31923_;
  assign new_n31925_ = ~new_n31920_ & ~new_n31924_;
  assign new_n31926_ = ~ys__n602 & ~new_n31925_;
  assign new_n31927_ = new_n17849_ & ~new_n31925_;
  assign new_n31928_ = ys__n26455 & new_n17846_;
  assign new_n31929_ = ys__n26455 & new_n17848_;
  assign new_n31930_ = ~new_n31928_ & ~new_n31929_;
  assign new_n31931_ = ~new_n17849_ & ~new_n31930_;
  assign new_n31932_ = ~new_n31927_ & ~new_n31931_;
  assign new_n31933_ = ys__n602 & ~new_n31932_;
  assign ys__n26689 = new_n31926_ | new_n31933_;
  assign new_n31935_ = ~ys__n778 & ys__n26455;
  assign new_n31936_ = ys__n778 & ys__n26455;
  assign new_n31937_ = new_n17849_ & new_n31936_;
  assign new_n31938_ = ~new_n31935_ & ~new_n31937_;
  assign new_n31939_ = ~ys__n602 & ~new_n31938_;
  assign new_n31940_ = new_n17849_ & ~new_n31938_;
  assign new_n31941_ = ys__n26285 & new_n17846_;
  assign new_n31942_ = ys__n26285 & new_n17848_;
  assign new_n31943_ = ~new_n31941_ & ~new_n31942_;
  assign new_n31944_ = ~new_n17849_ & ~new_n31943_;
  assign new_n31945_ = ~new_n31940_ & ~new_n31944_;
  assign new_n31946_ = ys__n602 & ~new_n31945_;
  assign ys__n26691 = new_n31939_ | new_n31946_;
  assign new_n31948_ = ~ys__n778 & ys__n26285;
  assign new_n31949_ = ys__n26285 & new_n17849_;
  assign new_n31950_ = ys__n26560 & ~new_n17849_;
  assign new_n31951_ = ~new_n31949_ & ~new_n31950_;
  assign new_n31952_ = ys__n778 & ~new_n31951_;
  assign new_n31953_ = ~new_n31948_ & ~new_n31952_;
  assign new_n31954_ = ~ys__n602 & ~new_n31953_;
  assign new_n31955_ = new_n17849_ & ~new_n31953_;
  assign new_n31956_ = ys__n26460 & new_n17846_;
  assign new_n31957_ = ys__n26460 & new_n17848_;
  assign new_n31958_ = ~new_n31956_ & ~new_n31957_;
  assign new_n31959_ = ~new_n17849_ & ~new_n31958_;
  assign new_n31960_ = ~new_n31955_ & ~new_n31959_;
  assign new_n31961_ = ys__n602 & ~new_n31960_;
  assign ys__n26693 = new_n31954_ | new_n31961_;
  assign new_n31963_ = ~ys__n778 & ys__n26460;
  assign new_n31964_ = ys__n26460 & new_n17849_;
  assign new_n31965_ = ys__n26561 & ~new_n17849_;
  assign new_n31966_ = ~new_n31964_ & ~new_n31965_;
  assign new_n31967_ = ys__n778 & ~new_n31966_;
  assign new_n31968_ = ~new_n31963_ & ~new_n31967_;
  assign new_n31969_ = ~ys__n602 & ~new_n31968_;
  assign new_n31970_ = new_n17849_ & ~new_n31968_;
  assign new_n31971_ = ys__n26463 & new_n17846_;
  assign new_n31972_ = ys__n26463 & new_n17848_;
  assign new_n31973_ = ~new_n31971_ & ~new_n31972_;
  assign new_n31974_ = ~new_n17849_ & ~new_n31973_;
  assign new_n31975_ = ~new_n31970_ & ~new_n31974_;
  assign new_n31976_ = ys__n602 & ~new_n31975_;
  assign ys__n26695 = new_n31969_ | new_n31976_;
  assign new_n31978_ = ~ys__n778 & ys__n26463;
  assign new_n31979_ = ys__n778 & ys__n26463;
  assign new_n31980_ = new_n17849_ & new_n31979_;
  assign new_n31981_ = ~new_n31978_ & ~new_n31980_;
  assign new_n31982_ = ~ys__n602 & ~new_n31981_;
  assign new_n31983_ = new_n17849_ & ~new_n31981_;
  assign new_n31984_ = ys__n26466 & new_n17846_;
  assign new_n31985_ = ys__n26466 & new_n17848_;
  assign new_n31986_ = ~new_n31984_ & ~new_n31985_;
  assign new_n31987_ = ~new_n17849_ & ~new_n31986_;
  assign new_n31988_ = ~new_n31983_ & ~new_n31987_;
  assign new_n31989_ = ys__n602 & ~new_n31988_;
  assign ys__n26697 = new_n31982_ | new_n31989_;
  assign new_n31991_ = ~ys__n778 & ys__n26466;
  assign new_n31992_ = ys__n26466 & new_n17849_;
  assign new_n31993_ = ys__n26562 & ~new_n17849_;
  assign new_n31994_ = ~new_n31992_ & ~new_n31993_;
  assign new_n31995_ = ys__n778 & ~new_n31994_;
  assign new_n31996_ = ~new_n31991_ & ~new_n31995_;
  assign new_n31997_ = ~ys__n602 & ~new_n31996_;
  assign new_n31998_ = new_n17849_ & ~new_n31996_;
  assign new_n31999_ = ys__n26469 & new_n17846_;
  assign new_n32000_ = ys__n26469 & new_n17848_;
  assign new_n32001_ = ~new_n31999_ & ~new_n32000_;
  assign new_n32002_ = ~new_n17849_ & ~new_n32001_;
  assign new_n32003_ = ~new_n31998_ & ~new_n32002_;
  assign new_n32004_ = ys__n602 & ~new_n32003_;
  assign ys__n26699 = new_n31997_ | new_n32004_;
  assign new_n32006_ = ~ys__n778 & ys__n26469;
  assign new_n32007_ = ys__n26469 & new_n17849_;
  assign new_n32008_ = ys__n26563 & ~new_n17849_;
  assign new_n32009_ = ~new_n32007_ & ~new_n32008_;
  assign new_n32010_ = ys__n778 & ~new_n32009_;
  assign new_n32011_ = ~new_n32006_ & ~new_n32010_;
  assign new_n32012_ = ~ys__n602 & ~new_n32011_;
  assign new_n32013_ = new_n17849_ & ~new_n32011_;
  assign new_n32014_ = ys__n26472 & new_n17846_;
  assign new_n32015_ = ys__n26472 & new_n17848_;
  assign new_n32016_ = ~new_n32014_ & ~new_n32015_;
  assign new_n32017_ = ~new_n17849_ & ~new_n32016_;
  assign new_n32018_ = ~new_n32013_ & ~new_n32017_;
  assign new_n32019_ = ys__n602 & ~new_n32018_;
  assign ys__n26701 = new_n32012_ | new_n32019_;
  assign new_n32021_ = ~ys__n778 & ys__n26472;
  assign new_n32022_ = ys__n26472 & new_n17849_;
  assign new_n32023_ = ys__n26564 & ~new_n17849_;
  assign new_n32024_ = ~new_n32022_ & ~new_n32023_;
  assign new_n32025_ = ys__n778 & ~new_n32024_;
  assign new_n32026_ = ~new_n32021_ & ~new_n32025_;
  assign new_n32027_ = ~ys__n602 & ~new_n32026_;
  assign new_n32028_ = new_n17849_ & ~new_n32026_;
  assign new_n32029_ = ys__n26475 & new_n17846_;
  assign new_n32030_ = ys__n26475 & new_n17848_;
  assign new_n32031_ = ~new_n32029_ & ~new_n32030_;
  assign new_n32032_ = ~new_n17849_ & ~new_n32031_;
  assign new_n32033_ = ~new_n32028_ & ~new_n32032_;
  assign new_n32034_ = ys__n602 & ~new_n32033_;
  assign ys__n26703 = new_n32027_ | new_n32034_;
  assign new_n32036_ = ~ys__n778 & ys__n26475;
  assign new_n32037_ = ys__n26475 & new_n17849_;
  assign new_n32038_ = ys__n18173 & ~new_n17849_;
  assign new_n32039_ = ~new_n32037_ & ~new_n32038_;
  assign new_n32040_ = ys__n778 & ~new_n32039_;
  assign new_n32041_ = ~new_n32036_ & ~new_n32040_;
  assign new_n32042_ = ~ys__n602 & ~new_n32041_;
  assign new_n32043_ = new_n17849_ & ~new_n32041_;
  assign new_n32044_ = ys__n26478 & new_n17846_;
  assign new_n32045_ = ys__n26478 & new_n17848_;
  assign new_n32046_ = ~new_n32044_ & ~new_n32045_;
  assign new_n32047_ = ~new_n17849_ & ~new_n32046_;
  assign new_n32048_ = ~new_n32043_ & ~new_n32047_;
  assign new_n32049_ = ys__n602 & ~new_n32048_;
  assign ys__n26705 = new_n32042_ | new_n32049_;
  assign new_n32051_ = ~ys__n778 & ys__n26478;
  assign new_n32052_ = ys__n26478 & new_n17849_;
  assign new_n32053_ = ys__n26565 & ~new_n17849_;
  assign new_n32054_ = ~new_n32052_ & ~new_n32053_;
  assign new_n32055_ = ys__n778 & ~new_n32054_;
  assign new_n32056_ = ~new_n32051_ & ~new_n32055_;
  assign new_n32057_ = ~ys__n602 & ~new_n32056_;
  assign new_n32058_ = new_n17849_ & ~new_n32056_;
  assign new_n32059_ = ys__n26481 & new_n17846_;
  assign new_n32060_ = ys__n26481 & new_n17848_;
  assign new_n32061_ = ~new_n32059_ & ~new_n32060_;
  assign new_n32062_ = ~new_n17849_ & ~new_n32061_;
  assign new_n32063_ = ~new_n32058_ & ~new_n32062_;
  assign new_n32064_ = ys__n602 & ~new_n32063_;
  assign ys__n26707 = new_n32057_ | new_n32064_;
  assign new_n32066_ = ~ys__n778 & ys__n26481;
  assign new_n32067_ = ys__n26481 & new_n17849_;
  assign new_n32068_ = ~new_n17849_ & ys__n26566;
  assign new_n32069_ = ~new_n32067_ & ~new_n32068_;
  assign new_n32070_ = ys__n778 & ~new_n32069_;
  assign new_n32071_ = ~new_n32066_ & ~new_n32070_;
  assign new_n32072_ = ~ys__n602 & ~new_n32071_;
  assign new_n32073_ = new_n17849_ & ~new_n32071_;
  assign new_n32074_ = ys__n26484 & new_n17846_;
  assign new_n32075_ = ys__n26484 & new_n17848_;
  assign new_n32076_ = ~new_n32074_ & ~new_n32075_;
  assign new_n32077_ = ~new_n17849_ & ~new_n32076_;
  assign new_n32078_ = ~new_n32073_ & ~new_n32077_;
  assign new_n32079_ = ys__n602 & ~new_n32078_;
  assign ys__n26709 = new_n32072_ | new_n32079_;
  assign new_n32081_ = ~ys__n778 & ys__n26484;
  assign new_n32082_ = ys__n26484 & new_n17849_;
  assign new_n32083_ = ys__n26567 & ~new_n17849_;
  assign new_n32084_ = ~new_n32082_ & ~new_n32083_;
  assign new_n32085_ = ys__n778 & ~new_n32084_;
  assign new_n32086_ = ~new_n32081_ & ~new_n32085_;
  assign new_n32087_ = ~ys__n602 & ~new_n32086_;
  assign new_n32088_ = new_n17849_ & ~new_n32086_;
  assign new_n32089_ = ys__n26487 & new_n17846_;
  assign new_n32090_ = ys__n26487 & new_n17848_;
  assign new_n32091_ = ~new_n32089_ & ~new_n32090_;
  assign new_n32092_ = ~new_n17849_ & ~new_n32091_;
  assign new_n32093_ = ~new_n32088_ & ~new_n32092_;
  assign new_n32094_ = ys__n602 & ~new_n32093_;
  assign ys__n26711 = new_n32087_ | new_n32094_;
  assign new_n32096_ = ~ys__n778 & ys__n26487;
  assign new_n32097_ = ys__n26487 & new_n17849_;
  assign new_n32098_ = new_n17849_ & ~new_n32097_;
  assign new_n32099_ = ys__n778 & ~new_n32098_;
  assign new_n32100_ = ~new_n32096_ & ~new_n32099_;
  assign new_n32101_ = ~ys__n602 & ~new_n32100_;
  assign new_n32102_ = new_n17849_ & ~new_n32100_;
  assign new_n32103_ = ys__n26490 & new_n17846_;
  assign new_n32104_ = ys__n26490 & new_n17848_;
  assign new_n32105_ = ~new_n32103_ & ~new_n32104_;
  assign new_n32106_ = ~new_n17849_ & ~new_n32105_;
  assign new_n32107_ = ~new_n32102_ & ~new_n32106_;
  assign new_n32108_ = ys__n602 & ~new_n32107_;
  assign ys__n26713 = new_n32101_ | new_n32108_;
  assign new_n32110_ = ~ys__n778 & ys__n26490;
  assign new_n32111_ = ys__n26490 & new_n17849_;
  assign new_n32112_ = ys__n26568 & ~new_n17849_;
  assign new_n32113_ = ~new_n32111_ & ~new_n32112_;
  assign new_n32114_ = ys__n778 & ~new_n32113_;
  assign new_n32115_ = ~new_n32110_ & ~new_n32114_;
  assign new_n32116_ = ~ys__n602 & ~new_n32115_;
  assign new_n32117_ = new_n17849_ & ~new_n32115_;
  assign new_n32118_ = ys__n26493 & new_n17846_;
  assign new_n32119_ = ys__n26493 & new_n17848_;
  assign new_n32120_ = ~new_n32118_ & ~new_n32119_;
  assign new_n32121_ = ~new_n17849_ & ~new_n32120_;
  assign new_n32122_ = ~new_n32117_ & ~new_n32121_;
  assign new_n32123_ = ys__n602 & ~new_n32122_;
  assign ys__n26715 = new_n32116_ | new_n32123_;
  assign new_n32125_ = ~ys__n778 & ys__n26493;
  assign new_n32126_ = ys__n26493 & new_n17849_;
  assign new_n32127_ = ys__n26569 & ~new_n17849_;
  assign new_n32128_ = ~new_n32126_ & ~new_n32127_;
  assign new_n32129_ = ys__n778 & ~new_n32128_;
  assign new_n32130_ = ~new_n32125_ & ~new_n32129_;
  assign new_n32131_ = ~ys__n602 & ~new_n32130_;
  assign new_n32132_ = new_n17849_ & ~new_n32130_;
  assign new_n32133_ = ys__n26496 & new_n17846_;
  assign new_n32134_ = ys__n26496 & new_n17848_;
  assign new_n32135_ = ~new_n32133_ & ~new_n32134_;
  assign new_n32136_ = ~new_n17849_ & ~new_n32135_;
  assign new_n32137_ = ~new_n32132_ & ~new_n32136_;
  assign new_n32138_ = ys__n602 & ~new_n32137_;
  assign ys__n26717 = new_n32131_ | new_n32138_;
  assign new_n32140_ = ~ys__n778 & ys__n26496;
  assign new_n32141_ = ys__n26496 & new_n17849_;
  assign new_n32142_ = ys__n26570 & ~new_n17849_;
  assign new_n32143_ = ~new_n32141_ & ~new_n32142_;
  assign new_n32144_ = ys__n778 & ~new_n32143_;
  assign new_n32145_ = ~new_n32140_ & ~new_n32144_;
  assign new_n32146_ = ~ys__n602 & ~new_n32145_;
  assign new_n32147_ = new_n17849_ & ~new_n32145_;
  assign new_n32148_ = ys__n26499 & new_n17846_;
  assign new_n32149_ = ys__n26499 & new_n17848_;
  assign new_n32150_ = ~new_n32148_ & ~new_n32149_;
  assign new_n32151_ = ~new_n17849_ & ~new_n32150_;
  assign new_n32152_ = ~new_n32147_ & ~new_n32151_;
  assign new_n32153_ = ys__n602 & ~new_n32152_;
  assign ys__n26719 = new_n32146_ | new_n32153_;
  assign new_n32155_ = ~ys__n778 & ys__n26499;
  assign new_n32156_ = ys__n26499 & new_n17849_;
  assign new_n32157_ = ys__n26571 & ~new_n17849_;
  assign new_n32158_ = ~new_n32156_ & ~new_n32157_;
  assign new_n32159_ = ys__n778 & ~new_n32158_;
  assign new_n32160_ = ~new_n32155_ & ~new_n32159_;
  assign new_n32161_ = ~ys__n602 & ~new_n32160_;
  assign new_n32162_ = new_n17849_ & ~new_n32160_;
  assign new_n32163_ = ys__n26502 & new_n17846_;
  assign new_n32164_ = ys__n26502 & new_n17848_;
  assign new_n32165_ = ~new_n32163_ & ~new_n32164_;
  assign new_n32166_ = ~new_n17849_ & ~new_n32165_;
  assign new_n32167_ = ~new_n32162_ & ~new_n32166_;
  assign new_n32168_ = ys__n602 & ~new_n32167_;
  assign ys__n26721 = new_n32161_ | new_n32168_;
  assign new_n32170_ = ~ys__n778 & ys__n26502;
  assign new_n32171_ = ys__n778 & ys__n26502;
  assign new_n32172_ = new_n17849_ & new_n32171_;
  assign new_n32173_ = ~new_n32170_ & ~new_n32172_;
  assign new_n32174_ = ~ys__n602 & ~new_n32173_;
  assign new_n32175_ = new_n17849_ & ~new_n32173_;
  assign new_n32176_ = ys__n26505 & new_n17846_;
  assign new_n32177_ = ys__n26505 & new_n17848_;
  assign new_n32178_ = ~new_n32176_ & ~new_n32177_;
  assign new_n32179_ = ~new_n17849_ & ~new_n32178_;
  assign new_n32180_ = ~new_n32175_ & ~new_n32179_;
  assign new_n32181_ = ys__n602 & ~new_n32180_;
  assign ys__n26723 = new_n32174_ | new_n32181_;
  assign new_n32183_ = ~ys__n778 & ys__n26505;
  assign new_n32184_ = ys__n778 & ys__n26505;
  assign new_n32185_ = new_n17849_ & new_n32184_;
  assign new_n32186_ = ~new_n32183_ & ~new_n32185_;
  assign new_n32187_ = ~ys__n602 & ~new_n32186_;
  assign new_n32188_ = new_n17849_ & ~new_n32186_;
  assign new_n32189_ = ys__n26508 & new_n17846_;
  assign new_n32190_ = ys__n26508 & new_n17848_;
  assign new_n32191_ = ~new_n32189_ & ~new_n32190_;
  assign new_n32192_ = ~new_n17849_ & ~new_n32191_;
  assign new_n32193_ = ~new_n32188_ & ~new_n32192_;
  assign new_n32194_ = ys__n602 & ~new_n32193_;
  assign ys__n26725 = new_n32187_ | new_n32194_;
  assign new_n32196_ = ~ys__n778 & ys__n26508;
  assign new_n32197_ = ys__n778 & ys__n26508;
  assign new_n32198_ = new_n17849_ & new_n32197_;
  assign new_n32199_ = ~new_n32196_ & ~new_n32198_;
  assign new_n32200_ = ~ys__n602 & ~new_n32199_;
  assign new_n32201_ = new_n17849_ & ~new_n32199_;
  assign new_n32202_ = ys__n26511 & new_n17846_;
  assign new_n32203_ = ys__n26511 & new_n17848_;
  assign new_n32204_ = ~new_n32202_ & ~new_n32203_;
  assign new_n32205_ = ~new_n17849_ & ~new_n32204_;
  assign new_n32206_ = ~new_n32201_ & ~new_n32205_;
  assign new_n32207_ = ys__n602 & ~new_n32206_;
  assign ys__n26727 = new_n32200_ | new_n32207_;
  assign new_n32209_ = ~ys__n778 & ys__n26511;
  assign new_n32210_ = ys__n778 & ys__n26511;
  assign new_n32211_ = new_n17849_ & new_n32210_;
  assign new_n32212_ = ~new_n32209_ & ~new_n32211_;
  assign new_n32213_ = ~ys__n602 & ~new_n32212_;
  assign new_n32214_ = new_n17849_ & ~new_n32212_;
  assign new_n32215_ = ys__n26514 & new_n17846_;
  assign new_n32216_ = ys__n26514 & new_n17848_;
  assign new_n32217_ = ~new_n32215_ & ~new_n32216_;
  assign new_n32218_ = ~new_n17849_ & ~new_n32217_;
  assign new_n32219_ = ~new_n32214_ & ~new_n32218_;
  assign new_n32220_ = ys__n602 & ~new_n32219_;
  assign ys__n26729 = new_n32213_ | new_n32220_;
  assign new_n32222_ = ~ys__n778 & ys__n26514;
  assign new_n32223_ = ys__n778 & ys__n26514;
  assign new_n32224_ = new_n17849_ & new_n32223_;
  assign new_n32225_ = ~new_n32222_ & ~new_n32224_;
  assign new_n32226_ = ~ys__n602 & ~new_n32225_;
  assign new_n32227_ = new_n17849_ & ~new_n32225_;
  assign new_n32228_ = ys__n26517 & new_n17846_;
  assign new_n32229_ = ys__n26517 & new_n17848_;
  assign new_n32230_ = ~new_n32228_ & ~new_n32229_;
  assign new_n32231_ = ~new_n17849_ & ~new_n32230_;
  assign new_n32232_ = ~new_n32227_ & ~new_n32231_;
  assign new_n32233_ = ys__n602 & ~new_n32232_;
  assign ys__n26731 = new_n32226_ | new_n32233_;
  assign new_n32235_ = ~ys__n778 & ys__n26517;
  assign new_n32236_ = ys__n26517 & new_n17849_;
  assign new_n32237_ = ys__n26572 & ~new_n17849_;
  assign new_n32238_ = ~new_n32236_ & ~new_n32237_;
  assign new_n32239_ = ys__n778 & ~new_n32238_;
  assign new_n32240_ = ~new_n32235_ & ~new_n32239_;
  assign new_n32241_ = ~ys__n602 & ~new_n32240_;
  assign new_n32242_ = new_n17849_ & ~new_n32240_;
  assign new_n32243_ = ys__n25980 & new_n17846_;
  assign new_n32244_ = new_n17848_ & new_n31780_;
  assign new_n32245_ = ~new_n32243_ & ~new_n32244_;
  assign new_n32246_ = ~new_n17849_ & ~new_n32245_;
  assign new_n32247_ = ~new_n32242_ & ~new_n32246_;
  assign new_n32248_ = ys__n602 & ~new_n32247_;
  assign ys__n26733 = new_n32241_ | new_n32248_;
  assign new_n32250_ = ~ys__n778 & ys__n26359;
  assign new_n32251_ = ys__n26359 & new_n17857_;
  assign new_n32252_ = ys__n6112 & ~ys__n18173;
  assign new_n32253_ = ys__n18173 & ys__n18829;
  assign new_n32254_ = ~new_n32252_ & ~new_n32253_;
  assign new_n32255_ = ~new_n17857_ & ~new_n32254_;
  assign new_n32256_ = ~new_n32251_ & ~new_n32255_;
  assign new_n32257_ = ys__n778 & ~new_n32256_;
  assign new_n32258_ = ~new_n32250_ & ~new_n32257_;
  assign new_n32259_ = ~ys__n602 & ~new_n32258_;
  assign new_n32260_ = new_n17857_ & ~new_n32258_;
  assign new_n32261_ = ys__n26362 & ~new_n17857_;
  assign new_n32262_ = ~new_n32260_ & ~new_n32261_;
  assign new_n32263_ = ys__n602 & ~new_n32262_;
  assign ys__n26734 = new_n32259_ | new_n32263_;
  assign new_n32265_ = ~ys__n778 & ys__n26362;
  assign new_n32266_ = ys__n26362 & new_n17857_;
  assign new_n32267_ = ys__n6113 & ~ys__n18173;
  assign new_n32268_ = ys__n18173 & ys__n18831;
  assign new_n32269_ = ~new_n32267_ & ~new_n32268_;
  assign new_n32270_ = ~new_n17857_ & ~new_n32269_;
  assign new_n32271_ = ~new_n32266_ & ~new_n32270_;
  assign new_n32272_ = ys__n778 & ~new_n32271_;
  assign new_n32273_ = ~new_n32265_ & ~new_n32272_;
  assign new_n32274_ = ~ys__n602 & ~new_n32273_;
  assign new_n32275_ = new_n17857_ & ~new_n32273_;
  assign new_n32276_ = ys__n26161 & ~new_n17857_;
  assign new_n32277_ = ~new_n32275_ & ~new_n32276_;
  assign new_n32278_ = ys__n602 & ~new_n32277_;
  assign ys__n26735 = new_n32274_ | new_n32278_;
  assign new_n32280_ = ~ys__n778 & ys__n26161;
  assign new_n32281_ = ys__n26161 & new_n17857_;
  assign new_n32282_ = ys__n172 & ~ys__n18173;
  assign new_n32283_ = ys__n18173 & ys__n18833;
  assign new_n32284_ = ~new_n32282_ & ~new_n32283_;
  assign new_n32285_ = ~new_n17857_ & ~new_n32284_;
  assign new_n32286_ = ~new_n32281_ & ~new_n32285_;
  assign new_n32287_ = ys__n778 & ~new_n32286_;
  assign new_n32288_ = ~new_n32280_ & ~new_n32287_;
  assign new_n32289_ = ~ys__n602 & ~new_n32288_;
  assign new_n32290_ = new_n17857_ & ~new_n32288_;
  assign new_n32291_ = ys__n26162 & ~new_n17857_;
  assign new_n32292_ = ~new_n32290_ & ~new_n32291_;
  assign new_n32293_ = ys__n602 & ~new_n32292_;
  assign ys__n26736 = new_n32289_ | new_n32293_;
  assign new_n32295_ = ~ys__n778 & ys__n26162;
  assign new_n32296_ = ys__n26162 & new_n17857_;
  assign new_n32297_ = ys__n338 & ~ys__n18173;
  assign new_n32298_ = ys__n18173 & ys__n18835;
  assign new_n32299_ = ~new_n32297_ & ~new_n32298_;
  assign new_n32300_ = ~new_n17857_ & ~new_n32299_;
  assign new_n32301_ = ~new_n32296_ & ~new_n32300_;
  assign new_n32302_ = ys__n778 & ~new_n32301_;
  assign new_n32303_ = ~new_n32295_ & ~new_n32302_;
  assign new_n32304_ = ~ys__n602 & ~new_n32303_;
  assign new_n32305_ = new_n17857_ & ~new_n32303_;
  assign new_n32306_ = ys__n26164 & ~new_n17857_;
  assign new_n32307_ = ~new_n32305_ & ~new_n32306_;
  assign new_n32308_ = ys__n602 & ~new_n32307_;
  assign ys__n26737 = new_n32304_ | new_n32308_;
  assign new_n32310_ = ~ys__n778 & ys__n26164;
  assign new_n32311_ = ys__n26164 & new_n17857_;
  assign new_n32312_ = ys__n22 & ~ys__n18173;
  assign new_n32313_ = ys__n18173 & ys__n18837;
  assign new_n32314_ = ~new_n32312_ & ~new_n32313_;
  assign new_n32315_ = ~new_n17857_ & ~new_n32314_;
  assign new_n32316_ = ~new_n32311_ & ~new_n32315_;
  assign new_n32317_ = ys__n778 & ~new_n32316_;
  assign new_n32318_ = ~new_n32310_ & ~new_n32317_;
  assign new_n32319_ = ~ys__n602 & ~new_n32318_;
  assign new_n32320_ = new_n17857_ & ~new_n32318_;
  assign new_n32321_ = ys__n26166 & ~new_n17857_;
  assign new_n32322_ = ~new_n32320_ & ~new_n32321_;
  assign new_n32323_ = ys__n602 & ~new_n32322_;
  assign ys__n26738 = new_n32319_ | new_n32323_;
  assign new_n32325_ = ~ys__n778 & ys__n26166;
  assign new_n32326_ = ys__n26166 & new_n17857_;
  assign new_n32327_ = ys__n316 & ~ys__n18173;
  assign new_n32328_ = ys__n18173 & ys__n18839;
  assign new_n32329_ = ~new_n32327_ & ~new_n32328_;
  assign new_n32330_ = ~new_n17857_ & ~new_n32329_;
  assign new_n32331_ = ~new_n32326_ & ~new_n32330_;
  assign new_n32332_ = ys__n778 & ~new_n32331_;
  assign new_n32333_ = ~new_n32325_ & ~new_n32332_;
  assign new_n32334_ = ~ys__n602 & ~new_n32333_;
  assign new_n32335_ = new_n17857_ & ~new_n32333_;
  assign new_n32336_ = ys__n26168 & ~new_n17857_;
  assign new_n32337_ = ~new_n32335_ & ~new_n32336_;
  assign new_n32338_ = ys__n602 & ~new_n32337_;
  assign ys__n26739 = new_n32334_ | new_n32338_;
  assign new_n32340_ = ~ys__n778 & ys__n26168;
  assign new_n32341_ = ys__n26168 & new_n17857_;
  assign new_n32342_ = ys__n6115 & ~ys__n18173;
  assign new_n32343_ = ys__n18173 & ys__n18841;
  assign new_n32344_ = ~new_n32342_ & ~new_n32343_;
  assign new_n32345_ = ~new_n17857_ & ~new_n32344_;
  assign new_n32346_ = ~new_n32341_ & ~new_n32345_;
  assign new_n32347_ = ys__n778 & ~new_n32346_;
  assign new_n32348_ = ~new_n32340_ & ~new_n32347_;
  assign new_n32349_ = ~ys__n602 & ~new_n32348_;
  assign new_n32350_ = new_n17857_ & ~new_n32348_;
  assign new_n32351_ = ys__n26170 & ~new_n17857_;
  assign new_n32352_ = ~new_n32350_ & ~new_n32351_;
  assign new_n32353_ = ys__n602 & ~new_n32352_;
  assign ys__n26740 = new_n32349_ | new_n32353_;
  assign new_n32355_ = ~ys__n778 & ys__n26170;
  assign new_n32356_ = ys__n26170 & new_n17857_;
  assign new_n32357_ = ys__n44 & ~ys__n18173;
  assign new_n32358_ = ys__n18173 & ys__n18843;
  assign new_n32359_ = ~new_n32357_ & ~new_n32358_;
  assign new_n32360_ = ~new_n17857_ & ~new_n32359_;
  assign new_n32361_ = ~new_n32356_ & ~new_n32360_;
  assign new_n32362_ = ys__n778 & ~new_n32361_;
  assign new_n32363_ = ~new_n32355_ & ~new_n32362_;
  assign new_n32364_ = ~ys__n602 & ~new_n32363_;
  assign new_n32365_ = new_n17857_ & ~new_n32363_;
  assign new_n32366_ = ys__n26172 & ~new_n17857_;
  assign new_n32367_ = ~new_n32365_ & ~new_n32366_;
  assign new_n32368_ = ys__n602 & ~new_n32367_;
  assign ys__n26741 = new_n32364_ | new_n32368_;
  assign new_n32370_ = ~ys__n778 & ys__n26172;
  assign new_n32371_ = ys__n26172 & new_n17857_;
  assign new_n32372_ = ys__n340 & ~ys__n18173;
  assign new_n32373_ = ys__n18173 & ys__n18845;
  assign new_n32374_ = ~new_n32372_ & ~new_n32373_;
  assign new_n32375_ = ~new_n17857_ & ~new_n32374_;
  assign new_n32376_ = ~new_n32371_ & ~new_n32375_;
  assign new_n32377_ = ys__n778 & ~new_n32376_;
  assign new_n32378_ = ~new_n32370_ & ~new_n32377_;
  assign new_n32379_ = ~ys__n602 & ~new_n32378_;
  assign new_n32380_ = new_n17857_ & ~new_n32378_;
  assign new_n32381_ = ys__n26174 & ~new_n17857_;
  assign new_n32382_ = ~new_n32380_ & ~new_n32381_;
  assign new_n32383_ = ys__n602 & ~new_n32382_;
  assign ys__n26742 = new_n32379_ | new_n32383_;
  assign new_n32385_ = ~ys__n778 & ys__n26174;
  assign new_n32386_ = ys__n26174 & new_n17857_;
  assign new_n32387_ = ys__n46 & ~ys__n18173;
  assign new_n32388_ = ys__n18173 & ys__n18847;
  assign new_n32389_ = ~new_n32387_ & ~new_n32388_;
  assign new_n32390_ = ~new_n17857_ & ~new_n32389_;
  assign new_n32391_ = ~new_n32386_ & ~new_n32390_;
  assign new_n32392_ = ys__n778 & ~new_n32391_;
  assign new_n32393_ = ~new_n32385_ & ~new_n32392_;
  assign new_n32394_ = ~ys__n602 & ~new_n32393_;
  assign new_n32395_ = new_n17857_ & ~new_n32393_;
  assign new_n32396_ = ys__n26176 & ~new_n17857_;
  assign new_n32397_ = ~new_n32395_ & ~new_n32396_;
  assign new_n32398_ = ys__n602 & ~new_n32397_;
  assign ys__n26743 = new_n32394_ | new_n32398_;
  assign new_n32400_ = ~ys__n778 & ys__n26176;
  assign new_n32401_ = ys__n26176 & new_n17857_;
  assign new_n32402_ = ys__n6118 & ~ys__n18173;
  assign new_n32403_ = ys__n18173 & ys__n18849;
  assign new_n32404_ = ~new_n32402_ & ~new_n32403_;
  assign new_n32405_ = ~new_n17857_ & ~new_n32404_;
  assign new_n32406_ = ~new_n32401_ & ~new_n32405_;
  assign new_n32407_ = ys__n778 & ~new_n32406_;
  assign new_n32408_ = ~new_n32400_ & ~new_n32407_;
  assign new_n32409_ = ~ys__n602 & ~new_n32408_;
  assign new_n32410_ = new_n17857_ & ~new_n32408_;
  assign new_n32411_ = ys__n26178 & ~new_n17857_;
  assign new_n32412_ = ~new_n32410_ & ~new_n32411_;
  assign new_n32413_ = ys__n602 & ~new_n32412_;
  assign ys__n26744 = new_n32409_ | new_n32413_;
  assign new_n32415_ = ~ys__n778 & ys__n26178;
  assign new_n32416_ = ys__n26178 & new_n17857_;
  assign new_n32417_ = ys__n6119 & ~ys__n18173;
  assign new_n32418_ = ys__n18173 & ys__n18851;
  assign new_n32419_ = ~new_n32417_ & ~new_n32418_;
  assign new_n32420_ = ~new_n17857_ & ~new_n32419_;
  assign new_n32421_ = ~new_n32416_ & ~new_n32420_;
  assign new_n32422_ = ys__n778 & ~new_n32421_;
  assign new_n32423_ = ~new_n32415_ & ~new_n32422_;
  assign new_n32424_ = ~ys__n602 & ~new_n32423_;
  assign new_n32425_ = new_n17857_ & ~new_n32423_;
  assign new_n32426_ = ys__n26180 & ~new_n17857_;
  assign new_n32427_ = ~new_n32425_ & ~new_n32426_;
  assign new_n32428_ = ys__n602 & ~new_n32427_;
  assign ys__n26745 = new_n32424_ | new_n32428_;
  assign new_n32430_ = ~ys__n778 & ys__n26180;
  assign new_n32431_ = ys__n26180 & new_n17857_;
  assign new_n32432_ = ys__n6120 & ~ys__n18173;
  assign new_n32433_ = ys__n18173 & ys__n18853;
  assign new_n32434_ = ~new_n32432_ & ~new_n32433_;
  assign new_n32435_ = ~new_n17857_ & ~new_n32434_;
  assign new_n32436_ = ~new_n32431_ & ~new_n32435_;
  assign new_n32437_ = ys__n778 & ~new_n32436_;
  assign new_n32438_ = ~new_n32430_ & ~new_n32437_;
  assign new_n32439_ = ~ys__n602 & ~new_n32438_;
  assign new_n32440_ = new_n17857_ & ~new_n32438_;
  assign new_n32441_ = ys__n26182 & ~new_n17857_;
  assign new_n32442_ = ~new_n32440_ & ~new_n32441_;
  assign new_n32443_ = ys__n602 & ~new_n32442_;
  assign ys__n26746 = new_n32439_ | new_n32443_;
  assign new_n32445_ = ~ys__n778 & ys__n26182;
  assign new_n32446_ = ys__n26182 & new_n17857_;
  assign new_n32447_ = ys__n6121 & ~ys__n18173;
  assign new_n32448_ = ys__n18173 & ys__n18855;
  assign new_n32449_ = ~new_n32447_ & ~new_n32448_;
  assign new_n32450_ = ~new_n17857_ & ~new_n32449_;
  assign new_n32451_ = ~new_n32446_ & ~new_n32450_;
  assign new_n32452_ = ys__n778 & ~new_n32451_;
  assign new_n32453_ = ~new_n32445_ & ~new_n32452_;
  assign new_n32454_ = ~ys__n602 & ~new_n32453_;
  assign new_n32455_ = new_n17857_ & ~new_n32453_;
  assign new_n32456_ = ys__n26184 & ~new_n17857_;
  assign new_n32457_ = ~new_n32455_ & ~new_n32456_;
  assign new_n32458_ = ys__n602 & ~new_n32457_;
  assign ys__n26747 = new_n32454_ | new_n32458_;
  assign new_n32460_ = ~ys__n778 & ys__n26184;
  assign new_n32461_ = ys__n26184 & new_n17857_;
  assign new_n32462_ = ys__n6123 & ~ys__n18173;
  assign new_n32463_ = ys__n18173 & ys__n18857;
  assign new_n32464_ = ~new_n32462_ & ~new_n32463_;
  assign new_n32465_ = ~new_n17857_ & ~new_n32464_;
  assign new_n32466_ = ~new_n32461_ & ~new_n32465_;
  assign new_n32467_ = ys__n778 & ~new_n32466_;
  assign new_n32468_ = ~new_n32460_ & ~new_n32467_;
  assign new_n32469_ = ~ys__n602 & ~new_n32468_;
  assign new_n32470_ = new_n17857_ & ~new_n32468_;
  assign new_n32471_ = ys__n26186 & ~new_n17857_;
  assign new_n32472_ = ~new_n32470_ & ~new_n32471_;
  assign new_n32473_ = ys__n602 & ~new_n32472_;
  assign ys__n26748 = new_n32469_ | new_n32473_;
  assign new_n32475_ = ~ys__n778 & ys__n26186;
  assign new_n32476_ = ys__n26186 & new_n17857_;
  assign new_n32477_ = ys__n6124 & ~ys__n18173;
  assign new_n32478_ = ys__n18173 & ys__n18859;
  assign new_n32479_ = ~new_n32477_ & ~new_n32478_;
  assign new_n32480_ = ~new_n17857_ & ~new_n32479_;
  assign new_n32481_ = ~new_n32476_ & ~new_n32480_;
  assign new_n32482_ = ys__n778 & ~new_n32481_;
  assign new_n32483_ = ~new_n32475_ & ~new_n32482_;
  assign new_n32484_ = ~ys__n602 & ~new_n32483_;
  assign new_n32485_ = new_n17857_ & ~new_n32483_;
  assign new_n32486_ = ys__n26188 & ~new_n17857_;
  assign new_n32487_ = ~new_n32485_ & ~new_n32486_;
  assign new_n32488_ = ys__n602 & ~new_n32487_;
  assign ys__n26749 = new_n32484_ | new_n32488_;
  assign new_n32490_ = ~ys__n778 & ys__n26188;
  assign new_n32491_ = ys__n26188 & new_n17857_;
  assign new_n32492_ = ys__n6126 & ~ys__n18173;
  assign new_n32493_ = ys__n18173 & ys__n18861;
  assign new_n32494_ = ~new_n32492_ & ~new_n32493_;
  assign new_n32495_ = ~new_n17857_ & ~new_n32494_;
  assign new_n32496_ = ~new_n32491_ & ~new_n32495_;
  assign new_n32497_ = ys__n778 & ~new_n32496_;
  assign new_n32498_ = ~new_n32490_ & ~new_n32497_;
  assign new_n32499_ = ~ys__n602 & ~new_n32498_;
  assign new_n32500_ = new_n17857_ & ~new_n32498_;
  assign new_n32501_ = ys__n26190 & ~new_n17857_;
  assign new_n32502_ = ~new_n32500_ & ~new_n32501_;
  assign new_n32503_ = ys__n602 & ~new_n32502_;
  assign ys__n26750 = new_n32499_ | new_n32503_;
  assign new_n32505_ = ~ys__n778 & ys__n26190;
  assign new_n32506_ = ys__n26190 & new_n17857_;
  assign new_n32507_ = ys__n6127 & ~ys__n18173;
  assign new_n32508_ = ys__n18173 & ys__n18863;
  assign new_n32509_ = ~new_n32507_ & ~new_n32508_;
  assign new_n32510_ = ~new_n17857_ & ~new_n32509_;
  assign new_n32511_ = ~new_n32506_ & ~new_n32510_;
  assign new_n32512_ = ys__n778 & ~new_n32511_;
  assign new_n32513_ = ~new_n32505_ & ~new_n32512_;
  assign new_n32514_ = ~ys__n602 & ~new_n32513_;
  assign new_n32515_ = new_n17857_ & ~new_n32513_;
  assign new_n32516_ = ys__n26192 & ~new_n17857_;
  assign new_n32517_ = ~new_n32515_ & ~new_n32516_;
  assign new_n32518_ = ys__n602 & ~new_n32517_;
  assign ys__n26751 = new_n32514_ | new_n32518_;
  assign new_n32520_ = ~ys__n778 & ys__n26192;
  assign new_n32521_ = ys__n26192 & new_n17857_;
  assign new_n32522_ = ys__n6129 & ~ys__n18173;
  assign new_n32523_ = ys__n18173 & ys__n18865;
  assign new_n32524_ = ~new_n32522_ & ~new_n32523_;
  assign new_n32525_ = ~new_n17857_ & ~new_n32524_;
  assign new_n32526_ = ~new_n32521_ & ~new_n32525_;
  assign new_n32527_ = ys__n778 & ~new_n32526_;
  assign new_n32528_ = ~new_n32520_ & ~new_n32527_;
  assign new_n32529_ = ~ys__n602 & ~new_n32528_;
  assign new_n32530_ = new_n17857_ & ~new_n32528_;
  assign new_n32531_ = ys__n26194 & ~new_n17857_;
  assign new_n32532_ = ~new_n32530_ & ~new_n32531_;
  assign new_n32533_ = ys__n602 & ~new_n32532_;
  assign ys__n26752 = new_n32529_ | new_n32533_;
  assign new_n32535_ = ~ys__n778 & ys__n26194;
  assign new_n32536_ = ys__n26194 & new_n17857_;
  assign new_n32537_ = ys__n6130 & ~ys__n18173;
  assign new_n32538_ = ys__n18173 & ys__n18867;
  assign new_n32539_ = ~new_n32537_ & ~new_n32538_;
  assign new_n32540_ = ~new_n17857_ & ~new_n32539_;
  assign new_n32541_ = ~new_n32536_ & ~new_n32540_;
  assign new_n32542_ = ys__n778 & ~new_n32541_;
  assign new_n32543_ = ~new_n32535_ & ~new_n32542_;
  assign new_n32544_ = ~ys__n602 & ~new_n32543_;
  assign new_n32545_ = new_n17857_ & ~new_n32543_;
  assign new_n32546_ = ys__n26196 & ~new_n17857_;
  assign new_n32547_ = ~new_n32545_ & ~new_n32546_;
  assign new_n32548_ = ys__n602 & ~new_n32547_;
  assign ys__n26753 = new_n32544_ | new_n32548_;
  assign new_n32550_ = ~ys__n778 & ys__n26196;
  assign new_n32551_ = ys__n26196 & new_n17857_;
  assign new_n32552_ = ys__n42 & ~ys__n18173;
  assign new_n32553_ = ys__n18173 & ys__n18869;
  assign new_n32554_ = ~new_n32552_ & ~new_n32553_;
  assign new_n32555_ = ~new_n17857_ & ~new_n32554_;
  assign new_n32556_ = ~new_n32551_ & ~new_n32555_;
  assign new_n32557_ = ys__n778 & ~new_n32556_;
  assign new_n32558_ = ~new_n32550_ & ~new_n32557_;
  assign new_n32559_ = ~ys__n602 & ~new_n32558_;
  assign new_n32560_ = new_n17857_ & ~new_n32558_;
  assign new_n32561_ = ys__n26198 & ~new_n17857_;
  assign new_n32562_ = ~new_n32560_ & ~new_n32561_;
  assign new_n32563_ = ys__n602 & ~new_n32562_;
  assign ys__n26754 = new_n32559_ | new_n32563_;
  assign new_n32565_ = ~ys__n778 & ys__n26198;
  assign new_n32566_ = ys__n26198 & new_n17857_;
  assign new_n32567_ = ys__n40 & ~ys__n18173;
  assign new_n32568_ = ys__n18173 & ys__n18871;
  assign new_n32569_ = ~new_n32567_ & ~new_n32568_;
  assign new_n32570_ = ~new_n17857_ & ~new_n32569_;
  assign new_n32571_ = ~new_n32566_ & ~new_n32570_;
  assign new_n32572_ = ys__n778 & ~new_n32571_;
  assign new_n32573_ = ~new_n32565_ & ~new_n32572_;
  assign new_n32574_ = ~ys__n602 & ~new_n32573_;
  assign new_n32575_ = new_n17857_ & ~new_n32573_;
  assign new_n32576_ = ys__n26200 & ~new_n17857_;
  assign new_n32577_ = ~new_n32575_ & ~new_n32576_;
  assign new_n32578_ = ys__n602 & ~new_n32577_;
  assign ys__n26755 = new_n32574_ | new_n32578_;
  assign new_n32580_ = ~ys__n778 & ys__n26200;
  assign new_n32581_ = ys__n26200 & new_n17857_;
  assign new_n32582_ = ys__n6133 & ~ys__n18173;
  assign new_n32583_ = ys__n18173 & ys__n18873;
  assign new_n32584_ = ~new_n32582_ & ~new_n32583_;
  assign new_n32585_ = ~new_n17857_ & ~new_n32584_;
  assign new_n32586_ = ~new_n32581_ & ~new_n32585_;
  assign new_n32587_ = ys__n778 & ~new_n32586_;
  assign new_n32588_ = ~new_n32580_ & ~new_n32587_;
  assign new_n32589_ = ~ys__n602 & ~new_n32588_;
  assign new_n32590_ = new_n17857_ & ~new_n32588_;
  assign new_n32591_ = ys__n26202 & ~new_n17857_;
  assign new_n32592_ = ~new_n32590_ & ~new_n32591_;
  assign new_n32593_ = ys__n602 & ~new_n32592_;
  assign ys__n26756 = new_n32589_ | new_n32593_;
  assign new_n32595_ = ~ys__n778 & ys__n26202;
  assign new_n32596_ = ys__n26202 & new_n17857_;
  assign new_n32597_ = ys__n6134 & ~ys__n18173;
  assign new_n32598_ = ys__n18173 & ys__n18875;
  assign new_n32599_ = ~new_n32597_ & ~new_n32598_;
  assign new_n32600_ = ~new_n17857_ & ~new_n32599_;
  assign new_n32601_ = ~new_n32596_ & ~new_n32600_;
  assign new_n32602_ = ys__n778 & ~new_n32601_;
  assign new_n32603_ = ~new_n32595_ & ~new_n32602_;
  assign new_n32604_ = ~ys__n602 & ~new_n32603_;
  assign new_n32605_ = new_n17857_ & ~new_n32603_;
  assign new_n32606_ = ys__n26204 & ~new_n17857_;
  assign new_n32607_ = ~new_n32605_ & ~new_n32606_;
  assign new_n32608_ = ys__n602 & ~new_n32607_;
  assign ys__n26757 = new_n32604_ | new_n32608_;
  assign new_n32610_ = ~ys__n778 & ys__n26204;
  assign new_n32611_ = ys__n26204 & new_n17857_;
  assign new_n32612_ = ys__n38 & ~ys__n18173;
  assign new_n32613_ = ys__n18173 & ys__n18877;
  assign new_n32614_ = ~new_n32612_ & ~new_n32613_;
  assign new_n32615_ = ~new_n17857_ & ~new_n32614_;
  assign new_n32616_ = ~new_n32611_ & ~new_n32615_;
  assign new_n32617_ = ys__n778 & ~new_n32616_;
  assign new_n32618_ = ~new_n32610_ & ~new_n32617_;
  assign new_n32619_ = ~ys__n602 & ~new_n32618_;
  assign new_n32620_ = new_n17857_ & ~new_n32618_;
  assign new_n32621_ = ys__n26206 & ~new_n17857_;
  assign new_n32622_ = ~new_n32620_ & ~new_n32621_;
  assign new_n32623_ = ys__n602 & ~new_n32622_;
  assign ys__n26758 = new_n32619_ | new_n32623_;
  assign new_n32625_ = ~ys__n778 & ys__n26206;
  assign new_n32626_ = ys__n26206 & new_n17857_;
  assign new_n32627_ = ys__n36 & ~ys__n18173;
  assign new_n32628_ = ys__n18173 & ys__n18879;
  assign new_n32629_ = ~new_n32627_ & ~new_n32628_;
  assign new_n32630_ = ~new_n17857_ & ~new_n32629_;
  assign new_n32631_ = ~new_n32626_ & ~new_n32630_;
  assign new_n32632_ = ys__n778 & ~new_n32631_;
  assign new_n32633_ = ~new_n32625_ & ~new_n32632_;
  assign new_n32634_ = ~ys__n602 & ~new_n32633_;
  assign new_n32635_ = new_n17857_ & ~new_n32633_;
  assign new_n32636_ = ys__n26208 & ~new_n17857_;
  assign new_n32637_ = ~new_n32635_ & ~new_n32636_;
  assign new_n32638_ = ys__n602 & ~new_n32637_;
  assign ys__n26759 = new_n32634_ | new_n32638_;
  assign new_n32640_ = ~ys__n778 & ys__n26208;
  assign new_n32641_ = ys__n26208 & new_n17857_;
  assign new_n32642_ = ys__n34 & ~ys__n18173;
  assign new_n32643_ = ys__n18173 & ys__n18881;
  assign new_n32644_ = ~new_n32642_ & ~new_n32643_;
  assign new_n32645_ = ~new_n17857_ & ~new_n32644_;
  assign new_n32646_ = ~new_n32641_ & ~new_n32645_;
  assign new_n32647_ = ys__n778 & ~new_n32646_;
  assign new_n32648_ = ~new_n32640_ & ~new_n32647_;
  assign new_n32649_ = ~ys__n602 & ~new_n32648_;
  assign new_n32650_ = new_n17857_ & ~new_n32648_;
  assign new_n32651_ = ys__n26210 & ~new_n17857_;
  assign new_n32652_ = ~new_n32650_ & ~new_n32651_;
  assign new_n32653_ = ys__n602 & ~new_n32652_;
  assign ys__n26760 = new_n32649_ | new_n32653_;
  assign new_n32655_ = ~ys__n778 & ys__n26210;
  assign new_n32656_ = ys__n26210 & new_n17857_;
  assign new_n32657_ = ys__n32 & ~ys__n18173;
  assign new_n32658_ = ys__n18173 & ys__n18883;
  assign new_n32659_ = ~new_n32657_ & ~new_n32658_;
  assign new_n32660_ = ~new_n17857_ & ~new_n32659_;
  assign new_n32661_ = ~new_n32656_ & ~new_n32660_;
  assign new_n32662_ = ys__n778 & ~new_n32661_;
  assign new_n32663_ = ~new_n32655_ & ~new_n32662_;
  assign new_n32664_ = ~ys__n602 & ~new_n32663_;
  assign new_n32665_ = new_n17857_ & ~new_n32663_;
  assign new_n32666_ = ys__n26212 & ~new_n17857_;
  assign new_n32667_ = ~new_n32665_ & ~new_n32666_;
  assign new_n32668_ = ys__n602 & ~new_n32667_;
  assign ys__n26761 = new_n32664_ | new_n32668_;
  assign new_n32670_ = ~ys__n778 & ys__n26212;
  assign new_n32671_ = ys__n26212 & new_n17857_;
  assign new_n32672_ = ys__n30 & ~ys__n18173;
  assign new_n32673_ = ys__n18173 & ys__n18885;
  assign new_n32674_ = ~new_n32672_ & ~new_n32673_;
  assign new_n32675_ = ~new_n17857_ & ~new_n32674_;
  assign new_n32676_ = ~new_n32671_ & ~new_n32675_;
  assign new_n32677_ = ys__n778 & ~new_n32676_;
  assign new_n32678_ = ~new_n32670_ & ~new_n32677_;
  assign new_n32679_ = ~ys__n602 & ~new_n32678_;
  assign new_n32680_ = new_n17857_ & ~new_n32678_;
  assign new_n32681_ = ys__n26214 & ~new_n17857_;
  assign new_n32682_ = ~new_n32680_ & ~new_n32681_;
  assign new_n32683_ = ys__n602 & ~new_n32682_;
  assign ys__n26762 = new_n32679_ | new_n32683_;
  assign new_n32685_ = ~ys__n778 & ys__n26214;
  assign new_n32686_ = ys__n26214 & new_n17857_;
  assign new_n32687_ = ys__n28 & ~ys__n18173;
  assign new_n32688_ = ys__n18173 & ys__n18887;
  assign new_n32689_ = ~new_n32687_ & ~new_n32688_;
  assign new_n32690_ = ~new_n17857_ & ~new_n32689_;
  assign new_n32691_ = ~new_n32686_ & ~new_n32690_;
  assign new_n32692_ = ys__n778 & ~new_n32691_;
  assign new_n32693_ = ~new_n32685_ & ~new_n32692_;
  assign new_n32694_ = ~ys__n602 & ~new_n32693_;
  assign new_n32695_ = new_n17857_ & ~new_n32693_;
  assign new_n32696_ = ys__n26216 & ~new_n17857_;
  assign new_n32697_ = ~new_n32695_ & ~new_n32696_;
  assign new_n32698_ = ys__n602 & ~new_n32697_;
  assign ys__n26763 = new_n32694_ | new_n32698_;
  assign new_n32700_ = ~ys__n778 & ys__n26216;
  assign new_n32701_ = ys__n26216 & new_n17857_;
  assign new_n32702_ = ys__n26 & ~ys__n18173;
  assign new_n32703_ = ys__n18173 & ys__n18889;
  assign new_n32704_ = ~new_n32702_ & ~new_n32703_;
  assign new_n32705_ = ~new_n17857_ & ~new_n32704_;
  assign new_n32706_ = ~new_n32701_ & ~new_n32705_;
  assign new_n32707_ = ys__n778 & ~new_n32706_;
  assign new_n32708_ = ~new_n32700_ & ~new_n32707_;
  assign new_n32709_ = ~ys__n602 & ~new_n32708_;
  assign new_n32710_ = new_n17857_ & ~new_n32708_;
  assign new_n32711_ = ys__n26218 & ~new_n17857_;
  assign new_n32712_ = ~new_n32710_ & ~new_n32711_;
  assign new_n32713_ = ys__n602 & ~new_n32712_;
  assign ys__n26764 = new_n32709_ | new_n32713_;
  assign new_n32715_ = ~ys__n778 & ys__n26218;
  assign new_n32716_ = ys__n26218 & new_n17857_;
  assign new_n32717_ = ys__n24 & ~ys__n18173;
  assign new_n32718_ = ys__n18173 & ys__n18891;
  assign new_n32719_ = ~new_n32717_ & ~new_n32718_;
  assign new_n32720_ = ~new_n17857_ & ~new_n32719_;
  assign new_n32721_ = ~new_n32716_ & ~new_n32720_;
  assign new_n32722_ = ys__n778 & ~new_n32721_;
  assign new_n32723_ = ~new_n32715_ & ~new_n32722_;
  assign new_n32724_ = ~ys__n602 & ~new_n32723_;
  assign new_n32725_ = new_n17857_ & ~new_n32723_;
  assign new_n32726_ = ~new_n17857_ & new_n31780_;
  assign new_n32727_ = ~new_n32725_ & ~new_n32726_;
  assign new_n32728_ = ys__n602 & ~new_n32727_;
  assign ys__n26765 = new_n32724_ | new_n32728_;
  assign ys__n26802 = ys__n18448 & new_n13380_;
  assign ys__n26803 = new_n13384_ & ys__n26802;
  assign ys__n26804 = ys__n18451 & new_n13380_;
  assign ys__n26805 = new_n13384_ & ys__n26804;
  assign ys__n26806 = ys__n18454 & new_n13380_;
  assign ys__n26807 = new_n13384_ & ys__n26806;
  assign ys__n26808 = ys__n18457 & new_n13380_;
  assign ys__n26809 = new_n13384_ & ys__n26808;
  assign ys__n26810 = ys__n18460 & new_n13380_;
  assign ys__n26811 = new_n13384_ & ys__n26810;
  assign ys__n26812 = ys__n18463 & new_n13380_;
  assign ys__n26813 = new_n13384_ & ys__n26812;
  assign ys__n26814 = ys__n18466 & new_n13380_;
  assign ys__n26815 = new_n13384_ & ys__n26814;
  assign ys__n26816 = ys__n18469 & new_n13380_;
  assign ys__n26817 = new_n13384_ & ys__n26816;
  assign ys__n26818 = ys__n18472 & new_n13380_;
  assign ys__n26819 = new_n13384_ & ys__n26818;
  assign ys__n26820 = ys__n18475 & new_n13380_;
  assign ys__n26821 = new_n13384_ & ys__n26820;
  assign ys__n26822 = ys__n18478 & new_n13380_;
  assign ys__n26823 = new_n13384_ & ys__n26822;
  assign ys__n26824 = ys__n18481 & new_n13380_;
  assign ys__n26825 = new_n13384_ & ys__n26824;
  assign ys__n26826 = ys__n18484 & new_n13380_;
  assign ys__n26827 = new_n13384_ & ys__n26826;
  assign ys__n26828 = ys__n18487 & new_n13380_;
  assign ys__n26829 = new_n13384_ & ys__n26828;
  assign ys__n26830 = ys__n18490 & new_n13380_;
  assign ys__n26831 = new_n13384_ & ys__n26830;
  assign ys__n26832 = ys__n18493 & new_n13380_;
  assign ys__n26833 = new_n13384_ & ys__n26832;
  assign ys__n26834 = ys__n18496 & new_n13380_;
  assign ys__n26835 = new_n13384_ & ys__n26834;
  assign ys__n26836 = ys__n18499 & new_n13380_;
  assign ys__n26837 = new_n13384_ & ys__n26836;
  assign ys__n26838 = ys__n18502 & new_n13380_;
  assign ys__n26839 = new_n13384_ & ys__n26838;
  assign ys__n26840 = ys__n18505 & new_n13380_;
  assign ys__n26841 = new_n13384_ & ys__n26840;
  assign ys__n26842 = ys__n18508 & new_n13380_;
  assign ys__n26843 = new_n13384_ & ys__n26842;
  assign ys__n26844 = ys__n18511 & new_n13380_;
  assign ys__n26845 = new_n13384_ & ys__n26844;
  assign ys__n26846 = ys__n18514 & new_n13380_;
  assign ys__n26847 = new_n13384_ & ys__n26846;
  assign ys__n26848 = ys__n18517 & new_n13380_;
  assign ys__n26849 = new_n13384_ & ys__n26848;
  assign ys__n26850 = ys__n18520 & new_n13380_;
  assign ys__n26851 = new_n13384_ & ys__n26850;
  assign ys__n26852 = ys__n18523 & new_n13380_;
  assign ys__n26853 = new_n13384_ & ys__n26852;
  assign ys__n26854 = ys__n18526 & new_n13380_;
  assign ys__n26855 = new_n13384_ & ys__n26854;
  assign ys__n26856 = ys__n18529 & new_n13380_;
  assign ys__n26857 = new_n13384_ & ys__n26856;
  assign ys__n26858 = ys__n18532 & new_n13380_;
  assign ys__n26859 = new_n13384_ & ys__n26858;
  assign ys__n26860 = ys__n18535 & new_n13380_;
  assign ys__n26861 = new_n13384_ & ys__n26860;
  assign ys__n26862 = ys__n18538 & new_n13380_;
  assign ys__n26863 = new_n13384_ & ys__n26862;
  assign ys__n26864 = ys__n18541 & new_n13380_;
  assign ys__n26865 = new_n13384_ & ys__n26864;
  assign ys__n26866 = ys__n18448 & new_n13379_;
  assign ys__n26867 = new_n13384_ & ys__n26866;
  assign ys__n26868 = ys__n18451 & new_n13379_;
  assign ys__n26869 = new_n13384_ & ys__n26868;
  assign ys__n26870 = ys__n18454 & new_n13379_;
  assign ys__n26871 = new_n13384_ & ys__n26870;
  assign ys__n26872 = ys__n18457 & new_n13379_;
  assign ys__n26873 = new_n13384_ & ys__n26872;
  assign ys__n26874 = ys__n18460 & new_n13379_;
  assign ys__n26875 = new_n13384_ & ys__n26874;
  assign ys__n26876 = ys__n18463 & new_n13379_;
  assign ys__n26877 = new_n13384_ & ys__n26876;
  assign ys__n26878 = ys__n18466 & new_n13379_;
  assign ys__n26879 = new_n13384_ & ys__n26878;
  assign ys__n26880 = ys__n18469 & new_n13379_;
  assign ys__n26881 = new_n13384_ & ys__n26880;
  assign ys__n26882 = ys__n18472 & new_n13379_;
  assign ys__n26883 = new_n13384_ & ys__n26882;
  assign ys__n26884 = ys__n18475 & new_n13379_;
  assign ys__n26885 = new_n13384_ & ys__n26884;
  assign ys__n26886 = ys__n18478 & new_n13379_;
  assign ys__n26887 = new_n13384_ & ys__n26886;
  assign ys__n26888 = ys__n18481 & new_n13379_;
  assign ys__n26889 = new_n13384_ & ys__n26888;
  assign ys__n26890 = ys__n18484 & new_n13379_;
  assign ys__n26891 = new_n13384_ & ys__n26890;
  assign ys__n26892 = ys__n18487 & new_n13379_;
  assign ys__n26893 = new_n13384_ & ys__n26892;
  assign ys__n26894 = ys__n18490 & new_n13379_;
  assign ys__n26895 = new_n13384_ & ys__n26894;
  assign ys__n26896 = ys__n18493 & new_n13379_;
  assign ys__n26897 = new_n13384_ & ys__n26896;
  assign ys__n26898 = ys__n18496 & new_n13379_;
  assign ys__n26899 = new_n13384_ & ys__n26898;
  assign ys__n26900 = ys__n18499 & new_n13379_;
  assign ys__n26901 = new_n13384_ & ys__n26900;
  assign ys__n26902 = ys__n18502 & new_n13379_;
  assign ys__n26903 = new_n13384_ & ys__n26902;
  assign ys__n26904 = ys__n18505 & new_n13379_;
  assign ys__n26905 = new_n13384_ & ys__n26904;
  assign ys__n26906 = ys__n18508 & new_n13379_;
  assign ys__n26907 = new_n13384_ & ys__n26906;
  assign ys__n26908 = ys__n18511 & new_n13379_;
  assign ys__n26909 = new_n13384_ & ys__n26908;
  assign ys__n26910 = ys__n18514 & new_n13379_;
  assign ys__n26911 = new_n13384_ & ys__n26910;
  assign ys__n26912 = ys__n18517 & new_n13379_;
  assign ys__n26913 = new_n13384_ & ys__n26912;
  assign ys__n26914 = ys__n18520 & new_n13379_;
  assign ys__n26915 = new_n13384_ & ys__n26914;
  assign ys__n26916 = ys__n18523 & new_n13379_;
  assign ys__n26917 = new_n13384_ & ys__n26916;
  assign ys__n26918 = ys__n18526 & new_n13379_;
  assign ys__n26919 = new_n13384_ & ys__n26918;
  assign ys__n26920 = ys__n18529 & new_n13379_;
  assign ys__n26921 = new_n13384_ & ys__n26920;
  assign ys__n26922 = ys__n18532 & new_n13379_;
  assign ys__n26923 = new_n13384_ & ys__n26922;
  assign ys__n26924 = ys__n18535 & new_n13379_;
  assign ys__n26925 = new_n13384_ & ys__n26924;
  assign ys__n26926 = ys__n18538 & new_n13379_;
  assign ys__n26927 = new_n13384_ & ys__n26926;
  assign ys__n26928 = ys__n18541 & new_n13379_;
  assign ys__n26929 = new_n13384_ & ys__n26928;
  assign ys__n26930 = ys__n18448 & new_n13382_;
  assign ys__n26931 = new_n13384_ & ys__n26930;
  assign ys__n26932 = ys__n18451 & new_n13382_;
  assign ys__n26933 = new_n13384_ & ys__n26932;
  assign ys__n26934 = ys__n18454 & new_n13382_;
  assign ys__n26935 = new_n13384_ & ys__n26934;
  assign ys__n26936 = ys__n18457 & new_n13382_;
  assign ys__n26937 = new_n13384_ & ys__n26936;
  assign ys__n26938 = ys__n18460 & new_n13382_;
  assign ys__n26939 = new_n13384_ & ys__n26938;
  assign ys__n26940 = ys__n18463 & new_n13382_;
  assign ys__n26941 = new_n13384_ & ys__n26940;
  assign ys__n26942 = ys__n18466 & new_n13382_;
  assign ys__n26943 = new_n13384_ & ys__n26942;
  assign ys__n26944 = ys__n18469 & new_n13382_;
  assign ys__n26945 = new_n13384_ & ys__n26944;
  assign ys__n26946 = ys__n18472 & new_n13382_;
  assign ys__n26947 = new_n13384_ & ys__n26946;
  assign ys__n26948 = ys__n18475 & new_n13382_;
  assign ys__n26949 = new_n13384_ & ys__n26948;
  assign ys__n26950 = ys__n18478 & new_n13382_;
  assign ys__n26951 = new_n13384_ & ys__n26950;
  assign ys__n26952 = ys__n18481 & new_n13382_;
  assign ys__n26953 = new_n13384_ & ys__n26952;
  assign ys__n26954 = ys__n18484 & new_n13382_;
  assign ys__n26955 = new_n13384_ & ys__n26954;
  assign ys__n26956 = ys__n18487 & new_n13382_;
  assign ys__n26957 = new_n13384_ & ys__n26956;
  assign ys__n26958 = ys__n18490 & new_n13382_;
  assign ys__n26959 = new_n13384_ & ys__n26958;
  assign ys__n26960 = ys__n18493 & new_n13382_;
  assign ys__n26961 = new_n13384_ & ys__n26960;
  assign ys__n26962 = ys__n18496 & new_n13382_;
  assign ys__n26963 = new_n13384_ & ys__n26962;
  assign ys__n26964 = ys__n18499 & new_n13382_;
  assign ys__n26965 = new_n13384_ & ys__n26964;
  assign ys__n26966 = ys__n18502 & new_n13382_;
  assign ys__n26967 = new_n13384_ & ys__n26966;
  assign ys__n26968 = ys__n18505 & new_n13382_;
  assign ys__n26969 = new_n13384_ & ys__n26968;
  assign ys__n26970 = ys__n18508 & new_n13382_;
  assign ys__n26971 = new_n13384_ & ys__n26970;
  assign ys__n26972 = ys__n18511 & new_n13382_;
  assign ys__n26973 = new_n13384_ & ys__n26972;
  assign ys__n26974 = ys__n18514 & new_n13382_;
  assign ys__n26975 = new_n13384_ & ys__n26974;
  assign ys__n26976 = ys__n18517 & new_n13382_;
  assign ys__n26977 = new_n13384_ & ys__n26976;
  assign ys__n26978 = ys__n18520 & new_n13382_;
  assign ys__n26979 = new_n13384_ & ys__n26978;
  assign ys__n26980 = ys__n18523 & new_n13382_;
  assign ys__n26981 = new_n13384_ & ys__n26980;
  assign ys__n26982 = ys__n18526 & new_n13382_;
  assign ys__n26983 = new_n13384_ & ys__n26982;
  assign ys__n26984 = ys__n18529 & new_n13382_;
  assign ys__n26985 = new_n13384_ & ys__n26984;
  assign ys__n26986 = ys__n18532 & new_n13382_;
  assign ys__n26987 = new_n13384_ & ys__n26986;
  assign ys__n26988 = ys__n18535 & new_n13382_;
  assign ys__n26989 = new_n13384_ & ys__n26988;
  assign ys__n26990 = ys__n18538 & new_n13382_;
  assign ys__n26991 = new_n13384_ & ys__n26990;
  assign ys__n26992 = ys__n18541 & new_n13382_;
  assign ys__n26993 = new_n13384_ & ys__n26992;
  assign ys__n26994 = ys__n18448 & new_n13490_;
  assign ys__n26995 = new_n13384_ & ys__n26994;
  assign ys__n26996 = ys__n18451 & new_n13490_;
  assign ys__n26997 = new_n13384_ & ys__n26996;
  assign ys__n26998 = ys__n18454 & new_n13490_;
  assign ys__n26999 = new_n13384_ & ys__n26998;
  assign ys__n27000 = ys__n18457 & new_n13490_;
  assign ys__n27001 = new_n13384_ & ys__n27000;
  assign ys__n27002 = ys__n18460 & new_n13490_;
  assign ys__n27003 = new_n13384_ & ys__n27002;
  assign ys__n27004 = ys__n18463 & new_n13490_;
  assign ys__n27005 = new_n13384_ & ys__n27004;
  assign ys__n27006 = ys__n18466 & new_n13490_;
  assign ys__n27007 = new_n13384_ & ys__n27006;
  assign ys__n27008 = ys__n18469 & new_n13490_;
  assign ys__n27009 = new_n13384_ & ys__n27008;
  assign ys__n27010 = ys__n18472 & new_n13490_;
  assign ys__n27011 = new_n13384_ & ys__n27010;
  assign ys__n27012 = ys__n18475 & new_n13490_;
  assign ys__n27013 = new_n13384_ & ys__n27012;
  assign ys__n27014 = ys__n18478 & new_n13490_;
  assign ys__n27015 = new_n13384_ & ys__n27014;
  assign ys__n27016 = ys__n18481 & new_n13490_;
  assign ys__n27017 = new_n13384_ & ys__n27016;
  assign ys__n27018 = ys__n18484 & new_n13490_;
  assign ys__n27019 = new_n13384_ & ys__n27018;
  assign ys__n27020 = ys__n18487 & new_n13490_;
  assign ys__n27021 = new_n13384_ & ys__n27020;
  assign ys__n27022 = ys__n18490 & new_n13490_;
  assign ys__n27023 = new_n13384_ & ys__n27022;
  assign ys__n27024 = ys__n18493 & new_n13490_;
  assign ys__n27025 = new_n13384_ & ys__n27024;
  assign ys__n27026 = ys__n18496 & new_n13490_;
  assign ys__n27027 = new_n13384_ & ys__n27026;
  assign ys__n27028 = ys__n18499 & new_n13490_;
  assign ys__n27029 = new_n13384_ & ys__n27028;
  assign ys__n27030 = ys__n18502 & new_n13490_;
  assign ys__n27031 = new_n13384_ & ys__n27030;
  assign ys__n27032 = ys__n18505 & new_n13490_;
  assign ys__n27033 = new_n13384_ & ys__n27032;
  assign ys__n27034 = ys__n18508 & new_n13490_;
  assign ys__n27035 = new_n13384_ & ys__n27034;
  assign ys__n27036 = ys__n18511 & new_n13490_;
  assign ys__n27037 = new_n13384_ & ys__n27036;
  assign ys__n27038 = ys__n18514 & new_n13490_;
  assign ys__n27039 = new_n13384_ & ys__n27038;
  assign ys__n27040 = ys__n18517 & new_n13490_;
  assign ys__n27041 = new_n13384_ & ys__n27040;
  assign ys__n27042 = ys__n18520 & new_n13490_;
  assign ys__n27043 = new_n13384_ & ys__n27042;
  assign ys__n27044 = ys__n18523 & new_n13490_;
  assign ys__n27045 = new_n13384_ & ys__n27044;
  assign ys__n27046 = ys__n18526 & new_n13490_;
  assign ys__n27047 = new_n13384_ & ys__n27046;
  assign ys__n27048 = ys__n18529 & new_n13490_;
  assign ys__n27049 = new_n13384_ & ys__n27048;
  assign ys__n27050 = ys__n18532 & new_n13490_;
  assign ys__n27051 = new_n13384_ & ys__n27050;
  assign ys__n27052 = ys__n18535 & new_n13490_;
  assign ys__n27053 = new_n13384_ & ys__n27052;
  assign ys__n27054 = ys__n18538 & new_n13490_;
  assign ys__n27055 = new_n13384_ & ys__n27054;
  assign ys__n27056 = ys__n18541 & new_n13490_;
  assign ys__n27057 = new_n13384_ & ys__n27056;
  assign ys__n27058 = new_n13376_ & ys__n26802;
  assign ys__n27059 = new_n13376_ & ys__n26804;
  assign ys__n27060 = new_n13376_ & ys__n26806;
  assign ys__n27061 = new_n13376_ & ys__n26808;
  assign ys__n27062 = new_n13376_ & ys__n26810;
  assign ys__n27063 = new_n13376_ & ys__n26812;
  assign ys__n27064 = new_n13376_ & ys__n26814;
  assign ys__n27065 = new_n13376_ & ys__n26816;
  assign ys__n27066 = new_n13376_ & ys__n26818;
  assign ys__n27067 = new_n13376_ & ys__n26820;
  assign ys__n27068 = new_n13376_ & ys__n26822;
  assign ys__n27069 = new_n13376_ & ys__n26824;
  assign ys__n27070 = new_n13376_ & ys__n26826;
  assign ys__n27071 = new_n13376_ & ys__n26828;
  assign ys__n27072 = new_n13376_ & ys__n26830;
  assign ys__n27073 = new_n13376_ & ys__n26832;
  assign ys__n27074 = new_n13376_ & ys__n26834;
  assign ys__n27075 = new_n13376_ & ys__n26836;
  assign ys__n27076 = new_n13376_ & ys__n26838;
  assign ys__n27077 = new_n13376_ & ys__n26840;
  assign ys__n27078 = new_n13376_ & ys__n26842;
  assign ys__n27079 = new_n13376_ & ys__n26844;
  assign ys__n27080 = new_n13376_ & ys__n26846;
  assign ys__n27081 = new_n13376_ & ys__n26848;
  assign ys__n27082 = new_n13376_ & ys__n26850;
  assign ys__n27083 = new_n13376_ & ys__n26852;
  assign ys__n27084 = new_n13376_ & ys__n26854;
  assign ys__n27085 = new_n13376_ & ys__n26856;
  assign ys__n27086 = new_n13376_ & ys__n26858;
  assign ys__n27087 = new_n13376_ & ys__n26860;
  assign ys__n27088 = new_n13376_ & ys__n26862;
  assign ys__n27089 = new_n13376_ & ys__n26864;
  assign ys__n27090 = new_n13376_ & ys__n26866;
  assign ys__n27091 = new_n13376_ & ys__n26868;
  assign ys__n27092 = new_n13376_ & ys__n26870;
  assign ys__n27093 = new_n13376_ & ys__n26872;
  assign ys__n27094 = new_n13376_ & ys__n26874;
  assign ys__n27095 = new_n13376_ & ys__n26876;
  assign ys__n27096 = new_n13376_ & ys__n26878;
  assign ys__n27097 = new_n13376_ & ys__n26880;
  assign ys__n27098 = new_n13376_ & ys__n26882;
  assign ys__n27099 = new_n13376_ & ys__n26884;
  assign ys__n27100 = new_n13376_ & ys__n26886;
  assign ys__n27101 = new_n13376_ & ys__n26888;
  assign ys__n27102 = new_n13376_ & ys__n26890;
  assign ys__n27103 = new_n13376_ & ys__n26892;
  assign ys__n27104 = new_n13376_ & ys__n26894;
  assign ys__n27105 = new_n13376_ & ys__n26896;
  assign ys__n27106 = new_n13376_ & ys__n26898;
  assign ys__n27107 = new_n13376_ & ys__n26900;
  assign ys__n27108 = new_n13376_ & ys__n26902;
  assign ys__n27109 = new_n13376_ & ys__n26904;
  assign ys__n27110 = new_n13376_ & ys__n26906;
  assign ys__n27111 = new_n13376_ & ys__n26908;
  assign ys__n27112 = new_n13376_ & ys__n26910;
  assign ys__n27113 = new_n13376_ & ys__n26912;
  assign ys__n27114 = new_n13376_ & ys__n26914;
  assign ys__n27115 = new_n13376_ & ys__n26916;
  assign ys__n27116 = new_n13376_ & ys__n26918;
  assign ys__n27117 = new_n13376_ & ys__n26920;
  assign ys__n27118 = new_n13376_ & ys__n26922;
  assign ys__n27119 = new_n13376_ & ys__n26924;
  assign ys__n27120 = new_n13376_ & ys__n26926;
  assign ys__n27121 = new_n13376_ & ys__n26928;
  assign ys__n27122 = new_n13376_ & ys__n26930;
  assign ys__n27123 = new_n13376_ & ys__n26932;
  assign ys__n27124 = new_n13376_ & ys__n26934;
  assign ys__n27125 = new_n13376_ & ys__n26936;
  assign ys__n27126 = new_n13376_ & ys__n26938;
  assign ys__n27127 = new_n13376_ & ys__n26940;
  assign ys__n27128 = new_n13376_ & ys__n26942;
  assign ys__n27129 = new_n13376_ & ys__n26944;
  assign ys__n27130 = new_n13376_ & ys__n26946;
  assign ys__n27131 = new_n13376_ & ys__n26948;
  assign ys__n27132 = new_n13376_ & ys__n26950;
  assign ys__n27133 = new_n13376_ & ys__n26952;
  assign ys__n27134 = new_n13376_ & ys__n26954;
  assign ys__n27135 = new_n13376_ & ys__n26956;
  assign ys__n27136 = new_n13376_ & ys__n26958;
  assign ys__n27137 = new_n13376_ & ys__n26960;
  assign ys__n27138 = new_n13376_ & ys__n26962;
  assign ys__n27139 = new_n13376_ & ys__n26964;
  assign ys__n27140 = new_n13376_ & ys__n26966;
  assign ys__n27141 = new_n13376_ & ys__n26968;
  assign ys__n27142 = new_n13376_ & ys__n26970;
  assign ys__n27143 = new_n13376_ & ys__n26972;
  assign ys__n27144 = new_n13376_ & ys__n26974;
  assign ys__n27145 = new_n13376_ & ys__n26976;
  assign ys__n27146 = new_n13376_ & ys__n26978;
  assign ys__n27147 = new_n13376_ & ys__n26980;
  assign ys__n27148 = new_n13376_ & ys__n26982;
  assign ys__n27149 = new_n13376_ & ys__n26984;
  assign ys__n27150 = new_n13376_ & ys__n26986;
  assign ys__n27151 = new_n13376_ & ys__n26988;
  assign ys__n27152 = new_n13376_ & ys__n26990;
  assign ys__n27153 = new_n13376_ & ys__n26992;
  assign ys__n27154 = new_n13376_ & ys__n26994;
  assign ys__n27155 = new_n13376_ & ys__n26996;
  assign ys__n27156 = new_n13376_ & ys__n26998;
  assign ys__n27157 = new_n13376_ & ys__n27000;
  assign ys__n27158 = new_n13376_ & ys__n27002;
  assign ys__n27159 = new_n13376_ & ys__n27004;
  assign ys__n27160 = new_n13376_ & ys__n27006;
  assign ys__n27161 = new_n13376_ & ys__n27008;
  assign ys__n27162 = new_n13376_ & ys__n27010;
  assign ys__n27163 = new_n13376_ & ys__n27012;
  assign ys__n27164 = new_n13376_ & ys__n27014;
  assign ys__n27165 = new_n13376_ & ys__n27016;
  assign ys__n27166 = new_n13376_ & ys__n27018;
  assign ys__n27167 = new_n13376_ & ys__n27020;
  assign ys__n27168 = new_n13376_ & ys__n27022;
  assign ys__n27169 = new_n13376_ & ys__n27024;
  assign ys__n27170 = new_n13376_ & ys__n27026;
  assign ys__n27171 = new_n13376_ & ys__n27028;
  assign ys__n27172 = new_n13376_ & ys__n27030;
  assign ys__n27173 = new_n13376_ & ys__n27032;
  assign ys__n27174 = new_n13376_ & ys__n27034;
  assign ys__n27175 = new_n13376_ & ys__n27036;
  assign ys__n27176 = new_n13376_ & ys__n27038;
  assign ys__n27177 = new_n13376_ & ys__n27040;
  assign ys__n27178 = new_n13376_ & ys__n27042;
  assign ys__n27179 = new_n13376_ & ys__n27044;
  assign ys__n27180 = new_n13376_ & ys__n27046;
  assign ys__n27181 = new_n13376_ & ys__n27048;
  assign ys__n27182 = new_n13376_ & ys__n27050;
  assign ys__n27183 = new_n13376_ & ys__n27052;
  assign ys__n27184 = new_n13376_ & ys__n27054;
  assign ys__n27185 = new_n13376_ & ys__n27056;
  assign ys__n27186 = new_n13374_ & ys__n26802;
  assign ys__n27187 = new_n13374_ & ys__n26804;
  assign ys__n27188 = new_n13374_ & ys__n26806;
  assign ys__n27189 = new_n13374_ & ys__n26808;
  assign ys__n27190 = new_n13374_ & ys__n26810;
  assign ys__n27191 = new_n13374_ & ys__n26812;
  assign ys__n27192 = new_n13374_ & ys__n26814;
  assign ys__n27193 = new_n13374_ & ys__n26816;
  assign ys__n27194 = new_n13374_ & ys__n26818;
  assign ys__n27195 = new_n13374_ & ys__n26820;
  assign ys__n27196 = new_n13374_ & ys__n26822;
  assign ys__n27197 = new_n13374_ & ys__n26824;
  assign ys__n27198 = new_n13374_ & ys__n26826;
  assign ys__n27199 = new_n13374_ & ys__n26828;
  assign ys__n27200 = new_n13374_ & ys__n26830;
  assign ys__n27201 = new_n13374_ & ys__n26832;
  assign ys__n27202 = new_n13374_ & ys__n26834;
  assign ys__n27203 = new_n13374_ & ys__n26836;
  assign ys__n27204 = new_n13374_ & ys__n26838;
  assign ys__n27205 = new_n13374_ & ys__n26840;
  assign ys__n27206 = new_n13374_ & ys__n26842;
  assign ys__n27207 = new_n13374_ & ys__n26844;
  assign ys__n27208 = new_n13374_ & ys__n26846;
  assign ys__n27209 = new_n13374_ & ys__n26848;
  assign ys__n27210 = new_n13374_ & ys__n26850;
  assign ys__n27211 = new_n13374_ & ys__n26852;
  assign ys__n27212 = new_n13374_ & ys__n26854;
  assign ys__n27213 = new_n13374_ & ys__n26856;
  assign ys__n27214 = new_n13374_ & ys__n26858;
  assign ys__n27215 = new_n13374_ & ys__n26860;
  assign ys__n27216 = new_n13374_ & ys__n26862;
  assign ys__n27217 = new_n13374_ & ys__n26864;
  assign ys__n27218 = new_n13374_ & ys__n26866;
  assign ys__n27219 = new_n13374_ & ys__n26868;
  assign ys__n27220 = new_n13374_ & ys__n26870;
  assign ys__n27221 = new_n13374_ & ys__n26872;
  assign ys__n27222 = new_n13374_ & ys__n26874;
  assign ys__n27223 = new_n13374_ & ys__n26876;
  assign ys__n27224 = new_n13374_ & ys__n26878;
  assign ys__n27225 = new_n13374_ & ys__n26880;
  assign ys__n27226 = new_n13374_ & ys__n26882;
  assign ys__n27227 = new_n13374_ & ys__n26884;
  assign ys__n27228 = new_n13374_ & ys__n26886;
  assign ys__n27229 = new_n13374_ & ys__n26888;
  assign ys__n27230 = new_n13374_ & ys__n26890;
  assign ys__n27231 = new_n13374_ & ys__n26892;
  assign ys__n27232 = new_n13374_ & ys__n26894;
  assign ys__n27233 = new_n13374_ & ys__n26896;
  assign ys__n27234 = new_n13374_ & ys__n26898;
  assign ys__n27235 = new_n13374_ & ys__n26900;
  assign ys__n27236 = new_n13374_ & ys__n26902;
  assign ys__n27237 = new_n13374_ & ys__n26904;
  assign ys__n27238 = new_n13374_ & ys__n26906;
  assign ys__n27239 = new_n13374_ & ys__n26908;
  assign ys__n27240 = new_n13374_ & ys__n26910;
  assign ys__n27241 = new_n13374_ & ys__n26912;
  assign ys__n27242 = new_n13374_ & ys__n26914;
  assign ys__n27243 = new_n13374_ & ys__n26916;
  assign ys__n27244 = new_n13374_ & ys__n26918;
  assign ys__n27245 = new_n13374_ & ys__n26920;
  assign ys__n27246 = new_n13374_ & ys__n26922;
  assign ys__n27247 = new_n13374_ & ys__n26924;
  assign ys__n27248 = new_n13374_ & ys__n26926;
  assign ys__n27249 = new_n13374_ & ys__n26928;
  assign ys__n27250 = new_n13374_ & ys__n26930;
  assign ys__n27251 = new_n13374_ & ys__n26932;
  assign ys__n27252 = new_n13374_ & ys__n26934;
  assign ys__n27253 = new_n13374_ & ys__n26936;
  assign ys__n27254 = new_n13374_ & ys__n26938;
  assign ys__n27255 = new_n13374_ & ys__n26940;
  assign ys__n27256 = new_n13374_ & ys__n26942;
  assign ys__n27257 = new_n13374_ & ys__n26944;
  assign ys__n27258 = new_n13374_ & ys__n26946;
  assign ys__n27259 = new_n13374_ & ys__n26948;
  assign ys__n27260 = new_n13374_ & ys__n26950;
  assign ys__n27261 = new_n13374_ & ys__n26952;
  assign ys__n27262 = new_n13374_ & ys__n26954;
  assign ys__n27263 = new_n13374_ & ys__n26956;
  assign ys__n27264 = new_n13374_ & ys__n26958;
  assign ys__n27265 = new_n13374_ & ys__n26960;
  assign ys__n27266 = new_n13374_ & ys__n26962;
  assign ys__n27267 = new_n13374_ & ys__n26964;
  assign ys__n27268 = new_n13374_ & ys__n26966;
  assign ys__n27269 = new_n13374_ & ys__n26968;
  assign ys__n27270 = new_n13374_ & ys__n26970;
  assign ys__n27271 = new_n13374_ & ys__n26972;
  assign ys__n27272 = new_n13374_ & ys__n26974;
  assign ys__n27273 = new_n13374_ & ys__n26976;
  assign ys__n27274 = new_n13374_ & ys__n26978;
  assign ys__n27275 = new_n13374_ & ys__n26980;
  assign ys__n27276 = new_n13374_ & ys__n26982;
  assign ys__n27277 = new_n13374_ & ys__n26984;
  assign ys__n27278 = new_n13374_ & ys__n26986;
  assign ys__n27279 = new_n13374_ & ys__n26988;
  assign ys__n27280 = new_n13374_ & ys__n26990;
  assign ys__n27281 = new_n13374_ & ys__n26992;
  assign ys__n27282 = new_n13374_ & ys__n26994;
  assign ys__n27283 = new_n13374_ & ys__n26996;
  assign ys__n27284 = new_n13374_ & ys__n26998;
  assign ys__n27285 = new_n13374_ & ys__n27000;
  assign ys__n27286 = new_n13374_ & ys__n27002;
  assign ys__n27287 = new_n13374_ & ys__n27004;
  assign ys__n27288 = new_n13374_ & ys__n27006;
  assign ys__n27289 = new_n13374_ & ys__n27008;
  assign ys__n27290 = new_n13374_ & ys__n27010;
  assign ys__n27291 = new_n13374_ & ys__n27012;
  assign ys__n27292 = new_n13374_ & ys__n27014;
  assign ys__n27293 = new_n13374_ & ys__n27016;
  assign ys__n27294 = new_n13374_ & ys__n27018;
  assign ys__n27295 = new_n13374_ & ys__n27020;
  assign ys__n27296 = new_n13374_ & ys__n27022;
  assign ys__n27297 = new_n13374_ & ys__n27024;
  assign ys__n27298 = new_n13374_ & ys__n27026;
  assign ys__n27299 = new_n13374_ & ys__n27028;
  assign ys__n27300 = new_n13374_ & ys__n27030;
  assign ys__n27301 = new_n13374_ & ys__n27032;
  assign ys__n27302 = new_n13374_ & ys__n27034;
  assign ys__n27303 = new_n13374_ & ys__n27036;
  assign ys__n27304 = new_n13374_ & ys__n27038;
  assign ys__n27305 = new_n13374_ & ys__n27040;
  assign ys__n27306 = new_n13374_ & ys__n27042;
  assign ys__n27307 = new_n13374_ & ys__n27044;
  assign ys__n27308 = new_n13374_ & ys__n27046;
  assign ys__n27309 = new_n13374_ & ys__n27048;
  assign ys__n27310 = new_n13374_ & ys__n27050;
  assign ys__n27311 = new_n13374_ & ys__n27052;
  assign ys__n27312 = new_n13374_ & ys__n27054;
  assign ys__n27313 = new_n13374_ & ys__n27056;
  assign ys__n27314 = new_n13375_ & ys__n26804;
  assign ys__n27315 = new_n13375_ & ys__n26806;
  assign ys__n27316 = new_n13375_ & ys__n26808;
  assign ys__n27317 = new_n13375_ & ys__n26810;
  assign ys__n27318 = new_n13375_ & ys__n26812;
  assign ys__n27319 = new_n13375_ & ys__n26814;
  assign ys__n27320 = new_n13375_ & ys__n26816;
  assign ys__n27321 = new_n13375_ & ys__n26818;
  assign ys__n27322 = new_n13375_ & ys__n26820;
  assign ys__n27323 = new_n13375_ & ys__n26822;
  assign ys__n27324 = new_n13375_ & ys__n26824;
  assign ys__n27325 = new_n13375_ & ys__n26826;
  assign ys__n27326 = new_n13375_ & ys__n26828;
  assign ys__n27327 = new_n13375_ & ys__n26830;
  assign ys__n27328 = new_n13375_ & ys__n26832;
  assign ys__n27329 = new_n13375_ & ys__n26834;
  assign ys__n27330 = new_n13375_ & ys__n26836;
  assign ys__n27331 = new_n13375_ & ys__n26838;
  assign ys__n27332 = new_n13375_ & ys__n26840;
  assign ys__n27333 = new_n13375_ & ys__n26842;
  assign ys__n27334 = new_n13375_ & ys__n26844;
  assign ys__n27335 = new_n13375_ & ys__n26846;
  assign ys__n27336 = new_n13375_ & ys__n26848;
  assign ys__n27337 = new_n13375_ & ys__n26850;
  assign ys__n27338 = new_n13375_ & ys__n26852;
  assign ys__n27339 = new_n13375_ & ys__n26854;
  assign ys__n27340 = new_n13375_ & ys__n26856;
  assign ys__n27341 = new_n13375_ & ys__n26858;
  assign ys__n27342 = new_n13375_ & ys__n26860;
  assign ys__n27343 = new_n13375_ & ys__n26862;
  assign ys__n27344 = new_n13375_ & ys__n26864;
  assign ys__n27345 = new_n13375_ & ys__n26868;
  assign ys__n27346 = new_n13375_ & ys__n26870;
  assign ys__n27347 = new_n13375_ & ys__n26872;
  assign ys__n27348 = new_n13375_ & ys__n26874;
  assign ys__n27349 = new_n13375_ & ys__n26876;
  assign ys__n27350 = new_n13375_ & ys__n26878;
  assign ys__n27351 = new_n13375_ & ys__n26880;
  assign ys__n27352 = new_n13375_ & ys__n26882;
  assign ys__n27353 = new_n13375_ & ys__n26884;
  assign ys__n27354 = new_n13375_ & ys__n26886;
  assign ys__n27355 = new_n13375_ & ys__n26888;
  assign ys__n27356 = new_n13375_ & ys__n26890;
  assign ys__n27357 = new_n13375_ & ys__n26892;
  assign ys__n27358 = new_n13375_ & ys__n26894;
  assign ys__n27359 = new_n13375_ & ys__n26896;
  assign ys__n27360 = new_n13375_ & ys__n26898;
  assign ys__n27361 = new_n13375_ & ys__n26900;
  assign ys__n27362 = new_n13375_ & ys__n26902;
  assign ys__n27363 = new_n13375_ & ys__n26904;
  assign ys__n27364 = new_n13375_ & ys__n26906;
  assign ys__n27365 = new_n13375_ & ys__n26908;
  assign ys__n27366 = new_n13375_ & ys__n26910;
  assign ys__n27367 = new_n13375_ & ys__n26912;
  assign ys__n27368 = new_n13375_ & ys__n26914;
  assign ys__n27369 = new_n13375_ & ys__n26916;
  assign ys__n27370 = new_n13375_ & ys__n26918;
  assign ys__n27371 = new_n13375_ & ys__n26920;
  assign ys__n27372 = new_n13375_ & ys__n26922;
  assign ys__n27373 = new_n13375_ & ys__n26924;
  assign ys__n27374 = new_n13375_ & ys__n26926;
  assign ys__n27375 = new_n13375_ & ys__n26928;
  assign ys__n27376 = new_n13375_ & ys__n26932;
  assign ys__n27377 = new_n13375_ & ys__n26934;
  assign ys__n27378 = new_n13375_ & ys__n26936;
  assign ys__n27379 = new_n13375_ & ys__n26938;
  assign ys__n27380 = new_n13375_ & ys__n26940;
  assign ys__n27381 = new_n13375_ & ys__n26942;
  assign ys__n27382 = new_n13375_ & ys__n26944;
  assign ys__n27383 = new_n13375_ & ys__n26946;
  assign ys__n27384 = new_n13375_ & ys__n26948;
  assign ys__n27385 = new_n13375_ & ys__n26950;
  assign ys__n27386 = new_n13375_ & ys__n26952;
  assign ys__n27387 = new_n13375_ & ys__n26954;
  assign ys__n27388 = new_n13375_ & ys__n26956;
  assign ys__n27389 = new_n13375_ & ys__n26958;
  assign ys__n27390 = new_n13375_ & ys__n26960;
  assign ys__n27391 = new_n13375_ & ys__n26962;
  assign ys__n27392 = new_n13375_ & ys__n26964;
  assign ys__n27393 = new_n13375_ & ys__n26966;
  assign ys__n27394 = new_n13375_ & ys__n26968;
  assign ys__n27395 = new_n13375_ & ys__n26970;
  assign ys__n27396 = new_n13375_ & ys__n26972;
  assign ys__n27397 = new_n13375_ & ys__n26974;
  assign ys__n27398 = new_n13375_ & ys__n26976;
  assign ys__n27399 = new_n13375_ & ys__n26978;
  assign ys__n27400 = new_n13375_ & ys__n26980;
  assign ys__n27401 = new_n13375_ & ys__n26982;
  assign ys__n27402 = new_n13375_ & ys__n26984;
  assign ys__n27403 = new_n13375_ & ys__n26986;
  assign ys__n27404 = new_n13375_ & ys__n26988;
  assign ys__n27405 = new_n13375_ & ys__n26990;
  assign ys__n27406 = new_n13375_ & ys__n26992;
  assign ys__n27407 = new_n13375_ & ys__n26996;
  assign ys__n27408 = new_n13375_ & ys__n26998;
  assign ys__n27409 = new_n13375_ & ys__n27000;
  assign ys__n27410 = new_n13375_ & ys__n27002;
  assign ys__n27411 = new_n13375_ & ys__n27004;
  assign ys__n27412 = new_n13375_ & ys__n27006;
  assign ys__n27413 = new_n13375_ & ys__n27008;
  assign ys__n27414 = new_n13375_ & ys__n27010;
  assign ys__n27415 = new_n13375_ & ys__n27012;
  assign ys__n27416 = new_n13375_ & ys__n27014;
  assign ys__n27417 = new_n13375_ & ys__n27016;
  assign ys__n27418 = new_n13375_ & ys__n27018;
  assign ys__n27419 = new_n13375_ & ys__n27020;
  assign ys__n27420 = new_n13375_ & ys__n27022;
  assign ys__n27421 = new_n13375_ & ys__n27024;
  assign ys__n27422 = new_n13375_ & ys__n27026;
  assign ys__n27423 = new_n13375_ & ys__n27028;
  assign ys__n27424 = new_n13375_ & ys__n27030;
  assign ys__n27425 = new_n13375_ & ys__n27032;
  assign ys__n27426 = new_n13375_ & ys__n27034;
  assign ys__n27427 = new_n13375_ & ys__n27036;
  assign ys__n27428 = new_n13375_ & ys__n27038;
  assign ys__n27429 = new_n13375_ & ys__n27040;
  assign ys__n27430 = new_n13375_ & ys__n27042;
  assign ys__n27431 = new_n13375_ & ys__n27044;
  assign ys__n27432 = new_n13375_ & ys__n27046;
  assign ys__n27433 = new_n13375_ & ys__n27048;
  assign ys__n27434 = new_n13375_ & ys__n27050;
  assign ys__n27435 = new_n13375_ & ys__n27052;
  assign ys__n27436 = new_n13375_ & ys__n27054;
  assign ys__n27437 = new_n13375_ & ys__n27056;
  assign new_n33366_ = ys__n26766 & ~new_n27901_;
  assign new_n33367_ = ys__n26766 & ~new_n27837_;
  assign new_n33368_ = ~new_n27839_ & ~new_n33367_;
  assign new_n33369_ = new_n27901_ & ~new_n33368_;
  assign new_n33370_ = ~new_n33366_ & ~new_n33369_;
  assign new_n33371_ = ys__n6126 & ys__n46936;
  assign new_n33372_ = ~ys__n6126 & ~ys__n46936;
  assign new_n33373_ = ~ys__n46906 & ~new_n33372_;
  assign new_n33374_ = ~new_n33371_ & new_n33373_;
  assign new_n33375_ = ys__n6127 & ys__n46937;
  assign new_n33376_ = ~ys__n6127 & ~ys__n46937;
  assign new_n33377_ = ~ys__n46908 & ~new_n33376_;
  assign new_n33378_ = ~new_n33375_ & new_n33377_;
  assign new_n33379_ = ~new_n33374_ & ~new_n33378_;
  assign new_n33380_ = ys__n6129 & ys__n46938;
  assign new_n33381_ = ~ys__n6129 & ~ys__n46938;
  assign new_n33382_ = ~ys__n46910 & ~new_n33381_;
  assign new_n33383_ = ~new_n33380_ & new_n33382_;
  assign new_n33384_ = ys__n6130 & ys__n46939;
  assign new_n33385_ = ~ys__n6130 & ~ys__n46939;
  assign new_n33386_ = ~ys__n46912 & ~new_n33385_;
  assign new_n33387_ = ~new_n33384_ & new_n33386_;
  assign new_n33388_ = ~new_n33383_ & ~new_n33387_;
  assign new_n33389_ = new_n33379_ & new_n33388_;
  assign new_n33390_ = ys__n6120 & ys__n46932;
  assign new_n33391_ = ~ys__n6120 & ~ys__n46932;
  assign new_n33392_ = ~ys__n46898 & ~new_n33391_;
  assign new_n33393_ = ~new_n33390_ & new_n33392_;
  assign new_n33394_ = ys__n6121 & ys__n46933;
  assign new_n33395_ = ~ys__n6121 & ~ys__n46933;
  assign new_n33396_ = ~ys__n46900 & ~new_n33395_;
  assign new_n33397_ = ~new_n33394_ & new_n33396_;
  assign new_n33398_ = ~new_n33393_ & ~new_n33397_;
  assign new_n33399_ = ys__n6123 & ys__n46934;
  assign new_n33400_ = ~ys__n6123 & ~ys__n46934;
  assign new_n33401_ = ~ys__n46902 & ~new_n33400_;
  assign new_n33402_ = ~new_n33399_ & new_n33401_;
  assign new_n33403_ = ys__n6124 & ys__n46935;
  assign new_n33404_ = ~ys__n6124 & ~ys__n46935;
  assign new_n33405_ = ~ys__n46904 & ~new_n33404_;
  assign new_n33406_ = ~new_n33403_ & new_n33405_;
  assign new_n33407_ = ~new_n33402_ & ~new_n33406_;
  assign new_n33408_ = new_n33398_ & new_n33407_;
  assign new_n33409_ = new_n33389_ & new_n33408_;
  assign new_n33410_ = ys__n18448 & ys__n46843;
  assign new_n33411_ = ~ys__n18448 & ~ys__n46843;
  assign new_n33412_ = ~ys__n46780 & ~new_n33411_;
  assign new_n33413_ = ~new_n33410_ & new_n33412_;
  assign new_n33414_ = ys__n18451 & ys__n46844;
  assign new_n33415_ = ~ys__n18451 & ~ys__n46844;
  assign new_n33416_ = ~ys__n46782 & ~new_n33415_;
  assign new_n33417_ = ~new_n33414_ & new_n33416_;
  assign new_n33418_ = ~new_n33413_ & ~new_n33417_;
  assign new_n33419_ = ys__n18454 & ys__n46845;
  assign new_n33420_ = ~ys__n18454 & ~ys__n46845;
  assign new_n33421_ = ~ys__n46784 & ~new_n33420_;
  assign new_n33422_ = ~new_n33419_ & new_n33421_;
  assign new_n33423_ = ys__n18457 & ys__n46846;
  assign new_n33424_ = ~ys__n18457 & ~ys__n46846;
  assign new_n33425_ = ~ys__n46786 & ~new_n33424_;
  assign new_n33426_ = ~new_n33423_ & new_n33425_;
  assign new_n33427_ = ~new_n33422_ & ~new_n33426_;
  assign new_n33428_ = new_n33418_ & new_n33427_;
  assign new_n33429_ = ys__n42 & ys__n46940;
  assign new_n33430_ = ~ys__n42 & ~ys__n46940;
  assign new_n33431_ = ~ys__n46914 & ~new_n33430_;
  assign new_n33432_ = ~new_n33429_ & new_n33431_;
  assign new_n33433_ = ys__n40 & ys__n46941;
  assign new_n33434_ = ~ys__n40 & ~ys__n46941;
  assign new_n33435_ = ~ys__n46916 & ~new_n33434_;
  assign new_n33436_ = ~new_n33433_ & new_n33435_;
  assign new_n33437_ = ~new_n33432_ & ~new_n33436_;
  assign new_n33438_ = ys__n6133 & ys__n46942;
  assign new_n33439_ = ~ys__n6133 & ~ys__n46942;
  assign new_n33440_ = ~ys__n46918 & ~new_n33439_;
  assign new_n33441_ = ~new_n33438_ & new_n33440_;
  assign new_n33442_ = ys__n6134 & ys__n46943;
  assign new_n33443_ = ~ys__n6134 & ~ys__n46943;
  assign new_n33444_ = ~ys__n46920 & ~new_n33443_;
  assign new_n33445_ = ~new_n33442_ & new_n33444_;
  assign new_n33446_ = ~new_n33441_ & ~new_n33445_;
  assign new_n33447_ = new_n33437_ & new_n33446_;
  assign new_n33448_ = new_n33428_ & new_n33447_;
  assign new_n33449_ = new_n33409_ & new_n33448_;
  assign new_n33450_ = ys__n6113 & ys__n46921;
  assign new_n33451_ = ~ys__n6113 & ~ys__n46921;
  assign new_n33452_ = ~ys__n46876 & ~new_n33451_;
  assign new_n33453_ = ~new_n33450_ & new_n33452_;
  assign new_n33454_ = ~ys__n38 & ~ys__n46944;
  assign new_n33455_ = ys__n38 & ys__n46944;
  assign new_n33456_ = ~new_n33454_ & ~new_n33455_;
  assign new_n33457_ = ~ys__n36 & ~ys__n46945;
  assign new_n33458_ = ys__n36 & ys__n46945;
  assign new_n33459_ = ~new_n33457_ & ~new_n33458_;
  assign new_n33460_ = ~new_n33456_ & ~new_n33459_;
  assign new_n33461_ = ~new_n33453_ & new_n33460_;
  assign new_n33462_ = ys__n172 & ys__n46922;
  assign new_n33463_ = ~ys__n172 & ~ys__n46922;
  assign new_n33464_ = ~ys__n46878 & ~new_n33463_;
  assign new_n33465_ = ~new_n33462_ & new_n33464_;
  assign new_n33466_ = ys__n338 & ys__n46923;
  assign new_n33467_ = ~ys__n338 & ~ys__n46923;
  assign new_n33468_ = ~ys__n46880 & ~new_n33467_;
  assign new_n33469_ = ~new_n33466_ & new_n33468_;
  assign new_n33470_ = ~new_n33465_ & ~new_n33469_;
  assign new_n33471_ = new_n33461_ & new_n33470_;
  assign new_n33472_ = ~ys__n26 & ~ys__n46950;
  assign new_n33473_ = ys__n26 & ys__n46950;
  assign new_n33474_ = ~new_n33472_ & ~new_n33473_;
  assign new_n33475_ = ~ys__n24 & ~ys__n46951;
  assign new_n33476_ = ys__n24 & ys__n46951;
  assign new_n33477_ = ~new_n33475_ & ~new_n33476_;
  assign new_n33478_ = ~new_n33474_ & ~new_n33477_;
  assign new_n33479_ = ~ys__n46230 & ys__n46231;
  assign new_n33480_ = ys__n46230 & ~ys__n46231;
  assign new_n33481_ = ~new_n33479_ & ~new_n33480_;
  assign new_n33482_ = ys__n18059 & ys__n18065;
  assign new_n33483_ = ~ys__n27479 & new_n33482_;
  assign new_n33484_ = ~new_n33481_ & ~new_n33483_;
  assign new_n33485_ = new_n33478_ & new_n33484_;
  assign new_n33486_ = ~ys__n34 & ~ys__n46946;
  assign new_n33487_ = ys__n34 & ys__n46946;
  assign new_n33488_ = ~new_n33486_ & ~new_n33487_;
  assign new_n33489_ = ~ys__n32 & ~ys__n46947;
  assign new_n33490_ = ys__n32 & ys__n46947;
  assign new_n33491_ = ~new_n33489_ & ~new_n33490_;
  assign new_n33492_ = ~new_n33488_ & ~new_n33491_;
  assign new_n33493_ = ~ys__n30 & ~ys__n46948;
  assign new_n33494_ = ys__n30 & ys__n46948;
  assign new_n33495_ = ~new_n33493_ & ~new_n33494_;
  assign new_n33496_ = ~ys__n28 & ~ys__n46949;
  assign new_n33497_ = ys__n28 & ys__n46949;
  assign new_n33498_ = ~new_n33496_ & ~new_n33497_;
  assign new_n33499_ = ~new_n33495_ & ~new_n33498_;
  assign new_n33500_ = new_n33492_ & new_n33499_;
  assign new_n33501_ = new_n33485_ & new_n33500_;
  assign new_n33502_ = new_n33471_ & new_n33501_;
  assign new_n33503_ = ys__n340 & ys__n46928;
  assign new_n33504_ = ~ys__n340 & ~ys__n46928;
  assign new_n33505_ = ~ys__n46890 & ~new_n33504_;
  assign new_n33506_ = ~new_n33503_ & new_n33505_;
  assign new_n33507_ = ys__n46 & ys__n46929;
  assign new_n33508_ = ~ys__n46 & ~ys__n46929;
  assign new_n33509_ = ~ys__n46892 & ~new_n33508_;
  assign new_n33510_ = ~new_n33507_ & new_n33509_;
  assign new_n33511_ = ~new_n33506_ & ~new_n33510_;
  assign new_n33512_ = ys__n6118 & ys__n46930;
  assign new_n33513_ = ~ys__n6118 & ~ys__n46930;
  assign new_n33514_ = ~ys__n46894 & ~new_n33513_;
  assign new_n33515_ = ~new_n33512_ & new_n33514_;
  assign new_n33516_ = ys__n6119 & ys__n46931;
  assign new_n33517_ = ~ys__n6119 & ~ys__n46931;
  assign new_n33518_ = ~ys__n46896 & ~new_n33517_;
  assign new_n33519_ = ~new_n33516_ & new_n33518_;
  assign new_n33520_ = ~new_n33515_ & ~new_n33519_;
  assign new_n33521_ = new_n33511_ & new_n33520_;
  assign new_n33522_ = ys__n22 & ys__n46924;
  assign new_n33523_ = ~ys__n22 & ~ys__n46924;
  assign new_n33524_ = ~ys__n46882 & ~new_n33523_;
  assign new_n33525_ = ~new_n33522_ & new_n33524_;
  assign new_n33526_ = ys__n316 & ys__n46925;
  assign new_n33527_ = ~ys__n316 & ~ys__n46925;
  assign new_n33528_ = ~ys__n46884 & ~new_n33527_;
  assign new_n33529_ = ~new_n33526_ & new_n33528_;
  assign new_n33530_ = ~new_n33525_ & ~new_n33529_;
  assign new_n33531_ = ys__n6115 & ys__n46926;
  assign new_n33532_ = ~ys__n6115 & ~ys__n46926;
  assign new_n33533_ = ~ys__n46886 & ~new_n33532_;
  assign new_n33534_ = ~new_n33531_ & new_n33533_;
  assign new_n33535_ = ys__n44 & ys__n46927;
  assign new_n33536_ = ~ys__n44 & ~ys__n46927;
  assign new_n33537_ = ~ys__n46888 & ~new_n33536_;
  assign new_n33538_ = ~new_n33535_ & new_n33537_;
  assign new_n33539_ = ~new_n33534_ & ~new_n33538_;
  assign new_n33540_ = new_n33530_ & new_n33539_;
  assign new_n33541_ = new_n33521_ & new_n33540_;
  assign new_n33542_ = new_n33502_ & new_n33541_;
  assign new_n33543_ = new_n33449_ & new_n33542_;
  assign new_n33544_ = ys__n18520 & ys__n46867;
  assign new_n33545_ = ~ys__n18520 & ~ys__n46867;
  assign new_n33546_ = ~ys__n46828 & ~new_n33545_;
  assign new_n33547_ = ~new_n33544_ & new_n33546_;
  assign new_n33548_ = ys__n18523 & ys__n46868;
  assign new_n33549_ = ~ys__n18523 & ~ys__n46868;
  assign new_n33550_ = ~ys__n46830 & ~new_n33549_;
  assign new_n33551_ = ~new_n33548_ & new_n33550_;
  assign new_n33552_ = ~new_n33547_ & ~new_n33551_;
  assign new_n33553_ = ys__n18526 & ys__n46869;
  assign new_n33554_ = ~ys__n18526 & ~ys__n46869;
  assign new_n33555_ = ~ys__n46832 & ~new_n33554_;
  assign new_n33556_ = ~new_n33553_ & new_n33555_;
  assign new_n33557_ = ys__n18529 & ys__n46870;
  assign new_n33558_ = ~ys__n18529 & ~ys__n46870;
  assign new_n33559_ = ~ys__n46834 & ~new_n33558_;
  assign new_n33560_ = ~new_n33557_ & new_n33559_;
  assign new_n33561_ = ~new_n33556_ & ~new_n33560_;
  assign new_n33562_ = new_n33552_ & new_n33561_;
  assign new_n33563_ = ys__n18508 & ys__n46863;
  assign new_n33564_ = ~ys__n18508 & ~ys__n46863;
  assign new_n33565_ = ~ys__n46820 & ~new_n33564_;
  assign new_n33566_ = ~new_n33563_ & new_n33565_;
  assign new_n33567_ = ys__n18511 & ys__n46864;
  assign new_n33568_ = ~ys__n18511 & ~ys__n46864;
  assign new_n33569_ = ~ys__n46822 & ~new_n33568_;
  assign new_n33570_ = ~new_n33567_ & new_n33569_;
  assign new_n33571_ = ~new_n33566_ & ~new_n33570_;
  assign new_n33572_ = ys__n18514 & ys__n46865;
  assign new_n33573_ = ~ys__n18514 & ~ys__n46865;
  assign new_n33574_ = ~ys__n46824 & ~new_n33573_;
  assign new_n33575_ = ~new_n33572_ & new_n33574_;
  assign new_n33576_ = ys__n18517 & ys__n46866;
  assign new_n33577_ = ~ys__n18517 & ~ys__n46866;
  assign new_n33578_ = ~ys__n46826 & ~new_n33577_;
  assign new_n33579_ = ~new_n33576_ & new_n33578_;
  assign new_n33580_ = ~new_n33575_ & ~new_n33579_;
  assign new_n33581_ = new_n33571_ & new_n33580_;
  assign new_n33582_ = new_n33562_ & new_n33581_;
  assign new_n33583_ = ~ys__n18059 & ~ys__n18065;
  assign new_n33584_ = ~ys__n18208 & new_n33583_;
  assign new_n33585_ = ~ys__n18061 & new_n33584_;
  assign new_n33586_ = ys__n18059 & ~ys__n18065;
  assign new_n33587_ = ys__n18208 & new_n33586_;
  assign new_n33588_ = ~ys__n18067 & new_n33587_;
  assign new_n33589_ = ~ys__n18208 & new_n33586_;
  assign new_n33590_ = ~ys__n18063 & new_n33589_;
  assign new_n33591_ = ~new_n33588_ & ~new_n33590_;
  assign new_n33592_ = ~new_n33585_ & new_n33591_;
  assign new_n33593_ = ys__n18532 & ys__n46871;
  assign new_n33594_ = ~ys__n18532 & ~ys__n46871;
  assign new_n33595_ = ~ys__n46836 & ~new_n33594_;
  assign new_n33596_ = ~new_n33593_ & new_n33595_;
  assign new_n33597_ = ys__n18535 & ys__n46872;
  assign new_n33598_ = ~ys__n18535 & ~ys__n46872;
  assign new_n33599_ = ~ys__n46838 & ~new_n33598_;
  assign new_n33600_ = ~new_n33597_ & new_n33599_;
  assign new_n33601_ = ~new_n33596_ & ~new_n33600_;
  assign new_n33602_ = ys__n18538 & ys__n46873;
  assign new_n33603_ = ~ys__n18538 & ~ys__n46873;
  assign new_n33604_ = ~ys__n46840 & ~new_n33603_;
  assign new_n33605_ = ~new_n33602_ & new_n33604_;
  assign new_n33606_ = ys__n18541 & ys__n46874;
  assign new_n33607_ = ~ys__n18541 & ~ys__n46874;
  assign new_n33608_ = ~ys__n46842 & ~new_n33607_;
  assign new_n33609_ = ~new_n33606_ & new_n33608_;
  assign new_n33610_ = ~new_n33605_ & ~new_n33609_;
  assign new_n33611_ = new_n33601_ & new_n33610_;
  assign new_n33612_ = new_n33592_ & new_n33611_;
  assign new_n33613_ = new_n33582_ & new_n33612_;
  assign new_n33614_ = ys__n18472 & ys__n46851;
  assign new_n33615_ = ~ys__n18472 & ~ys__n46851;
  assign new_n33616_ = ~ys__n46796 & ~new_n33615_;
  assign new_n33617_ = ~new_n33614_ & new_n33616_;
  assign new_n33618_ = ys__n18475 & ys__n46852;
  assign new_n33619_ = ~ys__n18475 & ~ys__n46852;
  assign new_n33620_ = ~ys__n46798 & ~new_n33619_;
  assign new_n33621_ = ~new_n33618_ & new_n33620_;
  assign new_n33622_ = ~new_n33617_ & ~new_n33621_;
  assign new_n33623_ = ys__n18478 & ys__n46853;
  assign new_n33624_ = ~ys__n18478 & ~ys__n46853;
  assign new_n33625_ = ~ys__n46800 & ~new_n33624_;
  assign new_n33626_ = ~new_n33623_ & new_n33625_;
  assign new_n33627_ = ys__n18481 & ys__n46854;
  assign new_n33628_ = ~ys__n18481 & ~ys__n46854;
  assign new_n33629_ = ~ys__n46802 & ~new_n33628_;
  assign new_n33630_ = ~new_n33627_ & new_n33629_;
  assign new_n33631_ = ~new_n33626_ & ~new_n33630_;
  assign new_n33632_ = new_n33622_ & new_n33631_;
  assign new_n33633_ = ys__n18460 & ys__n46847;
  assign new_n33634_ = ~ys__n18460 & ~ys__n46847;
  assign new_n33635_ = ~ys__n46788 & ~new_n33634_;
  assign new_n33636_ = ~new_n33633_ & new_n33635_;
  assign new_n33637_ = ys__n18463 & ys__n46848;
  assign new_n33638_ = ~ys__n18463 & ~ys__n46848;
  assign new_n33639_ = ~ys__n46790 & ~new_n33638_;
  assign new_n33640_ = ~new_n33637_ & new_n33639_;
  assign new_n33641_ = ~new_n33636_ & ~new_n33640_;
  assign new_n33642_ = ys__n18466 & ys__n46849;
  assign new_n33643_ = ~ys__n18466 & ~ys__n46849;
  assign new_n33644_ = ~ys__n46792 & ~new_n33643_;
  assign new_n33645_ = ~new_n33642_ & new_n33644_;
  assign new_n33646_ = ys__n18469 & ys__n46850;
  assign new_n33647_ = ~ys__n18469 & ~ys__n46850;
  assign new_n33648_ = ~ys__n46794 & ~new_n33647_;
  assign new_n33649_ = ~new_n33646_ & new_n33648_;
  assign new_n33650_ = ~new_n33645_ & ~new_n33649_;
  assign new_n33651_ = new_n33641_ & new_n33650_;
  assign new_n33652_ = new_n33632_ & new_n33651_;
  assign new_n33653_ = ys__n18496 & ys__n46859;
  assign new_n33654_ = ~ys__n18496 & ~ys__n46859;
  assign new_n33655_ = ~ys__n46812 & ~new_n33654_;
  assign new_n33656_ = ~new_n33653_ & new_n33655_;
  assign new_n33657_ = ys__n18499 & ys__n46860;
  assign new_n33658_ = ~ys__n18499 & ~ys__n46860;
  assign new_n33659_ = ~ys__n46814 & ~new_n33658_;
  assign new_n33660_ = ~new_n33657_ & new_n33659_;
  assign new_n33661_ = ~new_n33656_ & ~new_n33660_;
  assign new_n33662_ = ys__n18502 & ys__n46861;
  assign new_n33663_ = ~ys__n18502 & ~ys__n46861;
  assign new_n33664_ = ~ys__n46816 & ~new_n33663_;
  assign new_n33665_ = ~new_n33662_ & new_n33664_;
  assign new_n33666_ = ys__n18505 & ys__n46862;
  assign new_n33667_ = ~ys__n18505 & ~ys__n46862;
  assign new_n33668_ = ~ys__n46818 & ~new_n33667_;
  assign new_n33669_ = ~new_n33666_ & new_n33668_;
  assign new_n33670_ = ~new_n33665_ & ~new_n33669_;
  assign new_n33671_ = new_n33661_ & new_n33670_;
  assign new_n33672_ = ys__n18484 & ys__n46855;
  assign new_n33673_ = ~ys__n18484 & ~ys__n46855;
  assign new_n33674_ = ~ys__n46804 & ~new_n33673_;
  assign new_n33675_ = ~new_n33672_ & new_n33674_;
  assign new_n33676_ = ys__n18487 & ys__n46856;
  assign new_n33677_ = ~ys__n18487 & ~ys__n46856;
  assign new_n33678_ = ~ys__n46806 & ~new_n33677_;
  assign new_n33679_ = ~new_n33676_ & new_n33678_;
  assign new_n33680_ = ~new_n33675_ & ~new_n33679_;
  assign new_n33681_ = ys__n18490 & ys__n46857;
  assign new_n33682_ = ~ys__n18490 & ~ys__n46857;
  assign new_n33683_ = ~ys__n46808 & ~new_n33682_;
  assign new_n33684_ = ~new_n33681_ & new_n33683_;
  assign new_n33685_ = ys__n18493 & ys__n46858;
  assign new_n33686_ = ~ys__n18493 & ~ys__n46858;
  assign new_n33687_ = ~ys__n46810 & ~new_n33686_;
  assign new_n33688_ = ~new_n33685_ & new_n33687_;
  assign new_n33689_ = ~new_n33684_ & ~new_n33688_;
  assign new_n33690_ = new_n33680_ & new_n33689_;
  assign new_n33691_ = new_n33671_ & new_n33690_;
  assign new_n33692_ = new_n33652_ & new_n33691_;
  assign new_n33693_ = new_n33613_ & new_n33692_;
  assign new_n33694_ = new_n33543_ & new_n33693_;
  assign new_n33695_ = ~new_n33370_ & ~new_n33694_;
  assign new_n33696_ = ~ys__n27481 & ~new_n33370_;
  assign new_n33697_ = ~ys__n27481 & ~new_n33696_;
  assign new_n33698_ = ~ys__n27485 & ~new_n33697_;
  assign new_n33699_ = ~ys__n27485 & ~new_n33698_;
  assign new_n33700_ = new_n33694_ & ~new_n33699_;
  assign ys__n27484 = new_n33695_ | new_n33700_;
  assign new_n33702_ = ys__n26768 & ~new_n27901_;
  assign new_n33703_ = ys__n26768 & ~new_n27837_;
  assign new_n33704_ = ~new_n27846_ & ~new_n33703_;
  assign new_n33705_ = new_n27901_ & ~new_n33704_;
  assign new_n33706_ = ~new_n33702_ & ~new_n33705_;
  assign new_n33707_ = ys__n6126 & ys__n46760;
  assign new_n33708_ = ~ys__n6126 & ~ys__n46760;
  assign new_n33709_ = ~ys__n46730 & ~new_n33708_;
  assign new_n33710_ = ~new_n33707_ & new_n33709_;
  assign new_n33711_ = ys__n6127 & ys__n46761;
  assign new_n33712_ = ~ys__n6127 & ~ys__n46761;
  assign new_n33713_ = ~ys__n46732 & ~new_n33712_;
  assign new_n33714_ = ~new_n33711_ & new_n33713_;
  assign new_n33715_ = ~new_n33710_ & ~new_n33714_;
  assign new_n33716_ = ys__n6129 & ys__n46762;
  assign new_n33717_ = ~ys__n6129 & ~ys__n46762;
  assign new_n33718_ = ~ys__n46734 & ~new_n33717_;
  assign new_n33719_ = ~new_n33716_ & new_n33718_;
  assign new_n33720_ = ys__n6130 & ys__n46763;
  assign new_n33721_ = ~ys__n6130 & ~ys__n46763;
  assign new_n33722_ = ~ys__n46736 & ~new_n33721_;
  assign new_n33723_ = ~new_n33720_ & new_n33722_;
  assign new_n33724_ = ~new_n33719_ & ~new_n33723_;
  assign new_n33725_ = new_n33715_ & new_n33724_;
  assign new_n33726_ = ys__n6120 & ys__n46756;
  assign new_n33727_ = ~ys__n6120 & ~ys__n46756;
  assign new_n33728_ = ~ys__n46722 & ~new_n33727_;
  assign new_n33729_ = ~new_n33726_ & new_n33728_;
  assign new_n33730_ = ys__n6121 & ys__n46757;
  assign new_n33731_ = ~ys__n6121 & ~ys__n46757;
  assign new_n33732_ = ~ys__n46724 & ~new_n33731_;
  assign new_n33733_ = ~new_n33730_ & new_n33732_;
  assign new_n33734_ = ~new_n33729_ & ~new_n33733_;
  assign new_n33735_ = ys__n6123 & ys__n46758;
  assign new_n33736_ = ~ys__n6123 & ~ys__n46758;
  assign new_n33737_ = ~ys__n46726 & ~new_n33736_;
  assign new_n33738_ = ~new_n33735_ & new_n33737_;
  assign new_n33739_ = ys__n6124 & ys__n46759;
  assign new_n33740_ = ~ys__n6124 & ~ys__n46759;
  assign new_n33741_ = ~ys__n46728 & ~new_n33740_;
  assign new_n33742_ = ~new_n33739_ & new_n33741_;
  assign new_n33743_ = ~new_n33738_ & ~new_n33742_;
  assign new_n33744_ = new_n33734_ & new_n33743_;
  assign new_n33745_ = new_n33725_ & new_n33744_;
  assign new_n33746_ = ys__n18448 & ys__n46667;
  assign new_n33747_ = ~ys__n18448 & ~ys__n46667;
  assign new_n33748_ = ~ys__n46604 & ~new_n33747_;
  assign new_n33749_ = ~new_n33746_ & new_n33748_;
  assign new_n33750_ = ys__n18451 & ys__n46668;
  assign new_n33751_ = ~ys__n18451 & ~ys__n46668;
  assign new_n33752_ = ~ys__n46606 & ~new_n33751_;
  assign new_n33753_ = ~new_n33750_ & new_n33752_;
  assign new_n33754_ = ~new_n33749_ & ~new_n33753_;
  assign new_n33755_ = ys__n18454 & ys__n46669;
  assign new_n33756_ = ~ys__n18454 & ~ys__n46669;
  assign new_n33757_ = ~ys__n46608 & ~new_n33756_;
  assign new_n33758_ = ~new_n33755_ & new_n33757_;
  assign new_n33759_ = ys__n18457 & ys__n46670;
  assign new_n33760_ = ~ys__n18457 & ~ys__n46670;
  assign new_n33761_ = ~ys__n46610 & ~new_n33760_;
  assign new_n33762_ = ~new_n33759_ & new_n33761_;
  assign new_n33763_ = ~new_n33758_ & ~new_n33762_;
  assign new_n33764_ = new_n33754_ & new_n33763_;
  assign new_n33765_ = ys__n42 & ys__n46764;
  assign new_n33766_ = ~ys__n42 & ~ys__n46764;
  assign new_n33767_ = ~ys__n46738 & ~new_n33766_;
  assign new_n33768_ = ~new_n33765_ & new_n33767_;
  assign new_n33769_ = ys__n40 & ys__n46765;
  assign new_n33770_ = ~ys__n40 & ~ys__n46765;
  assign new_n33771_ = ~ys__n46740 & ~new_n33770_;
  assign new_n33772_ = ~new_n33769_ & new_n33771_;
  assign new_n33773_ = ~new_n33768_ & ~new_n33772_;
  assign new_n33774_ = ys__n6133 & ys__n46766;
  assign new_n33775_ = ~ys__n6133 & ~ys__n46766;
  assign new_n33776_ = ~ys__n46742 & ~new_n33775_;
  assign new_n33777_ = ~new_n33774_ & new_n33776_;
  assign new_n33778_ = ys__n6134 & ys__n46767;
  assign new_n33779_ = ~ys__n6134 & ~ys__n46767;
  assign new_n33780_ = ~ys__n46744 & ~new_n33779_;
  assign new_n33781_ = ~new_n33778_ & new_n33780_;
  assign new_n33782_ = ~new_n33777_ & ~new_n33781_;
  assign new_n33783_ = new_n33773_ & new_n33782_;
  assign new_n33784_ = new_n33764_ & new_n33783_;
  assign new_n33785_ = new_n33745_ & new_n33784_;
  assign new_n33786_ = ys__n6113 & ys__n46745;
  assign new_n33787_ = ~ys__n6113 & ~ys__n46745;
  assign new_n33788_ = ~ys__n46700 & ~new_n33787_;
  assign new_n33789_ = ~new_n33786_ & new_n33788_;
  assign new_n33790_ = ~ys__n38 & ~ys__n46768;
  assign new_n33791_ = ys__n38 & ys__n46768;
  assign new_n33792_ = ~new_n33790_ & ~new_n33791_;
  assign new_n33793_ = ~new_n33481_ & ~new_n33792_;
  assign new_n33794_ = ~new_n33789_ & new_n33793_;
  assign new_n33795_ = ys__n172 & ys__n46746;
  assign new_n33796_ = ~ys__n172 & ~ys__n46746;
  assign new_n33797_ = ~ys__n46702 & ~new_n33796_;
  assign new_n33798_ = ~new_n33795_ & new_n33797_;
  assign new_n33799_ = ys__n338 & ys__n46747;
  assign new_n33800_ = ~ys__n338 & ~ys__n46747;
  assign new_n33801_ = ~ys__n46704 & ~new_n33800_;
  assign new_n33802_ = ~new_n33799_ & new_n33801_;
  assign new_n33803_ = ~new_n33798_ & ~new_n33802_;
  assign new_n33804_ = new_n33794_ & new_n33803_;
  assign new_n33805_ = ~ys__n28 & ~ys__n46773;
  assign new_n33806_ = ys__n28 & ys__n46773;
  assign new_n33807_ = ~new_n33805_ & ~new_n33806_;
  assign new_n33808_ = ~ys__n26 & ~ys__n46774;
  assign new_n33809_ = ys__n26 & ys__n46774;
  assign new_n33810_ = ~new_n33808_ & ~new_n33809_;
  assign new_n33811_ = ~new_n33807_ & ~new_n33810_;
  assign new_n33812_ = ~ys__n24 & ~ys__n46775;
  assign new_n33813_ = ys__n24 & ys__n46775;
  assign new_n33814_ = ~new_n33812_ & ~new_n33813_;
  assign new_n33815_ = ~ys__n27488 & new_n33482_;
  assign new_n33816_ = ~new_n33814_ & ~new_n33815_;
  assign new_n33817_ = new_n33811_ & new_n33816_;
  assign new_n33818_ = ~ys__n36 & ~ys__n46769;
  assign new_n33819_ = ys__n36 & ys__n46769;
  assign new_n33820_ = ~new_n33818_ & ~new_n33819_;
  assign new_n33821_ = ~ys__n34 & ~ys__n46770;
  assign new_n33822_ = ys__n34 & ys__n46770;
  assign new_n33823_ = ~new_n33821_ & ~new_n33822_;
  assign new_n33824_ = ~new_n33820_ & ~new_n33823_;
  assign new_n33825_ = ~ys__n32 & ~ys__n46771;
  assign new_n33826_ = ys__n32 & ys__n46771;
  assign new_n33827_ = ~new_n33825_ & ~new_n33826_;
  assign new_n33828_ = ~ys__n30 & ~ys__n46772;
  assign new_n33829_ = ys__n30 & ys__n46772;
  assign new_n33830_ = ~new_n33828_ & ~new_n33829_;
  assign new_n33831_ = ~new_n33827_ & ~new_n33830_;
  assign new_n33832_ = new_n33824_ & new_n33831_;
  assign new_n33833_ = new_n33817_ & new_n33832_;
  assign new_n33834_ = new_n33804_ & new_n33833_;
  assign new_n33835_ = ys__n340 & ys__n46752;
  assign new_n33836_ = ~ys__n340 & ~ys__n46752;
  assign new_n33837_ = ~ys__n46714 & ~new_n33836_;
  assign new_n33838_ = ~new_n33835_ & new_n33837_;
  assign new_n33839_ = ys__n46 & ys__n46753;
  assign new_n33840_ = ~ys__n46 & ~ys__n46753;
  assign new_n33841_ = ~ys__n46716 & ~new_n33840_;
  assign new_n33842_ = ~new_n33839_ & new_n33841_;
  assign new_n33843_ = ~new_n33838_ & ~new_n33842_;
  assign new_n33844_ = ys__n6118 & ys__n46754;
  assign new_n33845_ = ~ys__n6118 & ~ys__n46754;
  assign new_n33846_ = ~ys__n46718 & ~new_n33845_;
  assign new_n33847_ = ~new_n33844_ & new_n33846_;
  assign new_n33848_ = ys__n6119 & ys__n46755;
  assign new_n33849_ = ~ys__n6119 & ~ys__n46755;
  assign new_n33850_ = ~ys__n46720 & ~new_n33849_;
  assign new_n33851_ = ~new_n33848_ & new_n33850_;
  assign new_n33852_ = ~new_n33847_ & ~new_n33851_;
  assign new_n33853_ = new_n33843_ & new_n33852_;
  assign new_n33854_ = ys__n22 & ys__n46748;
  assign new_n33855_ = ~ys__n22 & ~ys__n46748;
  assign new_n33856_ = ~ys__n46706 & ~new_n33855_;
  assign new_n33857_ = ~new_n33854_ & new_n33856_;
  assign new_n33858_ = ys__n316 & ys__n46749;
  assign new_n33859_ = ~ys__n316 & ~ys__n46749;
  assign new_n33860_ = ~ys__n46708 & ~new_n33859_;
  assign new_n33861_ = ~new_n33858_ & new_n33860_;
  assign new_n33862_ = ~new_n33857_ & ~new_n33861_;
  assign new_n33863_ = ys__n6115 & ys__n46750;
  assign new_n33864_ = ~ys__n6115 & ~ys__n46750;
  assign new_n33865_ = ~ys__n46710 & ~new_n33864_;
  assign new_n33866_ = ~new_n33863_ & new_n33865_;
  assign new_n33867_ = ys__n44 & ys__n46751;
  assign new_n33868_ = ~ys__n44 & ~ys__n46751;
  assign new_n33869_ = ~ys__n46712 & ~new_n33868_;
  assign new_n33870_ = ~new_n33867_ & new_n33869_;
  assign new_n33871_ = ~new_n33866_ & ~new_n33870_;
  assign new_n33872_ = new_n33862_ & new_n33871_;
  assign new_n33873_ = new_n33853_ & new_n33872_;
  assign new_n33874_ = new_n33834_ & new_n33873_;
  assign new_n33875_ = new_n33785_ & new_n33874_;
  assign new_n33876_ = ys__n18520 & ys__n46691;
  assign new_n33877_ = ~ys__n18520 & ~ys__n46691;
  assign new_n33878_ = ~ys__n46652 & ~new_n33877_;
  assign new_n33879_ = ~new_n33876_ & new_n33878_;
  assign new_n33880_ = ys__n18523 & ys__n46692;
  assign new_n33881_ = ~ys__n18523 & ~ys__n46692;
  assign new_n33882_ = ~ys__n46654 & ~new_n33881_;
  assign new_n33883_ = ~new_n33880_ & new_n33882_;
  assign new_n33884_ = ~new_n33879_ & ~new_n33883_;
  assign new_n33885_ = ys__n18526 & ys__n46693;
  assign new_n33886_ = ~ys__n18526 & ~ys__n46693;
  assign new_n33887_ = ~ys__n46656 & ~new_n33886_;
  assign new_n33888_ = ~new_n33885_ & new_n33887_;
  assign new_n33889_ = ys__n18529 & ys__n46694;
  assign new_n33890_ = ~ys__n18529 & ~ys__n46694;
  assign new_n33891_ = ~ys__n46658 & ~new_n33890_;
  assign new_n33892_ = ~new_n33889_ & new_n33891_;
  assign new_n33893_ = ~new_n33888_ & ~new_n33892_;
  assign new_n33894_ = new_n33884_ & new_n33893_;
  assign new_n33895_ = ys__n18508 & ys__n46687;
  assign new_n33896_ = ~ys__n18508 & ~ys__n46687;
  assign new_n33897_ = ~ys__n46644 & ~new_n33896_;
  assign new_n33898_ = ~new_n33895_ & new_n33897_;
  assign new_n33899_ = ys__n18511 & ys__n46688;
  assign new_n33900_ = ~ys__n18511 & ~ys__n46688;
  assign new_n33901_ = ~ys__n46646 & ~new_n33900_;
  assign new_n33902_ = ~new_n33899_ & new_n33901_;
  assign new_n33903_ = ~new_n33898_ & ~new_n33902_;
  assign new_n33904_ = ys__n18514 & ys__n46689;
  assign new_n33905_ = ~ys__n18514 & ~ys__n46689;
  assign new_n33906_ = ~ys__n46648 & ~new_n33905_;
  assign new_n33907_ = ~new_n33904_ & new_n33906_;
  assign new_n33908_ = ys__n18517 & ys__n46690;
  assign new_n33909_ = ~ys__n18517 & ~ys__n46690;
  assign new_n33910_ = ~ys__n46650 & ~new_n33909_;
  assign new_n33911_ = ~new_n33908_ & new_n33910_;
  assign new_n33912_ = ~new_n33907_ & ~new_n33911_;
  assign new_n33913_ = new_n33903_ & new_n33912_;
  assign new_n33914_ = new_n33894_ & new_n33913_;
  assign new_n33915_ = ~ys__n18053 & new_n33584_;
  assign new_n33916_ = ~ys__n18057 & new_n33587_;
  assign new_n33917_ = ~ys__n18055 & new_n33589_;
  assign new_n33918_ = ~new_n33916_ & ~new_n33917_;
  assign new_n33919_ = ~new_n33915_ & new_n33918_;
  assign new_n33920_ = ys__n18532 & ys__n46695;
  assign new_n33921_ = ~ys__n18532 & ~ys__n46695;
  assign new_n33922_ = ~ys__n46660 & ~new_n33921_;
  assign new_n33923_ = ~new_n33920_ & new_n33922_;
  assign new_n33924_ = ys__n18535 & ys__n46696;
  assign new_n33925_ = ~ys__n18535 & ~ys__n46696;
  assign new_n33926_ = ~ys__n46662 & ~new_n33925_;
  assign new_n33927_ = ~new_n33924_ & new_n33926_;
  assign new_n33928_ = ~new_n33923_ & ~new_n33927_;
  assign new_n33929_ = ys__n18538 & ys__n46697;
  assign new_n33930_ = ~ys__n18538 & ~ys__n46697;
  assign new_n33931_ = ~ys__n46664 & ~new_n33930_;
  assign new_n33932_ = ~new_n33929_ & new_n33931_;
  assign new_n33933_ = ys__n18541 & ys__n46698;
  assign new_n33934_ = ~ys__n18541 & ~ys__n46698;
  assign new_n33935_ = ~ys__n46666 & ~new_n33934_;
  assign new_n33936_ = ~new_n33933_ & new_n33935_;
  assign new_n33937_ = ~new_n33932_ & ~new_n33936_;
  assign new_n33938_ = new_n33928_ & new_n33937_;
  assign new_n33939_ = new_n33919_ & new_n33938_;
  assign new_n33940_ = new_n33914_ & new_n33939_;
  assign new_n33941_ = ys__n18472 & ys__n46675;
  assign new_n33942_ = ~ys__n18472 & ~ys__n46675;
  assign new_n33943_ = ~ys__n46620 & ~new_n33942_;
  assign new_n33944_ = ~new_n33941_ & new_n33943_;
  assign new_n33945_ = ys__n18475 & ys__n46676;
  assign new_n33946_ = ~ys__n18475 & ~ys__n46676;
  assign new_n33947_ = ~ys__n46622 & ~new_n33946_;
  assign new_n33948_ = ~new_n33945_ & new_n33947_;
  assign new_n33949_ = ~new_n33944_ & ~new_n33948_;
  assign new_n33950_ = ys__n18478 & ys__n46677;
  assign new_n33951_ = ~ys__n18478 & ~ys__n46677;
  assign new_n33952_ = ~ys__n46624 & ~new_n33951_;
  assign new_n33953_ = ~new_n33950_ & new_n33952_;
  assign new_n33954_ = ys__n18481 & ys__n46678;
  assign new_n33955_ = ~ys__n18481 & ~ys__n46678;
  assign new_n33956_ = ~ys__n46626 & ~new_n33955_;
  assign new_n33957_ = ~new_n33954_ & new_n33956_;
  assign new_n33958_ = ~new_n33953_ & ~new_n33957_;
  assign new_n33959_ = new_n33949_ & new_n33958_;
  assign new_n33960_ = ys__n18460 & ys__n46671;
  assign new_n33961_ = ~ys__n18460 & ~ys__n46671;
  assign new_n33962_ = ~ys__n46612 & ~new_n33961_;
  assign new_n33963_ = ~new_n33960_ & new_n33962_;
  assign new_n33964_ = ys__n18463 & ys__n46672;
  assign new_n33965_ = ~ys__n18463 & ~ys__n46672;
  assign new_n33966_ = ~ys__n46614 & ~new_n33965_;
  assign new_n33967_ = ~new_n33964_ & new_n33966_;
  assign new_n33968_ = ~new_n33963_ & ~new_n33967_;
  assign new_n33969_ = ys__n18466 & ys__n46673;
  assign new_n33970_ = ~ys__n18466 & ~ys__n46673;
  assign new_n33971_ = ~ys__n46616 & ~new_n33970_;
  assign new_n33972_ = ~new_n33969_ & new_n33971_;
  assign new_n33973_ = ys__n18469 & ys__n46674;
  assign new_n33974_ = ~ys__n18469 & ~ys__n46674;
  assign new_n33975_ = ~ys__n46618 & ~new_n33974_;
  assign new_n33976_ = ~new_n33973_ & new_n33975_;
  assign new_n33977_ = ~new_n33972_ & ~new_n33976_;
  assign new_n33978_ = new_n33968_ & new_n33977_;
  assign new_n33979_ = new_n33959_ & new_n33978_;
  assign new_n33980_ = ys__n18496 & ys__n46683;
  assign new_n33981_ = ~ys__n18496 & ~ys__n46683;
  assign new_n33982_ = ~ys__n46636 & ~new_n33981_;
  assign new_n33983_ = ~new_n33980_ & new_n33982_;
  assign new_n33984_ = ys__n18499 & ys__n46684;
  assign new_n33985_ = ~ys__n18499 & ~ys__n46684;
  assign new_n33986_ = ~ys__n46638 & ~new_n33985_;
  assign new_n33987_ = ~new_n33984_ & new_n33986_;
  assign new_n33988_ = ~new_n33983_ & ~new_n33987_;
  assign new_n33989_ = ys__n18502 & ys__n46685;
  assign new_n33990_ = ~ys__n18502 & ~ys__n46685;
  assign new_n33991_ = ~ys__n46640 & ~new_n33990_;
  assign new_n33992_ = ~new_n33989_ & new_n33991_;
  assign new_n33993_ = ys__n18505 & ys__n46686;
  assign new_n33994_ = ~ys__n18505 & ~ys__n46686;
  assign new_n33995_ = ~ys__n46642 & ~new_n33994_;
  assign new_n33996_ = ~new_n33993_ & new_n33995_;
  assign new_n33997_ = ~new_n33992_ & ~new_n33996_;
  assign new_n33998_ = new_n33988_ & new_n33997_;
  assign new_n33999_ = ys__n18484 & ys__n46679;
  assign new_n34000_ = ~ys__n18484 & ~ys__n46679;
  assign new_n34001_ = ~ys__n46628 & ~new_n34000_;
  assign new_n34002_ = ~new_n33999_ & new_n34001_;
  assign new_n34003_ = ys__n18487 & ys__n46680;
  assign new_n34004_ = ~ys__n18487 & ~ys__n46680;
  assign new_n34005_ = ~ys__n46630 & ~new_n34004_;
  assign new_n34006_ = ~new_n34003_ & new_n34005_;
  assign new_n34007_ = ~new_n34002_ & ~new_n34006_;
  assign new_n34008_ = ys__n18490 & ys__n46681;
  assign new_n34009_ = ~ys__n18490 & ~ys__n46681;
  assign new_n34010_ = ~ys__n46632 & ~new_n34009_;
  assign new_n34011_ = ~new_n34008_ & new_n34010_;
  assign new_n34012_ = ys__n18493 & ys__n46682;
  assign new_n34013_ = ~ys__n18493 & ~ys__n46682;
  assign new_n34014_ = ~ys__n46634 & ~new_n34013_;
  assign new_n34015_ = ~new_n34012_ & new_n34014_;
  assign new_n34016_ = ~new_n34011_ & ~new_n34015_;
  assign new_n34017_ = new_n34007_ & new_n34016_;
  assign new_n34018_ = new_n33998_ & new_n34017_;
  assign new_n34019_ = new_n33979_ & new_n34018_;
  assign new_n34020_ = new_n33940_ & new_n34019_;
  assign new_n34021_ = new_n33875_ & new_n34020_;
  assign new_n34022_ = ~new_n33706_ & ~new_n34021_;
  assign new_n34023_ = ~ys__n27496 & ~new_n33706_;
  assign new_n34024_ = ~ys__n27496 & ~new_n34023_;
  assign new_n34025_ = ~ys__n27498 & ~new_n34024_;
  assign new_n34026_ = ~ys__n27498 & ~new_n34025_;
  assign new_n34027_ = new_n34021_ & ~new_n34026_;
  assign ys__n27493 = new_n34022_ | new_n34027_;
  assign new_n34029_ = ys__n26770 & ~new_n27901_;
  assign new_n34030_ = ys__n26770 & ~new_n27837_;
  assign new_n34031_ = ~new_n27853_ & ~new_n34030_;
  assign new_n34032_ = new_n27901_ & ~new_n34031_;
  assign new_n34033_ = ~new_n34029_ & ~new_n34032_;
  assign new_n34034_ = ys__n6126 & ys__n46584;
  assign new_n34035_ = ~ys__n6126 & ~ys__n46584;
  assign new_n34036_ = ~ys__n46554 & ~new_n34035_;
  assign new_n34037_ = ~new_n34034_ & new_n34036_;
  assign new_n34038_ = ys__n6127 & ys__n46585;
  assign new_n34039_ = ~ys__n6127 & ~ys__n46585;
  assign new_n34040_ = ~ys__n46556 & ~new_n34039_;
  assign new_n34041_ = ~new_n34038_ & new_n34040_;
  assign new_n34042_ = ~new_n34037_ & ~new_n34041_;
  assign new_n34043_ = ys__n6129 & ys__n46586;
  assign new_n34044_ = ~ys__n6129 & ~ys__n46586;
  assign new_n34045_ = ~ys__n46558 & ~new_n34044_;
  assign new_n34046_ = ~new_n34043_ & new_n34045_;
  assign new_n34047_ = ys__n6130 & ys__n46587;
  assign new_n34048_ = ~ys__n6130 & ~ys__n46587;
  assign new_n34049_ = ~ys__n46560 & ~new_n34048_;
  assign new_n34050_ = ~new_n34047_ & new_n34049_;
  assign new_n34051_ = ~new_n34046_ & ~new_n34050_;
  assign new_n34052_ = new_n34042_ & new_n34051_;
  assign new_n34053_ = ys__n6120 & ys__n46580;
  assign new_n34054_ = ~ys__n6120 & ~ys__n46580;
  assign new_n34055_ = ~ys__n46546 & ~new_n34054_;
  assign new_n34056_ = ~new_n34053_ & new_n34055_;
  assign new_n34057_ = ys__n6121 & ys__n46581;
  assign new_n34058_ = ~ys__n6121 & ~ys__n46581;
  assign new_n34059_ = ~ys__n46548 & ~new_n34058_;
  assign new_n34060_ = ~new_n34057_ & new_n34059_;
  assign new_n34061_ = ~new_n34056_ & ~new_n34060_;
  assign new_n34062_ = ys__n6123 & ys__n46582;
  assign new_n34063_ = ~ys__n6123 & ~ys__n46582;
  assign new_n34064_ = ~ys__n46550 & ~new_n34063_;
  assign new_n34065_ = ~new_n34062_ & new_n34064_;
  assign new_n34066_ = ys__n6124 & ys__n46583;
  assign new_n34067_ = ~ys__n6124 & ~ys__n46583;
  assign new_n34068_ = ~ys__n46552 & ~new_n34067_;
  assign new_n34069_ = ~new_n34066_ & new_n34068_;
  assign new_n34070_ = ~new_n34065_ & ~new_n34069_;
  assign new_n34071_ = new_n34061_ & new_n34070_;
  assign new_n34072_ = new_n34052_ & new_n34071_;
  assign new_n34073_ = ys__n18448 & ys__n46491;
  assign new_n34074_ = ~ys__n18448 & ~ys__n46491;
  assign new_n34075_ = ~ys__n46428 & ~new_n34074_;
  assign new_n34076_ = ~new_n34073_ & new_n34075_;
  assign new_n34077_ = ys__n18451 & ys__n46492;
  assign new_n34078_ = ~ys__n18451 & ~ys__n46492;
  assign new_n34079_ = ~ys__n46430 & ~new_n34078_;
  assign new_n34080_ = ~new_n34077_ & new_n34079_;
  assign new_n34081_ = ~new_n34076_ & ~new_n34080_;
  assign new_n34082_ = ys__n18454 & ys__n46493;
  assign new_n34083_ = ~ys__n18454 & ~ys__n46493;
  assign new_n34084_ = ~ys__n46432 & ~new_n34083_;
  assign new_n34085_ = ~new_n34082_ & new_n34084_;
  assign new_n34086_ = ys__n18457 & ys__n46494;
  assign new_n34087_ = ~ys__n18457 & ~ys__n46494;
  assign new_n34088_ = ~ys__n46434 & ~new_n34087_;
  assign new_n34089_ = ~new_n34086_ & new_n34088_;
  assign new_n34090_ = ~new_n34085_ & ~new_n34089_;
  assign new_n34091_ = new_n34081_ & new_n34090_;
  assign new_n34092_ = ys__n42 & ys__n46588;
  assign new_n34093_ = ~ys__n42 & ~ys__n46588;
  assign new_n34094_ = ~ys__n46562 & ~new_n34093_;
  assign new_n34095_ = ~new_n34092_ & new_n34094_;
  assign new_n34096_ = ys__n40 & ys__n46589;
  assign new_n34097_ = ~ys__n40 & ~ys__n46589;
  assign new_n34098_ = ~ys__n46564 & ~new_n34097_;
  assign new_n34099_ = ~new_n34096_ & new_n34098_;
  assign new_n34100_ = ~new_n34095_ & ~new_n34099_;
  assign new_n34101_ = ys__n6133 & ys__n46590;
  assign new_n34102_ = ~ys__n6133 & ~ys__n46590;
  assign new_n34103_ = ~ys__n46566 & ~new_n34102_;
  assign new_n34104_ = ~new_n34101_ & new_n34103_;
  assign new_n34105_ = ys__n6134 & ys__n46591;
  assign new_n34106_ = ~ys__n6134 & ~ys__n46591;
  assign new_n34107_ = ~ys__n46568 & ~new_n34106_;
  assign new_n34108_ = ~new_n34105_ & new_n34107_;
  assign new_n34109_ = ~new_n34104_ & ~new_n34108_;
  assign new_n34110_ = new_n34100_ & new_n34109_;
  assign new_n34111_ = new_n34091_ & new_n34110_;
  assign new_n34112_ = new_n34072_ & new_n34111_;
  assign new_n34113_ = ys__n6113 & ys__n46569;
  assign new_n34114_ = ~ys__n6113 & ~ys__n46569;
  assign new_n34115_ = ~ys__n46524 & ~new_n34114_;
  assign new_n34116_ = ~new_n34113_ & new_n34115_;
  assign new_n34117_ = ~ys__n38 & ~ys__n46592;
  assign new_n34118_ = ys__n38 & ys__n46592;
  assign new_n34119_ = ~new_n34117_ & ~new_n34118_;
  assign new_n34120_ = ~new_n33481_ & ~new_n34119_;
  assign new_n34121_ = ~new_n34116_ & new_n34120_;
  assign new_n34122_ = ys__n172 & ys__n46570;
  assign new_n34123_ = ~ys__n172 & ~ys__n46570;
  assign new_n34124_ = ~ys__n46526 & ~new_n34123_;
  assign new_n34125_ = ~new_n34122_ & new_n34124_;
  assign new_n34126_ = ys__n338 & ys__n46571;
  assign new_n34127_ = ~ys__n338 & ~ys__n46571;
  assign new_n34128_ = ~ys__n46528 & ~new_n34127_;
  assign new_n34129_ = ~new_n34126_ & new_n34128_;
  assign new_n34130_ = ~new_n34125_ & ~new_n34129_;
  assign new_n34131_ = new_n34121_ & new_n34130_;
  assign new_n34132_ = ~ys__n28 & ~ys__n46597;
  assign new_n34133_ = ys__n28 & ys__n46597;
  assign new_n34134_ = ~new_n34132_ & ~new_n34133_;
  assign new_n34135_ = ~ys__n26 & ~ys__n46598;
  assign new_n34136_ = ys__n26 & ys__n46598;
  assign new_n34137_ = ~new_n34135_ & ~new_n34136_;
  assign new_n34138_ = ~new_n34134_ & ~new_n34137_;
  assign new_n34139_ = ~ys__n24 & ~ys__n46599;
  assign new_n34140_ = ys__n24 & ys__n46599;
  assign new_n34141_ = ~new_n34139_ & ~new_n34140_;
  assign new_n34142_ = ~ys__n27499 & new_n33482_;
  assign new_n34143_ = ~new_n34141_ & ~new_n34142_;
  assign new_n34144_ = new_n34138_ & new_n34143_;
  assign new_n34145_ = ~ys__n36 & ~ys__n46593;
  assign new_n34146_ = ys__n36 & ys__n46593;
  assign new_n34147_ = ~new_n34145_ & ~new_n34146_;
  assign new_n34148_ = ~ys__n34 & ~ys__n46594;
  assign new_n34149_ = ys__n34 & ys__n46594;
  assign new_n34150_ = ~new_n34148_ & ~new_n34149_;
  assign new_n34151_ = ~new_n34147_ & ~new_n34150_;
  assign new_n34152_ = ~ys__n32 & ~ys__n46595;
  assign new_n34153_ = ys__n32 & ys__n46595;
  assign new_n34154_ = ~new_n34152_ & ~new_n34153_;
  assign new_n34155_ = ~ys__n30 & ~ys__n46596;
  assign new_n34156_ = ys__n30 & ys__n46596;
  assign new_n34157_ = ~new_n34155_ & ~new_n34156_;
  assign new_n34158_ = ~new_n34154_ & ~new_n34157_;
  assign new_n34159_ = new_n34151_ & new_n34158_;
  assign new_n34160_ = new_n34144_ & new_n34159_;
  assign new_n34161_ = new_n34131_ & new_n34160_;
  assign new_n34162_ = ys__n340 & ys__n46576;
  assign new_n34163_ = ~ys__n340 & ~ys__n46576;
  assign new_n34164_ = ~ys__n46538 & ~new_n34163_;
  assign new_n34165_ = ~new_n34162_ & new_n34164_;
  assign new_n34166_ = ys__n46 & ys__n46577;
  assign new_n34167_ = ~ys__n46 & ~ys__n46577;
  assign new_n34168_ = ~ys__n46540 & ~new_n34167_;
  assign new_n34169_ = ~new_n34166_ & new_n34168_;
  assign new_n34170_ = ~new_n34165_ & ~new_n34169_;
  assign new_n34171_ = ys__n6118 & ys__n46578;
  assign new_n34172_ = ~ys__n6118 & ~ys__n46578;
  assign new_n34173_ = ~ys__n46542 & ~new_n34172_;
  assign new_n34174_ = ~new_n34171_ & new_n34173_;
  assign new_n34175_ = ys__n6119 & ys__n46579;
  assign new_n34176_ = ~ys__n6119 & ~ys__n46579;
  assign new_n34177_ = ~ys__n46544 & ~new_n34176_;
  assign new_n34178_ = ~new_n34175_ & new_n34177_;
  assign new_n34179_ = ~new_n34174_ & ~new_n34178_;
  assign new_n34180_ = new_n34170_ & new_n34179_;
  assign new_n34181_ = ys__n22 & ys__n46572;
  assign new_n34182_ = ~ys__n22 & ~ys__n46572;
  assign new_n34183_ = ~ys__n46530 & ~new_n34182_;
  assign new_n34184_ = ~new_n34181_ & new_n34183_;
  assign new_n34185_ = ys__n316 & ys__n46573;
  assign new_n34186_ = ~ys__n316 & ~ys__n46573;
  assign new_n34187_ = ~ys__n46532 & ~new_n34186_;
  assign new_n34188_ = ~new_n34185_ & new_n34187_;
  assign new_n34189_ = ~new_n34184_ & ~new_n34188_;
  assign new_n34190_ = ys__n6115 & ys__n46574;
  assign new_n34191_ = ~ys__n6115 & ~ys__n46574;
  assign new_n34192_ = ~ys__n46534 & ~new_n34191_;
  assign new_n34193_ = ~new_n34190_ & new_n34192_;
  assign new_n34194_ = ys__n44 & ys__n46575;
  assign new_n34195_ = ~ys__n44 & ~ys__n46575;
  assign new_n34196_ = ~ys__n46536 & ~new_n34195_;
  assign new_n34197_ = ~new_n34194_ & new_n34196_;
  assign new_n34198_ = ~new_n34193_ & ~new_n34197_;
  assign new_n34199_ = new_n34189_ & new_n34198_;
  assign new_n34200_ = new_n34180_ & new_n34199_;
  assign new_n34201_ = new_n34161_ & new_n34200_;
  assign new_n34202_ = new_n34112_ & new_n34201_;
  assign new_n34203_ = ys__n18520 & ys__n46515;
  assign new_n34204_ = ~ys__n18520 & ~ys__n46515;
  assign new_n34205_ = ~ys__n46476 & ~new_n34204_;
  assign new_n34206_ = ~new_n34203_ & new_n34205_;
  assign new_n34207_ = ys__n18523 & ys__n46516;
  assign new_n34208_ = ~ys__n18523 & ~ys__n46516;
  assign new_n34209_ = ~ys__n46478 & ~new_n34208_;
  assign new_n34210_ = ~new_n34207_ & new_n34209_;
  assign new_n34211_ = ~new_n34206_ & ~new_n34210_;
  assign new_n34212_ = ys__n18526 & ys__n46517;
  assign new_n34213_ = ~ys__n18526 & ~ys__n46517;
  assign new_n34214_ = ~ys__n46480 & ~new_n34213_;
  assign new_n34215_ = ~new_n34212_ & new_n34214_;
  assign new_n34216_ = ys__n18529 & ys__n46518;
  assign new_n34217_ = ~ys__n18529 & ~ys__n46518;
  assign new_n34218_ = ~ys__n46482 & ~new_n34217_;
  assign new_n34219_ = ~new_n34216_ & new_n34218_;
  assign new_n34220_ = ~new_n34215_ & ~new_n34219_;
  assign new_n34221_ = new_n34211_ & new_n34220_;
  assign new_n34222_ = ys__n18508 & ys__n46511;
  assign new_n34223_ = ~ys__n18508 & ~ys__n46511;
  assign new_n34224_ = ~ys__n46468 & ~new_n34223_;
  assign new_n34225_ = ~new_n34222_ & new_n34224_;
  assign new_n34226_ = ys__n18511 & ys__n46512;
  assign new_n34227_ = ~ys__n18511 & ~ys__n46512;
  assign new_n34228_ = ~ys__n46470 & ~new_n34227_;
  assign new_n34229_ = ~new_n34226_ & new_n34228_;
  assign new_n34230_ = ~new_n34225_ & ~new_n34229_;
  assign new_n34231_ = ys__n18514 & ys__n46513;
  assign new_n34232_ = ~ys__n18514 & ~ys__n46513;
  assign new_n34233_ = ~ys__n46472 & ~new_n34232_;
  assign new_n34234_ = ~new_n34231_ & new_n34233_;
  assign new_n34235_ = ys__n18517 & ys__n46514;
  assign new_n34236_ = ~ys__n18517 & ~ys__n46514;
  assign new_n34237_ = ~ys__n46474 & ~new_n34236_;
  assign new_n34238_ = ~new_n34235_ & new_n34237_;
  assign new_n34239_ = ~new_n34234_ & ~new_n34238_;
  assign new_n34240_ = new_n34230_ & new_n34239_;
  assign new_n34241_ = new_n34221_ & new_n34240_;
  assign new_n34242_ = ~ys__n18047 & new_n33584_;
  assign new_n34243_ = ~ys__n18051 & new_n33587_;
  assign new_n34244_ = ~ys__n18049 & new_n33589_;
  assign new_n34245_ = ~new_n34243_ & ~new_n34244_;
  assign new_n34246_ = ~new_n34242_ & new_n34245_;
  assign new_n34247_ = ys__n18532 & ys__n46519;
  assign new_n34248_ = ~ys__n18532 & ~ys__n46519;
  assign new_n34249_ = ~ys__n46484 & ~new_n34248_;
  assign new_n34250_ = ~new_n34247_ & new_n34249_;
  assign new_n34251_ = ys__n18535 & ys__n46520;
  assign new_n34252_ = ~ys__n18535 & ~ys__n46520;
  assign new_n34253_ = ~ys__n46486 & ~new_n34252_;
  assign new_n34254_ = ~new_n34251_ & new_n34253_;
  assign new_n34255_ = ~new_n34250_ & ~new_n34254_;
  assign new_n34256_ = ys__n18538 & ys__n46521;
  assign new_n34257_ = ~ys__n18538 & ~ys__n46521;
  assign new_n34258_ = ~ys__n46488 & ~new_n34257_;
  assign new_n34259_ = ~new_n34256_ & new_n34258_;
  assign new_n34260_ = ys__n18541 & ys__n46522;
  assign new_n34261_ = ~ys__n18541 & ~ys__n46522;
  assign new_n34262_ = ~ys__n46490 & ~new_n34261_;
  assign new_n34263_ = ~new_n34260_ & new_n34262_;
  assign new_n34264_ = ~new_n34259_ & ~new_n34263_;
  assign new_n34265_ = new_n34255_ & new_n34264_;
  assign new_n34266_ = new_n34246_ & new_n34265_;
  assign new_n34267_ = new_n34241_ & new_n34266_;
  assign new_n34268_ = ys__n18472 & ys__n46499;
  assign new_n34269_ = ~ys__n18472 & ~ys__n46499;
  assign new_n34270_ = ~ys__n46444 & ~new_n34269_;
  assign new_n34271_ = ~new_n34268_ & new_n34270_;
  assign new_n34272_ = ys__n18475 & ys__n46500;
  assign new_n34273_ = ~ys__n18475 & ~ys__n46500;
  assign new_n34274_ = ~ys__n46446 & ~new_n34273_;
  assign new_n34275_ = ~new_n34272_ & new_n34274_;
  assign new_n34276_ = ~new_n34271_ & ~new_n34275_;
  assign new_n34277_ = ys__n18478 & ys__n46501;
  assign new_n34278_ = ~ys__n18478 & ~ys__n46501;
  assign new_n34279_ = ~ys__n46448 & ~new_n34278_;
  assign new_n34280_ = ~new_n34277_ & new_n34279_;
  assign new_n34281_ = ys__n18481 & ys__n46502;
  assign new_n34282_ = ~ys__n18481 & ~ys__n46502;
  assign new_n34283_ = ~ys__n46450 & ~new_n34282_;
  assign new_n34284_ = ~new_n34281_ & new_n34283_;
  assign new_n34285_ = ~new_n34280_ & ~new_n34284_;
  assign new_n34286_ = new_n34276_ & new_n34285_;
  assign new_n34287_ = ys__n18460 & ys__n46495;
  assign new_n34288_ = ~ys__n18460 & ~ys__n46495;
  assign new_n34289_ = ~ys__n46436 & ~new_n34288_;
  assign new_n34290_ = ~new_n34287_ & new_n34289_;
  assign new_n34291_ = ys__n18463 & ys__n46496;
  assign new_n34292_ = ~ys__n18463 & ~ys__n46496;
  assign new_n34293_ = ~ys__n46438 & ~new_n34292_;
  assign new_n34294_ = ~new_n34291_ & new_n34293_;
  assign new_n34295_ = ~new_n34290_ & ~new_n34294_;
  assign new_n34296_ = ys__n18466 & ys__n46497;
  assign new_n34297_ = ~ys__n18466 & ~ys__n46497;
  assign new_n34298_ = ~ys__n46440 & ~new_n34297_;
  assign new_n34299_ = ~new_n34296_ & new_n34298_;
  assign new_n34300_ = ys__n18469 & ys__n46498;
  assign new_n34301_ = ~ys__n18469 & ~ys__n46498;
  assign new_n34302_ = ~ys__n46442 & ~new_n34301_;
  assign new_n34303_ = ~new_n34300_ & new_n34302_;
  assign new_n34304_ = ~new_n34299_ & ~new_n34303_;
  assign new_n34305_ = new_n34295_ & new_n34304_;
  assign new_n34306_ = new_n34286_ & new_n34305_;
  assign new_n34307_ = ys__n18496 & ys__n46507;
  assign new_n34308_ = ~ys__n18496 & ~ys__n46507;
  assign new_n34309_ = ~ys__n46460 & ~new_n34308_;
  assign new_n34310_ = ~new_n34307_ & new_n34309_;
  assign new_n34311_ = ys__n18499 & ys__n46508;
  assign new_n34312_ = ~ys__n18499 & ~ys__n46508;
  assign new_n34313_ = ~ys__n46462 & ~new_n34312_;
  assign new_n34314_ = ~new_n34311_ & new_n34313_;
  assign new_n34315_ = ~new_n34310_ & ~new_n34314_;
  assign new_n34316_ = ys__n18502 & ys__n46509;
  assign new_n34317_ = ~ys__n18502 & ~ys__n46509;
  assign new_n34318_ = ~ys__n46464 & ~new_n34317_;
  assign new_n34319_ = ~new_n34316_ & new_n34318_;
  assign new_n34320_ = ys__n18505 & ys__n46510;
  assign new_n34321_ = ~ys__n18505 & ~ys__n46510;
  assign new_n34322_ = ~ys__n46466 & ~new_n34321_;
  assign new_n34323_ = ~new_n34320_ & new_n34322_;
  assign new_n34324_ = ~new_n34319_ & ~new_n34323_;
  assign new_n34325_ = new_n34315_ & new_n34324_;
  assign new_n34326_ = ys__n18484 & ys__n46503;
  assign new_n34327_ = ~ys__n18484 & ~ys__n46503;
  assign new_n34328_ = ~ys__n46452 & ~new_n34327_;
  assign new_n34329_ = ~new_n34326_ & new_n34328_;
  assign new_n34330_ = ys__n18487 & ys__n46504;
  assign new_n34331_ = ~ys__n18487 & ~ys__n46504;
  assign new_n34332_ = ~ys__n46454 & ~new_n34331_;
  assign new_n34333_ = ~new_n34330_ & new_n34332_;
  assign new_n34334_ = ~new_n34329_ & ~new_n34333_;
  assign new_n34335_ = ys__n18490 & ys__n46505;
  assign new_n34336_ = ~ys__n18490 & ~ys__n46505;
  assign new_n34337_ = ~ys__n46456 & ~new_n34336_;
  assign new_n34338_ = ~new_n34335_ & new_n34337_;
  assign new_n34339_ = ys__n18493 & ys__n46506;
  assign new_n34340_ = ~ys__n18493 & ~ys__n46506;
  assign new_n34341_ = ~ys__n46458 & ~new_n34340_;
  assign new_n34342_ = ~new_n34339_ & new_n34341_;
  assign new_n34343_ = ~new_n34338_ & ~new_n34342_;
  assign new_n34344_ = new_n34334_ & new_n34343_;
  assign new_n34345_ = new_n34325_ & new_n34344_;
  assign new_n34346_ = new_n34306_ & new_n34345_;
  assign new_n34347_ = new_n34267_ & new_n34346_;
  assign new_n34348_ = new_n34202_ & new_n34347_;
  assign new_n34349_ = ~new_n34033_ & ~new_n34348_;
  assign new_n34350_ = ~ys__n27507 & ~new_n34033_;
  assign new_n34351_ = ~ys__n27507 & ~new_n34350_;
  assign new_n34352_ = ~ys__n27509 & ~new_n34351_;
  assign new_n34353_ = ~ys__n27509 & ~new_n34352_;
  assign new_n34354_ = new_n34348_ & ~new_n34353_;
  assign ys__n27504 = new_n34349_ | new_n34354_;
  assign new_n34356_ = ys__n27481 & new_n33694_;
  assign new_n34357_ = ~new_n34021_ & new_n34356_;
  assign new_n34358_ = ~ys__n27496 & new_n34356_;
  assign new_n34359_ = ~ys__n27496 & ~new_n34358_;
  assign new_n34360_ = new_n34021_ & ~new_n34359_;
  assign new_n34361_ = ~new_n34357_ & ~new_n34360_;
  assign new_n34362_ = ~new_n34348_ & ~new_n34361_;
  assign new_n34363_ = ~ys__n27507 & ~new_n34361_;
  assign new_n34364_ = ~ys__n27507 & ~new_n34363_;
  assign new_n34365_ = new_n34348_ & ~new_n34364_;
  assign new_n34366_ = ~new_n34362_ & ~new_n34365_;
  assign new_n34367_ = ys__n6126 & ys__n46408;
  assign new_n34368_ = ~ys__n6126 & ~ys__n46408;
  assign new_n34369_ = ~ys__n46378 & ~new_n34368_;
  assign new_n34370_ = ~new_n34367_ & new_n34369_;
  assign new_n34371_ = ys__n6127 & ys__n46409;
  assign new_n34372_ = ~ys__n6127 & ~ys__n46409;
  assign new_n34373_ = ~ys__n46380 & ~new_n34372_;
  assign new_n34374_ = ~new_n34371_ & new_n34373_;
  assign new_n34375_ = ~new_n34370_ & ~new_n34374_;
  assign new_n34376_ = ys__n6129 & ys__n46410;
  assign new_n34377_ = ~ys__n6129 & ~ys__n46410;
  assign new_n34378_ = ~ys__n46382 & ~new_n34377_;
  assign new_n34379_ = ~new_n34376_ & new_n34378_;
  assign new_n34380_ = ys__n6130 & ys__n46411;
  assign new_n34381_ = ~ys__n6130 & ~ys__n46411;
  assign new_n34382_ = ~ys__n46384 & ~new_n34381_;
  assign new_n34383_ = ~new_n34380_ & new_n34382_;
  assign new_n34384_ = ~new_n34379_ & ~new_n34383_;
  assign new_n34385_ = new_n34375_ & new_n34384_;
  assign new_n34386_ = ys__n6120 & ys__n46404;
  assign new_n34387_ = ~ys__n6120 & ~ys__n46404;
  assign new_n34388_ = ~ys__n46370 & ~new_n34387_;
  assign new_n34389_ = ~new_n34386_ & new_n34388_;
  assign new_n34390_ = ys__n6121 & ys__n46405;
  assign new_n34391_ = ~ys__n6121 & ~ys__n46405;
  assign new_n34392_ = ~ys__n46372 & ~new_n34391_;
  assign new_n34393_ = ~new_n34390_ & new_n34392_;
  assign new_n34394_ = ~new_n34389_ & ~new_n34393_;
  assign new_n34395_ = ys__n6123 & ys__n46406;
  assign new_n34396_ = ~ys__n6123 & ~ys__n46406;
  assign new_n34397_ = ~ys__n46374 & ~new_n34396_;
  assign new_n34398_ = ~new_n34395_ & new_n34397_;
  assign new_n34399_ = ys__n6124 & ys__n46407;
  assign new_n34400_ = ~ys__n6124 & ~ys__n46407;
  assign new_n34401_ = ~ys__n46376 & ~new_n34400_;
  assign new_n34402_ = ~new_n34399_ & new_n34401_;
  assign new_n34403_ = ~new_n34398_ & ~new_n34402_;
  assign new_n34404_ = new_n34394_ & new_n34403_;
  assign new_n34405_ = new_n34385_ & new_n34404_;
  assign new_n34406_ = ys__n18448 & ys__n46315;
  assign new_n34407_ = ~ys__n18448 & ~ys__n46315;
  assign new_n34408_ = ~ys__n46252 & ~new_n34407_;
  assign new_n34409_ = ~new_n34406_ & new_n34408_;
  assign new_n34410_ = ys__n18451 & ys__n46316;
  assign new_n34411_ = ~ys__n18451 & ~ys__n46316;
  assign new_n34412_ = ~ys__n46254 & ~new_n34411_;
  assign new_n34413_ = ~new_n34410_ & new_n34412_;
  assign new_n34414_ = ~new_n34409_ & ~new_n34413_;
  assign new_n34415_ = ys__n18454 & ys__n46317;
  assign new_n34416_ = ~ys__n18454 & ~ys__n46317;
  assign new_n34417_ = ~ys__n46256 & ~new_n34416_;
  assign new_n34418_ = ~new_n34415_ & new_n34417_;
  assign new_n34419_ = ys__n18457 & ys__n46318;
  assign new_n34420_ = ~ys__n18457 & ~ys__n46318;
  assign new_n34421_ = ~ys__n46258 & ~new_n34420_;
  assign new_n34422_ = ~new_n34419_ & new_n34421_;
  assign new_n34423_ = ~new_n34418_ & ~new_n34422_;
  assign new_n34424_ = new_n34414_ & new_n34423_;
  assign new_n34425_ = ys__n42 & ys__n46412;
  assign new_n34426_ = ~ys__n42 & ~ys__n46412;
  assign new_n34427_ = ~ys__n46386 & ~new_n34426_;
  assign new_n34428_ = ~new_n34425_ & new_n34427_;
  assign new_n34429_ = ys__n40 & ys__n46413;
  assign new_n34430_ = ~ys__n40 & ~ys__n46413;
  assign new_n34431_ = ~ys__n46388 & ~new_n34430_;
  assign new_n34432_ = ~new_n34429_ & new_n34431_;
  assign new_n34433_ = ~new_n34428_ & ~new_n34432_;
  assign new_n34434_ = ys__n6133 & ys__n46414;
  assign new_n34435_ = ~ys__n6133 & ~ys__n46414;
  assign new_n34436_ = ~ys__n46390 & ~new_n34435_;
  assign new_n34437_ = ~new_n34434_ & new_n34436_;
  assign new_n34438_ = ys__n6134 & ys__n46415;
  assign new_n34439_ = ~ys__n6134 & ~ys__n46415;
  assign new_n34440_ = ~ys__n46392 & ~new_n34439_;
  assign new_n34441_ = ~new_n34438_ & new_n34440_;
  assign new_n34442_ = ~new_n34437_ & ~new_n34441_;
  assign new_n34443_ = new_n34433_ & new_n34442_;
  assign new_n34444_ = new_n34424_ & new_n34443_;
  assign new_n34445_ = new_n34405_ & new_n34444_;
  assign new_n34446_ = ys__n6113 & ys__n46393;
  assign new_n34447_ = ~ys__n6113 & ~ys__n46393;
  assign new_n34448_ = ~ys__n46348 & ~new_n34447_;
  assign new_n34449_ = ~new_n34446_ & new_n34448_;
  assign new_n34450_ = ~ys__n38 & ~ys__n46416;
  assign new_n34451_ = ys__n38 & ys__n46416;
  assign new_n34452_ = ~new_n34450_ & ~new_n34451_;
  assign new_n34453_ = ~new_n33481_ & ~new_n34452_;
  assign new_n34454_ = ~new_n34449_ & new_n34453_;
  assign new_n34455_ = ys__n172 & ys__n46394;
  assign new_n34456_ = ~ys__n172 & ~ys__n46394;
  assign new_n34457_ = ~ys__n46350 & ~new_n34456_;
  assign new_n34458_ = ~new_n34455_ & new_n34457_;
  assign new_n34459_ = ys__n338 & ys__n46395;
  assign new_n34460_ = ~ys__n338 & ~ys__n46395;
  assign new_n34461_ = ~ys__n46352 & ~new_n34460_;
  assign new_n34462_ = ~new_n34459_ & new_n34461_;
  assign new_n34463_ = ~new_n34458_ & ~new_n34462_;
  assign new_n34464_ = new_n34454_ & new_n34463_;
  assign new_n34465_ = ~ys__n28 & ~ys__n46421;
  assign new_n34466_ = ys__n28 & ys__n46421;
  assign new_n34467_ = ~new_n34465_ & ~new_n34466_;
  assign new_n34468_ = ~ys__n26 & ~ys__n46422;
  assign new_n34469_ = ys__n26 & ys__n46422;
  assign new_n34470_ = ~new_n34468_ & ~new_n34469_;
  assign new_n34471_ = ~new_n34467_ & ~new_n34470_;
  assign new_n34472_ = ~ys__n24 & ~ys__n46423;
  assign new_n34473_ = ys__n24 & ys__n46423;
  assign new_n34474_ = ~new_n34472_ & ~new_n34473_;
  assign new_n34475_ = ~ys__n27510 & new_n33482_;
  assign new_n34476_ = ~new_n34474_ & ~new_n34475_;
  assign new_n34477_ = new_n34471_ & new_n34476_;
  assign new_n34478_ = ~ys__n36 & ~ys__n46417;
  assign new_n34479_ = ys__n36 & ys__n46417;
  assign new_n34480_ = ~new_n34478_ & ~new_n34479_;
  assign new_n34481_ = ~ys__n34 & ~ys__n46418;
  assign new_n34482_ = ys__n34 & ys__n46418;
  assign new_n34483_ = ~new_n34481_ & ~new_n34482_;
  assign new_n34484_ = ~new_n34480_ & ~new_n34483_;
  assign new_n34485_ = ~ys__n32 & ~ys__n46419;
  assign new_n34486_ = ys__n32 & ys__n46419;
  assign new_n34487_ = ~new_n34485_ & ~new_n34486_;
  assign new_n34488_ = ~ys__n30 & ~ys__n46420;
  assign new_n34489_ = ys__n30 & ys__n46420;
  assign new_n34490_ = ~new_n34488_ & ~new_n34489_;
  assign new_n34491_ = ~new_n34487_ & ~new_n34490_;
  assign new_n34492_ = new_n34484_ & new_n34491_;
  assign new_n34493_ = new_n34477_ & new_n34492_;
  assign new_n34494_ = new_n34464_ & new_n34493_;
  assign new_n34495_ = ys__n340 & ys__n46400;
  assign new_n34496_ = ~ys__n340 & ~ys__n46400;
  assign new_n34497_ = ~ys__n46362 & ~new_n34496_;
  assign new_n34498_ = ~new_n34495_ & new_n34497_;
  assign new_n34499_ = ys__n46 & ys__n46401;
  assign new_n34500_ = ~ys__n46 & ~ys__n46401;
  assign new_n34501_ = ~ys__n46364 & ~new_n34500_;
  assign new_n34502_ = ~new_n34499_ & new_n34501_;
  assign new_n34503_ = ~new_n34498_ & ~new_n34502_;
  assign new_n34504_ = ys__n6118 & ys__n46402;
  assign new_n34505_ = ~ys__n6118 & ~ys__n46402;
  assign new_n34506_ = ~ys__n46366 & ~new_n34505_;
  assign new_n34507_ = ~new_n34504_ & new_n34506_;
  assign new_n34508_ = ys__n6119 & ys__n46403;
  assign new_n34509_ = ~ys__n6119 & ~ys__n46403;
  assign new_n34510_ = ~ys__n46368 & ~new_n34509_;
  assign new_n34511_ = ~new_n34508_ & new_n34510_;
  assign new_n34512_ = ~new_n34507_ & ~new_n34511_;
  assign new_n34513_ = new_n34503_ & new_n34512_;
  assign new_n34514_ = ys__n22 & ys__n46396;
  assign new_n34515_ = ~ys__n22 & ~ys__n46396;
  assign new_n34516_ = ~ys__n46354 & ~new_n34515_;
  assign new_n34517_ = ~new_n34514_ & new_n34516_;
  assign new_n34518_ = ys__n316 & ys__n46397;
  assign new_n34519_ = ~ys__n316 & ~ys__n46397;
  assign new_n34520_ = ~ys__n46356 & ~new_n34519_;
  assign new_n34521_ = ~new_n34518_ & new_n34520_;
  assign new_n34522_ = ~new_n34517_ & ~new_n34521_;
  assign new_n34523_ = ys__n6115 & ys__n46398;
  assign new_n34524_ = ~ys__n6115 & ~ys__n46398;
  assign new_n34525_ = ~ys__n46358 & ~new_n34524_;
  assign new_n34526_ = ~new_n34523_ & new_n34525_;
  assign new_n34527_ = ys__n44 & ys__n46399;
  assign new_n34528_ = ~ys__n44 & ~ys__n46399;
  assign new_n34529_ = ~ys__n46360 & ~new_n34528_;
  assign new_n34530_ = ~new_n34527_ & new_n34529_;
  assign new_n34531_ = ~new_n34526_ & ~new_n34530_;
  assign new_n34532_ = new_n34522_ & new_n34531_;
  assign new_n34533_ = new_n34513_ & new_n34532_;
  assign new_n34534_ = new_n34494_ & new_n34533_;
  assign new_n34535_ = new_n34445_ & new_n34534_;
  assign new_n34536_ = ys__n18520 & ys__n46339;
  assign new_n34537_ = ~ys__n18520 & ~ys__n46339;
  assign new_n34538_ = ~ys__n46300 & ~new_n34537_;
  assign new_n34539_ = ~new_n34536_ & new_n34538_;
  assign new_n34540_ = ys__n18523 & ys__n46340;
  assign new_n34541_ = ~ys__n18523 & ~ys__n46340;
  assign new_n34542_ = ~ys__n46302 & ~new_n34541_;
  assign new_n34543_ = ~new_n34540_ & new_n34542_;
  assign new_n34544_ = ~new_n34539_ & ~new_n34543_;
  assign new_n34545_ = ys__n18526 & ys__n46341;
  assign new_n34546_ = ~ys__n18526 & ~ys__n46341;
  assign new_n34547_ = ~ys__n46304 & ~new_n34546_;
  assign new_n34548_ = ~new_n34545_ & new_n34547_;
  assign new_n34549_ = ys__n18529 & ys__n46342;
  assign new_n34550_ = ~ys__n18529 & ~ys__n46342;
  assign new_n34551_ = ~ys__n46306 & ~new_n34550_;
  assign new_n34552_ = ~new_n34549_ & new_n34551_;
  assign new_n34553_ = ~new_n34548_ & ~new_n34552_;
  assign new_n34554_ = new_n34544_ & new_n34553_;
  assign new_n34555_ = ys__n18508 & ys__n46335;
  assign new_n34556_ = ~ys__n18508 & ~ys__n46335;
  assign new_n34557_ = ~ys__n46292 & ~new_n34556_;
  assign new_n34558_ = ~new_n34555_ & new_n34557_;
  assign new_n34559_ = ys__n18511 & ys__n46336;
  assign new_n34560_ = ~ys__n18511 & ~ys__n46336;
  assign new_n34561_ = ~ys__n46294 & ~new_n34560_;
  assign new_n34562_ = ~new_n34559_ & new_n34561_;
  assign new_n34563_ = ~new_n34558_ & ~new_n34562_;
  assign new_n34564_ = ys__n18514 & ys__n46337;
  assign new_n34565_ = ~ys__n18514 & ~ys__n46337;
  assign new_n34566_ = ~ys__n46296 & ~new_n34565_;
  assign new_n34567_ = ~new_n34564_ & new_n34566_;
  assign new_n34568_ = ys__n18517 & ys__n46338;
  assign new_n34569_ = ~ys__n18517 & ~ys__n46338;
  assign new_n34570_ = ~ys__n46298 & ~new_n34569_;
  assign new_n34571_ = ~new_n34568_ & new_n34570_;
  assign new_n34572_ = ~new_n34567_ & ~new_n34571_;
  assign new_n34573_ = new_n34563_ & new_n34572_;
  assign new_n34574_ = new_n34554_ & new_n34573_;
  assign new_n34575_ = ~ys__n18041 & new_n33584_;
  assign new_n34576_ = ~ys__n18045 & new_n33587_;
  assign new_n34577_ = ~ys__n18043 & new_n33589_;
  assign new_n34578_ = ~new_n34576_ & ~new_n34577_;
  assign new_n34579_ = ~new_n34575_ & new_n34578_;
  assign new_n34580_ = ys__n18532 & ys__n46343;
  assign new_n34581_ = ~ys__n18532 & ~ys__n46343;
  assign new_n34582_ = ~ys__n46308 & ~new_n34581_;
  assign new_n34583_ = ~new_n34580_ & new_n34582_;
  assign new_n34584_ = ys__n18535 & ys__n46344;
  assign new_n34585_ = ~ys__n18535 & ~ys__n46344;
  assign new_n34586_ = ~ys__n46310 & ~new_n34585_;
  assign new_n34587_ = ~new_n34584_ & new_n34586_;
  assign new_n34588_ = ~new_n34583_ & ~new_n34587_;
  assign new_n34589_ = ys__n18538 & ys__n46345;
  assign new_n34590_ = ~ys__n18538 & ~ys__n46345;
  assign new_n34591_ = ~ys__n46312 & ~new_n34590_;
  assign new_n34592_ = ~new_n34589_ & new_n34591_;
  assign new_n34593_ = ys__n18541 & ys__n46346;
  assign new_n34594_ = ~ys__n18541 & ~ys__n46346;
  assign new_n34595_ = ~ys__n46314 & ~new_n34594_;
  assign new_n34596_ = ~new_n34593_ & new_n34595_;
  assign new_n34597_ = ~new_n34592_ & ~new_n34596_;
  assign new_n34598_ = new_n34588_ & new_n34597_;
  assign new_n34599_ = new_n34579_ & new_n34598_;
  assign new_n34600_ = new_n34574_ & new_n34599_;
  assign new_n34601_ = ys__n18472 & ys__n46323;
  assign new_n34602_ = ~ys__n18472 & ~ys__n46323;
  assign new_n34603_ = ~ys__n46268 & ~new_n34602_;
  assign new_n34604_ = ~new_n34601_ & new_n34603_;
  assign new_n34605_ = ys__n18475 & ys__n46324;
  assign new_n34606_ = ~ys__n18475 & ~ys__n46324;
  assign new_n34607_ = ~ys__n46270 & ~new_n34606_;
  assign new_n34608_ = ~new_n34605_ & new_n34607_;
  assign new_n34609_ = ~new_n34604_ & ~new_n34608_;
  assign new_n34610_ = ys__n18478 & ys__n46325;
  assign new_n34611_ = ~ys__n18478 & ~ys__n46325;
  assign new_n34612_ = ~ys__n46272 & ~new_n34611_;
  assign new_n34613_ = ~new_n34610_ & new_n34612_;
  assign new_n34614_ = ys__n18481 & ys__n46326;
  assign new_n34615_ = ~ys__n18481 & ~ys__n46326;
  assign new_n34616_ = ~ys__n46274 & ~new_n34615_;
  assign new_n34617_ = ~new_n34614_ & new_n34616_;
  assign new_n34618_ = ~new_n34613_ & ~new_n34617_;
  assign new_n34619_ = new_n34609_ & new_n34618_;
  assign new_n34620_ = ys__n18460 & ys__n46319;
  assign new_n34621_ = ~ys__n18460 & ~ys__n46319;
  assign new_n34622_ = ~ys__n46260 & ~new_n34621_;
  assign new_n34623_ = ~new_n34620_ & new_n34622_;
  assign new_n34624_ = ys__n18463 & ys__n46320;
  assign new_n34625_ = ~ys__n18463 & ~ys__n46320;
  assign new_n34626_ = ~ys__n46262 & ~new_n34625_;
  assign new_n34627_ = ~new_n34624_ & new_n34626_;
  assign new_n34628_ = ~new_n34623_ & ~new_n34627_;
  assign new_n34629_ = ys__n18466 & ys__n46321;
  assign new_n34630_ = ~ys__n18466 & ~ys__n46321;
  assign new_n34631_ = ~ys__n46264 & ~new_n34630_;
  assign new_n34632_ = ~new_n34629_ & new_n34631_;
  assign new_n34633_ = ys__n18469 & ys__n46322;
  assign new_n34634_ = ~ys__n18469 & ~ys__n46322;
  assign new_n34635_ = ~ys__n46266 & ~new_n34634_;
  assign new_n34636_ = ~new_n34633_ & new_n34635_;
  assign new_n34637_ = ~new_n34632_ & ~new_n34636_;
  assign new_n34638_ = new_n34628_ & new_n34637_;
  assign new_n34639_ = new_n34619_ & new_n34638_;
  assign new_n34640_ = ys__n18496 & ys__n46331;
  assign new_n34641_ = ~ys__n18496 & ~ys__n46331;
  assign new_n34642_ = ~ys__n46284 & ~new_n34641_;
  assign new_n34643_ = ~new_n34640_ & new_n34642_;
  assign new_n34644_ = ys__n18499 & ys__n46332;
  assign new_n34645_ = ~ys__n18499 & ~ys__n46332;
  assign new_n34646_ = ~ys__n46286 & ~new_n34645_;
  assign new_n34647_ = ~new_n34644_ & new_n34646_;
  assign new_n34648_ = ~new_n34643_ & ~new_n34647_;
  assign new_n34649_ = ys__n18502 & ys__n46333;
  assign new_n34650_ = ~ys__n18502 & ~ys__n46333;
  assign new_n34651_ = ~ys__n46288 & ~new_n34650_;
  assign new_n34652_ = ~new_n34649_ & new_n34651_;
  assign new_n34653_ = ys__n18505 & ys__n46334;
  assign new_n34654_ = ~ys__n18505 & ~ys__n46334;
  assign new_n34655_ = ~ys__n46290 & ~new_n34654_;
  assign new_n34656_ = ~new_n34653_ & new_n34655_;
  assign new_n34657_ = ~new_n34652_ & ~new_n34656_;
  assign new_n34658_ = new_n34648_ & new_n34657_;
  assign new_n34659_ = ys__n18484 & ys__n46327;
  assign new_n34660_ = ~ys__n18484 & ~ys__n46327;
  assign new_n34661_ = ~ys__n46276 & ~new_n34660_;
  assign new_n34662_ = ~new_n34659_ & new_n34661_;
  assign new_n34663_ = ys__n18487 & ys__n46328;
  assign new_n34664_ = ~ys__n18487 & ~ys__n46328;
  assign new_n34665_ = ~ys__n46278 & ~new_n34664_;
  assign new_n34666_ = ~new_n34663_ & new_n34665_;
  assign new_n34667_ = ~new_n34662_ & ~new_n34666_;
  assign new_n34668_ = ys__n18490 & ys__n46329;
  assign new_n34669_ = ~ys__n18490 & ~ys__n46329;
  assign new_n34670_ = ~ys__n46280 & ~new_n34669_;
  assign new_n34671_ = ~new_n34668_ & new_n34670_;
  assign new_n34672_ = ys__n18493 & ys__n46330;
  assign new_n34673_ = ~ys__n18493 & ~ys__n46330;
  assign new_n34674_ = ~ys__n46282 & ~new_n34673_;
  assign new_n34675_ = ~new_n34672_ & new_n34674_;
  assign new_n34676_ = ~new_n34671_ & ~new_n34675_;
  assign new_n34677_ = new_n34667_ & new_n34676_;
  assign new_n34678_ = new_n34658_ & new_n34677_;
  assign new_n34679_ = new_n34639_ & new_n34678_;
  assign new_n34680_ = new_n34600_ & new_n34679_;
  assign new_n34681_ = new_n34535_ & new_n34680_;
  assign new_n34682_ = ~new_n34366_ & ~new_n34681_;
  assign new_n34683_ = ~ys__n27518 & ~new_n34366_;
  assign new_n34684_ = ~ys__n27518 & ~new_n34683_;
  assign new_n34685_ = new_n34681_ & ~new_n34684_;
  assign ys__n27513 = new_n34682_ | new_n34685_;
  assign new_n34687_ = ys__n26772 & ~new_n27901_;
  assign new_n34688_ = ys__n26772 & ~new_n27837_;
  assign new_n34689_ = ~new_n27860_ & ~new_n34688_;
  assign new_n34690_ = new_n27901_ & ~new_n34689_;
  assign new_n34691_ = ~new_n34687_ & ~new_n34690_;
  assign new_n34692_ = ~new_n34681_ & ~new_n34691_;
  assign new_n34693_ = ~ys__n27518 & ~new_n34691_;
  assign new_n34694_ = ~ys__n27518 & ~new_n34693_;
  assign new_n34695_ = ~ys__n27520 & ~new_n34694_;
  assign new_n34696_ = ~ys__n27520 & ~new_n34695_;
  assign new_n34697_ = new_n34681_ & ~new_n34696_;
  assign ys__n27515 = new_n34692_ | new_n34697_;
  assign new_n34699_ = ys__n27485 & new_n33694_;
  assign new_n34700_ = ~new_n34021_ & new_n34699_;
  assign new_n34701_ = ~ys__n27498 & new_n34699_;
  assign new_n34702_ = ~ys__n27498 & ~new_n34701_;
  assign new_n34703_ = new_n34021_ & ~new_n34702_;
  assign new_n34704_ = ~new_n34700_ & ~new_n34703_;
  assign new_n34705_ = ~new_n34348_ & ~new_n34704_;
  assign new_n34706_ = ~ys__n27509 & ~new_n34704_;
  assign new_n34707_ = ~ys__n27509 & ~new_n34706_;
  assign new_n34708_ = new_n34348_ & ~new_n34707_;
  assign new_n34709_ = ~new_n34705_ & ~new_n34708_;
  assign new_n34710_ = ~new_n34681_ & ~new_n34709_;
  assign new_n34711_ = ~ys__n27520 & ~new_n34709_;
  assign new_n34712_ = ~ys__n27520 & ~new_n34711_;
  assign new_n34713_ = new_n34681_ & ~new_n34712_;
  assign ys__n27517 = new_n34710_ | new_n34713_;
  assign new_n34715_ = ys__n874 & ys__n18214;
  assign new_n34716_ = ys__n874 & ys__n18218;
  assign new_n34717_ = new_n34715_ & ~new_n34716_;
  assign new_n34718_ = ys__n18217 & new_n34715_;
  assign new_n34719_ = new_n34716_ & new_n34718_;
  assign ys__n27550 = new_n34717_ | new_n34719_;
  assign new_n34721_ = ~ys__n18217 & ~new_n34716_;
  assign new_n34722_ = ys__n18217 & new_n34716_;
  assign ys__n27551 = new_n34721_ | new_n34722_;
  assign new_n34724_ = ~ys__n18393 & ys__n27737;
  assign new_n34725_ = ys__n828 & ys__n18393;
  assign ys__n27598 = new_n34724_ | new_n34725_;
  assign new_n34727_ = ~ys__n18317 & new_n13228_;
  assign new_n34728_ = ys__n18317 & new_n13233_;
  assign new_n34729_ = ~new_n34727_ & ~new_n34728_;
  assign new_n34730_ = ys__n18065 & ~new_n34729_;
  assign new_n34731_ = ys__n27607 & ~new_n34730_;
  assign new_n34732_ = ys__n27608 & new_n34730_;
  assign ys__n27610 = new_n34731_ | new_n34732_;
  assign new_n34734_ = ys__n27611 & ~new_n34730_;
  assign new_n34735_ = ys__n27612 & new_n34730_;
  assign ys__n27613 = new_n34734_ | new_n34735_;
  assign new_n34737_ = ys__n27614 & ~new_n34730_;
  assign new_n34738_ = ys__n27615 & new_n34730_;
  assign ys__n27616 = new_n34737_ | new_n34738_;
  assign new_n34740_ = ys__n27617 & ~new_n34730_;
  assign new_n34741_ = ys__n27618 & new_n34730_;
  assign ys__n27619 = new_n34740_ | new_n34741_;
  assign new_n34743_ = ys__n27620 & ~new_n34730_;
  assign new_n34744_ = ys__n27621 & new_n34730_;
  assign ys__n27622 = new_n34743_ | new_n34744_;
  assign new_n34746_ = ys__n27623 & ~new_n34730_;
  assign new_n34747_ = ys__n27624 & new_n34730_;
  assign ys__n27625 = new_n34746_ | new_n34747_;
  assign new_n34749_ = ys__n27626 & ~new_n34730_;
  assign new_n34750_ = ys__n27627 & new_n34730_;
  assign ys__n27628 = new_n34749_ | new_n34750_;
  assign new_n34752_ = ys__n27629 & ~new_n34730_;
  assign new_n34753_ = ys__n27630 & new_n34730_;
  assign ys__n27631 = new_n34752_ | new_n34753_;
  assign new_n34755_ = ys__n27632 & ~new_n34730_;
  assign new_n34756_ = ys__n27633 & new_n34730_;
  assign ys__n27634 = new_n34755_ | new_n34756_;
  assign new_n34758_ = ys__n27635 & ~new_n34730_;
  assign new_n34759_ = ys__n27636 & new_n34730_;
  assign ys__n27637 = new_n34758_ | new_n34759_;
  assign new_n34761_ = ys__n27638 & ~new_n34730_;
  assign new_n34762_ = ys__n27639 & new_n34730_;
  assign ys__n27640 = new_n34761_ | new_n34762_;
  assign new_n34764_ = ys__n27641 & ~new_n34730_;
  assign new_n34765_ = ys__n27642 & new_n34730_;
  assign ys__n27643 = new_n34764_ | new_n34765_;
  assign new_n34767_ = ys__n27644 & ~new_n34730_;
  assign new_n34768_ = ys__n27645 & new_n34730_;
  assign ys__n27646 = new_n34767_ | new_n34768_;
  assign new_n34770_ = ys__n27647 & ~new_n34730_;
  assign new_n34771_ = ys__n27648 & new_n34730_;
  assign ys__n27649 = new_n34770_ | new_n34771_;
  assign new_n34773_ = ys__n27650 & ~new_n34730_;
  assign new_n34774_ = ys__n27651 & new_n34730_;
  assign ys__n27652 = new_n34773_ | new_n34774_;
  assign new_n34776_ = ys__n27653 & ~new_n34730_;
  assign new_n34777_ = ys__n27654 & new_n34730_;
  assign ys__n27655 = new_n34776_ | new_n34777_;
  assign new_n34779_ = ys__n27656 & ~new_n34730_;
  assign new_n34780_ = ys__n27657 & new_n34730_;
  assign ys__n27658 = new_n34779_ | new_n34780_;
  assign new_n34782_ = ys__n27659 & ~new_n34730_;
  assign new_n34783_ = ys__n27660 & new_n34730_;
  assign ys__n27661 = new_n34782_ | new_n34783_;
  assign new_n34785_ = ys__n27662 & ~new_n34730_;
  assign new_n34786_ = ys__n27663 & new_n34730_;
  assign ys__n27664 = new_n34785_ | new_n34786_;
  assign new_n34788_ = ys__n27665 & ~new_n34730_;
  assign new_n34789_ = ys__n27666 & new_n34730_;
  assign ys__n27667 = new_n34788_ | new_n34789_;
  assign new_n34791_ = ys__n27668 & ~new_n34730_;
  assign new_n34792_ = ys__n27669 & new_n34730_;
  assign ys__n27670 = new_n34791_ | new_n34792_;
  assign new_n34794_ = ys__n27671 & ~new_n34730_;
  assign new_n34795_ = ys__n27672 & new_n34730_;
  assign ys__n27673 = new_n34794_ | new_n34795_;
  assign new_n34797_ = ys__n27674 & ~new_n34730_;
  assign new_n34798_ = ys__n27675 & new_n34730_;
  assign ys__n27676 = new_n34797_ | new_n34798_;
  assign new_n34800_ = ys__n27677 & ~new_n34730_;
  assign new_n34801_ = ys__n27678 & new_n34730_;
  assign ys__n27679 = new_n34800_ | new_n34801_;
  assign new_n34803_ = ys__n27680 & ~new_n34730_;
  assign new_n34804_ = ys__n27681 & new_n34730_;
  assign ys__n27682 = new_n34803_ | new_n34804_;
  assign new_n34806_ = ys__n27683 & ~new_n34730_;
  assign new_n34807_ = ys__n27684 & new_n34730_;
  assign ys__n27685 = new_n34806_ | new_n34807_;
  assign new_n34809_ = ys__n27686 & ~new_n34730_;
  assign new_n34810_ = ys__n27687 & new_n34730_;
  assign ys__n27688 = new_n34809_ | new_n34810_;
  assign new_n34812_ = ys__n27689 & ~new_n34730_;
  assign new_n34813_ = ys__n27690 & new_n34730_;
  assign ys__n27691 = new_n34812_ | new_n34813_;
  assign new_n34815_ = ys__n27692 & ~new_n34730_;
  assign new_n34816_ = ys__n27693 & new_n34730_;
  assign ys__n27694 = new_n34815_ | new_n34816_;
  assign new_n34818_ = ys__n27695 & ~new_n34730_;
  assign new_n34819_ = ys__n27696 & new_n34730_;
  assign ys__n27697 = new_n34818_ | new_n34819_;
  assign new_n34821_ = ys__n27698 & ~new_n34730_;
  assign new_n34822_ = ys__n27699 & new_n34730_;
  assign ys__n27700 = new_n34821_ | new_n34822_;
  assign new_n34824_ = ys__n27701 & ~new_n34730_;
  assign new_n34825_ = ys__n27702 & new_n34730_;
  assign ys__n27703 = new_n34824_ | new_n34825_;
  assign new_n34827_ = ~ys__n18065 & ~new_n34729_;
  assign new_n34828_ = ys__n27607 & ~new_n34827_;
  assign new_n34829_ = ys__n27608 & new_n34827_;
  assign ys__n27705 = new_n34828_ | new_n34829_;
  assign new_n34831_ = ys__n27611 & ~new_n34827_;
  assign new_n34832_ = ys__n27612 & new_n34827_;
  assign ys__n27706 = new_n34831_ | new_n34832_;
  assign new_n34834_ = ys__n27614 & ~new_n34827_;
  assign new_n34835_ = ys__n27615 & new_n34827_;
  assign ys__n27707 = new_n34834_ | new_n34835_;
  assign new_n34837_ = ys__n27617 & ~new_n34827_;
  assign new_n34838_ = ys__n27618 & new_n34827_;
  assign ys__n27708 = new_n34837_ | new_n34838_;
  assign new_n34840_ = ys__n27620 & ~new_n34827_;
  assign new_n34841_ = ys__n27621 & new_n34827_;
  assign ys__n27709 = new_n34840_ | new_n34841_;
  assign new_n34843_ = ys__n27623 & ~new_n34827_;
  assign new_n34844_ = ys__n27624 & new_n34827_;
  assign ys__n27710 = new_n34843_ | new_n34844_;
  assign new_n34846_ = ys__n27626 & ~new_n34827_;
  assign new_n34847_ = ys__n27627 & new_n34827_;
  assign ys__n27711 = new_n34846_ | new_n34847_;
  assign new_n34849_ = ys__n27629 & ~new_n34827_;
  assign new_n34850_ = ys__n27630 & new_n34827_;
  assign ys__n27712 = new_n34849_ | new_n34850_;
  assign new_n34852_ = ys__n27632 & ~new_n34827_;
  assign new_n34853_ = ys__n27633 & new_n34827_;
  assign ys__n27713 = new_n34852_ | new_n34853_;
  assign new_n34855_ = ys__n27635 & ~new_n34827_;
  assign new_n34856_ = ys__n27636 & new_n34827_;
  assign ys__n27714 = new_n34855_ | new_n34856_;
  assign new_n34858_ = ys__n27638 & ~new_n34827_;
  assign new_n34859_ = ys__n27639 & new_n34827_;
  assign ys__n27715 = new_n34858_ | new_n34859_;
  assign new_n34861_ = ys__n27641 & ~new_n34827_;
  assign new_n34862_ = ys__n27642 & new_n34827_;
  assign ys__n27716 = new_n34861_ | new_n34862_;
  assign new_n34864_ = ys__n27644 & ~new_n34827_;
  assign new_n34865_ = ys__n27645 & new_n34827_;
  assign ys__n27717 = new_n34864_ | new_n34865_;
  assign new_n34867_ = ys__n27647 & ~new_n34827_;
  assign new_n34868_ = ys__n27648 & new_n34827_;
  assign ys__n27718 = new_n34867_ | new_n34868_;
  assign new_n34870_ = ys__n27650 & ~new_n34827_;
  assign new_n34871_ = ys__n27651 & new_n34827_;
  assign ys__n27719 = new_n34870_ | new_n34871_;
  assign new_n34873_ = ys__n27653 & ~new_n34827_;
  assign new_n34874_ = ys__n27654 & new_n34827_;
  assign ys__n27720 = new_n34873_ | new_n34874_;
  assign new_n34876_ = ys__n27656 & ~new_n34827_;
  assign new_n34877_ = ys__n27657 & new_n34827_;
  assign ys__n27721 = new_n34876_ | new_n34877_;
  assign new_n34879_ = ys__n27659 & ~new_n34827_;
  assign new_n34880_ = ys__n27660 & new_n34827_;
  assign ys__n27722 = new_n34879_ | new_n34880_;
  assign new_n34882_ = ys__n27662 & ~new_n34827_;
  assign new_n34883_ = ys__n27663 & new_n34827_;
  assign ys__n27723 = new_n34882_ | new_n34883_;
  assign new_n34885_ = ys__n27665 & ~new_n34827_;
  assign new_n34886_ = ys__n27666 & new_n34827_;
  assign ys__n27724 = new_n34885_ | new_n34886_;
  assign new_n34888_ = ys__n27668 & ~new_n34827_;
  assign new_n34889_ = ys__n27669 & new_n34827_;
  assign ys__n27725 = new_n34888_ | new_n34889_;
  assign new_n34891_ = ys__n27671 & ~new_n34827_;
  assign new_n34892_ = ys__n27672 & new_n34827_;
  assign ys__n27726 = new_n34891_ | new_n34892_;
  assign new_n34894_ = ys__n27674 & ~new_n34827_;
  assign new_n34895_ = ys__n27675 & new_n34827_;
  assign ys__n27727 = new_n34894_ | new_n34895_;
  assign new_n34897_ = ys__n27677 & ~new_n34827_;
  assign new_n34898_ = ys__n27678 & new_n34827_;
  assign ys__n27728 = new_n34897_ | new_n34898_;
  assign new_n34900_ = ys__n27680 & ~new_n34827_;
  assign new_n34901_ = ys__n27681 & new_n34827_;
  assign ys__n27729 = new_n34900_ | new_n34901_;
  assign new_n34903_ = ys__n27683 & ~new_n34827_;
  assign new_n34904_ = ys__n27684 & new_n34827_;
  assign ys__n27730 = new_n34903_ | new_n34904_;
  assign new_n34906_ = ys__n27686 & ~new_n34827_;
  assign new_n34907_ = ys__n27687 & new_n34827_;
  assign ys__n27731 = new_n34906_ | new_n34907_;
  assign new_n34909_ = ys__n27689 & ~new_n34827_;
  assign new_n34910_ = ys__n27690 & new_n34827_;
  assign ys__n27732 = new_n34909_ | new_n34910_;
  assign new_n34912_ = ys__n27692 & ~new_n34827_;
  assign new_n34913_ = ys__n27693 & new_n34827_;
  assign ys__n27733 = new_n34912_ | new_n34913_;
  assign new_n34915_ = ys__n27695 & ~new_n34827_;
  assign new_n34916_ = ys__n27696 & new_n34827_;
  assign ys__n27734 = new_n34915_ | new_n34916_;
  assign new_n34918_ = ys__n27698 & ~new_n34827_;
  assign new_n34919_ = ys__n27699 & new_n34827_;
  assign ys__n27735 = new_n34918_ | new_n34919_;
  assign new_n34921_ = ys__n27701 & ~new_n34827_;
  assign new_n34922_ = ys__n27702 & new_n34827_;
  assign ys__n27736 = new_n34921_ | new_n34922_;
  assign ys__n27739 = ~ys__n35065 & ~new_n12275_;
  assign new_n34925_ = ~ys__n18393 & ys__n27739;
  assign new_n34926_ = ys__n18393 & ys__n27740;
  assign ys__n27741 = new_n34925_ | new_n34926_;
  assign ys__n28258 = ~ys__n1535 & ys__n28243;
  assign ys__n28276 = ys__n1535 & ys__n28243;
  assign new_n34930_ = ys__n240 & ~ys__n1535;
  assign new_n34931_ = ~ys__n1535 & ~new_n34930_;
  assign ys__n28328 = ys__n28243 & ~new_n34931_;
  assign new_n34933_ = ys__n238 & ~ys__n1535;
  assign new_n34934_ = ~ys__n1535 & ~new_n34933_;
  assign ys__n28330 = ys__n28243 & ~new_n34934_;
  assign new_n34936_ = ys__n242 & ~ys__n1535;
  assign new_n34937_ = ~ys__n1535 & ~new_n34936_;
  assign ys__n28332 = ys__n28243 & ~new_n34937_;
  assign new_n34939_ = ~ys__n238 & ~ys__n242;
  assign new_n34940_ = ~ys__n1535 & new_n34939_;
  assign new_n34941_ = ~ys__n1535 & ~new_n34940_;
  assign ys__n28336 = ys__n28243 & ~new_n34941_;
  assign new_n34943_ = ys__n758 & ~ys__n760;
  assign new_n34944_ = ~ys__n762 & ~ys__n764;
  assign new_n34945_ = new_n34943_ & new_n34944_;
  assign new_n34946_ = ~ys__n766 & ys__n38198;
  assign new_n34947_ = new_n34945_ & new_n34946_;
  assign ys__n28343 = ~ys__n4566 & new_n34947_;
  assign new_n34949_ = ~ys__n758 & ys__n760;
  assign new_n34950_ = new_n34944_ & new_n34949_;
  assign new_n34951_ = new_n34946_ & new_n34950_;
  assign ys__n28345 = ~ys__n4566 & new_n34951_;
  assign new_n34953_ = ys__n758 & ys__n760;
  assign new_n34954_ = new_n34944_ & new_n34953_;
  assign new_n34955_ = new_n34946_ & new_n34954_;
  assign ys__n28347 = ~ys__n4566 & new_n34955_;
  assign new_n34957_ = ~ys__n758 & ~ys__n760;
  assign new_n34958_ = ys__n762 & ~ys__n764;
  assign new_n34959_ = new_n34957_ & new_n34958_;
  assign new_n34960_ = new_n34946_ & new_n34959_;
  assign ys__n28349 = ~ys__n4566 & new_n34960_;
  assign new_n34962_ = new_n34943_ & new_n34958_;
  assign new_n34963_ = new_n34946_ & new_n34962_;
  assign ys__n28351 = ~ys__n4566 & new_n34963_;
  assign new_n34965_ = new_n34949_ & new_n34958_;
  assign new_n34966_ = new_n34946_ & new_n34965_;
  assign ys__n28353 = ~ys__n4566 & new_n34966_;
  assign new_n34968_ = new_n34953_ & new_n34958_;
  assign new_n34969_ = new_n34946_ & new_n34968_;
  assign ys__n28355 = ~ys__n4566 & new_n34969_;
  assign new_n34971_ = ~ys__n762 & ys__n764;
  assign new_n34972_ = new_n34957_ & new_n34971_;
  assign new_n34973_ = new_n34946_ & new_n34972_;
  assign ys__n28357 = ~ys__n4566 & new_n34973_;
  assign new_n34975_ = new_n34943_ & new_n34971_;
  assign new_n34976_ = new_n34946_ & new_n34975_;
  assign ys__n28359 = ~ys__n4566 & new_n34976_;
  assign new_n34978_ = new_n34949_ & new_n34971_;
  assign new_n34979_ = new_n34946_ & new_n34978_;
  assign ys__n28361 = ~ys__n4566 & new_n34979_;
  assign new_n34981_ = new_n34953_ & new_n34971_;
  assign new_n34982_ = new_n34946_ & new_n34981_;
  assign ys__n28363 = ~ys__n4566 & new_n34982_;
  assign new_n34984_ = ys__n762 & ys__n764;
  assign new_n34985_ = new_n34957_ & new_n34984_;
  assign new_n34986_ = new_n34946_ & new_n34985_;
  assign ys__n28365 = ~ys__n4566 & new_n34986_;
  assign new_n34988_ = new_n34943_ & new_n34984_;
  assign new_n34989_ = new_n34946_ & new_n34988_;
  assign ys__n28367 = ~ys__n4566 & new_n34989_;
  assign new_n34991_ = new_n34949_ & new_n34984_;
  assign new_n34992_ = new_n34946_ & new_n34991_;
  assign ys__n28369 = ~ys__n4566 & new_n34992_;
  assign new_n34994_ = new_n34953_ & new_n34984_;
  assign new_n34995_ = new_n34946_ & new_n34994_;
  assign ys__n28371 = ~ys__n4566 & new_n34995_;
  assign new_n34997_ = ys__n766 & ys__n38198;
  assign new_n34998_ = new_n34944_ & new_n34997_;
  assign new_n34999_ = new_n34957_ & new_n34998_;
  assign ys__n28373 = ~ys__n4566 & new_n34999_;
  assign new_n35001_ = new_n34945_ & new_n34997_;
  assign ys__n28375 = ~ys__n4566 & new_n35001_;
  assign new_n35003_ = new_n34950_ & new_n34997_;
  assign ys__n28377 = ~ys__n4566 & new_n35003_;
  assign new_n35005_ = new_n34954_ & new_n34997_;
  assign ys__n28379 = ~ys__n4566 & new_n35005_;
  assign new_n35007_ = new_n34959_ & new_n34997_;
  assign ys__n28381 = ~ys__n4566 & new_n35007_;
  assign new_n35009_ = new_n34962_ & new_n34997_;
  assign ys__n28383 = ~ys__n4566 & new_n35009_;
  assign new_n35011_ = new_n34965_ & new_n34997_;
  assign ys__n28385 = ~ys__n4566 & new_n35011_;
  assign new_n35013_ = new_n34968_ & new_n34997_;
  assign ys__n28387 = ~ys__n4566 & new_n35013_;
  assign new_n35015_ = new_n34972_ & new_n34997_;
  assign ys__n28389 = ~ys__n4566 & new_n35015_;
  assign new_n35017_ = new_n34975_ & new_n34997_;
  assign ys__n28391 = ~ys__n4566 & new_n35017_;
  assign new_n35019_ = new_n34978_ & new_n34997_;
  assign ys__n28393 = ~ys__n4566 & new_n35019_;
  assign new_n35021_ = new_n34981_ & new_n34997_;
  assign ys__n28395 = ~ys__n4566 & new_n35021_;
  assign new_n35023_ = new_n34985_ & new_n34997_;
  assign ys__n28397 = ~ys__n4566 & new_n35023_;
  assign new_n35025_ = new_n34988_ & new_n34997_;
  assign ys__n28399 = ~ys__n4566 & new_n35025_;
  assign new_n35027_ = new_n34991_ & new_n34997_;
  assign ys__n28401 = ~ys__n4566 & new_n35027_;
  assign new_n35029_ = new_n34994_ & new_n34997_;
  assign ys__n28403 = ~ys__n4566 & new_n35029_;
  assign new_n35031_ = ~new_n15018_ & new_n15044_;
  assign new_n35032_ = new_n15018_ & new_n15051_;
  assign ys__n28406 = new_n35031_ | new_n35032_;
  assign new_n35034_ = ~ys__n738 & new_n15021_;
  assign new_n35035_ = new_n15036_ & new_n35034_;
  assign new_n35036_ = ~new_n15033_ & ~new_n35035_;
  assign new_n35037_ = ~new_n15018_ & new_n35036_;
  assign new_n35038_ = new_n15018_ & ~new_n15033_;
  assign ys__n28409 = new_n35037_ | new_n35038_;
  assign new_n35040_ = ys__n935 & ~ys__n478;
  assign new_n35041_ = ~ys__n232 & ~ys__n935;
  assign new_n35042_ = ~ys__n478 & new_n35041_;
  assign new_n35043_ = ~new_n35040_ & ~new_n35042_;
  assign new_n35044_ = ys__n38427 & ~new_n35043_;
  assign new_n35045_ = ys__n232 & ~ys__n935;
  assign new_n35046_ = ~ys__n478 & new_n35045_;
  assign new_n35047_ = ys__n47755 & new_n35046_;
  assign new_n35048_ = ~new_n35044_ & ~new_n35047_;
  assign new_n35049_ = ~ys__n478 & ~new_n35046_;
  assign new_n35050_ = new_n35043_ & new_n35049_;
  assign new_n35051_ = ~new_n13769_ & ~new_n35050_;
  assign new_n35052_ = ~new_n35048_ & new_n35051_;
  assign new_n35053_ = ys__n28462 & new_n13769_;
  assign ys__n28410 = new_n35052_ | new_n35053_;
  assign new_n35055_ = ~ys__n4454 & ys__n4455;
  assign new_n35056_ = ys__n22885 & new_n35055_;
  assign new_n35057_ = ys__n4454 & ys__n22822;
  assign new_n35058_ = ~new_n35056_ & ~new_n35057_;
  assign new_n35059_ = ~ys__n4452 & ~new_n35058_;
  assign new_n35060_ = ys__n4452 & ys__n22779;
  assign new_n35061_ = ~new_n35059_ & ~new_n35060_;
  assign new_n35062_ = ~ys__n4457 & ~new_n35061_;
  assign new_n35063_ = ys__n4457 & ys__n22715;
  assign new_n35064_ = ~new_n35062_ & ~new_n35063_;
  assign new_n35065_ = ~ys__n4451 & ~new_n35064_;
  assign new_n35066_ = ys__n4451 & ys__n22675;
  assign new_n35067_ = ~new_n35065_ & ~new_n35066_;
  assign new_n35068_ = ~ys__n4449 & ~ys__n4458;
  assign new_n35069_ = ~new_n35067_ & new_n35068_;
  assign new_n35070_ = ys__n4458 & ys__n22564;
  assign new_n35071_ = ~new_n35069_ & ~new_n35070_;
  assign new_n35072_ = ~ys__n4460 & ~ys__n4461;
  assign new_n35073_ = ~new_n35071_ & new_n35072_;
  assign new_n35074_ = ~ys__n4460 & ~new_n35073_;
  assign new_n35075_ = ~ys__n4448 & ~new_n35074_;
  assign new_n35076_ = ys__n4448 & ys__n28410;
  assign ys__n28411 = new_n35075_ | new_n35076_;
  assign new_n35078_ = ys__n38315 & ~new_n35043_;
  assign new_n35079_ = ys__n47756 & new_n35046_;
  assign new_n35080_ = ~new_n35078_ & ~new_n35079_;
  assign new_n35081_ = new_n35051_ & ~new_n35080_;
  assign new_n35082_ = ys__n28464 & new_n13769_;
  assign ys__n28412 = new_n35081_ | new_n35082_;
  assign new_n35084_ = ys__n22886 & new_n35055_;
  assign new_n35085_ = ys__n4454 & ys__n22824;
  assign new_n35086_ = ~new_n35084_ & ~new_n35085_;
  assign new_n35087_ = ~ys__n4452 & ~new_n35086_;
  assign new_n35088_ = ys__n4452 & ys__n22781;
  assign new_n35089_ = ~new_n35087_ & ~new_n35088_;
  assign new_n35090_ = ~ys__n4457 & ~new_n35089_;
  assign new_n35091_ = ys__n4457 & ys__n22717;
  assign new_n35092_ = ~new_n35090_ & ~new_n35091_;
  assign new_n35093_ = ~ys__n4451 & ~new_n35092_;
  assign new_n35094_ = ys__n4451 & ys__n22677;
  assign new_n35095_ = ~new_n35093_ & ~new_n35094_;
  assign new_n35096_ = new_n35068_ & ~new_n35095_;
  assign new_n35097_ = ys__n4458 & ys__n22566;
  assign new_n35098_ = ~new_n35096_ & ~new_n35097_;
  assign new_n35099_ = ~ys__n4448 & ~ys__n4460;
  assign new_n35100_ = ~ys__n4461 & new_n35099_;
  assign new_n35101_ = ~new_n35098_ & new_n35100_;
  assign new_n35102_ = ys__n4448 & ys__n28412;
  assign ys__n28413 = new_n35101_ | new_n35102_;
  assign new_n35104_ = ys__n47755 & ~new_n35043_;
  assign new_n35105_ = ys__n47757 & new_n35046_;
  assign new_n35106_ = ys__n38427 & ys__n478;
  assign new_n35107_ = ~new_n35105_ & ~new_n35106_;
  assign new_n35108_ = ~new_n35104_ & new_n35107_;
  assign new_n35109_ = new_n35051_ & ~new_n35108_;
  assign new_n35110_ = ys__n28466 & new_n13769_;
  assign ys__n28414 = new_n35109_ | new_n35110_;
  assign new_n35112_ = ys__n22887 & new_n35055_;
  assign new_n35113_ = ys__n4454 & ys__n22826;
  assign new_n35114_ = ~new_n35112_ & ~new_n35113_;
  assign new_n35115_ = ~ys__n4452 & ~new_n35114_;
  assign new_n35116_ = ys__n4452 & ys__n22783;
  assign new_n35117_ = ~new_n35115_ & ~new_n35116_;
  assign new_n35118_ = ~ys__n4457 & ~new_n35117_;
  assign new_n35119_ = ys__n4457 & ys__n22719;
  assign new_n35120_ = ~new_n35118_ & ~new_n35119_;
  assign new_n35121_ = ~ys__n4451 & ~new_n35120_;
  assign new_n35122_ = ys__n4451 & ys__n22679;
  assign new_n35123_ = ~new_n35121_ & ~new_n35122_;
  assign new_n35124_ = ~ys__n4449 & ~new_n35123_;
  assign new_n35125_ = ys__n4449 & ys__n22630;
  assign new_n35126_ = ~new_n35124_ & ~new_n35125_;
  assign new_n35127_ = ~ys__n4458 & ~new_n35126_;
  assign new_n35128_ = ys__n4458 & ys__n22568;
  assign new_n35129_ = ~new_n35127_ & ~new_n35128_;
  assign new_n35130_ = new_n35100_ & ~new_n35129_;
  assign new_n35131_ = ys__n4448 & ys__n28414;
  assign ys__n28415 = new_n35130_ | new_n35131_;
  assign new_n35133_ = ys__n47756 & ~new_n35043_;
  assign new_n35134_ = ys__n47758 & new_n35046_;
  assign new_n35135_ = ys__n38315 & ys__n478;
  assign new_n35136_ = ~new_n35134_ & ~new_n35135_;
  assign new_n35137_ = ~new_n35133_ & new_n35136_;
  assign new_n35138_ = new_n35051_ & ~new_n35137_;
  assign new_n35139_ = ys__n28468 & new_n13769_;
  assign ys__n28416 = new_n35138_ | new_n35139_;
  assign new_n35141_ = ys__n22888 & new_n35055_;
  assign new_n35142_ = ys__n4454 & ys__n22828;
  assign new_n35143_ = ~new_n35141_ & ~new_n35142_;
  assign new_n35144_ = ~ys__n4452 & ~new_n35143_;
  assign new_n35145_ = ys__n4452 & ys__n22785;
  assign new_n35146_ = ~new_n35144_ & ~new_n35145_;
  assign new_n35147_ = ~ys__n4457 & ~new_n35146_;
  assign new_n35148_ = ys__n4457 & ys__n22721;
  assign new_n35149_ = ~new_n35147_ & ~new_n35148_;
  assign new_n35150_ = ~ys__n4451 & ~new_n35149_;
  assign new_n35151_ = ys__n4451 & ys__n22681;
  assign new_n35152_ = ~new_n35150_ & ~new_n35151_;
  assign new_n35153_ = ~ys__n4449 & ~new_n35152_;
  assign new_n35154_ = ys__n4449 & ys__n22632;
  assign new_n35155_ = ~new_n35153_ & ~new_n35154_;
  assign new_n35156_ = ~ys__n4458 & ~new_n35155_;
  assign new_n35157_ = ys__n4458 & ys__n22570;
  assign new_n35158_ = ~new_n35156_ & ~new_n35157_;
  assign new_n35159_ = ~ys__n4461 & ~new_n35158_;
  assign new_n35160_ = ~ys__n4461 & ~new_n35159_;
  assign new_n35161_ = new_n35099_ & ~new_n35160_;
  assign new_n35162_ = ys__n4448 & ys__n28416;
  assign ys__n28417 = new_n35161_ | new_n35162_;
  assign new_n35164_ = ys__n47757 & ~new_n35043_;
  assign new_n35165_ = ys__n47755 & ys__n478;
  assign new_n35166_ = ~new_n35105_ & ~new_n35165_;
  assign new_n35167_ = ~new_n35164_ & new_n35166_;
  assign new_n35168_ = new_n35051_ & ~new_n35167_;
  assign new_n35169_ = ys__n28470 & new_n13769_;
  assign ys__n28418 = new_n35168_ | new_n35169_;
  assign new_n35171_ = ys__n22889 & new_n35055_;
  assign new_n35172_ = ys__n4454 & ys__n22830;
  assign new_n35173_ = ~new_n35171_ & ~new_n35172_;
  assign new_n35174_ = ~ys__n4452 & ~new_n35173_;
  assign new_n35175_ = ys__n4452 & ys__n22787;
  assign new_n35176_ = ~new_n35174_ & ~new_n35175_;
  assign new_n35177_ = ~ys__n4457 & ~new_n35176_;
  assign new_n35178_ = ys__n4457 & ys__n22723;
  assign new_n35179_ = ~new_n35177_ & ~new_n35178_;
  assign new_n35180_ = ~ys__n4451 & ~new_n35179_;
  assign new_n35181_ = ys__n4451 & ys__n22683;
  assign new_n35182_ = ~new_n35180_ & ~new_n35181_;
  assign new_n35183_ = ~ys__n4449 & ~new_n35182_;
  assign new_n35184_ = ys__n4449 & ys__n22634;
  assign new_n35185_ = ~new_n35183_ & ~new_n35184_;
  assign new_n35186_ = ~ys__n4458 & ~new_n35185_;
  assign new_n35187_ = ys__n4458 & ys__n22572;
  assign new_n35188_ = ~new_n35186_ & ~new_n35187_;
  assign new_n35189_ = new_n35100_ & ~new_n35188_;
  assign new_n35190_ = ys__n4448 & ys__n28418;
  assign ys__n28419 = new_n35189_ | new_n35190_;
  assign new_n35192_ = ys__n47758 & ~new_n35043_;
  assign new_n35193_ = ys__n47756 & ys__n478;
  assign new_n35194_ = ~new_n35134_ & ~new_n35193_;
  assign new_n35195_ = ~new_n35192_ & new_n35194_;
  assign new_n35196_ = new_n35051_ & ~new_n35195_;
  assign new_n35197_ = ys__n28472 & new_n13769_;
  assign ys__n28420 = new_n35196_ | new_n35197_;
  assign new_n35199_ = ys__n22890 & new_n35055_;
  assign new_n35200_ = ys__n4454 & ys__n22832;
  assign new_n35201_ = ~new_n35199_ & ~new_n35200_;
  assign new_n35202_ = ~ys__n4452 & ~new_n35201_;
  assign new_n35203_ = ys__n4452 & ys__n22789;
  assign new_n35204_ = ~new_n35202_ & ~new_n35203_;
  assign new_n35205_ = ~ys__n4457 & ~new_n35204_;
  assign new_n35206_ = ys__n4457 & ys__n22725;
  assign new_n35207_ = ~new_n35205_ & ~new_n35206_;
  assign new_n35208_ = ~ys__n4451 & ~new_n35207_;
  assign new_n35209_ = ys__n4451 & ys__n22685;
  assign new_n35210_ = ~new_n35208_ & ~new_n35209_;
  assign new_n35211_ = ~ys__n4449 & ~new_n35210_;
  assign new_n35212_ = ys__n4449 & ys__n22636;
  assign new_n35213_ = ~new_n35211_ & ~new_n35212_;
  assign new_n35214_ = ~ys__n4458 & ~new_n35213_;
  assign new_n35215_ = ys__n4458 & ys__n22574;
  assign new_n35216_ = ~new_n35214_ & ~new_n35215_;
  assign new_n35217_ = new_n35100_ & ~new_n35216_;
  assign new_n35218_ = ys__n4448 & ys__n28420;
  assign ys__n28421 = new_n35217_ | new_n35218_;
  assign new_n35220_ = ys__n22891 & new_n35055_;
  assign new_n35221_ = ys__n4454 & ys__n22834;
  assign new_n35222_ = ~new_n35220_ & ~new_n35221_;
  assign new_n35223_ = ~ys__n4452 & ~ys__n4457;
  assign new_n35224_ = ~new_n35222_ & new_n35223_;
  assign new_n35225_ = ys__n4457 & ys__n22727;
  assign new_n35226_ = ~new_n35224_ & ~new_n35225_;
  assign new_n35227_ = ~ys__n4451 & ~new_n35226_;
  assign new_n35228_ = ys__n4451 & ys__n22687;
  assign new_n35229_ = ~new_n35227_ & ~new_n35228_;
  assign new_n35230_ = new_n35068_ & ~new_n35229_;
  assign new_n35231_ = ys__n4458 & ys__n22576;
  assign new_n35232_ = ~new_n35230_ & ~new_n35231_;
  assign ys__n28422 = new_n35100_ & ~new_n35232_;
  assign new_n35234_ = ys__n22892 & new_n35055_;
  assign new_n35235_ = ys__n4454 & ys__n22836;
  assign new_n35236_ = ~new_n35234_ & ~new_n35235_;
  assign new_n35237_ = ~ys__n4452 & ~new_n35236_;
  assign new_n35238_ = ys__n4452 & ys__n22792;
  assign new_n35239_ = ~new_n35237_ & ~new_n35238_;
  assign new_n35240_ = ~ys__n4457 & ~new_n35239_;
  assign new_n35241_ = ys__n4457 & ys__n22729;
  assign new_n35242_ = ~new_n35240_ & ~new_n35241_;
  assign new_n35243_ = ~ys__n4451 & ~new_n35242_;
  assign new_n35244_ = ys__n4451 & ys__n22689;
  assign new_n35245_ = ~new_n35243_ & ~new_n35244_;
  assign new_n35246_ = new_n35068_ & ~new_n35245_;
  assign new_n35247_ = ys__n4458 & ys__n22578;
  assign new_n35248_ = ~new_n35246_ & ~new_n35247_;
  assign new_n35249_ = ~ys__n4461 & ~new_n35248_;
  assign new_n35250_ = ~ys__n4461 & ~new_n35249_;
  assign ys__n28423 = new_n35099_ & ~new_n35250_;
  assign new_n35252_ = ys__n22893 & new_n35055_;
  assign new_n35253_ = ys__n4454 & ys__n22838;
  assign new_n35254_ = ~new_n35252_ & ~new_n35253_;
  assign new_n35255_ = ~ys__n4452 & ~new_n35254_;
  assign new_n35256_ = ys__n4452 & ys__n22794;
  assign new_n35257_ = ~new_n35255_ & ~new_n35256_;
  assign new_n35258_ = ~ys__n4457 & ~new_n35257_;
  assign new_n35259_ = ys__n4457 & ys__n22731;
  assign new_n35260_ = ~new_n35258_ & ~new_n35259_;
  assign new_n35261_ = ~ys__n4449 & ~ys__n4451;
  assign new_n35262_ = ~new_n35260_ & new_n35261_;
  assign new_n35263_ = ys__n4449 & ys__n22640;
  assign new_n35264_ = ~new_n35262_ & ~new_n35263_;
  assign new_n35265_ = ~ys__n4458 & ~new_n35264_;
  assign new_n35266_ = ys__n4458 & ys__n22580;
  assign new_n35267_ = ~new_n35265_ & ~new_n35266_;
  assign new_n35268_ = ~ys__n4461 & ~new_n35267_;
  assign new_n35269_ = ~ys__n4461 & ~new_n35268_;
  assign new_n35270_ = ~ys__n4460 & ~new_n35269_;
  assign new_n35271_ = ~ys__n4460 & ~new_n35270_;
  assign new_n35272_ = ~ys__n4448 & ~new_n35271_;
  assign new_n35273_ = ys__n4448 & ys__n28424;
  assign ys__n28425 = new_n35272_ | new_n35273_;
  assign new_n35275_ = ys__n22894 & new_n35055_;
  assign new_n35276_ = ys__n4454 & ys__n22840;
  assign new_n35277_ = ~new_n35275_ & ~new_n35276_;
  assign new_n35278_ = new_n35223_ & ~new_n35277_;
  assign new_n35279_ = ys__n4457 & ys__n22733;
  assign new_n35280_ = ~new_n35278_ & ~new_n35279_;
  assign new_n35281_ = new_n35261_ & ~new_n35280_;
  assign new_n35282_ = ys__n4449 & ys__n22642;
  assign new_n35283_ = ~new_n35281_ & ~new_n35282_;
  assign new_n35284_ = ~ys__n4458 & ~new_n35283_;
  assign new_n35285_ = ys__n4458 & ys__n22582;
  assign new_n35286_ = ~new_n35284_ & ~new_n35285_;
  assign new_n35287_ = new_n35100_ & ~new_n35286_;
  assign new_n35288_ = ys__n4448 & ys__n28426;
  assign ys__n28427 = new_n35287_ | new_n35288_;
  assign new_n35290_ = ys__n22895 & new_n35055_;
  assign new_n35291_ = ys__n4454 & ys__n22842;
  assign new_n35292_ = ~new_n35290_ & ~new_n35291_;
  assign new_n35293_ = new_n35223_ & ~new_n35292_;
  assign new_n35294_ = ys__n4457 & ys__n22735;
  assign new_n35295_ = ~new_n35293_ & ~new_n35294_;
  assign new_n35296_ = new_n35261_ & ~new_n35295_;
  assign new_n35297_ = ys__n4449 & ys__n22644;
  assign new_n35298_ = ~new_n35296_ & ~new_n35297_;
  assign new_n35299_ = ~ys__n4458 & ~new_n35298_;
  assign new_n35300_ = ys__n4458 & ys__n22584;
  assign new_n35301_ = ~new_n35299_ & ~new_n35300_;
  assign new_n35302_ = new_n35100_ & ~new_n35301_;
  assign new_n35303_ = ys__n4448 & ys__n28428;
  assign ys__n28429 = new_n35302_ | new_n35303_;
  assign new_n35305_ = ys__n22896 & new_n35055_;
  assign new_n35306_ = ys__n4454 & ys__n22844;
  assign new_n35307_ = ~new_n35305_ & ~new_n35306_;
  assign new_n35308_ = new_n35223_ & ~new_n35307_;
  assign new_n35309_ = ys__n4457 & ys__n22737;
  assign new_n35310_ = ~new_n35308_ & ~new_n35309_;
  assign new_n35311_ = new_n35261_ & ~new_n35310_;
  assign new_n35312_ = ys__n4449 & ys__n22646;
  assign new_n35313_ = ~new_n35311_ & ~new_n35312_;
  assign new_n35314_ = ~ys__n4458 & ~new_n35313_;
  assign new_n35315_ = ys__n4458 & ys__n22586;
  assign new_n35316_ = ~new_n35314_ & ~new_n35315_;
  assign new_n35317_ = new_n35100_ & ~new_n35316_;
  assign new_n35318_ = ys__n4448 & ys__n28430;
  assign ys__n28431 = new_n35317_ | new_n35318_;
  assign new_n35320_ = ys__n22897 & new_n35055_;
  assign new_n35321_ = ys__n4454 & ys__n22846;
  assign new_n35322_ = ~new_n35320_ & ~new_n35321_;
  assign new_n35323_ = ~ys__n4452 & ~new_n35322_;
  assign new_n35324_ = ys__n4452 & ys__n22799;
  assign new_n35325_ = ~new_n35323_ & ~new_n35324_;
  assign new_n35326_ = ~ys__n4457 & ~new_n35325_;
  assign new_n35327_ = ys__n4457 & ys__n22739;
  assign new_n35328_ = ~new_n35326_ & ~new_n35327_;
  assign new_n35329_ = new_n35261_ & ~new_n35328_;
  assign new_n35330_ = ys__n4449 & ys__n22648;
  assign new_n35331_ = ~new_n35329_ & ~new_n35330_;
  assign new_n35332_ = ~ys__n4458 & ~new_n35331_;
  assign new_n35333_ = ys__n4458 & ys__n22588;
  assign new_n35334_ = ~new_n35332_ & ~new_n35333_;
  assign new_n35335_ = new_n35100_ & ~new_n35334_;
  assign new_n35336_ = ys__n4448 & ys__n28432;
  assign ys__n28433 = new_n35335_ | new_n35336_;
  assign new_n35338_ = ys__n22898 & new_n35055_;
  assign new_n35339_ = ys__n4454 & ys__n22848;
  assign new_n35340_ = ~new_n35338_ & ~new_n35339_;
  assign new_n35341_ = new_n35223_ & ~new_n35340_;
  assign new_n35342_ = ys__n4457 & ys__n22741;
  assign new_n35343_ = ~new_n35341_ & ~new_n35342_;
  assign new_n35344_ = new_n35261_ & ~new_n35343_;
  assign new_n35345_ = ys__n4449 & ys__n22650;
  assign new_n35346_ = ~new_n35344_ & ~new_n35345_;
  assign new_n35347_ = ~ys__n4458 & ~new_n35346_;
  assign new_n35348_ = ys__n4458 & ys__n22590;
  assign new_n35349_ = ~new_n35347_ & ~new_n35348_;
  assign new_n35350_ = new_n35100_ & ~new_n35349_;
  assign new_n35351_ = ys__n4448 & ys__n28434;
  assign ys__n28435 = new_n35350_ | new_n35351_;
  assign new_n35353_ = ys__n22899 & new_n35055_;
  assign new_n35354_ = ys__n4454 & ys__n22850;
  assign new_n35355_ = ~new_n35353_ & ~new_n35354_;
  assign new_n35356_ = new_n35223_ & ~new_n35355_;
  assign new_n35357_ = ys__n4457 & ys__n22743;
  assign new_n35358_ = ~new_n35356_ & ~new_n35357_;
  assign new_n35359_ = new_n35261_ & ~new_n35358_;
  assign new_n35360_ = ys__n4449 & ys__n22652;
  assign new_n35361_ = ~new_n35359_ & ~new_n35360_;
  assign new_n35362_ = ~ys__n4458 & ~new_n35361_;
  assign new_n35363_ = ys__n4458 & ys__n22592;
  assign new_n35364_ = ~new_n35362_ & ~new_n35363_;
  assign new_n35365_ = new_n35072_ & ~new_n35364_;
  assign new_n35366_ = ~ys__n4460 & ~new_n35365_;
  assign new_n35367_ = ~ys__n4448 & ~new_n35366_;
  assign new_n35368_ = ys__n4448 & ys__n28436;
  assign ys__n28437 = new_n35367_ | new_n35368_;
  assign new_n35370_ = ys__n22900 & new_n35055_;
  assign new_n35371_ = ys__n4454 & ys__n22852;
  assign new_n35372_ = ~new_n35370_ & ~new_n35371_;
  assign new_n35373_ = new_n35223_ & ~new_n35372_;
  assign new_n35374_ = ys__n4457 & ys__n22745;
  assign new_n35375_ = ~new_n35373_ & ~new_n35374_;
  assign new_n35376_ = new_n35261_ & ~new_n35375_;
  assign new_n35377_ = ys__n4449 & ys__n22654;
  assign new_n35378_ = ~new_n35376_ & ~new_n35377_;
  assign new_n35379_ = ~ys__n4458 & ~new_n35378_;
  assign new_n35380_ = ys__n4458 & ys__n22594;
  assign new_n35381_ = ~new_n35379_ & ~new_n35380_;
  assign new_n35382_ = new_n35072_ & ~new_n35381_;
  assign new_n35383_ = ~ys__n4460 & ~new_n35382_;
  assign new_n35384_ = ~ys__n4448 & ~new_n35383_;
  assign new_n35385_ = ys__n4448 & ys__n28438;
  assign ys__n28439 = new_n35384_ | new_n35385_;
  assign new_n35387_ = ys__n22901 & new_n35055_;
  assign new_n35388_ = ys__n4454 & ys__n22854;
  assign new_n35389_ = ~new_n35387_ & ~new_n35388_;
  assign new_n35390_ = new_n35223_ & ~new_n35389_;
  assign new_n35391_ = ys__n4457 & ys__n22747;
  assign new_n35392_ = ~new_n35390_ & ~new_n35391_;
  assign new_n35393_ = ~ys__n4458 & new_n35261_;
  assign new_n35394_ = ~new_n35392_ & new_n35393_;
  assign new_n35395_ = ys__n4458 & ys__n22596;
  assign new_n35396_ = ~new_n35394_ & ~new_n35395_;
  assign new_n35397_ = ~ys__n4461 & ~new_n35396_;
  assign new_n35398_ = ~ys__n4461 & ~new_n35397_;
  assign ys__n28440 = new_n35099_ & ~new_n35398_;
  assign new_n35400_ = ys__n22902 & new_n35055_;
  assign new_n35401_ = ys__n4454 & ys__n22856;
  assign new_n35402_ = ~new_n35400_ & ~new_n35401_;
  assign new_n35403_ = new_n35223_ & ~new_n35402_;
  assign new_n35404_ = ys__n4457 & ys__n22749;
  assign new_n35405_ = ~new_n35403_ & ~new_n35404_;
  assign new_n35406_ = new_n35393_ & ~new_n35405_;
  assign new_n35407_ = ys__n4458 & ys__n22598;
  assign new_n35408_ = ~new_n35406_ & ~new_n35407_;
  assign ys__n28441 = new_n35100_ & ~new_n35408_;
  assign new_n35410_ = ys__n22903 & new_n35055_;
  assign new_n35411_ = ys__n4454 & ys__n22858;
  assign new_n35412_ = ~new_n35410_ & ~new_n35411_;
  assign new_n35413_ = new_n35223_ & ~new_n35412_;
  assign new_n35414_ = ys__n4457 & ys__n22751;
  assign new_n35415_ = ~new_n35413_ & ~new_n35414_;
  assign new_n35416_ = new_n35393_ & ~new_n35415_;
  assign new_n35417_ = ys__n4458 & ys__n22600;
  assign new_n35418_ = ~new_n35416_ & ~new_n35417_;
  assign new_n35419_ = ~ys__n4461 & ~new_n35418_;
  assign new_n35420_ = ~ys__n4461 & ~new_n35419_;
  assign ys__n28442 = new_n35099_ & ~new_n35420_;
  assign new_n35422_ = ys__n22904 & new_n35055_;
  assign new_n35423_ = ys__n4454 & ys__n22860;
  assign new_n35424_ = ~new_n35422_ & ~new_n35423_;
  assign new_n35425_ = new_n35223_ & ~new_n35424_;
  assign new_n35426_ = ys__n4457 & ys__n22753;
  assign new_n35427_ = ~new_n35425_ & ~new_n35426_;
  assign new_n35428_ = new_n35393_ & ~new_n35427_;
  assign new_n35429_ = ys__n4458 & ys__n22602;
  assign new_n35430_ = ~new_n35428_ & ~new_n35429_;
  assign new_n35431_ = ~ys__n4461 & ~new_n35430_;
  assign new_n35432_ = ~ys__n4461 & ~new_n35431_;
  assign ys__n28443 = new_n35099_ & ~new_n35432_;
  assign new_n35434_ = ys__n22905 & new_n35055_;
  assign new_n35435_ = ys__n4454 & ys__n22862;
  assign new_n35436_ = ~new_n35434_ & ~new_n35435_;
  assign new_n35437_ = new_n35223_ & ~new_n35436_;
  assign new_n35438_ = ys__n4457 & ys__n22755;
  assign new_n35439_ = ~new_n35437_ & ~new_n35438_;
  assign new_n35440_ = new_n35393_ & ~new_n35439_;
  assign new_n35441_ = ys__n4458 & ys__n22604;
  assign new_n35442_ = ~new_n35440_ & ~new_n35441_;
  assign ys__n28444 = new_n35100_ & ~new_n35442_;
  assign new_n35444_ = ys__n22906 & new_n35055_;
  assign new_n35445_ = ys__n4454 & ys__n22864;
  assign new_n35446_ = ~new_n35444_ & ~new_n35445_;
  assign new_n35447_ = new_n35223_ & ~new_n35446_;
  assign new_n35448_ = ys__n4457 & ys__n22757;
  assign new_n35449_ = ~new_n35447_ & ~new_n35448_;
  assign new_n35450_ = new_n35393_ & ~new_n35449_;
  assign new_n35451_ = ys__n4458 & ys__n22606;
  assign new_n35452_ = ~new_n35450_ & ~new_n35451_;
  assign ys__n28445 = new_n35100_ & ~new_n35452_;
  assign new_n35454_ = ys__n22907 & new_n35055_;
  assign new_n35455_ = ys__n4454 & ys__n22866;
  assign new_n35456_ = ~new_n35454_ & ~new_n35455_;
  assign new_n35457_ = new_n35223_ & ~new_n35456_;
  assign new_n35458_ = ys__n4457 & ys__n22759;
  assign new_n35459_ = ~new_n35457_ & ~new_n35458_;
  assign new_n35460_ = new_n35393_ & ~new_n35459_;
  assign new_n35461_ = ys__n4458 & ys__n22608;
  assign new_n35462_ = ~new_n35460_ & ~new_n35461_;
  assign new_n35463_ = ~ys__n4461 & ~new_n35462_;
  assign new_n35464_ = ~ys__n4461 & ~new_n35463_;
  assign new_n35465_ = new_n35099_ & ~new_n35464_;
  assign new_n35466_ = ys__n4448 & ys__n28446;
  assign ys__n28447 = new_n35465_ | new_n35466_;
  assign new_n35468_ = ys__n22908 & new_n35055_;
  assign new_n35469_ = ys__n4454 & ys__n22868;
  assign new_n35470_ = ~new_n35468_ & ~new_n35469_;
  assign new_n35471_ = new_n35223_ & ~new_n35470_;
  assign new_n35472_ = ys__n4457 & ys__n22761;
  assign new_n35473_ = ~new_n35471_ & ~new_n35472_;
  assign new_n35474_ = new_n35393_ & ~new_n35473_;
  assign new_n35475_ = ys__n4458 & ys__n22610;
  assign new_n35476_ = ~new_n35474_ & ~new_n35475_;
  assign ys__n28448 = new_n35100_ & ~new_n35476_;
  assign new_n35478_ = ys__n22909 & new_n35055_;
  assign new_n35479_ = ys__n4454 & ys__n22870;
  assign new_n35480_ = ~new_n35478_ & ~new_n35479_;
  assign new_n35481_ = new_n35223_ & ~new_n35480_;
  assign new_n35482_ = ys__n4457 & ys__n22763;
  assign new_n35483_ = ~new_n35481_ & ~new_n35482_;
  assign new_n35484_ = new_n35393_ & ~new_n35483_;
  assign new_n35485_ = ys__n4458 & ys__n22612;
  assign new_n35486_ = ~new_n35484_ & ~new_n35485_;
  assign ys__n28449 = new_n35100_ & ~new_n35486_;
  assign new_n35488_ = ys__n22910 & new_n35055_;
  assign new_n35489_ = ys__n4454 & ys__n22872;
  assign new_n35490_ = ~new_n35488_ & ~new_n35489_;
  assign new_n35491_ = new_n35223_ & ~new_n35490_;
  assign new_n35492_ = ys__n4457 & ys__n22765;
  assign new_n35493_ = ~new_n35491_ & ~new_n35492_;
  assign new_n35494_ = new_n35393_ & ~new_n35493_;
  assign new_n35495_ = ys__n4458 & ys__n22614;
  assign new_n35496_ = ~new_n35494_ & ~new_n35495_;
  assign ys__n28450 = new_n35100_ & ~new_n35496_;
  assign new_n35498_ = ys__n22911 & new_n35055_;
  assign new_n35499_ = ys__n4454 & ys__n22874;
  assign new_n35500_ = ~new_n35498_ & ~new_n35499_;
  assign new_n35501_ = new_n35223_ & ~new_n35500_;
  assign new_n35502_ = ys__n4457 & ys__n22767;
  assign new_n35503_ = ~new_n35501_ & ~new_n35502_;
  assign new_n35504_ = new_n35393_ & ~new_n35503_;
  assign new_n35505_ = ys__n4458 & ys__n22616;
  assign new_n35506_ = ~new_n35504_ & ~new_n35505_;
  assign ys__n28451 = new_n35100_ & ~new_n35506_;
  assign new_n35508_ = ys__n22912 & new_n35055_;
  assign new_n35509_ = ys__n4454 & ys__n22876;
  assign new_n35510_ = ~new_n35508_ & ~new_n35509_;
  assign new_n35511_ = new_n35223_ & ~new_n35510_;
  assign new_n35512_ = ys__n4457 & ys__n22769;
  assign new_n35513_ = ~new_n35511_ & ~new_n35512_;
  assign new_n35514_ = new_n35393_ & ~new_n35513_;
  assign new_n35515_ = ys__n4458 & ys__n22618;
  assign new_n35516_ = ~new_n35514_ & ~new_n35515_;
  assign ys__n28452 = new_n35100_ & ~new_n35516_;
  assign new_n35518_ = ys__n22913 & new_n35055_;
  assign new_n35519_ = ys__n4454 & ys__n22878;
  assign new_n35520_ = ~new_n35518_ & ~new_n35519_;
  assign new_n35521_ = new_n35223_ & ~new_n35520_;
  assign new_n35522_ = ys__n4457 & ys__n22771;
  assign new_n35523_ = ~new_n35521_ & ~new_n35522_;
  assign new_n35524_ = new_n35261_ & ~new_n35523_;
  assign new_n35525_ = ys__n4449 & ys__n22668;
  assign new_n35526_ = ~new_n35524_ & ~new_n35525_;
  assign new_n35527_ = ~ys__n4458 & ~new_n35526_;
  assign new_n35528_ = ys__n4458 & ys__n22620;
  assign new_n35529_ = ~new_n35527_ & ~new_n35528_;
  assign new_n35530_ = new_n35100_ & ~new_n35529_;
  assign new_n35531_ = ys__n4448 & ys__n28453;
  assign ys__n28454 = new_n35530_ | new_n35531_;
  assign new_n35533_ = ys__n22914 & new_n35055_;
  assign new_n35534_ = ys__n4454 & ys__n22880;
  assign new_n35535_ = ~new_n35533_ & ~new_n35534_;
  assign new_n35536_ = new_n35223_ & ~new_n35535_;
  assign new_n35537_ = ys__n4457 & ys__n22773;
  assign new_n35538_ = ~new_n35536_ & ~new_n35537_;
  assign new_n35539_ = new_n35261_ & ~new_n35538_;
  assign new_n35540_ = ys__n4449 & ys__n22670;
  assign new_n35541_ = ~new_n35539_ & ~new_n35540_;
  assign new_n35542_ = ~ys__n4458 & ~new_n35541_;
  assign new_n35543_ = ys__n4458 & ys__n22622;
  assign new_n35544_ = ~new_n35542_ & ~new_n35543_;
  assign new_n35545_ = ~ys__n4461 & ~new_n35544_;
  assign new_n35546_ = ~ys__n4461 & ~new_n35545_;
  assign new_n35547_ = new_n35099_ & ~new_n35546_;
  assign new_n35548_ = ys__n4448 & ys__n28455;
  assign ys__n28456 = new_n35547_ | new_n35548_;
  assign new_n35550_ = ys__n22915 & new_n35055_;
  assign new_n35551_ = ys__n4454 & ys__n22882;
  assign new_n35552_ = ~new_n35550_ & ~new_n35551_;
  assign new_n35553_ = ~ys__n4452 & ~new_n35552_;
  assign new_n35554_ = ys__n4452 & ys__n22818;
  assign new_n35555_ = ~new_n35553_ & ~new_n35554_;
  assign new_n35556_ = ~ys__n4457 & ~new_n35555_;
  assign new_n35557_ = ys__n4457 & ys__n22775;
  assign new_n35558_ = ~new_n35556_ & ~new_n35557_;
  assign new_n35559_ = new_n35393_ & ~new_n35558_;
  assign new_n35560_ = ys__n4458 & ys__n22624;
  assign new_n35561_ = ~new_n35559_ & ~new_n35560_;
  assign new_n35562_ = new_n35100_ & ~new_n35561_;
  assign new_n35563_ = ys__n4448 & ys__n28457;
  assign ys__n28458 = new_n35562_ | new_n35563_;
  assign new_n35565_ = ys__n22916 & new_n35055_;
  assign new_n35566_ = ys__n4454 & ys__n22884;
  assign new_n35567_ = ~new_n35565_ & ~new_n35566_;
  assign new_n35568_ = ~ys__n4452 & ~new_n35567_;
  assign new_n35569_ = ys__n4452 & ys__n22820;
  assign new_n35570_ = ~new_n35568_ & ~new_n35569_;
  assign new_n35571_ = ~ys__n4457 & ~new_n35570_;
  assign new_n35572_ = ys__n4457 & ys__n22777;
  assign new_n35573_ = ~new_n35571_ & ~new_n35572_;
  assign new_n35574_ = new_n35261_ & ~new_n35573_;
  assign new_n35575_ = ys__n4449 & ys__n22673;
  assign new_n35576_ = ~new_n35574_ & ~new_n35575_;
  assign new_n35577_ = ~ys__n4458 & ~new_n35576_;
  assign new_n35578_ = ys__n4458 & ys__n22626;
  assign new_n35579_ = ~new_n35577_ & ~new_n35578_;
  assign new_n35580_ = new_n35100_ & ~new_n35579_;
  assign new_n35581_ = ys__n4448 & ys__n28459;
  assign ys__n28460 = new_n35580_ | new_n35581_;
  assign new_n35583_ = ~ys__n24256 & ~ys__n24260;
  assign new_n35584_ = ~ys__n28412 & ~new_n35583_;
  assign new_n35585_ = ys__n20053 & new_n35584_;
  assign new_n35586_ = ~ys__n33375 & ys__n18218;
  assign new_n35587_ = ~ys__n20053 & ~new_n35586_;
  assign new_n35588_ = ys__n28412 & ~new_n35583_;
  assign new_n35589_ = ~new_n35587_ & new_n35588_;
  assign ys__n28475 = new_n35585_ | new_n35589_;
  assign new_n35591_ = ~ys__n28243 & ys__n23483;
  assign new_n35592_ = ys__n22464 & ys__n28243;
  assign ys__n28476 = new_n35591_ | new_n35592_;
  assign new_n35594_ = ~ys__n28243 & ys__n23485;
  assign new_n35595_ = ys__n23548 & ys__n28243;
  assign ys__n28477 = new_n35594_ | new_n35595_;
  assign new_n35597_ = ~ys__n28243 & ys__n23487;
  assign new_n35598_ = ys__n23550 & ys__n28243;
  assign ys__n28478 = new_n35597_ | new_n35598_;
  assign new_n35600_ = ~ys__n28243 & ys__n23489;
  assign new_n35601_ = ys__n23552 & ys__n28243;
  assign ys__n28479 = new_n35600_ | new_n35601_;
  assign new_n35603_ = ~ys__n28243 & ys__n23491;
  assign new_n35604_ = ys__n23554 & ys__n28243;
  assign ys__n28480 = new_n35603_ | new_n35604_;
  assign new_n35606_ = ~ys__n28243 & ys__n23493;
  assign new_n35607_ = ys__n23556 & ys__n28243;
  assign ys__n28481 = new_n35606_ | new_n35607_;
  assign new_n35609_ = ~ys__n28243 & ys__n23495;
  assign new_n35610_ = ys__n23558 & ys__n28243;
  assign ys__n28482 = new_n35609_ | new_n35610_;
  assign new_n35612_ = ~ys__n28243 & ys__n23497;
  assign new_n35613_ = ys__n23560 & ys__n28243;
  assign ys__n28483 = new_n35612_ | new_n35613_;
  assign new_n35615_ = ~ys__n28243 & ys__n23499;
  assign new_n35616_ = ys__n23562 & ys__n28243;
  assign ys__n28484 = new_n35615_ | new_n35616_;
  assign new_n35618_ = ~ys__n28243 & ys__n23501;
  assign new_n35619_ = ys__n23564 & ys__n28243;
  assign ys__n28485 = new_n35618_ | new_n35619_;
  assign new_n35621_ = ~ys__n28243 & ys__n23503;
  assign new_n35622_ = ys__n23566 & ys__n28243;
  assign ys__n28486 = new_n35621_ | new_n35622_;
  assign new_n35624_ = ~ys__n28243 & ys__n23505;
  assign new_n35625_ = ys__n23568 & ys__n28243;
  assign ys__n28487 = new_n35624_ | new_n35625_;
  assign new_n35627_ = ~ys__n28243 & ys__n23507;
  assign new_n35628_ = ys__n23570 & ys__n28243;
  assign ys__n28488 = new_n35627_ | new_n35628_;
  assign new_n35630_ = ~ys__n28243 & ys__n23509;
  assign new_n35631_ = ys__n23572 & ys__n28243;
  assign ys__n28489 = new_n35630_ | new_n35631_;
  assign new_n35633_ = ~ys__n28243 & ys__n23511;
  assign new_n35634_ = ys__n23574 & ys__n28243;
  assign ys__n28490 = new_n35633_ | new_n35634_;
  assign new_n35636_ = ~ys__n28243 & ys__n23513;
  assign new_n35637_ = ys__n420 & ys__n28243;
  assign ys__n28491 = new_n35636_ | new_n35637_;
  assign new_n35639_ = ~ys__n28243 & ys__n23515;
  assign new_n35640_ = ys__n442 & ys__n28243;
  assign ys__n28492 = new_n35639_ | new_n35640_;
  assign new_n35642_ = ~ys__n28243 & ys__n23517;
  assign new_n35643_ = ys__n440 & ys__n28243;
  assign ys__n28493 = new_n35642_ | new_n35643_;
  assign new_n35645_ = ~ys__n28243 & ys__n23519;
  assign new_n35646_ = ys__n444 & ys__n28243;
  assign ys__n28494 = new_n35645_ | new_n35646_;
  assign new_n35648_ = ~ys__n28243 & ys__n23521;
  assign new_n35649_ = ys__n438 & ys__n28243;
  assign ys__n28495 = new_n35648_ | new_n35649_;
  assign new_n35651_ = ~ys__n28243 & ys__n23523;
  assign new_n35652_ = ys__n446 & ys__n28243;
  assign ys__n28496 = new_n35651_ | new_n35652_;
  assign new_n35654_ = ~ys__n28243 & ys__n23525;
  assign new_n35655_ = ys__n434 & ys__n28243;
  assign ys__n28497 = new_n35654_ | new_n35655_;
  assign new_n35657_ = ~ys__n28243 & ys__n23527;
  assign new_n35658_ = ys__n436 & ys__n28243;
  assign ys__n28498 = new_n35657_ | new_n35658_;
  assign new_n35660_ = ~ys__n28243 & ys__n23529;
  assign new_n35661_ = ys__n432 & ys__n28243;
  assign ys__n28499 = new_n35660_ | new_n35661_;
  assign new_n35663_ = ~ys__n28243 & ys__n23531;
  assign new_n35664_ = ys__n448 & ys__n28243;
  assign ys__n28500 = new_n35663_ | new_n35664_;
  assign new_n35666_ = ~ys__n28243 & ys__n23533;
  assign new_n35667_ = ys__n428 & ys__n28243;
  assign ys__n28501 = new_n35666_ | new_n35667_;
  assign new_n35669_ = ~ys__n28243 & ys__n23535;
  assign new_n35670_ = ys__n430 & ys__n28243;
  assign ys__n28502 = new_n35669_ | new_n35670_;
  assign new_n35672_ = ~ys__n28243 & ys__n23537;
  assign new_n35673_ = ys__n426 & ys__n28243;
  assign ys__n28503 = new_n35672_ | new_n35673_;
  assign new_n35675_ = ~ys__n28243 & ys__n23539;
  assign new_n35676_ = ys__n450 & ys__n28243;
  assign ys__n28504 = new_n35675_ | new_n35676_;
  assign new_n35678_ = ~ys__n28243 & ys__n23541;
  assign new_n35679_ = ys__n424 & ys__n28243;
  assign ys__n28505 = new_n35678_ | new_n35679_;
  assign new_n35681_ = ~ys__n28243 & ys__n23543;
  assign new_n35682_ = ys__n422 & ys__n28243;
  assign ys__n28506 = new_n35681_ | new_n35682_;
  assign new_n35684_ = ys__n47661 & new_n12768_;
  assign new_n35685_ = ys__n22822 & new_n12309_;
  assign new_n35686_ = ~new_n12314_ & new_n35685_;
  assign new_n35687_ = ~new_n12320_ & new_n35686_;
  assign new_n35688_ = ys__n23480 & new_n12320_;
  assign new_n35689_ = ~new_n35687_ & ~new_n35688_;
  assign new_n35690_ = ~new_n12404_ & ~new_n35689_;
  assign new_n35691_ = ys__n23480 & new_n12404_;
  assign new_n35692_ = ~new_n35690_ & ~new_n35691_;
  assign new_n35693_ = new_n12458_ & ~new_n12477_;
  assign new_n35694_ = ~new_n35692_ & new_n35693_;
  assign new_n35695_ = ys__n23480 & new_n12477_;
  assign new_n35696_ = ~new_n35694_ & ~new_n35695_;
  assign new_n35697_ = new_n12763_ & ~new_n35696_;
  assign new_n35698_ = ~new_n35684_ & ~new_n35697_;
  assign new_n35699_ = new_n12774_ & ~new_n35698_;
  assign new_n35700_ = ys__n47661 & new_n12778_;
  assign new_n35701_ = new_n12776_ & ~new_n35696_;
  assign new_n35702_ = ~new_n35700_ & ~new_n35701_;
  assign new_n35703_ = new_n12784_ & ~new_n35702_;
  assign ys__n28510 = new_n35699_ | new_n35703_;
  assign new_n35705_ = ys__n47662 & new_n12768_;
  assign new_n35706_ = ys__n22824 & ~new_n12314_;
  assign new_n35707_ = new_n12309_ & new_n35706_;
  assign new_n35708_ = ~new_n17411_ & ~new_n35707_;
  assign new_n35709_ = ~new_n12320_ & ~new_n35708_;
  assign new_n35710_ = ys__n22464 & new_n12320_;
  assign new_n35711_ = ~new_n35709_ & ~new_n35710_;
  assign new_n35712_ = ~new_n12404_ & ~new_n35711_;
  assign new_n35713_ = new_n12404_ & ys__n23483;
  assign new_n35714_ = ~new_n35712_ & ~new_n35713_;
  assign new_n35715_ = new_n35693_ & ~new_n35714_;
  assign new_n35716_ = ~ys__n22464 & new_n12523_;
  assign new_n35717_ = ys__n22464 & ~new_n12523_;
  assign new_n35718_ = ~new_n35716_ & ~new_n35717_;
  assign new_n35719_ = new_n12477_ & ~new_n35718_;
  assign new_n35720_ = ~new_n35715_ & ~new_n35719_;
  assign new_n35721_ = new_n12763_ & ~new_n35720_;
  assign new_n35722_ = ~new_n35705_ & ~new_n35721_;
  assign new_n35723_ = new_n12774_ & ~new_n35722_;
  assign new_n35724_ = ys__n47662 & new_n12778_;
  assign new_n35725_ = new_n12776_ & ~new_n35720_;
  assign new_n35726_ = ~new_n35724_ & ~new_n35725_;
  assign new_n35727_ = new_n12784_ & ~new_n35726_;
  assign ys__n28513 = new_n35723_ | new_n35727_;
  assign new_n35729_ = ys__n47664 & new_n12768_;
  assign new_n35730_ = ys__n22828 & ~new_n12314_;
  assign new_n35731_ = new_n12309_ & new_n35730_;
  assign new_n35732_ = ~new_n17423_ & ~new_n35731_;
  assign new_n35733_ = ~new_n12320_ & ~new_n35732_;
  assign new_n35734_ = ys__n23550 & new_n12320_;
  assign new_n35735_ = ~new_n35733_ & ~new_n35734_;
  assign new_n35736_ = ~new_n12404_ & ~new_n35735_;
  assign new_n35737_ = new_n12404_ & ys__n23487;
  assign new_n35738_ = ~new_n35736_ & ~new_n35737_;
  assign new_n35739_ = new_n12458_ & ~new_n35738_;
  assign new_n35740_ = ys__n526 & ~new_n12458_;
  assign new_n35741_ = ~new_n35739_ & ~new_n35740_;
  assign new_n35742_ = ~new_n12477_ & ~new_n35741_;
  assign new_n35743_ = ~new_n12506_ & new_n12524_;
  assign new_n35744_ = ~new_n12528_ & ~new_n35743_;
  assign new_n35745_ = new_n12517_ & ~new_n35744_;
  assign new_n35746_ = ~new_n12517_ & new_n35744_;
  assign new_n35747_ = ~new_n35745_ & ~new_n35746_;
  assign new_n35748_ = new_n12477_ & ~new_n35747_;
  assign new_n35749_ = ~new_n35742_ & ~new_n35748_;
  assign new_n35750_ = new_n12763_ & ~new_n35749_;
  assign new_n35751_ = ~new_n35729_ & ~new_n35750_;
  assign new_n35752_ = new_n12774_ & ~new_n35751_;
  assign new_n35753_ = ys__n47664 & new_n12778_;
  assign new_n35754_ = new_n12776_ & ~new_n35749_;
  assign new_n35755_ = ~new_n35753_ & ~new_n35754_;
  assign new_n35756_ = new_n12784_ & ~new_n35755_;
  assign ys__n28518 = new_n35752_ | new_n35756_;
  assign new_n35758_ = ys__n47671 & new_n12768_;
  assign new_n35759_ = ys__n22842 & ~new_n12314_;
  assign new_n35760_ = new_n12309_ & new_n35759_;
  assign new_n35761_ = ~new_n17465_ & ~new_n35760_;
  assign new_n35762_ = ~new_n12320_ & ~new_n35761_;
  assign new_n35763_ = ys__n23564 & new_n12320_;
  assign new_n35764_ = ~new_n35762_ & ~new_n35763_;
  assign new_n35765_ = ~new_n12404_ & ~new_n35764_;
  assign new_n35766_ = new_n12404_ & ys__n23501;
  assign new_n35767_ = ~new_n35765_ & ~new_n35766_;
  assign new_n35768_ = new_n12458_ & ~new_n35767_;
  assign new_n35769_ = ys__n518 & ~new_n12458_;
  assign new_n35770_ = ~new_n35768_ & ~new_n35769_;
  assign new_n35771_ = ~new_n12477_ & ~new_n35770_;
  assign new_n35772_ = ~new_n12590_ & new_n12670_;
  assign new_n35773_ = new_n12677_ & ~new_n35772_;
  assign new_n35774_ = new_n12648_ & ~new_n35773_;
  assign new_n35775_ = ~new_n12648_ & new_n35773_;
  assign new_n35776_ = ~new_n35774_ & ~new_n35775_;
  assign new_n35777_ = new_n12477_ & ~new_n35776_;
  assign new_n35778_ = ~new_n35771_ & ~new_n35777_;
  assign new_n35779_ = new_n12763_ & ~new_n35778_;
  assign new_n35780_ = ~new_n35758_ & ~new_n35779_;
  assign new_n35781_ = new_n12774_ & ~new_n35780_;
  assign new_n35782_ = ys__n47671 & new_n12778_;
  assign new_n35783_ = new_n12776_ & ~new_n35778_;
  assign new_n35784_ = ~new_n35782_ & ~new_n35783_;
  assign new_n35785_ = new_n12784_ & ~new_n35784_;
  assign ys__n28533 = new_n35781_ | new_n35785_;
  assign new_n35787_ = ys__n47672 & new_n12768_;
  assign new_n35788_ = ys__n22844 & ~new_n12314_;
  assign new_n35789_ = new_n12309_ & new_n35788_;
  assign new_n35790_ = ~new_n17471_ & ~new_n35789_;
  assign new_n35791_ = ~new_n12320_ & ~new_n35790_;
  assign new_n35792_ = ys__n23566 & new_n12320_;
  assign new_n35793_ = ~new_n35791_ & ~new_n35792_;
  assign new_n35794_ = ~new_n12404_ & ~new_n35793_;
  assign new_n35795_ = new_n12404_ & ys__n23503;
  assign new_n35796_ = ~new_n35794_ & ~new_n35795_;
  assign new_n35797_ = new_n12458_ & ~new_n35796_;
  assign new_n35798_ = ys__n548 & ~new_n12458_;
  assign new_n35799_ = ~new_n35797_ & ~new_n35798_;
  assign new_n35800_ = ~new_n12477_ & ~new_n35799_;
  assign new_n35801_ = ~new_n12648_ & ~new_n35773_;
  assign new_n35802_ = ~new_n12680_ & ~new_n35801_;
  assign new_n35803_ = new_n12638_ & ~new_n35802_;
  assign new_n35804_ = ~new_n12638_ & new_n35802_;
  assign new_n35805_ = ~new_n35803_ & ~new_n35804_;
  assign new_n35806_ = new_n12477_ & ~new_n35805_;
  assign new_n35807_ = ~new_n35800_ & ~new_n35806_;
  assign new_n35808_ = new_n12763_ & ~new_n35807_;
  assign new_n35809_ = ~new_n35787_ & ~new_n35808_;
  assign new_n35810_ = new_n12774_ & ~new_n35809_;
  assign new_n35811_ = ys__n47672 & new_n12778_;
  assign new_n35812_ = new_n12776_ & ~new_n35807_;
  assign new_n35813_ = ~new_n35811_ & ~new_n35812_;
  assign new_n35814_ = new_n12784_ & ~new_n35813_;
  assign ys__n28536 = new_n35810_ | new_n35814_;
  assign new_n35816_ = ys__n47673 & new_n12768_;
  assign new_n35817_ = ys__n22846 & ~new_n12314_;
  assign new_n35818_ = new_n12309_ & new_n35817_;
  assign new_n35819_ = ~new_n17477_ & ~new_n35818_;
  assign new_n35820_ = ~new_n12320_ & ~new_n35819_;
  assign new_n35821_ = ys__n23568 & new_n12320_;
  assign new_n35822_ = ~new_n35820_ & ~new_n35821_;
  assign new_n35823_ = ~new_n12404_ & ~new_n35822_;
  assign new_n35824_ = new_n12404_ & ys__n23505;
  assign new_n35825_ = ~new_n35823_ & ~new_n35824_;
  assign new_n35826_ = new_n12458_ & ~new_n35825_;
  assign new_n35827_ = ys__n550 & ~new_n12458_;
  assign new_n35828_ = ~new_n35826_ & ~new_n35827_;
  assign new_n35829_ = ~new_n12477_ & ~new_n35828_;
  assign new_n35830_ = ~new_n12590_ & new_n12671_;
  assign new_n35831_ = new_n12683_ & ~new_n35830_;
  assign new_n35832_ = new_n12627_ & ~new_n35831_;
  assign new_n35833_ = ~new_n12627_ & new_n35831_;
  assign new_n35834_ = ~new_n35832_ & ~new_n35833_;
  assign new_n35835_ = new_n12477_ & ~new_n35834_;
  assign new_n35836_ = ~new_n35829_ & ~new_n35835_;
  assign new_n35837_ = new_n12763_ & ~new_n35836_;
  assign new_n35838_ = ~new_n35816_ & ~new_n35837_;
  assign new_n35839_ = new_n12774_ & ~new_n35838_;
  assign new_n35840_ = ys__n47673 & new_n12778_;
  assign new_n35841_ = new_n12776_ & ~new_n35836_;
  assign new_n35842_ = ~new_n35840_ & ~new_n35841_;
  assign new_n35843_ = new_n12784_ & ~new_n35842_;
  assign ys__n28539 = new_n35839_ | new_n35843_;
  assign new_n35845_ = ys__n47674 & new_n12768_;
  assign new_n35846_ = ys__n22848 & ~new_n12314_;
  assign new_n35847_ = new_n12309_ & new_n35846_;
  assign new_n35848_ = ~new_n17483_ & ~new_n35847_;
  assign new_n35849_ = ~new_n12320_ & ~new_n35848_;
  assign new_n35850_ = ys__n23570 & new_n12320_;
  assign new_n35851_ = ~new_n35849_ & ~new_n35850_;
  assign new_n35852_ = ~new_n12404_ & ~new_n35851_;
  assign new_n35853_ = new_n12404_ & ys__n23507;
  assign new_n35854_ = ~new_n35852_ & ~new_n35853_;
  assign new_n35855_ = new_n12458_ & ~new_n35854_;
  assign new_n35856_ = ys__n640 & ~new_n12458_;
  assign new_n35857_ = ~new_n35855_ & ~new_n35856_;
  assign new_n35858_ = ~new_n12477_ & ~new_n35857_;
  assign new_n35859_ = ~new_n12627_ & ~new_n35831_;
  assign new_n35860_ = ~new_n12686_ & ~new_n35859_;
  assign new_n35861_ = new_n12618_ & ~new_n35860_;
  assign new_n35862_ = ~new_n12618_ & new_n35860_;
  assign new_n35863_ = ~new_n35861_ & ~new_n35862_;
  assign new_n35864_ = new_n12477_ & ~new_n35863_;
  assign new_n35865_ = ~new_n35858_ & ~new_n35864_;
  assign new_n35866_ = new_n12763_ & ~new_n35865_;
  assign new_n35867_ = ~new_n35845_ & ~new_n35866_;
  assign new_n35868_ = new_n12774_ & ~new_n35867_;
  assign new_n35869_ = ys__n47674 & new_n12778_;
  assign new_n35870_ = new_n12776_ & ~new_n35865_;
  assign new_n35871_ = ~new_n35869_ & ~new_n35870_;
  assign new_n35872_ = new_n12784_ & ~new_n35871_;
  assign ys__n28542 = new_n35868_ | new_n35872_;
  assign new_n35874_ = ys__n47675 & new_n12768_;
  assign new_n35875_ = ys__n22850 & ~new_n12314_;
  assign new_n35876_ = new_n12309_ & new_n35875_;
  assign new_n35877_ = ~new_n17489_ & ~new_n35876_;
  assign new_n35878_ = ~new_n12320_ & ~new_n35877_;
  assign new_n35879_ = ys__n23572 & new_n12320_;
  assign new_n35880_ = ~new_n35878_ & ~new_n35879_;
  assign new_n35881_ = ~new_n12404_ & ~new_n35880_;
  assign new_n35882_ = new_n12404_ & ys__n23509;
  assign new_n35883_ = ~new_n35881_ & ~new_n35882_;
  assign new_n35884_ = new_n12458_ & ~new_n35883_;
  assign new_n35885_ = ys__n638 & ~new_n12458_;
  assign new_n35886_ = ~new_n35884_ & ~new_n35885_;
  assign new_n35887_ = ~new_n12477_ & ~new_n35886_;
  assign new_n35888_ = new_n12628_ & ~new_n35831_;
  assign new_n35889_ = new_n12688_ & ~new_n35888_;
  assign new_n35890_ = new_n12608_ & ~new_n35889_;
  assign new_n35891_ = ~new_n12608_ & new_n35889_;
  assign new_n35892_ = ~new_n35890_ & ~new_n35891_;
  assign new_n35893_ = new_n12477_ & ~new_n35892_;
  assign new_n35894_ = ~new_n35887_ & ~new_n35893_;
  assign new_n35895_ = new_n12763_ & ~new_n35894_;
  assign new_n35896_ = ~new_n35874_ & ~new_n35895_;
  assign new_n35897_ = new_n12774_ & ~new_n35896_;
  assign new_n35898_ = ys__n47675 & new_n12778_;
  assign new_n35899_ = new_n12776_ & ~new_n35894_;
  assign new_n35900_ = ~new_n35898_ & ~new_n35899_;
  assign new_n35901_ = new_n12784_ & ~new_n35900_;
  assign ys__n28545 = new_n35897_ | new_n35901_;
  assign new_n35903_ = ys__n47676 & new_n12768_;
  assign new_n35904_ = ys__n22852 & ~new_n12314_;
  assign new_n35905_ = new_n12309_ & new_n35904_;
  assign new_n35906_ = ~new_n17495_ & ~new_n35905_;
  assign new_n35907_ = ~new_n12320_ & ~new_n35906_;
  assign new_n35908_ = ys__n23574 & new_n12320_;
  assign new_n35909_ = ~new_n35907_ & ~new_n35908_;
  assign new_n35910_ = ~new_n12404_ & ~new_n35909_;
  assign new_n35911_ = new_n12404_ & ys__n23511;
  assign new_n35912_ = ~new_n35910_ & ~new_n35911_;
  assign new_n35913_ = new_n12458_ & ~new_n35912_;
  assign new_n35914_ = ys__n636 & ~new_n12458_;
  assign new_n35915_ = ~new_n35913_ & ~new_n35914_;
  assign new_n35916_ = ~new_n12477_ & ~new_n35915_;
  assign new_n35917_ = ~new_n12608_ & ~new_n35889_;
  assign new_n35918_ = ~new_n12691_ & ~new_n35917_;
  assign new_n35919_ = new_n12599_ & ~new_n35918_;
  assign new_n35920_ = ~new_n12599_ & new_n35918_;
  assign new_n35921_ = ~new_n35919_ & ~new_n35920_;
  assign new_n35922_ = new_n12477_ & ~new_n35921_;
  assign new_n35923_ = ~new_n35916_ & ~new_n35922_;
  assign new_n35924_ = new_n12763_ & ~new_n35923_;
  assign new_n35925_ = ~new_n35903_ & ~new_n35924_;
  assign new_n35926_ = new_n12774_ & ~new_n35925_;
  assign new_n35927_ = ys__n47676 & new_n12778_;
  assign new_n35928_ = new_n12776_ & ~new_n35923_;
  assign new_n35929_ = ~new_n35927_ & ~new_n35928_;
  assign new_n35930_ = new_n12784_ & ~new_n35929_;
  assign ys__n28548 = new_n35926_ | new_n35930_;
  assign new_n35932_ = ys__n47677 & new_n12768_;
  assign new_n35933_ = ys__n22854 & ~new_n12314_;
  assign new_n35934_ = new_n12309_ & new_n35933_;
  assign new_n35935_ = ~new_n17501_ & ~new_n35934_;
  assign new_n35936_ = ~new_n12320_ & ~new_n35935_;
  assign new_n35937_ = ys__n420 & new_n12320_;
  assign new_n35938_ = ~new_n35936_ & ~new_n35937_;
  assign new_n35939_ = ~new_n12404_ & ~new_n35938_;
  assign new_n35940_ = new_n12404_ & ys__n23513;
  assign new_n35941_ = ~new_n35939_ & ~new_n35940_;
  assign new_n35942_ = new_n12458_ & ~new_n35941_;
  assign new_n35943_ = ys__n634 & ~new_n12458_;
  assign new_n35944_ = ~new_n35942_ & ~new_n35943_;
  assign new_n35945_ = ~new_n12477_ & ~new_n35944_;
  assign new_n35946_ = new_n12495_ & ~new_n12696_;
  assign new_n35947_ = ~new_n12495_ & new_n12696_;
  assign new_n35948_ = ~new_n35946_ & ~new_n35947_;
  assign new_n35949_ = new_n12477_ & ~new_n35948_;
  assign new_n35950_ = ~new_n35945_ & ~new_n35949_;
  assign new_n35951_ = new_n12763_ & ~new_n35950_;
  assign new_n35952_ = ~new_n35932_ & ~new_n35951_;
  assign new_n35953_ = new_n12774_ & ~new_n35952_;
  assign new_n35954_ = ys__n47677 & new_n12778_;
  assign new_n35955_ = new_n12776_ & ~new_n35950_;
  assign new_n35956_ = ~new_n35954_ & ~new_n35955_;
  assign new_n35957_ = new_n12784_ & ~new_n35956_;
  assign ys__n28551 = new_n35953_ | new_n35957_;
  assign new_n35959_ = ys__n47678 & new_n12768_;
  assign new_n35960_ = ys__n22856 & ~new_n12314_;
  assign new_n35961_ = new_n12309_ & new_n35960_;
  assign new_n35962_ = ~new_n17507_ & ~new_n35961_;
  assign new_n35963_ = ~new_n12320_ & ~new_n35962_;
  assign new_n35964_ = ys__n442 & new_n12320_;
  assign new_n35965_ = ~new_n35963_ & ~new_n35964_;
  assign new_n35966_ = ~new_n12404_ & ~new_n35965_;
  assign new_n35967_ = new_n12404_ & ys__n23515;
  assign new_n35968_ = ~new_n35966_ & ~new_n35967_;
  assign new_n35969_ = new_n12458_ & ~new_n35968_;
  assign new_n35970_ = ys__n642 & ~new_n12458_;
  assign new_n35971_ = ~new_n35969_ & ~new_n35970_;
  assign new_n35972_ = ~new_n12477_ & ~new_n35971_;
  assign new_n35973_ = ys__n442 & ~new_n12703_;
  assign new_n35974_ = ~ys__n442 & new_n12737_;
  assign new_n35975_ = ~ys__n442 & new_n12753_;
  assign new_n35976_ = ~new_n35974_ & ~new_n35975_;
  assign new_n35977_ = ~new_n35973_ & new_n35976_;
  assign new_n35978_ = new_n12759_ & ~new_n35977_;
  assign new_n35979_ = ~new_n35972_ & ~new_n35978_;
  assign new_n35980_ = new_n12763_ & ~new_n35979_;
  assign new_n35981_ = ~new_n35959_ & ~new_n35980_;
  assign new_n35982_ = new_n12774_ & ~new_n35981_;
  assign new_n35983_ = ys__n47678 & new_n12778_;
  assign new_n35984_ = new_n12776_ & ~new_n35979_;
  assign new_n35985_ = ~new_n35983_ & ~new_n35984_;
  assign new_n35986_ = new_n12784_ & ~new_n35985_;
  assign ys__n28554 = new_n35982_ | new_n35986_;
  assign new_n35988_ = ys__n47679 & new_n12768_;
  assign new_n35989_ = ys__n22858 & ~new_n12314_;
  assign new_n35990_ = new_n12309_ & new_n35989_;
  assign new_n35991_ = ~new_n17513_ & ~new_n35990_;
  assign new_n35992_ = ~new_n12320_ & ~new_n35991_;
  assign new_n35993_ = ys__n440 & new_n12320_;
  assign new_n35994_ = ~new_n35992_ & ~new_n35993_;
  assign new_n35995_ = ~new_n12404_ & ~new_n35994_;
  assign new_n35996_ = new_n12404_ & ys__n23517;
  assign new_n35997_ = ~new_n35995_ & ~new_n35996_;
  assign new_n35998_ = new_n12458_ & ~new_n35997_;
  assign new_n35999_ = ys__n514 & ~ys__n28243;
  assign new_n36000_ = ys__n28243 & ys__n28632;
  assign new_n36001_ = ~new_n35999_ & ~new_n36000_;
  assign new_n36002_ = ~new_n12458_ & ~new_n36001_;
  assign new_n36003_ = ~new_n35998_ & ~new_n36002_;
  assign new_n36004_ = ~new_n12477_ & ~new_n36003_;
  assign new_n36005_ = ys__n440 & ~new_n12703_;
  assign new_n36006_ = ~ys__n440 & ~ys__n442;
  assign new_n36007_ = ~new_n12742_ & ~new_n36006_;
  assign new_n36008_ = new_n12737_ & ~new_n36007_;
  assign new_n36009_ = ys__n440 & ~ys__n442;
  assign new_n36010_ = ~new_n12705_ & ~new_n36009_;
  assign new_n36011_ = new_n12753_ & ~new_n36010_;
  assign new_n36012_ = ~new_n36008_ & ~new_n36011_;
  assign new_n36013_ = ~new_n36005_ & new_n36012_;
  assign new_n36014_ = new_n12759_ & ~new_n36013_;
  assign new_n36015_ = ~new_n36004_ & ~new_n36014_;
  assign new_n36016_ = new_n12763_ & ~new_n36015_;
  assign new_n36017_ = ~new_n35988_ & ~new_n36016_;
  assign new_n36018_ = new_n12774_ & ~new_n36017_;
  assign new_n36019_ = ys__n47679 & new_n12778_;
  assign new_n36020_ = new_n12776_ & ~new_n36015_;
  assign new_n36021_ = ~new_n36019_ & ~new_n36020_;
  assign new_n36022_ = new_n12784_ & ~new_n36021_;
  assign ys__n28557 = new_n36018_ | new_n36022_;
  assign new_n36024_ = ys__n47680 & new_n12768_;
  assign new_n36025_ = ys__n22860 & ~new_n12314_;
  assign new_n36026_ = new_n12309_ & new_n36025_;
  assign new_n36027_ = ~new_n17519_ & ~new_n36026_;
  assign new_n36028_ = ~new_n12320_ & ~new_n36027_;
  assign new_n36029_ = ys__n444 & new_n12320_;
  assign new_n36030_ = ~new_n36028_ & ~new_n36029_;
  assign new_n36031_ = ~new_n12404_ & ~new_n36030_;
  assign new_n36032_ = new_n12404_ & ys__n23519;
  assign new_n36033_ = ~new_n36031_ & ~new_n36032_;
  assign new_n36034_ = new_n12458_ & ~new_n36033_;
  assign new_n36035_ = ys__n2024 & ~ys__n28243;
  assign new_n36036_ = ys__n28243 & ys__n28633;
  assign new_n36037_ = ~new_n36035_ & ~new_n36036_;
  assign new_n36038_ = ~new_n12458_ & ~new_n36037_;
  assign new_n36039_ = ~new_n36034_ & ~new_n36038_;
  assign new_n36040_ = ~new_n12477_ & ~new_n36039_;
  assign new_n36041_ = ys__n444 & ~new_n12703_;
  assign new_n36042_ = ys__n444 & ~new_n12706_;
  assign new_n36043_ = ~ys__n444 & new_n12706_;
  assign new_n36044_ = ~new_n36042_ & ~new_n36043_;
  assign new_n36045_ = new_n12737_ & ~new_n36044_;
  assign new_n36046_ = ~ys__n444 & new_n12742_;
  assign new_n36047_ = ys__n444 & ~new_n12742_;
  assign new_n36048_ = ~new_n36046_ & ~new_n36047_;
  assign new_n36049_ = new_n12753_ & ~new_n36048_;
  assign new_n36050_ = ~new_n36045_ & ~new_n36049_;
  assign new_n36051_ = ~new_n36041_ & new_n36050_;
  assign new_n36052_ = new_n12759_ & ~new_n36051_;
  assign new_n36053_ = ~new_n36040_ & ~new_n36052_;
  assign new_n36054_ = new_n12763_ & ~new_n36053_;
  assign new_n36055_ = ~new_n36024_ & ~new_n36054_;
  assign new_n36056_ = new_n12774_ & ~new_n36055_;
  assign new_n36057_ = ys__n47680 & new_n12778_;
  assign new_n36058_ = new_n12776_ & ~new_n36053_;
  assign new_n36059_ = ~new_n36057_ & ~new_n36058_;
  assign new_n36060_ = new_n12784_ & ~new_n36059_;
  assign ys__n28560 = new_n36056_ | new_n36060_;
  assign new_n36062_ = ys__n47681 & new_n12768_;
  assign new_n36063_ = ys__n22862 & ~new_n12314_;
  assign new_n36064_ = new_n12309_ & new_n36063_;
  assign new_n36065_ = ~new_n17525_ & ~new_n36064_;
  assign new_n36066_ = ~new_n12320_ & ~new_n36065_;
  assign new_n36067_ = ys__n438 & new_n12320_;
  assign new_n36068_ = ~new_n36066_ & ~new_n36067_;
  assign new_n36069_ = ~new_n12404_ & ~new_n36068_;
  assign new_n36070_ = new_n12404_ & ys__n23521;
  assign new_n36071_ = ~new_n36069_ & ~new_n36070_;
  assign new_n36072_ = new_n12458_ & ~new_n36071_;
  assign new_n36073_ = ys__n4478 & ~ys__n28243;
  assign new_n36074_ = ys__n28243 & ys__n28634;
  assign new_n36075_ = ~new_n36073_ & ~new_n36074_;
  assign new_n36076_ = ~new_n12458_ & ~new_n36075_;
  assign new_n36077_ = ~new_n36072_ & ~new_n36076_;
  assign new_n36078_ = ~new_n12477_ & ~new_n36077_;
  assign new_n36079_ = ys__n438 & ~new_n12703_;
  assign new_n36080_ = ~ys__n444 & ~new_n12706_;
  assign new_n36081_ = ~ys__n444 & ~new_n36080_;
  assign new_n36082_ = ys__n438 & ~new_n36081_;
  assign new_n36083_ = ~ys__n438 & new_n36081_;
  assign new_n36084_ = ~new_n36082_ & ~new_n36083_;
  assign new_n36085_ = new_n12737_ & ~new_n36084_;
  assign new_n36086_ = ys__n444 & new_n12742_;
  assign new_n36087_ = ~ys__n438 & new_n36086_;
  assign new_n36088_ = ys__n438 & ~new_n36086_;
  assign new_n36089_ = ~new_n36087_ & ~new_n36088_;
  assign new_n36090_ = new_n12753_ & ~new_n36089_;
  assign new_n36091_ = ~new_n36085_ & ~new_n36090_;
  assign new_n36092_ = ~new_n36079_ & new_n36091_;
  assign new_n36093_ = new_n12759_ & ~new_n36092_;
  assign new_n36094_ = ~new_n36078_ & ~new_n36093_;
  assign new_n36095_ = new_n12763_ & ~new_n36094_;
  assign new_n36096_ = ~new_n36062_ & ~new_n36095_;
  assign new_n36097_ = new_n12774_ & ~new_n36096_;
  assign new_n36098_ = ys__n47681 & new_n12778_;
  assign new_n36099_ = new_n12776_ & ~new_n36094_;
  assign new_n36100_ = ~new_n36098_ & ~new_n36099_;
  assign new_n36101_ = new_n12784_ & ~new_n36100_;
  assign ys__n28563 = new_n36097_ | new_n36101_;
  assign new_n36103_ = ys__n22864 & new_n12309_;
  assign new_n36104_ = ~new_n17115_ & ~new_n36103_;
  assign new_n36105_ = ~new_n12314_ & ~new_n36104_;
  assign new_n36106_ = ~new_n17531_ & ~new_n36105_;
  assign new_n36107_ = ~new_n12320_ & ~new_n36106_;
  assign new_n36108_ = ys__n446 & new_n12320_;
  assign new_n36109_ = ~new_n36107_ & ~new_n36108_;
  assign new_n36110_ = ~new_n12404_ & ~new_n36109_;
  assign new_n36111_ = new_n12404_ & ys__n23523;
  assign new_n36112_ = ~new_n36110_ & ~new_n36111_;
  assign new_n36113_ = new_n12458_ & ~new_n36112_;
  assign new_n36114_ = ys__n4480 & ~ys__n28243;
  assign new_n36115_ = ys__n28243 & ys__n28635;
  assign new_n36116_ = ~new_n36114_ & ~new_n36115_;
  assign new_n36117_ = ~new_n12458_ & ~new_n36116_;
  assign new_n36118_ = ~new_n36113_ & ~new_n36117_;
  assign new_n36119_ = ~new_n12477_ & ~new_n36118_;
  assign new_n36120_ = ys__n446 & ~new_n12703_;
  assign new_n36121_ = ys__n446 & ~new_n12711_;
  assign new_n36122_ = ~ys__n446 & new_n12711_;
  assign new_n36123_ = ~new_n36121_ & ~new_n36122_;
  assign new_n36124_ = new_n12737_ & ~new_n36123_;
  assign new_n36125_ = ~ys__n446 & new_n12744_;
  assign new_n36126_ = ys__n446 & ~new_n12744_;
  assign new_n36127_ = ~new_n36125_ & ~new_n36126_;
  assign new_n36128_ = new_n12753_ & ~new_n36127_;
  assign new_n36129_ = ~new_n36124_ & ~new_n36128_;
  assign new_n36130_ = ~new_n36120_ & new_n36129_;
  assign new_n36131_ = new_n12759_ & ~new_n36130_;
  assign new_n36132_ = ~new_n36119_ & ~new_n36131_;
  assign new_n36133_ = new_n12763_ & ~new_n36132_;
  assign new_n36134_ = ys__n47682 & new_n12768_;
  assign new_n36135_ = ~new_n17155_ & ~new_n36134_;
  assign new_n36136_ = ~new_n36133_ & new_n36135_;
  assign new_n36137_ = new_n12774_ & ~new_n36136_;
  assign new_n36138_ = new_n12776_ & ~new_n36132_;
  assign new_n36139_ = ys__n47682 & new_n12778_;
  assign new_n36140_ = ~new_n17155_ & ~new_n36139_;
  assign new_n36141_ = ~new_n36138_ & new_n36140_;
  assign new_n36142_ = new_n12784_ & ~new_n36141_;
  assign ys__n28566 = new_n36137_ | new_n36142_;
  assign new_n36144_ = ~ys__n23627 & ~ys__n23629;
  assign new_n36145_ = ~new_n12309_ & new_n36144_;
  assign new_n36146_ = ys__n22866 & new_n12309_;
  assign new_n36147_ = ~new_n36145_ & ~new_n36146_;
  assign new_n36148_ = ~new_n12314_ & ~new_n36147_;
  assign new_n36149_ = ~new_n17537_ & ~new_n36148_;
  assign new_n36150_ = ~new_n12320_ & ~new_n36149_;
  assign new_n36151_ = ys__n434 & new_n12320_;
  assign new_n36152_ = ~new_n36150_ & ~new_n36151_;
  assign new_n36153_ = ~new_n12404_ & ~new_n36152_;
  assign new_n36154_ = new_n12404_ & ys__n23525;
  assign new_n36155_ = ~new_n36153_ & ~new_n36154_;
  assign new_n36156_ = new_n12458_ & ~new_n36155_;
  assign new_n36157_ = ys__n516 & ~ys__n28243;
  assign new_n36158_ = ys__n28243 & ys__n28636;
  assign new_n36159_ = ~new_n36157_ & ~new_n36158_;
  assign new_n36160_ = ~new_n12458_ & ~new_n36159_;
  assign new_n36161_ = ~new_n36156_ & ~new_n36160_;
  assign new_n36162_ = ~new_n12477_ & ~new_n36161_;
  assign new_n36163_ = ys__n434 & ~new_n12703_;
  assign new_n36164_ = ~ys__n446 & ~new_n12711_;
  assign new_n36165_ = ~ys__n446 & ~new_n36164_;
  assign new_n36166_ = ys__n434 & ~new_n36165_;
  assign new_n36167_ = ~ys__n434 & new_n36165_;
  assign new_n36168_ = ~new_n36166_ & ~new_n36167_;
  assign new_n36169_ = new_n12737_ & ~new_n36168_;
  assign new_n36170_ = ys__n446 & new_n12744_;
  assign new_n36171_ = ~ys__n434 & new_n36170_;
  assign new_n36172_ = ys__n434 & ~new_n36170_;
  assign new_n36173_ = ~new_n36171_ & ~new_n36172_;
  assign new_n36174_ = new_n12753_ & ~new_n36173_;
  assign new_n36175_ = ~new_n36169_ & ~new_n36174_;
  assign new_n36176_ = ~new_n36163_ & new_n36175_;
  assign new_n36177_ = new_n12759_ & ~new_n36176_;
  assign new_n36178_ = ~new_n36162_ & ~new_n36177_;
  assign new_n36179_ = new_n12763_ & ~new_n36178_;
  assign new_n36180_ = ys__n935 & ~ys__n23629;
  assign new_n36181_ = ~new_n12765_ & ~new_n36180_;
  assign new_n36182_ = new_n12762_ & ~new_n36181_;
  assign new_n36183_ = ys__n47683 & new_n12768_;
  assign new_n36184_ = ~new_n36182_ & ~new_n36183_;
  assign new_n36185_ = ~new_n36179_ & new_n36184_;
  assign new_n36186_ = new_n12774_ & ~new_n36185_;
  assign new_n36187_ = new_n12776_ & ~new_n36178_;
  assign new_n36188_ = ys__n47683 & new_n12778_;
  assign new_n36189_ = ~new_n36182_ & ~new_n36188_;
  assign new_n36190_ = ~new_n36187_ & new_n36189_;
  assign new_n36191_ = new_n12784_ & ~new_n36190_;
  assign ys__n28569 = new_n36186_ | new_n36191_;
  assign new_n36193_ = ys__n22868 & new_n12309_;
  assign new_n36194_ = ~new_n36145_ & ~new_n36193_;
  assign new_n36195_ = ~new_n12314_ & ~new_n36194_;
  assign new_n36196_ = ~new_n17543_ & ~new_n36195_;
  assign new_n36197_ = ~new_n12320_ & ~new_n36196_;
  assign new_n36198_ = ys__n436 & new_n12320_;
  assign new_n36199_ = ~new_n36197_ & ~new_n36198_;
  assign new_n36200_ = ~new_n12404_ & ~new_n36199_;
  assign new_n36201_ = new_n12404_ & ys__n23527;
  assign new_n36202_ = ~new_n36200_ & ~new_n36201_;
  assign new_n36203_ = new_n12458_ & ~new_n36202_;
  assign new_n36204_ = ys__n4494 & ~ys__n28243;
  assign new_n36205_ = ys__n28243 & ys__n28637;
  assign new_n36206_ = ~new_n36204_ & ~new_n36205_;
  assign new_n36207_ = ~new_n12458_ & ~new_n36206_;
  assign new_n36208_ = ~new_n36203_ & ~new_n36207_;
  assign new_n36209_ = ~new_n12477_ & ~new_n36208_;
  assign new_n36210_ = ys__n436 & ~new_n12703_;
  assign new_n36211_ = ~new_n12711_ & new_n12713_;
  assign new_n36212_ = new_n12717_ & ~new_n36211_;
  assign new_n36213_ = ys__n436 & ~new_n36212_;
  assign new_n36214_ = ~ys__n436 & new_n36212_;
  assign new_n36215_ = ~new_n36213_ & ~new_n36214_;
  assign new_n36216_ = new_n12737_ & ~new_n36215_;
  assign new_n36217_ = new_n12744_ & new_n12745_;
  assign new_n36218_ = ~ys__n436 & new_n36217_;
  assign new_n36219_ = ys__n436 & ~new_n36217_;
  assign new_n36220_ = ~new_n36218_ & ~new_n36219_;
  assign new_n36221_ = new_n12753_ & ~new_n36220_;
  assign new_n36222_ = ~new_n36216_ & ~new_n36221_;
  assign new_n36223_ = ~new_n36210_ & new_n36222_;
  assign new_n36224_ = new_n12759_ & ~new_n36223_;
  assign new_n36225_ = ~new_n36209_ & ~new_n36224_;
  assign new_n36226_ = new_n12763_ & ~new_n36225_;
  assign new_n36227_ = ys__n47684 & new_n12768_;
  assign new_n36228_ = ~new_n36182_ & ~new_n36227_;
  assign new_n36229_ = ~new_n36226_ & new_n36228_;
  assign new_n36230_ = new_n12774_ & ~new_n36229_;
  assign new_n36231_ = new_n12776_ & ~new_n36225_;
  assign new_n36232_ = ys__n47684 & new_n12778_;
  assign new_n36233_ = ~new_n36182_ & ~new_n36232_;
  assign new_n36234_ = ~new_n36231_ & new_n36233_;
  assign new_n36235_ = new_n12784_ & ~new_n36234_;
  assign ys__n28572 = new_n36230_ | new_n36235_;
  assign new_n36237_ = ys__n22870 & new_n12309_;
  assign new_n36238_ = ~new_n12310_ & ~new_n36237_;
  assign new_n36239_ = ~new_n12314_ & ~new_n36238_;
  assign new_n36240_ = ~new_n17549_ & ~new_n36239_;
  assign new_n36241_ = ~new_n12320_ & ~new_n36240_;
  assign new_n36242_ = ys__n432 & new_n12320_;
  assign new_n36243_ = ~new_n36241_ & ~new_n36242_;
  assign new_n36244_ = ~new_n12404_ & ~new_n36243_;
  assign new_n36245_ = new_n12404_ & ys__n23529;
  assign new_n36246_ = ~new_n36244_ & ~new_n36245_;
  assign new_n36247_ = new_n12458_ & ~new_n36246_;
  assign new_n36248_ = ys__n4496 & ~ys__n28243;
  assign new_n36249_ = ys__n28243 & ys__n28638;
  assign new_n36250_ = ~new_n36248_ & ~new_n36249_;
  assign new_n36251_ = ~new_n12458_ & ~new_n36250_;
  assign new_n36252_ = ~new_n36247_ & ~new_n36251_;
  assign new_n36253_ = ~new_n12477_ & ~new_n36252_;
  assign new_n36254_ = ys__n432 & ~new_n12703_;
  assign new_n36255_ = ~ys__n436 & ~new_n36212_;
  assign new_n36256_ = ~ys__n436 & ~new_n36255_;
  assign new_n36257_ = ys__n432 & ~new_n36256_;
  assign new_n36258_ = ~ys__n432 & new_n36256_;
  assign new_n36259_ = ~new_n36257_ & ~new_n36258_;
  assign new_n36260_ = new_n12737_ & ~new_n36259_;
  assign new_n36261_ = ys__n436 & new_n36217_;
  assign new_n36262_ = ~ys__n432 & new_n36261_;
  assign new_n36263_ = ys__n432 & ~new_n36261_;
  assign new_n36264_ = ~new_n36262_ & ~new_n36263_;
  assign new_n36265_ = new_n12753_ & ~new_n36264_;
  assign new_n36266_ = ~new_n36260_ & ~new_n36265_;
  assign new_n36267_ = ~new_n36254_ & new_n36266_;
  assign new_n36268_ = new_n12759_ & ~new_n36267_;
  assign new_n36269_ = ~new_n36253_ & ~new_n36268_;
  assign new_n36270_ = new_n12763_ & ~new_n36269_;
  assign new_n36271_ = ys__n47685 & new_n12768_;
  assign new_n36272_ = ~new_n12767_ & ~new_n36271_;
  assign new_n36273_ = ~new_n36270_ & new_n36272_;
  assign new_n36274_ = new_n12774_ & ~new_n36273_;
  assign new_n36275_ = new_n12776_ & ~new_n36269_;
  assign new_n36276_ = ys__n47685 & new_n12778_;
  assign new_n36277_ = ~new_n12767_ & ~new_n36276_;
  assign new_n36278_ = ~new_n36275_ & new_n36277_;
  assign new_n36279_ = new_n12784_ & ~new_n36278_;
  assign ys__n28575 = new_n36274_ | new_n36279_;
  assign new_n36281_ = ys__n22872 & new_n12309_;
  assign new_n36282_ = ~new_n12310_ & ~new_n36281_;
  assign new_n36283_ = ~new_n12314_ & ~new_n36282_;
  assign new_n36284_ = ~new_n17555_ & ~new_n36283_;
  assign new_n36285_ = ~new_n12320_ & ~new_n36284_;
  assign new_n36286_ = ys__n448 & new_n12320_;
  assign new_n36287_ = ~new_n36285_ & ~new_n36286_;
  assign new_n36288_ = ~new_n12404_ & ~new_n36287_;
  assign new_n36289_ = new_n12404_ & ys__n23531;
  assign new_n36290_ = ~new_n36288_ & ~new_n36289_;
  assign new_n36291_ = new_n12458_ & ~new_n36290_;
  assign new_n36292_ = ys__n632 & ~ys__n28243;
  assign new_n36293_ = ys__n28243 & ys__n28639;
  assign new_n36294_ = ~new_n36292_ & ~new_n36293_;
  assign new_n36295_ = ~new_n12458_ & ~new_n36294_;
  assign new_n36296_ = ~new_n36291_ & ~new_n36295_;
  assign new_n36297_ = ~new_n12477_ & ~new_n36296_;
  assign new_n36298_ = ys__n448 & ~new_n12703_;
  assign new_n36299_ = ys__n448 & ~new_n12722_;
  assign new_n36300_ = ~ys__n448 & new_n12722_;
  assign new_n36301_ = ~new_n36299_ & ~new_n36300_;
  assign new_n36302_ = new_n12737_ & ~new_n36301_;
  assign new_n36303_ = ~ys__n448 & new_n12748_;
  assign new_n36304_ = ys__n448 & ~new_n12748_;
  assign new_n36305_ = ~new_n36303_ & ~new_n36304_;
  assign new_n36306_ = new_n12753_ & ~new_n36305_;
  assign new_n36307_ = ~new_n36302_ & ~new_n36306_;
  assign new_n36308_ = ~new_n36298_ & new_n36307_;
  assign new_n36309_ = new_n12759_ & ~new_n36308_;
  assign new_n36310_ = ~new_n36297_ & ~new_n36309_;
  assign new_n36311_ = new_n12763_ & ~new_n36310_;
  assign new_n36312_ = ys__n47686 & new_n12768_;
  assign new_n36313_ = ~new_n12767_ & ~new_n36312_;
  assign new_n36314_ = ~new_n36311_ & new_n36313_;
  assign new_n36315_ = new_n12774_ & ~new_n36314_;
  assign new_n36316_ = new_n12776_ & ~new_n36310_;
  assign new_n36317_ = ys__n47686 & new_n12778_;
  assign new_n36318_ = ~new_n12767_ & ~new_n36317_;
  assign new_n36319_ = ~new_n36316_ & new_n36318_;
  assign new_n36320_ = new_n12784_ & ~new_n36319_;
  assign ys__n28578 = new_n36315_ | new_n36320_;
  assign new_n36322_ = ys__n22874 & new_n12309_;
  assign new_n36323_ = ~new_n12310_ & ~new_n36322_;
  assign new_n36324_ = ~new_n12314_ & ~new_n36323_;
  assign new_n36325_ = ~new_n17561_ & ~new_n36324_;
  assign new_n36326_ = ~new_n12320_ & ~new_n36325_;
  assign new_n36327_ = ys__n428 & new_n12320_;
  assign new_n36328_ = ~new_n36326_ & ~new_n36327_;
  assign new_n36329_ = ~new_n12404_ & ~new_n36328_;
  assign new_n36330_ = new_n12404_ & ys__n23533;
  assign new_n36331_ = ~new_n36329_ & ~new_n36330_;
  assign new_n36332_ = new_n12458_ & ~new_n36331_;
  assign new_n36333_ = ys__n512 & ~ys__n28243;
  assign new_n36334_ = ys__n28243 & ys__n28640;
  assign new_n36335_ = ~new_n36333_ & ~new_n36334_;
  assign new_n36336_ = ~new_n12458_ & ~new_n36335_;
  assign new_n36337_ = ~new_n36332_ & ~new_n36336_;
  assign new_n36338_ = ~new_n12477_ & ~new_n36337_;
  assign new_n36339_ = ys__n428 & ~new_n12703_;
  assign new_n36340_ = ~ys__n448 & ~new_n12722_;
  assign new_n36341_ = ~ys__n448 & ~new_n36340_;
  assign new_n36342_ = ys__n428 & ~new_n36341_;
  assign new_n36343_ = ~ys__n428 & new_n36341_;
  assign new_n36344_ = ~new_n36342_ & ~new_n36343_;
  assign new_n36345_ = new_n12737_ & ~new_n36344_;
  assign new_n36346_ = ys__n448 & new_n12748_;
  assign new_n36347_ = ~ys__n428 & new_n36346_;
  assign new_n36348_ = ys__n428 & ~new_n36346_;
  assign new_n36349_ = ~new_n36347_ & ~new_n36348_;
  assign new_n36350_ = new_n12753_ & ~new_n36349_;
  assign new_n36351_ = ~new_n36345_ & ~new_n36350_;
  assign new_n36352_ = ~new_n36339_ & new_n36351_;
  assign new_n36353_ = new_n12759_ & ~new_n36352_;
  assign new_n36354_ = ~new_n36338_ & ~new_n36353_;
  assign new_n36355_ = new_n12763_ & ~new_n36354_;
  assign new_n36356_ = ys__n47687 & new_n12768_;
  assign new_n36357_ = ~new_n12767_ & ~new_n36356_;
  assign new_n36358_ = ~new_n36355_ & new_n36357_;
  assign new_n36359_ = new_n12774_ & ~new_n36358_;
  assign new_n36360_ = new_n12776_ & ~new_n36354_;
  assign new_n36361_ = ys__n47687 & new_n12778_;
  assign new_n36362_ = ~new_n12767_ & ~new_n36361_;
  assign new_n36363_ = ~new_n36360_ & new_n36362_;
  assign new_n36364_ = new_n12784_ & ~new_n36363_;
  assign ys__n28581 = new_n36359_ | new_n36364_;
  assign new_n36366_ = ys__n22876 & new_n12309_;
  assign new_n36367_ = ~new_n12310_ & ~new_n36366_;
  assign new_n36368_ = ~new_n12314_ & ~new_n36367_;
  assign new_n36369_ = ~new_n17567_ & ~new_n36368_;
  assign new_n36370_ = ~new_n12320_ & ~new_n36369_;
  assign new_n36371_ = ys__n430 & new_n12320_;
  assign new_n36372_ = ~new_n36370_ & ~new_n36371_;
  assign new_n36373_ = ~new_n12404_ & ~new_n36372_;
  assign new_n36374_ = new_n12404_ & ys__n23535;
  assign new_n36375_ = ~new_n36373_ & ~new_n36374_;
  assign new_n36376_ = new_n12458_ & ~new_n36375_;
  assign new_n36377_ = ys__n520 & ~ys__n28243;
  assign new_n36378_ = ys__n28243 & ys__n28641;
  assign new_n36379_ = ~new_n36377_ & ~new_n36378_;
  assign new_n36380_ = ~new_n12458_ & ~new_n36379_;
  assign new_n36381_ = ~new_n36376_ & ~new_n36380_;
  assign new_n36382_ = ~new_n12477_ & ~new_n36381_;
  assign new_n36383_ = ys__n430 & ~new_n12703_;
  assign new_n36384_ = ~new_n12722_ & new_n12724_;
  assign new_n36385_ = new_n12728_ & ~new_n36384_;
  assign new_n36386_ = ys__n430 & ~new_n36385_;
  assign new_n36387_ = ~ys__n430 & new_n36385_;
  assign new_n36388_ = ~new_n36386_ & ~new_n36387_;
  assign new_n36389_ = new_n12737_ & ~new_n36388_;
  assign new_n36390_ = new_n12739_ & new_n12748_;
  assign new_n36391_ = ~ys__n430 & new_n36390_;
  assign new_n36392_ = ys__n430 & ~new_n36390_;
  assign new_n36393_ = ~new_n36391_ & ~new_n36392_;
  assign new_n36394_ = new_n12753_ & ~new_n36393_;
  assign new_n36395_ = ~new_n36389_ & ~new_n36394_;
  assign new_n36396_ = ~new_n36383_ & new_n36395_;
  assign new_n36397_ = new_n12759_ & ~new_n36396_;
  assign new_n36398_ = ~new_n36382_ & ~new_n36397_;
  assign new_n36399_ = new_n12763_ & ~new_n36398_;
  assign new_n36400_ = ys__n47688 & new_n12768_;
  assign new_n36401_ = ~new_n12767_ & ~new_n36400_;
  assign new_n36402_ = ~new_n36399_ & new_n36401_;
  assign new_n36403_ = new_n12774_ & ~new_n36402_;
  assign new_n36404_ = new_n12776_ & ~new_n36398_;
  assign new_n36405_ = ys__n47688 & new_n12778_;
  assign new_n36406_ = ~new_n12767_ & ~new_n36405_;
  assign new_n36407_ = ~new_n36404_ & new_n36406_;
  assign new_n36408_ = new_n12784_ & ~new_n36407_;
  assign ys__n28584 = new_n36403_ | new_n36408_;
  assign new_n36410_ = ys__n22878 & new_n12309_;
  assign new_n36411_ = ~new_n12310_ & ~new_n36410_;
  assign new_n36412_ = ~new_n12314_ & ~new_n36411_;
  assign new_n36413_ = ~new_n17573_ & ~new_n36412_;
  assign new_n36414_ = ~new_n12320_ & ~new_n36413_;
  assign new_n36415_ = ys__n426 & new_n12320_;
  assign new_n36416_ = ~new_n36414_ & ~new_n36415_;
  assign new_n36417_ = ~new_n12404_ & ~new_n36416_;
  assign new_n36418_ = new_n12404_ & ys__n23537;
  assign new_n36419_ = ~new_n36417_ & ~new_n36418_;
  assign new_n36420_ = new_n12458_ & ~new_n36419_;
  assign new_n36421_ = ys__n426 & ~new_n12458_;
  assign new_n36422_ = ~new_n36420_ & ~new_n36421_;
  assign new_n36423_ = ~new_n12477_ & ~new_n36422_;
  assign new_n36424_ = ys__n426 & ~new_n12703_;
  assign new_n36425_ = ~ys__n430 & ~new_n36385_;
  assign new_n36426_ = ~ys__n430 & ~new_n36425_;
  assign new_n36427_ = ys__n426 & ~new_n36426_;
  assign new_n36428_ = ~ys__n426 & new_n36426_;
  assign new_n36429_ = ~new_n36427_ & ~new_n36428_;
  assign new_n36430_ = new_n12737_ & ~new_n36429_;
  assign new_n36431_ = ys__n430 & new_n36390_;
  assign new_n36432_ = ~ys__n426 & new_n36431_;
  assign new_n36433_ = ys__n426 & ~new_n36431_;
  assign new_n36434_ = ~new_n36432_ & ~new_n36433_;
  assign new_n36435_ = new_n12753_ & ~new_n36434_;
  assign new_n36436_ = ~new_n36430_ & ~new_n36435_;
  assign new_n36437_ = ~new_n36424_ & new_n36436_;
  assign new_n36438_ = new_n12759_ & ~new_n36437_;
  assign new_n36439_ = ~new_n36423_ & ~new_n36438_;
  assign new_n36440_ = new_n12763_ & ~new_n36439_;
  assign new_n36441_ = ys__n47689 & new_n12768_;
  assign new_n36442_ = ~new_n12767_ & ~new_n36441_;
  assign new_n36443_ = ~new_n36440_ & new_n36442_;
  assign new_n36444_ = new_n12774_ & ~new_n36443_;
  assign new_n36445_ = new_n12776_ & ~new_n36439_;
  assign new_n36446_ = ys__n47689 & new_n12778_;
  assign new_n36447_ = ~new_n12767_ & ~new_n36446_;
  assign new_n36448_ = ~new_n36445_ & new_n36447_;
  assign new_n36449_ = new_n12784_ & ~new_n36448_;
  assign ys__n28587 = new_n36444_ | new_n36449_;
  assign ys__n28661 = ys__n532 & ~ys__n28243;
  assign ys__n28662 = ys__n746 & ~ys__n28243;
  assign new_n36453_ = ~ys__n860 & new_n12120_;
  assign new_n36454_ = ~ys__n204 & new_n36453_;
  assign new_n36455_ = ~ys__n182 & ys__n192;
  assign new_n36456_ = new_n36454_ & new_n36455_;
  assign new_n36457_ = ys__n182 & ~ys__n184;
  assign new_n36458_ = ys__n204 & new_n36453_;
  assign new_n36459_ = new_n36457_ & new_n36458_;
  assign new_n36460_ = ~ys__n182 & ys__n204;
  assign new_n36461_ = new_n36453_ & new_n36460_;
  assign new_n36462_ = new_n36453_ & ~new_n36461_;
  assign new_n36463_ = ~new_n36459_ & new_n36462_;
  assign new_n36464_ = ~new_n36456_ & new_n36463_;
  assign new_n36465_ = ys__n182 & ys__n192;
  assign new_n36466_ = new_n36454_ & new_n36465_;
  assign new_n36467_ = ys__n182 & ys__n184;
  assign new_n36468_ = new_n36458_ & new_n36467_;
  assign new_n36469_ = ~ys__n192 & ~ys__n204;
  assign new_n36470_ = new_n36453_ & new_n36469_;
  assign new_n36471_ = ~new_n36468_ & ~new_n36470_;
  assign new_n36472_ = ~new_n36466_ & new_n36471_;
  assign new_n36473_ = new_n36464_ & new_n36472_;
  assign new_n36474_ = ys__n190 & new_n36467_;
  assign new_n36475_ = ys__n190 & new_n36457_;
  assign new_n36476_ = ~new_n36474_ & ~new_n36475_;
  assign new_n36477_ = ~ys__n182 & ys__n184;
  assign new_n36478_ = ys__n190 & new_n36477_;
  assign new_n36479_ = ~ys__n182 & ~ys__n184;
  assign new_n36480_ = ~ys__n190 & new_n36479_;
  assign new_n36481_ = ~new_n36478_ & ~new_n36480_;
  assign new_n36482_ = new_n36476_ & new_n36481_;
  assign new_n36483_ = ~new_n36457_ & ~new_n36467_;
  assign new_n36484_ = ~new_n36477_ & ~new_n36479_;
  assign new_n36485_ = new_n36483_ & new_n36484_;
  assign new_n36486_ = ~new_n36482_ & ~new_n36485_;
  assign new_n36487_ = ~new_n36464_ & new_n36486_;
  assign new_n36488_ = ~new_n36473_ & new_n36487_;
  assign new_n36489_ = ys__n4566 & new_n13716_;
  assign new_n36490_ = new_n36488_ & new_n36489_;
  assign new_n36491_ = ~new_n12139_ & new_n13713_;
  assign new_n36492_ = new_n36488_ & new_n36491_;
  assign new_n36493_ = ys__n186 & ~ys__n202;
  assign new_n36494_ = new_n36477_ & new_n36493_;
  assign new_n36495_ = ~ys__n38453 & new_n36494_;
  assign new_n36496_ = ~ys__n186 & ~ys__n202;
  assign new_n36497_ = new_n36477_ & new_n36496_;
  assign new_n36498_ = ~ys__n38453 & new_n36497_;
  assign new_n36499_ = ~new_n36495_ & ~new_n36498_;
  assign new_n36500_ = new_n36457_ & new_n36493_;
  assign new_n36501_ = ~ys__n38453 & new_n36500_;
  assign new_n36502_ = ~ys__n186 & ys__n202;
  assign new_n36503_ = new_n36457_ & new_n36502_;
  assign new_n36504_ = ~ys__n38453 & new_n36503_;
  assign new_n36505_ = ~new_n36501_ & ~new_n36504_;
  assign new_n36506_ = new_n36499_ & new_n36505_;
  assign new_n36507_ = ys__n38453 & new_n36502_;
  assign new_n36508_ = ys__n186 & ys__n202;
  assign new_n36509_ = new_n36467_ & new_n36508_;
  assign new_n36510_ = ~ys__n38453 & new_n36509_;
  assign new_n36511_ = ~new_n36507_ & ~new_n36510_;
  assign new_n36512_ = new_n36467_ & new_n36496_;
  assign new_n36513_ = ~ys__n38453 & new_n36512_;
  assign new_n36514_ = new_n36467_ & new_n36502_;
  assign new_n36515_ = ~ys__n38453 & new_n36514_;
  assign new_n36516_ = ~new_n36513_ & ~new_n36515_;
  assign new_n36517_ = new_n36511_ & new_n36516_;
  assign new_n36518_ = new_n36506_ & new_n36517_;
  assign new_n36519_ = new_n36467_ & new_n36493_;
  assign new_n36520_ = ~ys__n38453 & new_n36519_;
  assign new_n36521_ = ys__n38453 & new_n36496_;
  assign new_n36522_ = new_n36479_ & new_n36502_;
  assign new_n36523_ = ~ys__n38453 & new_n36522_;
  assign new_n36524_ = ~new_n36521_ & ~new_n36523_;
  assign new_n36525_ = ~new_n36520_ & new_n36524_;
  assign new_n36526_ = new_n36479_ & new_n36496_;
  assign new_n36527_ = ~ys__n38453 & new_n36526_;
  assign new_n36528_ = new_n36477_ & new_n36502_;
  assign new_n36529_ = ~ys__n38453 & new_n36528_;
  assign new_n36530_ = ~new_n36527_ & ~new_n36529_;
  assign new_n36531_ = new_n36457_ & new_n36508_;
  assign new_n36532_ = ~ys__n38453 & new_n36531_;
  assign new_n36533_ = new_n36530_ & ~new_n36532_;
  assign new_n36534_ = new_n36525_ & new_n36533_;
  assign new_n36535_ = new_n36457_ & new_n36496_;
  assign new_n36536_ = ~ys__n38453 & new_n36535_;
  assign new_n36537_ = new_n36479_ & new_n36493_;
  assign new_n36538_ = ~ys__n38453 & new_n36537_;
  assign new_n36539_ = new_n36477_ & new_n36508_;
  assign new_n36540_ = ~ys__n38453 & new_n36539_;
  assign new_n36541_ = ~new_n36538_ & ~new_n36540_;
  assign new_n36542_ = ~new_n36536_ & new_n36541_;
  assign new_n36543_ = ys__n38453 & new_n36493_;
  assign new_n36544_ = new_n36479_ & new_n36508_;
  assign new_n36545_ = ~ys__n38453 & new_n36544_;
  assign new_n36546_ = ~new_n36543_ & ~new_n36545_;
  assign new_n36547_ = ys__n38453 & new_n36508_;
  assign new_n36548_ = new_n36546_ & ~new_n36547_;
  assign new_n36549_ = new_n36542_ & new_n36548_;
  assign new_n36550_ = new_n36534_ & new_n36549_;
  assign new_n36551_ = new_n36518_ & new_n36550_;
  assign new_n36552_ = ~new_n36513_ & new_n36525_;
  assign new_n36553_ = ~new_n36501_ & ~new_n36536_;
  assign new_n36554_ = new_n36499_ & new_n36553_;
  assign new_n36555_ = new_n36546_ & new_n36554_;
  assign new_n36556_ = new_n36552_ & new_n36555_;
  assign new_n36557_ = new_n12139_ & ~new_n36556_;
  assign new_n36558_ = ~new_n36551_ & new_n36557_;
  assign new_n36559_ = ~new_n36492_ & ~new_n36558_;
  assign new_n36560_ = ~new_n12139_ & ~new_n36491_;
  assign new_n36561_ = ~ys__n4566 & ~new_n36560_;
  assign new_n36562_ = ~new_n36559_ & new_n36561_;
  assign new_n36563_ = ~new_n36490_ & ~new_n36562_;
  assign new_n36564_ = ~ys__n738 & ~new_n36563_;
  assign new_n36565_ = ys__n738 & new_n13713_;
  assign new_n36566_ = new_n36488_ & new_n36565_;
  assign ys__n28781 = new_n36564_ | new_n36566_;
  assign new_n36568_ = ys__n190 & ys__n192;
  assign new_n36569_ = ~new_n12121_ & ~new_n36568_;
  assign new_n36570_ = new_n36479_ & ~new_n36569_;
  assign new_n36571_ = ~ys__n192 & new_n36477_;
  assign new_n36572_ = ys__n192 & new_n36467_;
  assign new_n36573_ = ys__n192 & new_n36457_;
  assign new_n36574_ = ~new_n36572_ & ~new_n36573_;
  assign new_n36575_ = ~new_n36571_ & new_n36574_;
  assign new_n36576_ = ~new_n36570_ & new_n36575_;
  assign new_n36577_ = ~new_n36485_ & ~new_n36576_;
  assign new_n36578_ = ~new_n36464_ & new_n36577_;
  assign new_n36579_ = ~new_n36473_ & new_n36578_;
  assign new_n36580_ = new_n36489_ & new_n36579_;
  assign new_n36581_ = new_n36491_ & new_n36579_;
  assign new_n36582_ = ~new_n36501_ & new_n36546_;
  assign new_n36583_ = new_n36530_ & new_n36582_;
  assign new_n36584_ = new_n36542_ & new_n36583_;
  assign new_n36585_ = new_n36552_ & new_n36584_;
  assign new_n36586_ = new_n12139_ & ~new_n36551_;
  assign new_n36587_ = ~new_n36585_ & new_n36586_;
  assign new_n36588_ = ~new_n36581_ & ~new_n36587_;
  assign new_n36589_ = new_n36561_ & ~new_n36588_;
  assign new_n36590_ = ~new_n36580_ & ~new_n36589_;
  assign new_n36591_ = ~ys__n738 & ~new_n36590_;
  assign new_n36592_ = new_n36565_ & new_n36579_;
  assign ys__n28782 = new_n36591_ | new_n36592_;
  assign new_n36594_ = ys__n190 & ~ys__n192;
  assign new_n36595_ = ~ys__n192 & ~new_n36594_;
  assign new_n36596_ = ys__n204 & ~new_n36595_;
  assign new_n36597_ = ~ys__n204 & new_n36595_;
  assign new_n36598_ = ~new_n36596_ & ~new_n36597_;
  assign new_n36599_ = new_n36479_ & ~new_n36598_;
  assign new_n36600_ = ys__n192 & ys__n204;
  assign new_n36601_ = ~new_n36469_ & ~new_n36600_;
  assign new_n36602_ = new_n36477_ & ~new_n36601_;
  assign new_n36603_ = ys__n204 & new_n36467_;
  assign new_n36604_ = ~ys__n204 & new_n36457_;
  assign new_n36605_ = ~new_n36603_ & ~new_n36604_;
  assign new_n36606_ = ~new_n36602_ & new_n36605_;
  assign new_n36607_ = ~new_n36599_ & new_n36606_;
  assign new_n36608_ = ~new_n36464_ & ~new_n36485_;
  assign new_n36609_ = ~new_n36607_ & new_n36608_;
  assign new_n36610_ = ~new_n36473_ & new_n36609_;
  assign new_n36611_ = new_n36489_ & new_n36610_;
  assign new_n36612_ = new_n36491_ & new_n36610_;
  assign new_n36613_ = new_n36499_ & ~new_n36504_;
  assign new_n36614_ = new_n36541_ & new_n36546_;
  assign new_n36615_ = new_n36613_ & new_n36614_;
  assign new_n36616_ = new_n36533_ & new_n36615_;
  assign new_n36617_ = new_n36552_ & new_n36616_;
  assign new_n36618_ = new_n36586_ & ~new_n36617_;
  assign new_n36619_ = ~new_n36612_ & ~new_n36618_;
  assign new_n36620_ = new_n36561_ & ~new_n36619_;
  assign new_n36621_ = ~new_n36611_ & ~new_n36620_;
  assign new_n36622_ = ~ys__n738 & ~new_n36621_;
  assign new_n36623_ = new_n36565_ & new_n36610_;
  assign ys__n28783 = new_n36622_ | new_n36623_;
  assign new_n36625_ = ~ys__n204 & ~new_n36595_;
  assign new_n36626_ = ~ys__n204 & ~new_n36625_;
  assign new_n36627_ = ys__n860 & ~new_n36626_;
  assign new_n36628_ = ~ys__n860 & new_n36626_;
  assign new_n36629_ = ~new_n36627_ & ~new_n36628_;
  assign new_n36630_ = new_n36479_ & ~new_n36629_;
  assign new_n36631_ = ys__n192 & ~ys__n204;
  assign new_n36632_ = ~ys__n204 & ~new_n36631_;
  assign new_n36633_ = ys__n860 & ~new_n36632_;
  assign new_n36634_ = ~ys__n860 & new_n36632_;
  assign new_n36635_ = ~new_n36633_ & ~new_n36634_;
  assign new_n36636_ = new_n36477_ & ~new_n36635_;
  assign new_n36637_ = ~ys__n860 & new_n36467_;
  assign new_n36638_ = ys__n204 & ys__n860;
  assign new_n36639_ = ~new_n12122_ & ~new_n36638_;
  assign new_n36640_ = new_n36457_ & ~new_n36639_;
  assign new_n36641_ = ~new_n36637_ & ~new_n36640_;
  assign new_n36642_ = ~new_n36636_ & new_n36641_;
  assign new_n36643_ = ~new_n36630_ & new_n36642_;
  assign new_n36644_ = ~new_n36473_ & new_n36608_;
  assign new_n36645_ = ~new_n36643_ & new_n36644_;
  assign new_n36646_ = new_n36489_ & new_n36645_;
  assign new_n36647_ = new_n36491_ & new_n36645_;
  assign new_n36648_ = ~new_n36504_ & new_n36530_;
  assign new_n36649_ = ~new_n36498_ & ~new_n36536_;
  assign new_n36650_ = ~new_n36515_ & ~new_n36547_;
  assign new_n36651_ = new_n36649_ & new_n36650_;
  assign new_n36652_ = new_n36525_ & new_n36651_;
  assign new_n36653_ = new_n36648_ & new_n36652_;
  assign new_n36654_ = new_n12139_ & ~new_n36653_;
  assign new_n36655_ = ~new_n36551_ & new_n36654_;
  assign new_n36656_ = ~new_n36647_ & ~new_n36655_;
  assign new_n36657_ = new_n36561_ & ~new_n36656_;
  assign new_n36658_ = ~new_n36646_ & ~new_n36657_;
  assign new_n36659_ = ~ys__n738 & ~new_n36658_;
  assign new_n36660_ = new_n36565_ & new_n36645_;
  assign ys__n28784 = new_n36659_ | new_n36660_;
  assign new_n36662_ = ys__n204 & ~ys__n860;
  assign new_n36663_ = ~ys__n860 & ~new_n36662_;
  assign new_n36664_ = new_n12122_ & ~new_n36595_;
  assign new_n36665_ = new_n36663_ & ~new_n36664_;
  assign new_n36666_ = ys__n208 & ~new_n36665_;
  assign new_n36667_ = ~ys__n208 & new_n36665_;
  assign new_n36668_ = ~new_n36666_ & ~new_n36667_;
  assign new_n36669_ = new_n36479_ & ~new_n36668_;
  assign new_n36670_ = ys__n192 & new_n12122_;
  assign new_n36671_ = new_n36663_ & ~new_n36670_;
  assign new_n36672_ = ys__n208 & ~new_n36671_;
  assign new_n36673_ = ~ys__n208 & new_n36671_;
  assign new_n36674_ = ~new_n36672_ & ~new_n36673_;
  assign new_n36675_ = new_n36477_ & ~new_n36674_;
  assign new_n36676_ = ~ys__n204 & ys__n860;
  assign new_n36677_ = ~new_n36638_ & ~new_n36676_;
  assign new_n36678_ = ys__n208 & ~new_n36677_;
  assign new_n36679_ = ~ys__n208 & new_n36677_;
  assign new_n36680_ = ~new_n36678_ & ~new_n36679_;
  assign new_n36681_ = new_n36467_ & ~new_n36680_;
  assign new_n36682_ = ys__n208 & ~new_n36663_;
  assign new_n36683_ = ~ys__n208 & new_n36663_;
  assign new_n36684_ = ~new_n36682_ & ~new_n36683_;
  assign new_n36685_ = new_n36457_ & ~new_n36684_;
  assign new_n36686_ = ~new_n36681_ & ~new_n36685_;
  assign new_n36687_ = ~new_n36675_ & new_n36686_;
  assign new_n36688_ = ~new_n36669_ & new_n36687_;
  assign new_n36689_ = new_n36644_ & ~new_n36688_;
  assign new_n36690_ = new_n36489_ & new_n36689_;
  assign new_n36691_ = new_n36491_ & new_n36689_;
  assign new_n36692_ = new_n36516_ & new_n36649_;
  assign new_n36693_ = new_n36525_ & new_n36692_;
  assign new_n36694_ = new_n36648_ & new_n36693_;
  assign new_n36695_ = new_n12139_ & ~new_n36694_;
  assign new_n36696_ = ~new_n36551_ & new_n36695_;
  assign new_n36697_ = ~new_n36691_ & ~new_n36696_;
  assign new_n36698_ = new_n36561_ & ~new_n36697_;
  assign new_n36699_ = ~new_n36690_ & ~new_n36698_;
  assign new_n36700_ = ~ys__n738 & ~new_n36699_;
  assign new_n36701_ = new_n36565_ & new_n36689_;
  assign ys__n28785 = new_n36700_ | new_n36701_;
  assign new_n36703_ = ~ys__n208 & ~new_n36665_;
  assign new_n36704_ = ~ys__n208 & ~new_n36703_;
  assign new_n36705_ = ys__n206 & ~new_n36704_;
  assign new_n36706_ = ~ys__n206 & new_n36704_;
  assign new_n36707_ = ~new_n36705_ & ~new_n36706_;
  assign new_n36708_ = new_n36479_ & ~new_n36707_;
  assign new_n36709_ = ~ys__n208 & ~new_n36671_;
  assign new_n36710_ = ~ys__n208 & ~new_n36709_;
  assign new_n36711_ = ys__n206 & ~new_n36710_;
  assign new_n36712_ = ~ys__n206 & new_n36710_;
  assign new_n36713_ = ~new_n36711_ & ~new_n36712_;
  assign new_n36714_ = new_n36477_ & ~new_n36713_;
  assign new_n36715_ = ~ys__n208 & ~new_n36677_;
  assign new_n36716_ = ~ys__n208 & ~new_n36715_;
  assign new_n36717_ = ys__n206 & ~new_n36716_;
  assign new_n36718_ = ~ys__n206 & new_n36716_;
  assign new_n36719_ = ~new_n36717_ & ~new_n36718_;
  assign new_n36720_ = new_n36467_ & ~new_n36719_;
  assign new_n36721_ = ~ys__n208 & ~new_n36663_;
  assign new_n36722_ = ~ys__n208 & ~new_n36721_;
  assign new_n36723_ = ys__n206 & ~new_n36722_;
  assign new_n36724_ = ~ys__n206 & new_n36722_;
  assign new_n36725_ = ~new_n36723_ & ~new_n36724_;
  assign new_n36726_ = new_n36457_ & ~new_n36725_;
  assign new_n36727_ = ~new_n36720_ & ~new_n36726_;
  assign new_n36728_ = ~new_n36714_ & new_n36727_;
  assign new_n36729_ = ~new_n36708_ & new_n36728_;
  assign new_n36730_ = new_n36644_ & ~new_n36729_;
  assign new_n36731_ = new_n36489_ & new_n36730_;
  assign new_n36732_ = new_n36491_ & new_n36730_;
  assign new_n36733_ = ~new_n36495_ & ~new_n36501_;
  assign new_n36734_ = ~new_n36532_ & new_n36733_;
  assign new_n36735_ = new_n36511_ & new_n36541_;
  assign new_n36736_ = new_n36734_ & new_n36735_;
  assign new_n36737_ = new_n36548_ & new_n36736_;
  assign new_n36738_ = new_n12139_ & ~new_n36737_;
  assign new_n36739_ = ~new_n36551_ & new_n36738_;
  assign new_n36740_ = ~new_n36732_ & ~new_n36739_;
  assign new_n36741_ = new_n36561_ & ~new_n36740_;
  assign new_n36742_ = ~new_n36731_ & ~new_n36741_;
  assign new_n36743_ = ~ys__n738 & ~new_n36742_;
  assign new_n36744_ = new_n36565_ & new_n36730_;
  assign ys__n28786 = new_n36743_ | new_n36744_;
  assign new_n36746_ = ys__n47185 & ~new_n13716_;
  assign new_n36747_ = ys__n46962 & new_n36467_;
  assign new_n36748_ = ys__n46958 & new_n36457_;
  assign new_n36749_ = ~new_n36747_ & ~new_n36748_;
  assign new_n36750_ = ys__n46956 & new_n36477_;
  assign new_n36751_ = ys__n47184 & new_n36479_;
  assign new_n36752_ = ~new_n36750_ & ~new_n36751_;
  assign new_n36753_ = new_n36749_ & new_n36752_;
  assign new_n36754_ = ~new_n36485_ & ~new_n36753_;
  assign new_n36755_ = new_n13716_ & new_n36754_;
  assign new_n36756_ = ~new_n36746_ & ~new_n36755_;
  assign new_n36757_ = ys__n4566 & ~new_n36756_;
  assign new_n36758_ = new_n12127_ & ~new_n12138_;
  assign new_n36759_ = ys__n202 & new_n36758_;
  assign new_n36760_ = ys__n23339 & new_n36759_;
  assign new_n36761_ = ~ys__n202 & new_n36758_;
  assign new_n36762_ = ys__n22464 & new_n36761_;
  assign new_n36763_ = ~new_n36760_ & ~new_n36762_;
  assign new_n36764_ = ys__n202 & ~new_n36758_;
  assign new_n36765_ = ys__n28243 & new_n36764_;
  assign new_n36766_ = ~ys__n202 & ~new_n36758_;
  assign new_n36767_ = ys__n47106 & new_n36766_;
  assign new_n36768_ = ~new_n36765_ & ~new_n36767_;
  assign new_n36769_ = new_n36763_ & new_n36768_;
  assign new_n36770_ = ~new_n36759_ & ~new_n36761_;
  assign new_n36771_ = ~new_n36764_ & ~new_n36766_;
  assign new_n36772_ = new_n36770_ & new_n36771_;
  assign new_n36773_ = new_n12139_ & ~new_n36772_;
  assign new_n36774_ = ~new_n36769_ & new_n36773_;
  assign new_n36775_ = ys__n47185 & new_n13714_;
  assign new_n36776_ = new_n36491_ & new_n36754_;
  assign new_n36777_ = ~new_n36775_ & ~new_n36776_;
  assign new_n36778_ = ~new_n36774_ & new_n36777_;
  assign new_n36779_ = ~new_n13714_ & new_n36560_;
  assign new_n36780_ = ~ys__n4566 & ~new_n36779_;
  assign new_n36781_ = ~new_n36778_ & new_n36780_;
  assign new_n36782_ = ~new_n36757_ & ~new_n36781_;
  assign new_n36783_ = ~ys__n738 & ~new_n36782_;
  assign new_n36784_ = ys__n47185 & ~new_n13713_;
  assign new_n36785_ = new_n13713_ & new_n36754_;
  assign new_n36786_ = ~new_n36784_ & ~new_n36785_;
  assign new_n36787_ = ys__n738 & ~new_n36786_;
  assign ys__n28787 = new_n36783_ | new_n36787_;
  assign new_n36789_ = ys__n47184 & ~new_n13716_;
  assign new_n36790_ = ys__n46963 & new_n36467_;
  assign new_n36791_ = ys__n46959 & new_n36457_;
  assign new_n36792_ = ~new_n36790_ & ~new_n36791_;
  assign new_n36793_ = ys__n46957 & new_n36477_;
  assign new_n36794_ = ys__n46956 & new_n36479_;
  assign new_n36795_ = ~new_n36793_ & ~new_n36794_;
  assign new_n36796_ = new_n36792_ & new_n36795_;
  assign new_n36797_ = ~new_n36485_ & ~new_n36796_;
  assign new_n36798_ = new_n13716_ & new_n36797_;
  assign new_n36799_ = ~new_n36789_ & ~new_n36798_;
  assign new_n36800_ = ys__n4566 & ~new_n36799_;
  assign new_n36801_ = ys__n22464 & new_n36759_;
  assign new_n36802_ = ys__n23548 & new_n36761_;
  assign new_n36803_ = ~new_n36801_ & ~new_n36802_;
  assign new_n36804_ = ys__n47106 & new_n36764_;
  assign new_n36805_ = ys__n23111 & new_n36766_;
  assign new_n36806_ = ~new_n36804_ & ~new_n36805_;
  assign new_n36807_ = new_n36803_ & new_n36806_;
  assign new_n36808_ = new_n36773_ & ~new_n36807_;
  assign new_n36809_ = ys__n47184 & new_n13714_;
  assign new_n36810_ = new_n36491_ & new_n36797_;
  assign new_n36811_ = ~new_n36809_ & ~new_n36810_;
  assign new_n36812_ = ~new_n36808_ & new_n36811_;
  assign new_n36813_ = new_n36780_ & ~new_n36812_;
  assign new_n36814_ = ~new_n36800_ & ~new_n36813_;
  assign new_n36815_ = ~ys__n738 & ~new_n36814_;
  assign new_n36816_ = ys__n47184 & ~new_n13713_;
  assign new_n36817_ = new_n13713_ & new_n36797_;
  assign new_n36818_ = ~new_n36816_ & ~new_n36817_;
  assign new_n36819_ = ys__n738 & ~new_n36818_;
  assign ys__n28788 = new_n36815_ | new_n36819_;
  assign new_n36821_ = ys__n46956 & ~new_n13716_;
  assign new_n36822_ = ys__n46964 & new_n36467_;
  assign new_n36823_ = ys__n46960 & new_n36457_;
  assign new_n36824_ = ~new_n36822_ & ~new_n36823_;
  assign new_n36825_ = ys__n46958 & new_n36477_;
  assign new_n36826_ = ys__n46957 & new_n36479_;
  assign new_n36827_ = ~new_n36825_ & ~new_n36826_;
  assign new_n36828_ = new_n36824_ & new_n36827_;
  assign new_n36829_ = ~new_n36485_ & ~new_n36828_;
  assign new_n36830_ = new_n13716_ & new_n36829_;
  assign new_n36831_ = ~new_n36821_ & ~new_n36830_;
  assign new_n36832_ = ys__n4566 & ~new_n36831_;
  assign new_n36833_ = ys__n23548 & new_n36759_;
  assign new_n36834_ = ys__n23550 & new_n36761_;
  assign new_n36835_ = ~new_n36833_ & ~new_n36834_;
  assign new_n36836_ = ys__n23111 & new_n36764_;
  assign new_n36837_ = ys__n23114 & new_n36766_;
  assign new_n36838_ = ~new_n36836_ & ~new_n36837_;
  assign new_n36839_ = new_n36835_ & new_n36838_;
  assign new_n36840_ = new_n36773_ & ~new_n36839_;
  assign new_n36841_ = ys__n46956 & new_n13714_;
  assign new_n36842_ = new_n36491_ & new_n36829_;
  assign new_n36843_ = ~new_n36841_ & ~new_n36842_;
  assign new_n36844_ = ~new_n36840_ & new_n36843_;
  assign new_n36845_ = new_n36780_ & ~new_n36844_;
  assign new_n36846_ = ~new_n36832_ & ~new_n36845_;
  assign new_n36847_ = ~ys__n738 & ~new_n36846_;
  assign new_n36848_ = ys__n46956 & ~new_n13713_;
  assign new_n36849_ = new_n13713_ & new_n36829_;
  assign new_n36850_ = ~new_n36848_ & ~new_n36849_;
  assign new_n36851_ = ys__n738 & ~new_n36850_;
  assign ys__n28789 = new_n36847_ | new_n36851_;
  assign new_n36853_ = ys__n46957 & ~new_n13716_;
  assign new_n36854_ = ys__n46965 & new_n36467_;
  assign new_n36855_ = ys__n46961 & new_n36457_;
  assign new_n36856_ = ~new_n36854_ & ~new_n36855_;
  assign new_n36857_ = ys__n46959 & new_n36477_;
  assign new_n36858_ = ys__n46958 & new_n36479_;
  assign new_n36859_ = ~new_n36857_ & ~new_n36858_;
  assign new_n36860_ = new_n36856_ & new_n36859_;
  assign new_n36861_ = ~new_n36485_ & ~new_n36860_;
  assign new_n36862_ = new_n13716_ & new_n36861_;
  assign new_n36863_ = ~new_n36853_ & ~new_n36862_;
  assign new_n36864_ = ys__n4566 & ~new_n36863_;
  assign new_n36865_ = ys__n23550 & new_n36759_;
  assign new_n36866_ = ys__n23552 & new_n36761_;
  assign new_n36867_ = ~new_n36865_ & ~new_n36866_;
  assign new_n36868_ = ys__n23114 & new_n36764_;
  assign new_n36869_ = ys__n23117 & new_n36766_;
  assign new_n36870_ = ~new_n36868_ & ~new_n36869_;
  assign new_n36871_ = new_n36867_ & new_n36870_;
  assign new_n36872_ = new_n36773_ & ~new_n36871_;
  assign new_n36873_ = ys__n46957 & new_n13714_;
  assign new_n36874_ = new_n36491_ & new_n36861_;
  assign new_n36875_ = ~new_n36873_ & ~new_n36874_;
  assign new_n36876_ = ~new_n36872_ & new_n36875_;
  assign new_n36877_ = new_n36780_ & ~new_n36876_;
  assign new_n36878_ = ~new_n36864_ & ~new_n36877_;
  assign new_n36879_ = ~ys__n738 & ~new_n36878_;
  assign new_n36880_ = ys__n46957 & ~new_n13713_;
  assign new_n36881_ = new_n13713_ & new_n36861_;
  assign new_n36882_ = ~new_n36880_ & ~new_n36881_;
  assign new_n36883_ = ys__n738 & ~new_n36882_;
  assign ys__n28790 = new_n36879_ | new_n36883_;
  assign new_n36885_ = ys__n46958 & ~new_n13716_;
  assign new_n36886_ = ys__n46966 & new_n36467_;
  assign new_n36887_ = ys__n46962 & new_n36457_;
  assign new_n36888_ = ~new_n36886_ & ~new_n36887_;
  assign new_n36889_ = ys__n46960 & new_n36477_;
  assign new_n36890_ = ys__n46959 & new_n36479_;
  assign new_n36891_ = ~new_n36889_ & ~new_n36890_;
  assign new_n36892_ = new_n36888_ & new_n36891_;
  assign new_n36893_ = ~new_n36485_ & ~new_n36892_;
  assign new_n36894_ = new_n13716_ & new_n36893_;
  assign new_n36895_ = ~new_n36885_ & ~new_n36894_;
  assign new_n36896_ = ys__n4566 & ~new_n36895_;
  assign new_n36897_ = ys__n23552 & new_n36759_;
  assign new_n36898_ = ys__n23554 & new_n36761_;
  assign new_n36899_ = ~new_n36897_ & ~new_n36898_;
  assign new_n36900_ = ys__n23117 & new_n36764_;
  assign new_n36901_ = ys__n23120 & new_n36766_;
  assign new_n36902_ = ~new_n36900_ & ~new_n36901_;
  assign new_n36903_ = new_n36899_ & new_n36902_;
  assign new_n36904_ = new_n36773_ & ~new_n36903_;
  assign new_n36905_ = ys__n46958 & new_n13714_;
  assign new_n36906_ = new_n36491_ & new_n36893_;
  assign new_n36907_ = ~new_n36905_ & ~new_n36906_;
  assign new_n36908_ = ~new_n36904_ & new_n36907_;
  assign new_n36909_ = new_n36780_ & ~new_n36908_;
  assign new_n36910_ = ~new_n36896_ & ~new_n36909_;
  assign new_n36911_ = ~ys__n738 & ~new_n36910_;
  assign new_n36912_ = ys__n46958 & ~new_n13713_;
  assign new_n36913_ = new_n13713_ & new_n36893_;
  assign new_n36914_ = ~new_n36912_ & ~new_n36913_;
  assign new_n36915_ = ys__n738 & ~new_n36914_;
  assign ys__n28791 = new_n36911_ | new_n36915_;
  assign new_n36917_ = ys__n46959 & ~new_n13716_;
  assign new_n36918_ = ys__n46967 & new_n36467_;
  assign new_n36919_ = ys__n46963 & new_n36457_;
  assign new_n36920_ = ~new_n36918_ & ~new_n36919_;
  assign new_n36921_ = ys__n46961 & new_n36477_;
  assign new_n36922_ = ys__n46960 & new_n36479_;
  assign new_n36923_ = ~new_n36921_ & ~new_n36922_;
  assign new_n36924_ = new_n36920_ & new_n36923_;
  assign new_n36925_ = ~new_n36485_ & ~new_n36924_;
  assign new_n36926_ = new_n13716_ & new_n36925_;
  assign new_n36927_ = ~new_n36917_ & ~new_n36926_;
  assign new_n36928_ = ys__n4566 & ~new_n36927_;
  assign new_n36929_ = ys__n23554 & new_n36759_;
  assign new_n36930_ = ys__n23556 & new_n36761_;
  assign new_n36931_ = ~new_n36929_ & ~new_n36930_;
  assign new_n36932_ = ys__n23120 & new_n36764_;
  assign new_n36933_ = ys__n23123 & new_n36766_;
  assign new_n36934_ = ~new_n36932_ & ~new_n36933_;
  assign new_n36935_ = new_n36931_ & new_n36934_;
  assign new_n36936_ = new_n36773_ & ~new_n36935_;
  assign new_n36937_ = ys__n46959 & new_n13714_;
  assign new_n36938_ = new_n36491_ & new_n36925_;
  assign new_n36939_ = ~new_n36937_ & ~new_n36938_;
  assign new_n36940_ = ~new_n36936_ & new_n36939_;
  assign new_n36941_ = new_n36780_ & ~new_n36940_;
  assign new_n36942_ = ~new_n36928_ & ~new_n36941_;
  assign new_n36943_ = ~ys__n738 & ~new_n36942_;
  assign new_n36944_ = ys__n46959 & ~new_n13713_;
  assign new_n36945_ = new_n13713_ & new_n36925_;
  assign new_n36946_ = ~new_n36944_ & ~new_n36945_;
  assign new_n36947_ = ys__n738 & ~new_n36946_;
  assign ys__n28792 = new_n36943_ | new_n36947_;
  assign new_n36949_ = ys__n46960 & ~new_n13716_;
  assign new_n36950_ = ys__n46968 & new_n36467_;
  assign new_n36951_ = ys__n46964 & new_n36457_;
  assign new_n36952_ = ~new_n36950_ & ~new_n36951_;
  assign new_n36953_ = ys__n46962 & new_n36477_;
  assign new_n36954_ = ys__n46961 & new_n36479_;
  assign new_n36955_ = ~new_n36953_ & ~new_n36954_;
  assign new_n36956_ = new_n36952_ & new_n36955_;
  assign new_n36957_ = ~new_n36485_ & ~new_n36956_;
  assign new_n36958_ = new_n13716_ & new_n36957_;
  assign new_n36959_ = ~new_n36949_ & ~new_n36958_;
  assign new_n36960_ = ys__n4566 & ~new_n36959_;
  assign new_n36961_ = ys__n23556 & new_n36759_;
  assign new_n36962_ = ys__n23558 & new_n36761_;
  assign new_n36963_ = ~new_n36961_ & ~new_n36962_;
  assign new_n36964_ = ys__n23123 & new_n36764_;
  assign new_n36965_ = ys__n23126 & new_n36766_;
  assign new_n36966_ = ~new_n36964_ & ~new_n36965_;
  assign new_n36967_ = new_n36963_ & new_n36966_;
  assign new_n36968_ = new_n36773_ & ~new_n36967_;
  assign new_n36969_ = ys__n46960 & new_n13714_;
  assign new_n36970_ = new_n36491_ & new_n36957_;
  assign new_n36971_ = ~new_n36969_ & ~new_n36970_;
  assign new_n36972_ = ~new_n36968_ & new_n36971_;
  assign new_n36973_ = new_n36780_ & ~new_n36972_;
  assign new_n36974_ = ~new_n36960_ & ~new_n36973_;
  assign new_n36975_ = ~ys__n738 & ~new_n36974_;
  assign new_n36976_ = ys__n46960 & ~new_n13713_;
  assign new_n36977_ = new_n13713_ & new_n36957_;
  assign new_n36978_ = ~new_n36976_ & ~new_n36977_;
  assign new_n36979_ = ys__n738 & ~new_n36978_;
  assign ys__n28793 = new_n36975_ | new_n36979_;
  assign new_n36981_ = ys__n46961 & ~new_n13716_;
  assign new_n36982_ = ys__n46969 & new_n36467_;
  assign new_n36983_ = ys__n46965 & new_n36457_;
  assign new_n36984_ = ~new_n36982_ & ~new_n36983_;
  assign new_n36985_ = ys__n46963 & new_n36477_;
  assign new_n36986_ = ys__n46962 & new_n36479_;
  assign new_n36987_ = ~new_n36985_ & ~new_n36986_;
  assign new_n36988_ = new_n36984_ & new_n36987_;
  assign new_n36989_ = ~new_n36485_ & ~new_n36988_;
  assign new_n36990_ = new_n13716_ & new_n36989_;
  assign new_n36991_ = ~new_n36981_ & ~new_n36990_;
  assign new_n36992_ = ys__n4566 & ~new_n36991_;
  assign new_n36993_ = ys__n23558 & new_n36759_;
  assign new_n36994_ = ys__n23560 & new_n36761_;
  assign new_n36995_ = ~new_n36993_ & ~new_n36994_;
  assign new_n36996_ = ys__n23126 & new_n36764_;
  assign new_n36997_ = ys__n23129 & new_n36766_;
  assign new_n36998_ = ~new_n36996_ & ~new_n36997_;
  assign new_n36999_ = new_n36995_ & new_n36998_;
  assign new_n37000_ = new_n36773_ & ~new_n36999_;
  assign new_n37001_ = ys__n46961 & new_n13714_;
  assign new_n37002_ = new_n36491_ & new_n36989_;
  assign new_n37003_ = ~new_n37001_ & ~new_n37002_;
  assign new_n37004_ = ~new_n37000_ & new_n37003_;
  assign new_n37005_ = new_n36780_ & ~new_n37004_;
  assign new_n37006_ = ~new_n36992_ & ~new_n37005_;
  assign new_n37007_ = ~ys__n738 & ~new_n37006_;
  assign new_n37008_ = ys__n46961 & ~new_n13713_;
  assign new_n37009_ = new_n13713_ & new_n36989_;
  assign new_n37010_ = ~new_n37008_ & ~new_n37009_;
  assign new_n37011_ = ys__n738 & ~new_n37010_;
  assign ys__n28794 = new_n37007_ | new_n37011_;
  assign new_n37013_ = ys__n46970 & new_n36467_;
  assign new_n37014_ = ys__n46966 & new_n36457_;
  assign new_n37015_ = ~new_n37013_ & ~new_n37014_;
  assign new_n37016_ = ys__n46964 & new_n36477_;
  assign new_n37017_ = ys__n46963 & new_n36479_;
  assign new_n37018_ = ~new_n37016_ & ~new_n37017_;
  assign new_n37019_ = new_n37015_ & new_n37018_;
  assign new_n37020_ = ~new_n36485_ & ~new_n37019_;
  assign new_n37021_ = new_n36489_ & new_n37020_;
  assign new_n37022_ = new_n36491_ & new_n37020_;
  assign new_n37023_ = ys__n23560 & new_n36759_;
  assign new_n37024_ = ys__n23562 & new_n36761_;
  assign new_n37025_ = ~new_n37023_ & ~new_n37024_;
  assign new_n37026_ = ys__n23129 & new_n36764_;
  assign new_n37027_ = ys__n23132 & new_n36766_;
  assign new_n37028_ = ~new_n37026_ & ~new_n37027_;
  assign new_n37029_ = new_n37025_ & new_n37028_;
  assign new_n37030_ = new_n36773_ & ~new_n37029_;
  assign new_n37031_ = ~new_n37022_ & ~new_n37030_;
  assign new_n37032_ = new_n36780_ & ~new_n37031_;
  assign new_n37033_ = ~new_n37021_ & ~new_n37032_;
  assign new_n37034_ = ~ys__n738 & ~new_n37033_;
  assign new_n37035_ = new_n36565_ & new_n37020_;
  assign ys__n28796 = new_n37034_ | new_n37035_;
  assign new_n37037_ = ys__n46971 & new_n36467_;
  assign new_n37038_ = ys__n46967 & new_n36457_;
  assign new_n37039_ = ~new_n37037_ & ~new_n37038_;
  assign new_n37040_ = ys__n46965 & new_n36477_;
  assign new_n37041_ = ys__n46964 & new_n36479_;
  assign new_n37042_ = ~new_n37040_ & ~new_n37041_;
  assign new_n37043_ = new_n37039_ & new_n37042_;
  assign new_n37044_ = ~new_n36485_ & ~new_n37043_;
  assign new_n37045_ = new_n36489_ & new_n37044_;
  assign new_n37046_ = new_n36491_ & new_n37044_;
  assign new_n37047_ = ys__n23562 & new_n36759_;
  assign new_n37048_ = ys__n23564 & new_n36761_;
  assign new_n37049_ = ~new_n37047_ & ~new_n37048_;
  assign new_n37050_ = ys__n23132 & new_n36764_;
  assign new_n37051_ = ys__n23135 & new_n36766_;
  assign new_n37052_ = ~new_n37050_ & ~new_n37051_;
  assign new_n37053_ = new_n37049_ & new_n37052_;
  assign new_n37054_ = new_n36773_ & ~new_n37053_;
  assign new_n37055_ = ~new_n37046_ & ~new_n37054_;
  assign new_n37056_ = new_n36780_ & ~new_n37055_;
  assign new_n37057_ = ~new_n37045_ & ~new_n37056_;
  assign new_n37058_ = ~ys__n738 & ~new_n37057_;
  assign new_n37059_ = new_n36565_ & new_n37044_;
  assign ys__n28798 = new_n37058_ | new_n37059_;
  assign new_n37061_ = ys__n46972 & new_n36467_;
  assign new_n37062_ = ys__n46968 & new_n36457_;
  assign new_n37063_ = ~new_n37061_ & ~new_n37062_;
  assign new_n37064_ = ys__n46966 & new_n36477_;
  assign new_n37065_ = ys__n46965 & new_n36479_;
  assign new_n37066_ = ~new_n37064_ & ~new_n37065_;
  assign new_n37067_ = new_n37063_ & new_n37066_;
  assign new_n37068_ = ~new_n36485_ & ~new_n37067_;
  assign new_n37069_ = new_n36489_ & new_n37068_;
  assign new_n37070_ = new_n36491_ & new_n37068_;
  assign new_n37071_ = ys__n23564 & new_n36759_;
  assign new_n37072_ = ys__n23566 & new_n36761_;
  assign new_n37073_ = ~new_n37071_ & ~new_n37072_;
  assign new_n37074_ = ys__n23135 & new_n36764_;
  assign new_n37075_ = ys__n23138 & new_n36766_;
  assign new_n37076_ = ~new_n37074_ & ~new_n37075_;
  assign new_n37077_ = new_n37073_ & new_n37076_;
  assign new_n37078_ = new_n36773_ & ~new_n37077_;
  assign new_n37079_ = ~new_n37070_ & ~new_n37078_;
  assign new_n37080_ = new_n36780_ & ~new_n37079_;
  assign new_n37081_ = ~new_n37069_ & ~new_n37080_;
  assign new_n37082_ = ~ys__n738 & ~new_n37081_;
  assign new_n37083_ = new_n36565_ & new_n37068_;
  assign ys__n28800 = new_n37082_ | new_n37083_;
  assign new_n37085_ = ys__n46973 & new_n36467_;
  assign new_n37086_ = ys__n46969 & new_n36457_;
  assign new_n37087_ = ~new_n37085_ & ~new_n37086_;
  assign new_n37088_ = ys__n46967 & new_n36477_;
  assign new_n37089_ = ys__n46966 & new_n36479_;
  assign new_n37090_ = ~new_n37088_ & ~new_n37089_;
  assign new_n37091_ = new_n37087_ & new_n37090_;
  assign new_n37092_ = ~new_n36485_ & ~new_n37091_;
  assign new_n37093_ = new_n36489_ & new_n37092_;
  assign new_n37094_ = new_n36491_ & new_n37092_;
  assign new_n37095_ = ys__n23566 & new_n36759_;
  assign new_n37096_ = ys__n23568 & new_n36761_;
  assign new_n37097_ = ~new_n37095_ & ~new_n37096_;
  assign new_n37098_ = ys__n23138 & new_n36764_;
  assign new_n37099_ = ys__n23141 & new_n36766_;
  assign new_n37100_ = ~new_n37098_ & ~new_n37099_;
  assign new_n37101_ = new_n37097_ & new_n37100_;
  assign new_n37102_ = new_n36773_ & ~new_n37101_;
  assign new_n37103_ = ~new_n37094_ & ~new_n37102_;
  assign new_n37104_ = new_n36780_ & ~new_n37103_;
  assign new_n37105_ = ~new_n37093_ & ~new_n37104_;
  assign new_n37106_ = ~ys__n738 & ~new_n37105_;
  assign new_n37107_ = new_n36565_ & new_n37092_;
  assign ys__n28802 = new_n37106_ | new_n37107_;
  assign new_n37109_ = ys__n46974 & new_n36467_;
  assign new_n37110_ = ys__n46970 & new_n36457_;
  assign new_n37111_ = ~new_n37109_ & ~new_n37110_;
  assign new_n37112_ = ys__n46968 & new_n36477_;
  assign new_n37113_ = ys__n46967 & new_n36479_;
  assign new_n37114_ = ~new_n37112_ & ~new_n37113_;
  assign new_n37115_ = new_n37111_ & new_n37114_;
  assign new_n37116_ = ~new_n36485_ & ~new_n37115_;
  assign new_n37117_ = new_n36489_ & new_n37116_;
  assign new_n37118_ = new_n36491_ & new_n37116_;
  assign new_n37119_ = ys__n23568 & new_n36759_;
  assign new_n37120_ = ys__n23570 & new_n36761_;
  assign new_n37121_ = ~new_n37119_ & ~new_n37120_;
  assign new_n37122_ = ys__n23141 & new_n36764_;
  assign new_n37123_ = ys__n23144 & new_n36766_;
  assign new_n37124_ = ~new_n37122_ & ~new_n37123_;
  assign new_n37125_ = new_n37121_ & new_n37124_;
  assign new_n37126_ = new_n36773_ & ~new_n37125_;
  assign new_n37127_ = ~new_n37118_ & ~new_n37126_;
  assign new_n37128_ = new_n36780_ & ~new_n37127_;
  assign new_n37129_ = ~new_n37117_ & ~new_n37128_;
  assign new_n37130_ = ~ys__n738 & ~new_n37129_;
  assign new_n37131_ = new_n36565_ & new_n37116_;
  assign ys__n28804 = new_n37130_ | new_n37131_;
  assign new_n37133_ = ys__n46975 & new_n36467_;
  assign new_n37134_ = ys__n46971 & new_n36457_;
  assign new_n37135_ = ~new_n37133_ & ~new_n37134_;
  assign new_n37136_ = ys__n46969 & new_n36477_;
  assign new_n37137_ = ys__n46968 & new_n36479_;
  assign new_n37138_ = ~new_n37136_ & ~new_n37137_;
  assign new_n37139_ = new_n37135_ & new_n37138_;
  assign new_n37140_ = ~new_n36485_ & ~new_n37139_;
  assign new_n37141_ = new_n36489_ & new_n37140_;
  assign new_n37142_ = new_n36491_ & new_n37140_;
  assign new_n37143_ = ys__n23570 & new_n36759_;
  assign new_n37144_ = ys__n23572 & new_n36761_;
  assign new_n37145_ = ~new_n37143_ & ~new_n37144_;
  assign new_n37146_ = ys__n23144 & new_n36764_;
  assign new_n37147_ = ys__n23147 & new_n36766_;
  assign new_n37148_ = ~new_n37146_ & ~new_n37147_;
  assign new_n37149_ = new_n37145_ & new_n37148_;
  assign new_n37150_ = new_n36773_ & ~new_n37149_;
  assign new_n37151_ = ~new_n37142_ & ~new_n37150_;
  assign new_n37152_ = new_n36780_ & ~new_n37151_;
  assign new_n37153_ = ~new_n37141_ & ~new_n37152_;
  assign new_n37154_ = ~ys__n738 & ~new_n37153_;
  assign new_n37155_ = new_n36565_ & new_n37140_;
  assign ys__n28806 = new_n37154_ | new_n37155_;
  assign new_n37157_ = ys__n46976 & new_n36467_;
  assign new_n37158_ = ys__n46972 & new_n36457_;
  assign new_n37159_ = ~new_n37157_ & ~new_n37158_;
  assign new_n37160_ = ys__n46970 & new_n36477_;
  assign new_n37161_ = ys__n46969 & new_n36479_;
  assign new_n37162_ = ~new_n37160_ & ~new_n37161_;
  assign new_n37163_ = new_n37159_ & new_n37162_;
  assign new_n37164_ = ~new_n36485_ & ~new_n37163_;
  assign new_n37165_ = new_n36489_ & new_n37164_;
  assign new_n37166_ = new_n36491_ & new_n37164_;
  assign new_n37167_ = ys__n23572 & new_n36759_;
  assign new_n37168_ = ys__n23574 & new_n36761_;
  assign new_n37169_ = ~new_n37167_ & ~new_n37168_;
  assign new_n37170_ = ys__n23147 & new_n36764_;
  assign new_n37171_ = ys__n23150 & new_n36766_;
  assign new_n37172_ = ~new_n37170_ & ~new_n37171_;
  assign new_n37173_ = new_n37169_ & new_n37172_;
  assign new_n37174_ = new_n36773_ & ~new_n37173_;
  assign new_n37175_ = ~new_n37166_ & ~new_n37174_;
  assign new_n37176_ = new_n36780_ & ~new_n37175_;
  assign new_n37177_ = ~new_n37165_ & ~new_n37176_;
  assign new_n37178_ = ~ys__n738 & ~new_n37177_;
  assign new_n37179_ = new_n36565_ & new_n37164_;
  assign ys__n28808 = new_n37178_ | new_n37179_;
  assign new_n37181_ = ys__n46977 & new_n36467_;
  assign new_n37182_ = ys__n46973 & new_n36457_;
  assign new_n37183_ = ~new_n37181_ & ~new_n37182_;
  assign new_n37184_ = ys__n46971 & new_n36477_;
  assign new_n37185_ = ys__n46970 & new_n36479_;
  assign new_n37186_ = ~new_n37184_ & ~new_n37185_;
  assign new_n37187_ = new_n37183_ & new_n37186_;
  assign new_n37188_ = ~new_n36485_ & ~new_n37187_;
  assign new_n37189_ = new_n36489_ & new_n37188_;
  assign new_n37190_ = new_n36491_ & new_n37188_;
  assign new_n37191_ = ys__n23574 & new_n36759_;
  assign new_n37192_ = ys__n420 & new_n36761_;
  assign new_n37193_ = ~new_n37191_ & ~new_n37192_;
  assign new_n37194_ = ys__n23150 & new_n36764_;
  assign new_n37195_ = ys__n23153 & new_n36766_;
  assign new_n37196_ = ~new_n37194_ & ~new_n37195_;
  assign new_n37197_ = new_n37193_ & new_n37196_;
  assign new_n37198_ = new_n36773_ & ~new_n37197_;
  assign new_n37199_ = ~new_n37190_ & ~new_n37198_;
  assign new_n37200_ = new_n36780_ & ~new_n37199_;
  assign new_n37201_ = ~new_n37189_ & ~new_n37200_;
  assign new_n37202_ = ~ys__n738 & ~new_n37201_;
  assign new_n37203_ = new_n36565_ & new_n37188_;
  assign ys__n28810 = new_n37202_ | new_n37203_;
  assign new_n37205_ = ys__n46978 & new_n36467_;
  assign new_n37206_ = ys__n46974 & new_n36457_;
  assign new_n37207_ = ~new_n37205_ & ~new_n37206_;
  assign new_n37208_ = ys__n46972 & new_n36477_;
  assign new_n37209_ = ys__n46971 & new_n36479_;
  assign new_n37210_ = ~new_n37208_ & ~new_n37209_;
  assign new_n37211_ = new_n37207_ & new_n37210_;
  assign new_n37212_ = ~new_n36485_ & ~new_n37211_;
  assign new_n37213_ = new_n36489_ & new_n37212_;
  assign new_n37214_ = new_n36491_ & new_n37212_;
  assign new_n37215_ = ys__n420 & new_n36759_;
  assign new_n37216_ = ys__n442 & new_n36761_;
  assign new_n37217_ = ~new_n37215_ & ~new_n37216_;
  assign new_n37218_ = ys__n23153 & new_n36764_;
  assign new_n37219_ = ys__n23156 & new_n36766_;
  assign new_n37220_ = ~new_n37218_ & ~new_n37219_;
  assign new_n37221_ = new_n37217_ & new_n37220_;
  assign new_n37222_ = new_n36773_ & ~new_n37221_;
  assign new_n37223_ = ~new_n37214_ & ~new_n37222_;
  assign new_n37224_ = new_n36780_ & ~new_n37223_;
  assign new_n37225_ = ~new_n37213_ & ~new_n37224_;
  assign new_n37226_ = ~ys__n738 & ~new_n37225_;
  assign new_n37227_ = new_n36565_ & new_n37212_;
  assign ys__n28812 = new_n37226_ | new_n37227_;
  assign new_n37229_ = ys__n46979 & new_n36467_;
  assign new_n37230_ = ys__n46975 & new_n36457_;
  assign new_n37231_ = ~new_n37229_ & ~new_n37230_;
  assign new_n37232_ = ys__n46973 & new_n36477_;
  assign new_n37233_ = ys__n46972 & new_n36479_;
  assign new_n37234_ = ~new_n37232_ & ~new_n37233_;
  assign new_n37235_ = new_n37231_ & new_n37234_;
  assign new_n37236_ = ~new_n36485_ & ~new_n37235_;
  assign new_n37237_ = new_n36489_ & new_n37236_;
  assign new_n37238_ = new_n36491_ & new_n37236_;
  assign new_n37239_ = ys__n442 & new_n36759_;
  assign new_n37240_ = ys__n440 & new_n36761_;
  assign new_n37241_ = ~new_n37239_ & ~new_n37240_;
  assign new_n37242_ = ys__n23156 & new_n36764_;
  assign new_n37243_ = ys__n23159 & new_n36766_;
  assign new_n37244_ = ~new_n37242_ & ~new_n37243_;
  assign new_n37245_ = new_n37241_ & new_n37244_;
  assign new_n37246_ = new_n36773_ & ~new_n37245_;
  assign new_n37247_ = ~new_n37238_ & ~new_n37246_;
  assign new_n37248_ = new_n36780_ & ~new_n37247_;
  assign new_n37249_ = ~new_n37237_ & ~new_n37248_;
  assign new_n37250_ = ~ys__n738 & ~new_n37249_;
  assign new_n37251_ = new_n36565_ & new_n37236_;
  assign ys__n28814 = new_n37250_ | new_n37251_;
  assign new_n37253_ = ys__n46980 & new_n36467_;
  assign new_n37254_ = ys__n46976 & new_n36457_;
  assign new_n37255_ = ~new_n37253_ & ~new_n37254_;
  assign new_n37256_ = ys__n46974 & new_n36477_;
  assign new_n37257_ = ys__n46973 & new_n36479_;
  assign new_n37258_ = ~new_n37256_ & ~new_n37257_;
  assign new_n37259_ = new_n37255_ & new_n37258_;
  assign new_n37260_ = ~new_n36485_ & ~new_n37259_;
  assign new_n37261_ = new_n36489_ & new_n37260_;
  assign new_n37262_ = new_n36491_ & new_n37260_;
  assign new_n37263_ = ys__n440 & new_n36759_;
  assign new_n37264_ = ys__n444 & new_n36761_;
  assign new_n37265_ = ~new_n37263_ & ~new_n37264_;
  assign new_n37266_ = ys__n23159 & new_n36764_;
  assign new_n37267_ = ys__n23162 & new_n36766_;
  assign new_n37268_ = ~new_n37266_ & ~new_n37267_;
  assign new_n37269_ = new_n37265_ & new_n37268_;
  assign new_n37270_ = new_n36773_ & ~new_n37269_;
  assign new_n37271_ = ~new_n37262_ & ~new_n37270_;
  assign new_n37272_ = new_n36780_ & ~new_n37271_;
  assign new_n37273_ = ~new_n37261_ & ~new_n37272_;
  assign new_n37274_ = ~ys__n738 & ~new_n37273_;
  assign new_n37275_ = new_n36565_ & new_n37260_;
  assign ys__n28816 = new_n37274_ | new_n37275_;
  assign new_n37277_ = ys__n46981 & new_n36467_;
  assign new_n37278_ = ys__n46977 & new_n36457_;
  assign new_n37279_ = ~new_n37277_ & ~new_n37278_;
  assign new_n37280_ = ys__n46975 & new_n36477_;
  assign new_n37281_ = ys__n46974 & new_n36479_;
  assign new_n37282_ = ~new_n37280_ & ~new_n37281_;
  assign new_n37283_ = new_n37279_ & new_n37282_;
  assign new_n37284_ = ~new_n36485_ & ~new_n37283_;
  assign new_n37285_ = new_n36489_ & new_n37284_;
  assign new_n37286_ = new_n36491_ & new_n37284_;
  assign new_n37287_ = ys__n444 & new_n36759_;
  assign new_n37288_ = ys__n438 & new_n36761_;
  assign new_n37289_ = ~new_n37287_ & ~new_n37288_;
  assign new_n37290_ = ys__n23162 & new_n36764_;
  assign new_n37291_ = ys__n23165 & new_n36766_;
  assign new_n37292_ = ~new_n37290_ & ~new_n37291_;
  assign new_n37293_ = new_n37289_ & new_n37292_;
  assign new_n37294_ = new_n36773_ & ~new_n37293_;
  assign new_n37295_ = ~new_n37286_ & ~new_n37294_;
  assign new_n37296_ = new_n36780_ & ~new_n37295_;
  assign new_n37297_ = ~new_n37285_ & ~new_n37296_;
  assign new_n37298_ = ~ys__n738 & ~new_n37297_;
  assign new_n37299_ = new_n36565_ & new_n37284_;
  assign ys__n28818 = new_n37298_ | new_n37299_;
  assign new_n37301_ = ys__n46982 & new_n36467_;
  assign new_n37302_ = ys__n46978 & new_n36457_;
  assign new_n37303_ = ~new_n37301_ & ~new_n37302_;
  assign new_n37304_ = ys__n46976 & new_n36477_;
  assign new_n37305_ = ys__n46975 & new_n36479_;
  assign new_n37306_ = ~new_n37304_ & ~new_n37305_;
  assign new_n37307_ = new_n37303_ & new_n37306_;
  assign new_n37308_ = ~new_n36485_ & ~new_n37307_;
  assign new_n37309_ = new_n36489_ & new_n37308_;
  assign new_n37310_ = new_n36491_ & new_n37308_;
  assign new_n37311_ = ys__n438 & new_n36759_;
  assign new_n37312_ = ys__n446 & new_n36761_;
  assign new_n37313_ = ~new_n37311_ & ~new_n37312_;
  assign new_n37314_ = ys__n23165 & new_n36764_;
  assign new_n37315_ = ys__n23168 & new_n36766_;
  assign new_n37316_ = ~new_n37314_ & ~new_n37315_;
  assign new_n37317_ = new_n37313_ & new_n37316_;
  assign new_n37318_ = new_n36773_ & ~new_n37317_;
  assign new_n37319_ = ~new_n37310_ & ~new_n37318_;
  assign new_n37320_ = new_n36780_ & ~new_n37319_;
  assign new_n37321_ = ~new_n37309_ & ~new_n37320_;
  assign new_n37322_ = ~ys__n738 & ~new_n37321_;
  assign new_n37323_ = new_n36565_ & new_n37308_;
  assign ys__n28820 = new_n37322_ | new_n37323_;
  assign new_n37325_ = ys__n46983 & new_n36467_;
  assign new_n37326_ = ys__n46979 & new_n36457_;
  assign new_n37327_ = ~new_n37325_ & ~new_n37326_;
  assign new_n37328_ = ys__n46977 & new_n36477_;
  assign new_n37329_ = ys__n46976 & new_n36479_;
  assign new_n37330_ = ~new_n37328_ & ~new_n37329_;
  assign new_n37331_ = new_n37327_ & new_n37330_;
  assign new_n37332_ = ~new_n36485_ & ~new_n37331_;
  assign new_n37333_ = new_n36489_ & new_n37332_;
  assign new_n37334_ = new_n36491_ & new_n37332_;
  assign new_n37335_ = ys__n446 & new_n36759_;
  assign new_n37336_ = ys__n434 & new_n36761_;
  assign new_n37337_ = ~new_n37335_ & ~new_n37336_;
  assign new_n37338_ = ys__n23168 & new_n36764_;
  assign new_n37339_ = ys__n23171 & new_n36766_;
  assign new_n37340_ = ~new_n37338_ & ~new_n37339_;
  assign new_n37341_ = new_n37337_ & new_n37340_;
  assign new_n37342_ = new_n36773_ & ~new_n37341_;
  assign new_n37343_ = ~new_n37334_ & ~new_n37342_;
  assign new_n37344_ = new_n36780_ & ~new_n37343_;
  assign new_n37345_ = ~new_n37333_ & ~new_n37344_;
  assign new_n37346_ = ~ys__n738 & ~new_n37345_;
  assign new_n37347_ = new_n36565_ & new_n37332_;
  assign ys__n28822 = new_n37346_ | new_n37347_;
  assign new_n37349_ = ys__n46984 & new_n36467_;
  assign new_n37350_ = ys__n46980 & new_n36457_;
  assign new_n37351_ = ~new_n37349_ & ~new_n37350_;
  assign new_n37352_ = ys__n46978 & new_n36477_;
  assign new_n37353_ = ys__n46977 & new_n36479_;
  assign new_n37354_ = ~new_n37352_ & ~new_n37353_;
  assign new_n37355_ = new_n37351_ & new_n37354_;
  assign new_n37356_ = ~new_n36485_ & ~new_n37355_;
  assign new_n37357_ = new_n36489_ & new_n37356_;
  assign new_n37358_ = new_n36491_ & new_n37356_;
  assign new_n37359_ = ys__n434 & new_n36759_;
  assign new_n37360_ = ys__n436 & new_n36761_;
  assign new_n37361_ = ~new_n37359_ & ~new_n37360_;
  assign new_n37362_ = ys__n23171 & new_n36764_;
  assign new_n37363_ = ys__n23174 & new_n36766_;
  assign new_n37364_ = ~new_n37362_ & ~new_n37363_;
  assign new_n37365_ = new_n37361_ & new_n37364_;
  assign new_n37366_ = new_n36773_ & ~new_n37365_;
  assign new_n37367_ = ~new_n37358_ & ~new_n37366_;
  assign new_n37368_ = new_n36780_ & ~new_n37367_;
  assign new_n37369_ = ~new_n37357_ & ~new_n37368_;
  assign new_n37370_ = ~ys__n738 & ~new_n37369_;
  assign new_n37371_ = new_n36565_ & new_n37356_;
  assign ys__n28824 = new_n37370_ | new_n37371_;
  assign new_n37373_ = ys__n46985 & new_n36467_;
  assign new_n37374_ = ys__n46981 & new_n36457_;
  assign new_n37375_ = ~new_n37373_ & ~new_n37374_;
  assign new_n37376_ = ys__n46979 & new_n36477_;
  assign new_n37377_ = ys__n46978 & new_n36479_;
  assign new_n37378_ = ~new_n37376_ & ~new_n37377_;
  assign new_n37379_ = new_n37375_ & new_n37378_;
  assign new_n37380_ = ~new_n36485_ & ~new_n37379_;
  assign new_n37381_ = new_n36489_ & new_n37380_;
  assign new_n37382_ = new_n36491_ & new_n37380_;
  assign new_n37383_ = ys__n436 & new_n36759_;
  assign new_n37384_ = ys__n432 & new_n36761_;
  assign new_n37385_ = ~new_n37383_ & ~new_n37384_;
  assign new_n37386_ = ys__n23174 & new_n36764_;
  assign new_n37387_ = ys__n23177 & new_n36766_;
  assign new_n37388_ = ~new_n37386_ & ~new_n37387_;
  assign new_n37389_ = new_n37385_ & new_n37388_;
  assign new_n37390_ = new_n36773_ & ~new_n37389_;
  assign new_n37391_ = ~new_n37382_ & ~new_n37390_;
  assign new_n37392_ = new_n36780_ & ~new_n37391_;
  assign new_n37393_ = ~new_n37381_ & ~new_n37392_;
  assign new_n37394_ = ~ys__n738 & ~new_n37393_;
  assign new_n37395_ = new_n36565_ & new_n37380_;
  assign ys__n28826 = new_n37394_ | new_n37395_;
  assign new_n37397_ = ys__n46986 & new_n36467_;
  assign new_n37398_ = ys__n46982 & new_n36457_;
  assign new_n37399_ = ~new_n37397_ & ~new_n37398_;
  assign new_n37400_ = ys__n46980 & new_n36477_;
  assign new_n37401_ = ys__n46979 & new_n36479_;
  assign new_n37402_ = ~new_n37400_ & ~new_n37401_;
  assign new_n37403_ = new_n37399_ & new_n37402_;
  assign new_n37404_ = ~new_n36485_ & ~new_n37403_;
  assign new_n37405_ = new_n36489_ & new_n37404_;
  assign new_n37406_ = new_n36491_ & new_n37404_;
  assign new_n37407_ = ys__n432 & new_n36759_;
  assign new_n37408_ = ys__n448 & new_n36761_;
  assign new_n37409_ = ~new_n37407_ & ~new_n37408_;
  assign new_n37410_ = ys__n23177 & new_n36764_;
  assign new_n37411_ = ys__n23180 & new_n36766_;
  assign new_n37412_ = ~new_n37410_ & ~new_n37411_;
  assign new_n37413_ = new_n37409_ & new_n37412_;
  assign new_n37414_ = new_n36773_ & ~new_n37413_;
  assign new_n37415_ = ~new_n37406_ & ~new_n37414_;
  assign new_n37416_ = new_n36780_ & ~new_n37415_;
  assign new_n37417_ = ~new_n37405_ & ~new_n37416_;
  assign new_n37418_ = ~ys__n738 & ~new_n37417_;
  assign new_n37419_ = new_n36565_ & new_n37404_;
  assign ys__n28828 = new_n37418_ | new_n37419_;
  assign new_n37421_ = ys__n46987 & new_n36467_;
  assign new_n37422_ = ys__n46983 & new_n36457_;
  assign new_n37423_ = ~new_n37421_ & ~new_n37422_;
  assign new_n37424_ = ys__n46981 & new_n36477_;
  assign new_n37425_ = ys__n46980 & new_n36479_;
  assign new_n37426_ = ~new_n37424_ & ~new_n37425_;
  assign new_n37427_ = new_n37423_ & new_n37426_;
  assign new_n37428_ = ~new_n36485_ & ~new_n37427_;
  assign new_n37429_ = new_n36489_ & new_n37428_;
  assign new_n37430_ = new_n36491_ & new_n37428_;
  assign new_n37431_ = ys__n448 & new_n36759_;
  assign new_n37432_ = ys__n428 & new_n36761_;
  assign new_n37433_ = ~new_n37431_ & ~new_n37432_;
  assign new_n37434_ = ys__n23180 & new_n36764_;
  assign new_n37435_ = ys__n23183 & new_n36766_;
  assign new_n37436_ = ~new_n37434_ & ~new_n37435_;
  assign new_n37437_ = new_n37433_ & new_n37436_;
  assign new_n37438_ = new_n36773_ & ~new_n37437_;
  assign new_n37439_ = ~new_n37430_ & ~new_n37438_;
  assign new_n37440_ = new_n36780_ & ~new_n37439_;
  assign new_n37441_ = ~new_n37429_ & ~new_n37440_;
  assign new_n37442_ = ~ys__n738 & ~new_n37441_;
  assign new_n37443_ = new_n36565_ & new_n37428_;
  assign ys__n28830 = new_n37442_ | new_n37443_;
  assign new_n37445_ = ys__n46988 & new_n36467_;
  assign new_n37446_ = ys__n46984 & new_n36457_;
  assign new_n37447_ = ~new_n37445_ & ~new_n37446_;
  assign new_n37448_ = ys__n46982 & new_n36477_;
  assign new_n37449_ = ys__n46981 & new_n36479_;
  assign new_n37450_ = ~new_n37448_ & ~new_n37449_;
  assign new_n37451_ = new_n37447_ & new_n37450_;
  assign new_n37452_ = ~new_n36485_ & ~new_n37451_;
  assign new_n37453_ = new_n36489_ & new_n37452_;
  assign new_n37454_ = new_n36491_ & new_n37452_;
  assign new_n37455_ = ys__n428 & new_n36759_;
  assign new_n37456_ = ys__n430 & new_n36761_;
  assign new_n37457_ = ~new_n37455_ & ~new_n37456_;
  assign new_n37458_ = ys__n23183 & new_n36764_;
  assign new_n37459_ = ys__n23186 & new_n36766_;
  assign new_n37460_ = ~new_n37458_ & ~new_n37459_;
  assign new_n37461_ = new_n37457_ & new_n37460_;
  assign new_n37462_ = new_n36773_ & ~new_n37461_;
  assign new_n37463_ = ~new_n37454_ & ~new_n37462_;
  assign new_n37464_ = new_n36780_ & ~new_n37463_;
  assign new_n37465_ = ~new_n37453_ & ~new_n37464_;
  assign new_n37466_ = ~ys__n738 & ~new_n37465_;
  assign new_n37467_ = new_n36565_ & new_n37452_;
  assign ys__n28832 = new_n37466_ | new_n37467_;
  assign new_n37469_ = ys__n46989 & new_n36467_;
  assign new_n37470_ = ys__n46985 & new_n36457_;
  assign new_n37471_ = ~new_n37469_ & ~new_n37470_;
  assign new_n37472_ = ys__n46983 & new_n36477_;
  assign new_n37473_ = ys__n46982 & new_n36479_;
  assign new_n37474_ = ~new_n37472_ & ~new_n37473_;
  assign new_n37475_ = new_n37471_ & new_n37474_;
  assign new_n37476_ = ~new_n36485_ & ~new_n37475_;
  assign new_n37477_ = new_n36489_ & new_n37476_;
  assign new_n37478_ = new_n36491_ & new_n37476_;
  assign new_n37479_ = ys__n430 & new_n36759_;
  assign new_n37480_ = ys__n426 & new_n36761_;
  assign new_n37481_ = ~new_n37479_ & ~new_n37480_;
  assign new_n37482_ = ys__n23186 & new_n36764_;
  assign new_n37483_ = ys__n23189 & new_n36766_;
  assign new_n37484_ = ~new_n37482_ & ~new_n37483_;
  assign new_n37485_ = new_n37481_ & new_n37484_;
  assign new_n37486_ = new_n36773_ & ~new_n37485_;
  assign new_n37487_ = ~new_n37478_ & ~new_n37486_;
  assign new_n37488_ = new_n36780_ & ~new_n37487_;
  assign new_n37489_ = ~new_n37477_ & ~new_n37488_;
  assign new_n37490_ = ~ys__n738 & ~new_n37489_;
  assign new_n37491_ = new_n36565_ & new_n37476_;
  assign ys__n28834 = new_n37490_ | new_n37491_;
  assign new_n37493_ = ys__n46990 & new_n36467_;
  assign new_n37494_ = ys__n46986 & new_n36457_;
  assign new_n37495_ = ~new_n37493_ & ~new_n37494_;
  assign new_n37496_ = ys__n46984 & new_n36477_;
  assign new_n37497_ = ys__n46983 & new_n36479_;
  assign new_n37498_ = ~new_n37496_ & ~new_n37497_;
  assign new_n37499_ = new_n37495_ & new_n37498_;
  assign new_n37500_ = ~new_n36485_ & ~new_n37499_;
  assign new_n37501_ = new_n36489_ & new_n37500_;
  assign new_n37502_ = new_n36491_ & new_n37500_;
  assign new_n37503_ = ys__n426 & new_n36759_;
  assign new_n37504_ = ys__n450 & new_n36761_;
  assign new_n37505_ = ~new_n37503_ & ~new_n37504_;
  assign new_n37506_ = ys__n23189 & new_n36764_;
  assign new_n37507_ = ys__n23192 & new_n36766_;
  assign new_n37508_ = ~new_n37506_ & ~new_n37507_;
  assign new_n37509_ = new_n37505_ & new_n37508_;
  assign new_n37510_ = new_n36773_ & ~new_n37509_;
  assign new_n37511_ = ~new_n37502_ & ~new_n37510_;
  assign new_n37512_ = new_n36780_ & ~new_n37511_;
  assign new_n37513_ = ~new_n37501_ & ~new_n37512_;
  assign new_n37514_ = ~ys__n738 & ~new_n37513_;
  assign new_n37515_ = new_n36565_ & new_n37500_;
  assign ys__n28836 = new_n37514_ | new_n37515_;
  assign new_n37517_ = ys__n46991 & new_n36467_;
  assign new_n37518_ = ys__n46987 & new_n36457_;
  assign new_n37519_ = ~new_n37517_ & ~new_n37518_;
  assign new_n37520_ = ys__n46985 & new_n36477_;
  assign new_n37521_ = ys__n46984 & new_n36479_;
  assign new_n37522_ = ~new_n37520_ & ~new_n37521_;
  assign new_n37523_ = new_n37519_ & new_n37522_;
  assign new_n37524_ = ~new_n36485_ & ~new_n37523_;
  assign new_n37525_ = new_n36489_ & new_n37524_;
  assign new_n37526_ = new_n36491_ & new_n37524_;
  assign new_n37527_ = ys__n450 & new_n36759_;
  assign new_n37528_ = ys__n424 & new_n36761_;
  assign new_n37529_ = ~new_n37527_ & ~new_n37528_;
  assign new_n37530_ = ys__n23192 & new_n36764_;
  assign new_n37531_ = ys__n23195 & new_n36766_;
  assign new_n37532_ = ~new_n37530_ & ~new_n37531_;
  assign new_n37533_ = new_n37529_ & new_n37532_;
  assign new_n37534_ = new_n36773_ & ~new_n37533_;
  assign new_n37535_ = ~new_n37526_ & ~new_n37534_;
  assign new_n37536_ = new_n36780_ & ~new_n37535_;
  assign new_n37537_ = ~new_n37525_ & ~new_n37536_;
  assign new_n37538_ = ~ys__n738 & ~new_n37537_;
  assign new_n37539_ = new_n36565_ & new_n37524_;
  assign ys__n28838 = new_n37538_ | new_n37539_;
  assign new_n37541_ = ys__n46992 & new_n36467_;
  assign new_n37542_ = ys__n46988 & new_n36457_;
  assign new_n37543_ = ~new_n37541_ & ~new_n37542_;
  assign new_n37544_ = ys__n46986 & new_n36477_;
  assign new_n37545_ = ys__n46985 & new_n36479_;
  assign new_n37546_ = ~new_n37544_ & ~new_n37545_;
  assign new_n37547_ = new_n37543_ & new_n37546_;
  assign new_n37548_ = ~new_n36485_ & ~new_n37547_;
  assign new_n37549_ = new_n36489_ & new_n37548_;
  assign new_n37550_ = new_n36491_ & new_n37548_;
  assign new_n37551_ = ys__n424 & new_n36759_;
  assign new_n37552_ = ys__n422 & new_n36761_;
  assign new_n37553_ = ~new_n37551_ & ~new_n37552_;
  assign new_n37554_ = ys__n23195 & new_n36764_;
  assign new_n37555_ = ys__n23198 & new_n36766_;
  assign new_n37556_ = ~new_n37554_ & ~new_n37555_;
  assign new_n37557_ = new_n37553_ & new_n37556_;
  assign new_n37558_ = new_n36773_ & ~new_n37557_;
  assign new_n37559_ = ~new_n37550_ & ~new_n37558_;
  assign new_n37560_ = new_n36780_ & ~new_n37559_;
  assign new_n37561_ = ~new_n37549_ & ~new_n37560_;
  assign new_n37562_ = ~ys__n738 & ~new_n37561_;
  assign new_n37563_ = new_n36565_ & new_n37548_;
  assign ys__n28840 = new_n37562_ | new_n37563_;
  assign new_n37565_ = ys__n46993 & new_n36467_;
  assign new_n37566_ = ys__n46989 & new_n36457_;
  assign new_n37567_ = ~new_n37565_ & ~new_n37566_;
  assign new_n37568_ = ys__n46987 & new_n36477_;
  assign new_n37569_ = ys__n46986 & new_n36479_;
  assign new_n37570_ = ~new_n37568_ & ~new_n37569_;
  assign new_n37571_ = new_n37567_ & new_n37570_;
  assign new_n37572_ = ~new_n36485_ & ~new_n37571_;
  assign new_n37573_ = new_n36489_ & new_n37572_;
  assign new_n37574_ = new_n36491_ & new_n37572_;
  assign new_n37575_ = ys__n422 & new_n36759_;
  assign new_n37576_ = ys__n23198 & new_n36764_;
  assign new_n37577_ = ~new_n37575_ & ~new_n37576_;
  assign new_n37578_ = new_n36773_ & ~new_n37577_;
  assign new_n37579_ = ~new_n37574_ & ~new_n37578_;
  assign new_n37580_ = new_n36780_ & ~new_n37579_;
  assign new_n37581_ = ~new_n37573_ & ~new_n37580_;
  assign new_n37582_ = ~ys__n738 & ~new_n37581_;
  assign new_n37583_ = new_n36565_ & new_n37572_;
  assign ys__n28842 = new_n37582_ | new_n37583_;
  assign new_n37585_ = ys__n46987 & new_n36479_;
  assign new_n37586_ = ys__n46990 & new_n36457_;
  assign new_n37587_ = ys__n46988 & new_n36477_;
  assign new_n37588_ = ~new_n37586_ & ~new_n37587_;
  assign new_n37589_ = ~new_n37585_ & new_n37588_;
  assign new_n37590_ = ~new_n36485_ & ~new_n37589_;
  assign new_n37591_ = new_n36489_ & new_n37590_;
  assign new_n37592_ = ~ys__n4566 & new_n37590_;
  assign new_n37593_ = new_n36491_ & new_n37592_;
  assign new_n37594_ = ~new_n36779_ & new_n37593_;
  assign new_n37595_ = ~new_n37591_ & ~new_n37594_;
  assign new_n37596_ = ~ys__n738 & ~new_n37595_;
  assign new_n37597_ = new_n36565_ & new_n37590_;
  assign ys__n28844 = new_n37596_ | new_n37597_;
  assign new_n37599_ = ys__n46988 & new_n36479_;
  assign new_n37600_ = ys__n46991 & new_n36457_;
  assign new_n37601_ = ys__n46989 & new_n36477_;
  assign new_n37602_ = ~new_n37600_ & ~new_n37601_;
  assign new_n37603_ = ~new_n37599_ & new_n37602_;
  assign new_n37604_ = ~new_n36485_ & ~new_n37603_;
  assign new_n37605_ = new_n36489_ & new_n37604_;
  assign new_n37606_ = ~ys__n4566 & new_n37604_;
  assign new_n37607_ = new_n36491_ & new_n37606_;
  assign new_n37608_ = ~new_n36779_ & new_n37607_;
  assign new_n37609_ = ~new_n37605_ & ~new_n37608_;
  assign new_n37610_ = ~ys__n738 & ~new_n37609_;
  assign new_n37611_ = new_n36565_ & new_n37604_;
  assign ys__n28846 = new_n37610_ | new_n37611_;
  assign new_n37613_ = ys__n46989 & new_n36479_;
  assign new_n37614_ = ys__n46992 & new_n36457_;
  assign new_n37615_ = ys__n46990 & new_n36477_;
  assign new_n37616_ = ~new_n37614_ & ~new_n37615_;
  assign new_n37617_ = ~new_n37613_ & new_n37616_;
  assign new_n37618_ = ~new_n36485_ & ~new_n37617_;
  assign new_n37619_ = new_n36489_ & new_n37618_;
  assign new_n37620_ = ~ys__n4566 & new_n37618_;
  assign new_n37621_ = new_n36491_ & new_n37620_;
  assign new_n37622_ = ~new_n36779_ & new_n37621_;
  assign new_n37623_ = ~new_n37619_ & ~new_n37622_;
  assign new_n37624_ = ~ys__n738 & ~new_n37623_;
  assign new_n37625_ = new_n36565_ & new_n37618_;
  assign ys__n28848 = new_n37624_ | new_n37625_;
  assign new_n37627_ = ys__n46990 & new_n36479_;
  assign new_n37628_ = ys__n46993 & new_n36457_;
  assign new_n37629_ = ys__n46991 & new_n36477_;
  assign new_n37630_ = ~new_n37628_ & ~new_n37629_;
  assign new_n37631_ = ~new_n37627_ & new_n37630_;
  assign new_n37632_ = ~new_n36485_ & ~new_n37631_;
  assign new_n37633_ = new_n36489_ & new_n37632_;
  assign new_n37634_ = ~ys__n4566 & new_n37632_;
  assign new_n37635_ = new_n36491_ & new_n37634_;
  assign new_n37636_ = ~new_n36779_ & new_n37635_;
  assign new_n37637_ = ~new_n37633_ & ~new_n37636_;
  assign new_n37638_ = ~ys__n738 & ~new_n37637_;
  assign new_n37639_ = new_n36565_ & new_n37632_;
  assign ys__n28850 = new_n37638_ | new_n37639_;
  assign new_n37641_ = ys__n46992 & new_n36477_;
  assign new_n37642_ = ys__n46991 & new_n36479_;
  assign new_n37643_ = ~new_n37641_ & ~new_n37642_;
  assign new_n37644_ = ~new_n36485_ & ~new_n37643_;
  assign new_n37645_ = ys__n4566 & new_n37644_;
  assign new_n37646_ = new_n13716_ & new_n37645_;
  assign new_n37647_ = ~ys__n4566 & new_n37644_;
  assign new_n37648_ = new_n36491_ & new_n37647_;
  assign new_n37649_ = ~new_n36779_ & new_n37648_;
  assign new_n37650_ = ~new_n37646_ & ~new_n37649_;
  assign new_n37651_ = ~ys__n738 & ~new_n37650_;
  assign new_n37652_ = new_n36565_ & new_n37644_;
  assign ys__n28852 = new_n37651_ | new_n37652_;
  assign new_n37654_ = ys__n46993 & new_n36477_;
  assign new_n37655_ = ys__n46992 & new_n36479_;
  assign new_n37656_ = ~new_n37654_ & ~new_n37655_;
  assign new_n37657_ = ~new_n36485_ & ~new_n37656_;
  assign new_n37658_ = ys__n4566 & new_n37657_;
  assign new_n37659_ = new_n13716_ & new_n37658_;
  assign new_n37660_ = ~ys__n4566 & new_n37657_;
  assign new_n37661_ = new_n36491_ & new_n37660_;
  assign new_n37662_ = ~new_n36779_ & new_n37661_;
  assign new_n37663_ = ~new_n37659_ & ~new_n37662_;
  assign new_n37664_ = ~ys__n738 & ~new_n37663_;
  assign new_n37665_ = new_n36565_ & new_n37657_;
  assign ys__n28854 = new_n37664_ | new_n37665_;
  assign new_n37667_ = ys__n46993 & new_n36479_;
  assign new_n37668_ = ~new_n36485_ & new_n37667_;
  assign new_n37669_ = ys__n4566 & new_n37668_;
  assign new_n37670_ = new_n13716_ & new_n37669_;
  assign new_n37671_ = ~ys__n4566 & new_n37668_;
  assign new_n37672_ = new_n36491_ & new_n37671_;
  assign new_n37673_ = ~new_n36779_ & new_n37672_;
  assign new_n37674_ = ~new_n37670_ & ~new_n37673_;
  assign new_n37675_ = ~ys__n738 & ~new_n37674_;
  assign new_n37676_ = new_n36565_ & new_n37668_;
  assign ys__n28856 = new_n37675_ | new_n37676_;
  assign new_n37678_ = ~ys__n4625 & ~ys__n38494;
  assign new_n37679_ = new_n13359_ & new_n37678_;
  assign new_n37680_ = ~new_n24256_ & new_n37679_;
  assign new_n37681_ = ~new_n24248_ & ~new_n24576_;
  assign new_n37682_ = ~new_n24577_ & ~new_n37681_;
  assign new_n37683_ = ~new_n37679_ & ~new_n37682_;
  assign new_n37684_ = ~new_n37680_ & ~new_n37683_;
  assign new_n37685_ = new_n13344_ & ~new_n37684_;
  assign new_n37686_ = ~ys__n740 & ~new_n13344_;
  assign new_n37687_ = ~new_n37684_ & new_n37686_;
  assign ys__n29022 = new_n37685_ | new_n37687_;
  assign new_n37689_ = ~new_n24275_ & new_n37679_;
  assign new_n37690_ = ys__n30014 & ~new_n24549_;
  assign new_n37691_ = ys__n30046 & new_n24549_;
  assign new_n37692_ = ~new_n37690_ & ~new_n37691_;
  assign new_n37693_ = ~new_n24553_ & ~new_n37692_;
  assign new_n37694_ = ys__n30030 & ~new_n24549_;
  assign new_n37695_ = ys__n30062 & new_n24549_;
  assign new_n37696_ = ~new_n37694_ & ~new_n37695_;
  assign new_n37697_ = new_n24553_ & ~new_n37696_;
  assign new_n37698_ = ~new_n37693_ & ~new_n37697_;
  assign new_n37699_ = ~new_n24561_ & ~new_n37698_;
  assign new_n37700_ = ys__n30014 & new_n24561_;
  assign new_n37701_ = ~new_n37699_ & ~new_n37700_;
  assign new_n37702_ = ~new_n24565_ & ~new_n37701_;
  assign new_n37703_ = new_n24576_ & new_n37702_;
  assign new_n37704_ = new_n24267_ & ~new_n24576_;
  assign new_n37705_ = ~new_n37703_ & ~new_n37704_;
  assign new_n37706_ = ~new_n37679_ & ~new_n37705_;
  assign new_n37707_ = ~new_n37689_ & ~new_n37706_;
  assign new_n37708_ = new_n13344_ & ~new_n37707_;
  assign new_n37709_ = new_n37686_ & ~new_n37707_;
  assign ys__n29025 = new_n37708_ | new_n37709_;
  assign new_n37711_ = ~new_n24294_ & new_n37679_;
  assign new_n37712_ = ys__n30016 & ~new_n24549_;
  assign new_n37713_ = ys__n30048 & new_n24549_;
  assign new_n37714_ = ~new_n37712_ & ~new_n37713_;
  assign new_n37715_ = ~new_n24553_ & ~new_n37714_;
  assign new_n37716_ = ys__n30032 & ~new_n24549_;
  assign new_n37717_ = ys__n30064 & new_n24549_;
  assign new_n37718_ = ~new_n37716_ & ~new_n37717_;
  assign new_n37719_ = new_n24553_ & ~new_n37718_;
  assign new_n37720_ = ~new_n37715_ & ~new_n37719_;
  assign new_n37721_ = ~new_n24561_ & ~new_n37720_;
  assign new_n37722_ = ys__n30016 & new_n24561_;
  assign new_n37723_ = ~new_n37721_ & ~new_n37722_;
  assign new_n37724_ = ~new_n24565_ & ~new_n37723_;
  assign new_n37725_ = new_n24576_ & new_n37724_;
  assign new_n37726_ = new_n24286_ & ~new_n24576_;
  assign new_n37727_ = ~new_n37725_ & ~new_n37726_;
  assign new_n37728_ = ~new_n37679_ & ~new_n37727_;
  assign new_n37729_ = ~new_n37711_ & ~new_n37728_;
  assign new_n37730_ = new_n13344_ & ~new_n37729_;
  assign new_n37731_ = new_n37686_ & ~new_n37729_;
  assign ys__n29028 = new_n37730_ | new_n37731_;
  assign new_n37733_ = ~new_n24313_ & new_n37679_;
  assign new_n37734_ = ys__n30018 & ~new_n24549_;
  assign new_n37735_ = ys__n30050 & new_n24549_;
  assign new_n37736_ = ~new_n37734_ & ~new_n37735_;
  assign new_n37737_ = ~new_n24553_ & ~new_n37736_;
  assign new_n37738_ = ys__n30034 & ~new_n24549_;
  assign new_n37739_ = ys__n30066 & new_n24549_;
  assign new_n37740_ = ~new_n37738_ & ~new_n37739_;
  assign new_n37741_ = new_n24553_ & ~new_n37740_;
  assign new_n37742_ = ~new_n37737_ & ~new_n37741_;
  assign new_n37743_ = ~new_n24561_ & ~new_n37742_;
  assign new_n37744_ = ys__n30018 & new_n24561_;
  assign new_n37745_ = ~new_n37743_ & ~new_n37744_;
  assign new_n37746_ = ~new_n24565_ & ~new_n37745_;
  assign new_n37747_ = new_n24576_ & new_n37746_;
  assign new_n37748_ = new_n24305_ & ~new_n24576_;
  assign new_n37749_ = ~new_n37747_ & ~new_n37748_;
  assign new_n37750_ = ~new_n37679_ & ~new_n37749_;
  assign new_n37751_ = ~new_n37733_ & ~new_n37750_;
  assign new_n37752_ = new_n13344_ & ~new_n37751_;
  assign new_n37753_ = new_n37686_ & ~new_n37751_;
  assign ys__n29031 = new_n37752_ | new_n37753_;
  assign new_n37755_ = ~new_n24332_ & new_n37679_;
  assign new_n37756_ = ys__n30020 & ~new_n24549_;
  assign new_n37757_ = ys__n30052 & new_n24549_;
  assign new_n37758_ = ~new_n37756_ & ~new_n37757_;
  assign new_n37759_ = ~new_n24553_ & ~new_n37758_;
  assign new_n37760_ = ys__n30036 & ~new_n24549_;
  assign new_n37761_ = ys__n30068 & new_n24549_;
  assign new_n37762_ = ~new_n37760_ & ~new_n37761_;
  assign new_n37763_ = new_n24553_ & ~new_n37762_;
  assign new_n37764_ = ~new_n37759_ & ~new_n37763_;
  assign new_n37765_ = ~new_n24561_ & ~new_n37764_;
  assign new_n37766_ = ys__n30020 & new_n24561_;
  assign new_n37767_ = ~new_n37765_ & ~new_n37766_;
  assign new_n37768_ = ~new_n24565_ & ~new_n37767_;
  assign new_n37769_ = new_n24576_ & new_n37768_;
  assign new_n37770_ = new_n24324_ & ~new_n24576_;
  assign new_n37771_ = ~new_n37769_ & ~new_n37770_;
  assign new_n37772_ = ~new_n37679_ & ~new_n37771_;
  assign new_n37773_ = ~new_n37755_ & ~new_n37772_;
  assign new_n37774_ = new_n13344_ & ~new_n37773_;
  assign new_n37775_ = new_n37686_ & ~new_n37773_;
  assign ys__n29034 = new_n37774_ | new_n37775_;
  assign new_n37777_ = ~new_n24351_ & new_n37679_;
  assign new_n37778_ = ys__n30022 & ~new_n24549_;
  assign new_n37779_ = ys__n30054 & new_n24549_;
  assign new_n37780_ = ~new_n37778_ & ~new_n37779_;
  assign new_n37781_ = ~new_n24553_ & ~new_n37780_;
  assign new_n37782_ = ys__n30038 & ~new_n24549_;
  assign new_n37783_ = ys__n30070 & new_n24549_;
  assign new_n37784_ = ~new_n37782_ & ~new_n37783_;
  assign new_n37785_ = new_n24553_ & ~new_n37784_;
  assign new_n37786_ = ~new_n37781_ & ~new_n37785_;
  assign new_n37787_ = ~new_n24561_ & ~new_n37786_;
  assign new_n37788_ = ys__n30022 & new_n24561_;
  assign new_n37789_ = ~new_n37787_ & ~new_n37788_;
  assign new_n37790_ = ~new_n24565_ & ~new_n37789_;
  assign new_n37791_ = new_n24576_ & new_n37790_;
  assign new_n37792_ = new_n24343_ & ~new_n24576_;
  assign new_n37793_ = ~new_n37791_ & ~new_n37792_;
  assign new_n37794_ = ~new_n37679_ & ~new_n37793_;
  assign new_n37795_ = ~new_n37777_ & ~new_n37794_;
  assign new_n37796_ = new_n13344_ & ~new_n37795_;
  assign new_n37797_ = new_n37686_ & ~new_n37795_;
  assign ys__n29037 = new_n37796_ | new_n37797_;
  assign new_n37799_ = ~new_n24370_ & new_n37679_;
  assign new_n37800_ = ys__n30024 & ~new_n24549_;
  assign new_n37801_ = ys__n30056 & new_n24549_;
  assign new_n37802_ = ~new_n37800_ & ~new_n37801_;
  assign new_n37803_ = ~new_n24553_ & ~new_n37802_;
  assign new_n37804_ = ys__n30040 & ~new_n24549_;
  assign new_n37805_ = ys__n30072 & new_n24549_;
  assign new_n37806_ = ~new_n37804_ & ~new_n37805_;
  assign new_n37807_ = new_n24553_ & ~new_n37806_;
  assign new_n37808_ = ~new_n37803_ & ~new_n37807_;
  assign new_n37809_ = ~new_n24561_ & ~new_n37808_;
  assign new_n37810_ = ys__n30024 & new_n24561_;
  assign new_n37811_ = ~new_n37809_ & ~new_n37810_;
  assign new_n37812_ = ~new_n24565_ & ~new_n37811_;
  assign new_n37813_ = new_n24576_ & new_n37812_;
  assign new_n37814_ = new_n24362_ & ~new_n24576_;
  assign new_n37815_ = ~new_n37813_ & ~new_n37814_;
  assign new_n37816_ = ~new_n37679_ & ~new_n37815_;
  assign new_n37817_ = ~new_n37799_ & ~new_n37816_;
  assign new_n37818_ = new_n13344_ & ~new_n37817_;
  assign new_n37819_ = new_n37686_ & ~new_n37817_;
  assign ys__n29040 = new_n37818_ | new_n37819_;
  assign new_n37821_ = ~new_n24389_ & new_n37679_;
  assign new_n37822_ = ys__n30026 & ~new_n24549_;
  assign new_n37823_ = ys__n30058 & new_n24549_;
  assign new_n37824_ = ~new_n37822_ & ~new_n37823_;
  assign new_n37825_ = ~new_n24553_ & ~new_n37824_;
  assign new_n37826_ = ys__n30042 & ~new_n24549_;
  assign new_n37827_ = ys__n30074 & new_n24549_;
  assign new_n37828_ = ~new_n37826_ & ~new_n37827_;
  assign new_n37829_ = new_n24553_ & ~new_n37828_;
  assign new_n37830_ = ~new_n37825_ & ~new_n37829_;
  assign new_n37831_ = ~new_n24561_ & ~new_n37830_;
  assign new_n37832_ = ys__n30026 & new_n24561_;
  assign new_n37833_ = ~new_n37831_ & ~new_n37832_;
  assign new_n37834_ = ~new_n24565_ & ~new_n37833_;
  assign new_n37835_ = new_n24576_ & new_n37834_;
  assign new_n37836_ = new_n24381_ & ~new_n24576_;
  assign new_n37837_ = ~new_n37835_ & ~new_n37836_;
  assign new_n37838_ = ~new_n37679_ & ~new_n37837_;
  assign new_n37839_ = ~new_n37821_ & ~new_n37838_;
  assign new_n37840_ = new_n13344_ & ~new_n37839_;
  assign new_n37841_ = new_n37686_ & ~new_n37839_;
  assign ys__n29043 = new_n37840_ | new_n37841_;
  assign new_n37843_ = ~new_n24070_ & new_n37679_;
  assign new_n37844_ = ys__n14 & ~ys__n4688;
  assign new_n37845_ = ~ys__n14 & ys__n4688;
  assign new_n37846_ = ~new_n37844_ & ~new_n37845_;
  assign new_n37847_ = ~ys__n16 & ys__n2693;
  assign new_n37848_ = ys__n16 & ~ys__n2693;
  assign new_n37849_ = ~new_n37847_ & ~new_n37848_;
  assign new_n37850_ = new_n37846_ & ~new_n37849_;
  assign new_n37851_ = ~new_n37846_ & new_n37849_;
  assign new_n37852_ = ~new_n37850_ & ~new_n37851_;
  assign new_n37853_ = ~new_n24557_ & new_n37852_;
  assign new_n37854_ = ys__n14 & ~ys__n16;
  assign new_n37855_ = ~ys__n2693 & new_n37854_;
  assign new_n37856_ = ~ys__n2693 & ~new_n37855_;
  assign new_n37857_ = ~ys__n14 & ~ys__n16;
  assign new_n37858_ = ~ys__n2693 & new_n37857_;
  assign new_n37859_ = ~ys__n2693 & ~new_n37848_;
  assign new_n37860_ = ~new_n37855_ & new_n37859_;
  assign new_n37861_ = ~new_n37858_ & new_n37860_;
  assign new_n37862_ = ~new_n37856_ & ~new_n37861_;
  assign new_n37863_ = ~new_n37859_ & ~new_n37861_;
  assign new_n37864_ = new_n37862_ & new_n37863_;
  assign new_n37865_ = ys__n30074 & new_n37864_;
  assign new_n37866_ = ~new_n37862_ & new_n37863_;
  assign new_n37867_ = ys__n30058 & new_n37866_;
  assign new_n37868_ = ~new_n37865_ & ~new_n37867_;
  assign new_n37869_ = new_n37862_ & ~new_n37863_;
  assign new_n37870_ = ys__n30042 & new_n37869_;
  assign new_n37871_ = ~new_n37862_ & ~new_n37863_;
  assign new_n37872_ = ys__n30026 & new_n37871_;
  assign new_n37873_ = ~new_n37870_ & ~new_n37872_;
  assign new_n37874_ = new_n37868_ & new_n37873_;
  assign new_n37875_ = ~new_n37864_ & ~new_n37866_;
  assign new_n37876_ = ~new_n37869_ & ~new_n37871_;
  assign new_n37877_ = new_n37875_ & new_n37876_;
  assign new_n37878_ = ys__n38724 & ~new_n37877_;
  assign new_n37879_ = ~new_n37874_ & new_n37878_;
  assign new_n37880_ = ~new_n37852_ & new_n37879_;
  assign new_n37881_ = ~new_n37853_ & ~new_n37880_;
  assign new_n37882_ = ~new_n24561_ & ~new_n37881_;
  assign new_n37883_ = ys__n30028 & new_n24561_;
  assign new_n37884_ = ~new_n37882_ & ~new_n37883_;
  assign new_n37885_ = ~new_n24565_ & ~new_n37884_;
  assign new_n37886_ = new_n24576_ & new_n37885_;
  assign new_n37887_ = new_n24062_ & ~new_n24576_;
  assign new_n37888_ = ~new_n37886_ & ~new_n37887_;
  assign new_n37889_ = ~new_n37679_ & ~new_n37888_;
  assign new_n37890_ = ~new_n37843_ & ~new_n37889_;
  assign new_n37891_ = new_n13344_ & ~new_n37890_;
  assign new_n37892_ = new_n37686_ & ~new_n37890_;
  assign ys__n29046 = new_n37891_ | new_n37892_;
  assign new_n37894_ = ~new_n24088_ & new_n37679_;
  assign new_n37895_ = ~new_n37696_ & new_n37852_;
  assign new_n37896_ = ~new_n37880_ & ~new_n37895_;
  assign new_n37897_ = ~new_n24561_ & ~new_n37896_;
  assign new_n37898_ = ys__n30030 & new_n24561_;
  assign new_n37899_ = ~new_n37897_ & ~new_n37898_;
  assign new_n37900_ = ~new_n24565_ & ~new_n37899_;
  assign new_n37901_ = new_n24576_ & new_n37900_;
  assign new_n37902_ = new_n24080_ & ~new_n24576_;
  assign new_n37903_ = ~new_n37901_ & ~new_n37902_;
  assign new_n37904_ = ~new_n37679_ & ~new_n37903_;
  assign new_n37905_ = ~new_n37894_ & ~new_n37904_;
  assign new_n37906_ = new_n13344_ & ~new_n37905_;
  assign new_n37907_ = new_n37686_ & ~new_n37905_;
  assign ys__n29049 = new_n37906_ | new_n37907_;
  assign new_n37909_ = ~new_n24106_ & new_n37679_;
  assign new_n37910_ = ~new_n37718_ & new_n37852_;
  assign new_n37911_ = ~new_n37880_ & ~new_n37910_;
  assign new_n37912_ = ~new_n24561_ & ~new_n37911_;
  assign new_n37913_ = ys__n30032 & new_n24561_;
  assign new_n37914_ = ~new_n37912_ & ~new_n37913_;
  assign new_n37915_ = ~new_n24565_ & ~new_n37914_;
  assign new_n37916_ = new_n24576_ & new_n37915_;
  assign new_n37917_ = new_n24098_ & ~new_n24576_;
  assign new_n37918_ = ~new_n37916_ & ~new_n37917_;
  assign new_n37919_ = ~new_n37679_ & ~new_n37918_;
  assign new_n37920_ = ~new_n37909_ & ~new_n37919_;
  assign new_n37921_ = new_n13344_ & ~new_n37920_;
  assign new_n37922_ = new_n37686_ & ~new_n37920_;
  assign ys__n29052 = new_n37921_ | new_n37922_;
  assign new_n37924_ = ~new_n24124_ & new_n37679_;
  assign new_n37925_ = ~new_n37740_ & new_n37852_;
  assign new_n37926_ = ~new_n37880_ & ~new_n37925_;
  assign new_n37927_ = ~new_n24561_ & ~new_n37926_;
  assign new_n37928_ = ys__n30034 & new_n24561_;
  assign new_n37929_ = ~new_n37927_ & ~new_n37928_;
  assign new_n37930_ = ~new_n24565_ & ~new_n37929_;
  assign new_n37931_ = new_n24576_ & new_n37930_;
  assign new_n37932_ = new_n24116_ & ~new_n24576_;
  assign new_n37933_ = ~new_n37931_ & ~new_n37932_;
  assign new_n37934_ = ~new_n37679_ & ~new_n37933_;
  assign new_n37935_ = ~new_n37924_ & ~new_n37934_;
  assign new_n37936_ = new_n13344_ & ~new_n37935_;
  assign new_n37937_ = new_n37686_ & ~new_n37935_;
  assign ys__n29055 = new_n37936_ | new_n37937_;
  assign new_n37939_ = ~new_n24142_ & new_n37679_;
  assign new_n37940_ = ~new_n37762_ & new_n37852_;
  assign new_n37941_ = ~new_n37880_ & ~new_n37940_;
  assign new_n37942_ = ~new_n24561_ & ~new_n37941_;
  assign new_n37943_ = ys__n30036 & new_n24561_;
  assign new_n37944_ = ~new_n37942_ & ~new_n37943_;
  assign new_n37945_ = ~new_n24565_ & ~new_n37944_;
  assign new_n37946_ = new_n24576_ & new_n37945_;
  assign new_n37947_ = new_n24134_ & ~new_n24576_;
  assign new_n37948_ = ~new_n37946_ & ~new_n37947_;
  assign new_n37949_ = ~new_n37679_ & ~new_n37948_;
  assign new_n37950_ = ~new_n37939_ & ~new_n37949_;
  assign new_n37951_ = new_n13344_ & ~new_n37950_;
  assign new_n37952_ = new_n37686_ & ~new_n37950_;
  assign ys__n29058 = new_n37951_ | new_n37952_;
  assign new_n37954_ = ~new_n24160_ & new_n37679_;
  assign new_n37955_ = ~new_n37784_ & new_n37852_;
  assign new_n37956_ = ~new_n37880_ & ~new_n37955_;
  assign new_n37957_ = ~new_n24561_ & ~new_n37956_;
  assign new_n37958_ = ys__n30038 & new_n24561_;
  assign new_n37959_ = ~new_n37957_ & ~new_n37958_;
  assign new_n37960_ = ~new_n24565_ & ~new_n37959_;
  assign new_n37961_ = new_n24576_ & new_n37960_;
  assign new_n37962_ = new_n24152_ & ~new_n24576_;
  assign new_n37963_ = ~new_n37961_ & ~new_n37962_;
  assign new_n37964_ = ~new_n37679_ & ~new_n37963_;
  assign new_n37965_ = ~new_n37954_ & ~new_n37964_;
  assign new_n37966_ = new_n13344_ & ~new_n37965_;
  assign new_n37967_ = new_n37686_ & ~new_n37965_;
  assign ys__n29061 = new_n37966_ | new_n37967_;
  assign new_n37969_ = ~new_n24178_ & new_n37679_;
  assign new_n37970_ = ~new_n37806_ & new_n37852_;
  assign new_n37971_ = ~new_n37880_ & ~new_n37970_;
  assign new_n37972_ = ~new_n24561_ & ~new_n37971_;
  assign new_n37973_ = ys__n30040 & new_n24561_;
  assign new_n37974_ = ~new_n37972_ & ~new_n37973_;
  assign new_n37975_ = ~new_n24565_ & ~new_n37974_;
  assign new_n37976_ = new_n24576_ & new_n37975_;
  assign new_n37977_ = new_n24170_ & ~new_n24576_;
  assign new_n37978_ = ~new_n37976_ & ~new_n37977_;
  assign new_n37979_ = ~new_n37679_ & ~new_n37978_;
  assign new_n37980_ = ~new_n37969_ & ~new_n37979_;
  assign new_n37981_ = new_n13344_ & ~new_n37980_;
  assign new_n37982_ = new_n37686_ & ~new_n37980_;
  assign ys__n29064 = new_n37981_ | new_n37982_;
  assign new_n37984_ = ~new_n24196_ & new_n37679_;
  assign new_n37985_ = ~new_n37828_ & new_n37852_;
  assign new_n37986_ = ~new_n37880_ & ~new_n37985_;
  assign new_n37987_ = ~new_n24561_ & ~new_n37986_;
  assign new_n37988_ = ys__n30042 & new_n24561_;
  assign new_n37989_ = ~new_n37987_ & ~new_n37988_;
  assign new_n37990_ = ~new_n24565_ & ~new_n37989_;
  assign new_n37991_ = new_n24576_ & new_n37990_;
  assign new_n37992_ = new_n24188_ & ~new_n24576_;
  assign new_n37993_ = ~new_n37991_ & ~new_n37992_;
  assign new_n37994_ = ~new_n37679_ & ~new_n37993_;
  assign new_n37995_ = ~new_n37984_ & ~new_n37994_;
  assign new_n37996_ = new_n13344_ & ~new_n37995_;
  assign new_n37997_ = new_n37686_ & ~new_n37995_;
  assign ys__n29067 = new_n37996_ | new_n37997_;
  assign new_n37999_ = ~new_n23910_ & new_n37679_;
  assign new_n38000_ = ys__n14 & ys__n16;
  assign new_n38001_ = ys__n2693 & ys__n4688;
  assign new_n38002_ = new_n38000_ & new_n38001_;
  assign new_n38003_ = ys__n30044 & new_n38002_;
  assign new_n38004_ = new_n37879_ & ~new_n38002_;
  assign new_n38005_ = ~new_n38003_ & ~new_n38004_;
  assign new_n38006_ = ~new_n24561_ & ~new_n38005_;
  assign new_n38007_ = ys__n30044 & new_n24561_;
  assign new_n38008_ = ~new_n38006_ & ~new_n38007_;
  assign new_n38009_ = ~new_n24565_ & ~new_n38008_;
  assign new_n38010_ = new_n24576_ & new_n38009_;
  assign new_n38011_ = new_n23902_ & ~new_n24576_;
  assign new_n38012_ = ~new_n38010_ & ~new_n38011_;
  assign new_n38013_ = ~new_n37679_ & ~new_n38012_;
  assign new_n38014_ = ~new_n37999_ & ~new_n38013_;
  assign new_n38015_ = new_n13344_ & ~new_n38014_;
  assign new_n38016_ = new_n37686_ & ~new_n38014_;
  assign ys__n29070 = new_n38015_ | new_n38016_;
  assign new_n38018_ = ~new_n23925_ & new_n37679_;
  assign new_n38019_ = ys__n30046 & new_n38002_;
  assign new_n38020_ = ~new_n38004_ & ~new_n38019_;
  assign new_n38021_ = ~new_n24561_ & ~new_n38020_;
  assign new_n38022_ = ys__n30046 & new_n24561_;
  assign new_n38023_ = ~new_n38021_ & ~new_n38022_;
  assign new_n38024_ = ~new_n24565_ & ~new_n38023_;
  assign new_n38025_ = new_n24576_ & new_n38024_;
  assign new_n38026_ = new_n23917_ & ~new_n24576_;
  assign new_n38027_ = ~new_n38025_ & ~new_n38026_;
  assign new_n38028_ = ~new_n37679_ & ~new_n38027_;
  assign new_n38029_ = ~new_n38018_ & ~new_n38028_;
  assign new_n38030_ = new_n13344_ & ~new_n38029_;
  assign new_n38031_ = new_n37686_ & ~new_n38029_;
  assign ys__n29073 = new_n38030_ | new_n38031_;
  assign new_n38033_ = ~new_n23940_ & new_n37679_;
  assign new_n38034_ = ys__n30048 & new_n38002_;
  assign new_n38035_ = ~new_n38004_ & ~new_n38034_;
  assign new_n38036_ = ~new_n24561_ & ~new_n38035_;
  assign new_n38037_ = ys__n30048 & new_n24561_;
  assign new_n38038_ = ~new_n38036_ & ~new_n38037_;
  assign new_n38039_ = ~new_n24565_ & ~new_n38038_;
  assign new_n38040_ = new_n24576_ & new_n38039_;
  assign new_n38041_ = new_n23932_ & ~new_n24576_;
  assign new_n38042_ = ~new_n38040_ & ~new_n38041_;
  assign new_n38043_ = ~new_n37679_ & ~new_n38042_;
  assign new_n38044_ = ~new_n38033_ & ~new_n38043_;
  assign new_n38045_ = new_n13344_ & ~new_n38044_;
  assign new_n38046_ = new_n37686_ & ~new_n38044_;
  assign ys__n29076 = new_n38045_ | new_n38046_;
  assign new_n38048_ = ~new_n23955_ & new_n37679_;
  assign new_n38049_ = ys__n30050 & new_n38002_;
  assign new_n38050_ = ~new_n38004_ & ~new_n38049_;
  assign new_n38051_ = ~new_n24561_ & ~new_n38050_;
  assign new_n38052_ = ys__n30050 & new_n24561_;
  assign new_n38053_ = ~new_n38051_ & ~new_n38052_;
  assign new_n38054_ = ~new_n24565_ & ~new_n38053_;
  assign new_n38055_ = new_n24576_ & new_n38054_;
  assign new_n38056_ = new_n23947_ & ~new_n24576_;
  assign new_n38057_ = ~new_n38055_ & ~new_n38056_;
  assign new_n38058_ = ~new_n37679_ & ~new_n38057_;
  assign new_n38059_ = ~new_n38048_ & ~new_n38058_;
  assign new_n38060_ = new_n13344_ & ~new_n38059_;
  assign new_n38061_ = new_n37686_ & ~new_n38059_;
  assign ys__n29079 = new_n38060_ | new_n38061_;
  assign new_n38063_ = ~new_n23970_ & new_n37679_;
  assign new_n38064_ = ys__n30052 & new_n38002_;
  assign new_n38065_ = ~new_n38004_ & ~new_n38064_;
  assign new_n38066_ = ~new_n24561_ & ~new_n38065_;
  assign new_n38067_ = ys__n30052 & new_n24561_;
  assign new_n38068_ = ~new_n38066_ & ~new_n38067_;
  assign new_n38069_ = ~new_n24565_ & ~new_n38068_;
  assign new_n38070_ = new_n24576_ & new_n38069_;
  assign new_n38071_ = new_n23962_ & ~new_n24576_;
  assign new_n38072_ = ~new_n38070_ & ~new_n38071_;
  assign new_n38073_ = ~new_n37679_ & ~new_n38072_;
  assign new_n38074_ = ~new_n38063_ & ~new_n38073_;
  assign new_n38075_ = new_n13344_ & ~new_n38074_;
  assign new_n38076_ = new_n37686_ & ~new_n38074_;
  assign ys__n29082 = new_n38075_ | new_n38076_;
  assign new_n38078_ = ~new_n23985_ & new_n37679_;
  assign new_n38079_ = ys__n30054 & new_n38002_;
  assign new_n38080_ = ~new_n38004_ & ~new_n38079_;
  assign new_n38081_ = ~new_n24561_ & ~new_n38080_;
  assign new_n38082_ = ys__n30054 & new_n24561_;
  assign new_n38083_ = ~new_n38081_ & ~new_n38082_;
  assign new_n38084_ = ~new_n24565_ & ~new_n38083_;
  assign new_n38085_ = new_n24576_ & new_n38084_;
  assign new_n38086_ = new_n23977_ & ~new_n24576_;
  assign new_n38087_ = ~new_n38085_ & ~new_n38086_;
  assign new_n38088_ = ~new_n37679_ & ~new_n38087_;
  assign new_n38089_ = ~new_n38078_ & ~new_n38088_;
  assign new_n38090_ = new_n13344_ & ~new_n38089_;
  assign new_n38091_ = new_n37686_ & ~new_n38089_;
  assign ys__n29085 = new_n38090_ | new_n38091_;
  assign new_n38093_ = ~new_n24000_ & new_n37679_;
  assign new_n38094_ = ys__n30056 & new_n38002_;
  assign new_n38095_ = ~new_n38004_ & ~new_n38094_;
  assign new_n38096_ = ~new_n24561_ & ~new_n38095_;
  assign new_n38097_ = ys__n30056 & new_n24561_;
  assign new_n38098_ = ~new_n38096_ & ~new_n38097_;
  assign new_n38099_ = ~new_n24565_ & ~new_n38098_;
  assign new_n38100_ = new_n24576_ & new_n38099_;
  assign new_n38101_ = new_n23992_ & ~new_n24576_;
  assign new_n38102_ = ~new_n38100_ & ~new_n38101_;
  assign new_n38103_ = ~new_n37679_ & ~new_n38102_;
  assign new_n38104_ = ~new_n38093_ & ~new_n38103_;
  assign new_n38105_ = new_n13344_ & ~new_n38104_;
  assign new_n38106_ = new_n37686_ & ~new_n38104_;
  assign ys__n29088 = new_n38105_ | new_n38106_;
  assign new_n38108_ = ~new_n24015_ & new_n37679_;
  assign new_n38109_ = ys__n30058 & new_n38002_;
  assign new_n38110_ = ~new_n38004_ & ~new_n38109_;
  assign new_n38111_ = ~new_n24561_ & ~new_n38110_;
  assign new_n38112_ = ys__n30058 & new_n24561_;
  assign new_n38113_ = ~new_n38111_ & ~new_n38112_;
  assign new_n38114_ = ~new_n24565_ & ~new_n38113_;
  assign new_n38115_ = new_n24576_ & new_n38114_;
  assign new_n38116_ = new_n24007_ & ~new_n24576_;
  assign new_n38117_ = ~new_n38115_ & ~new_n38116_;
  assign new_n38118_ = ~new_n37679_ & ~new_n38117_;
  assign new_n38119_ = ~new_n38108_ & ~new_n38118_;
  assign new_n38120_ = new_n13344_ & ~new_n38119_;
  assign new_n38121_ = new_n37686_ & ~new_n38119_;
  assign ys__n29091 = new_n38120_ | new_n38121_;
  assign new_n38123_ = ~new_n23762_ & new_n37679_;
  assign new_n38124_ = ys__n30060 & new_n38002_;
  assign new_n38125_ = ~new_n38004_ & ~new_n38124_;
  assign new_n38126_ = ~new_n24561_ & ~new_n38125_;
  assign new_n38127_ = ys__n30060 & new_n24561_;
  assign new_n38128_ = ~new_n38126_ & ~new_n38127_;
  assign new_n38129_ = ~new_n24565_ & ~new_n38128_;
  assign new_n38130_ = new_n24576_ & new_n38129_;
  assign new_n38131_ = new_n23748_ & ~new_n24576_;
  assign new_n38132_ = ~new_n38130_ & ~new_n38131_;
  assign new_n38133_ = ~new_n37679_ & ~new_n38132_;
  assign new_n38134_ = ~new_n38123_ & ~new_n38133_;
  assign new_n38135_ = new_n13344_ & ~new_n38134_;
  assign new_n38136_ = new_n37686_ & ~new_n38134_;
  assign ys__n29094 = new_n38135_ | new_n38136_;
  assign new_n38138_ = ~new_n23777_ & new_n37679_;
  assign new_n38139_ = ys__n30062 & new_n38002_;
  assign new_n38140_ = ~new_n38004_ & ~new_n38139_;
  assign new_n38141_ = ~new_n24561_ & ~new_n38140_;
  assign new_n38142_ = ys__n30062 & new_n24561_;
  assign new_n38143_ = ~new_n38141_ & ~new_n38142_;
  assign new_n38144_ = ~new_n24565_ & ~new_n38143_;
  assign new_n38145_ = new_n24576_ & new_n38144_;
  assign new_n38146_ = new_n23769_ & ~new_n24576_;
  assign new_n38147_ = ~new_n38145_ & ~new_n38146_;
  assign new_n38148_ = ~new_n37679_ & ~new_n38147_;
  assign new_n38149_ = ~new_n38138_ & ~new_n38148_;
  assign new_n38150_ = new_n13344_ & ~new_n38149_;
  assign new_n38151_ = new_n37686_ & ~new_n38149_;
  assign ys__n29097 = new_n38150_ | new_n38151_;
  assign new_n38153_ = ~new_n23792_ & new_n37679_;
  assign new_n38154_ = ys__n30064 & new_n38002_;
  assign new_n38155_ = ~new_n38004_ & ~new_n38154_;
  assign new_n38156_ = ~new_n24561_ & ~new_n38155_;
  assign new_n38157_ = ys__n30064 & new_n24561_;
  assign new_n38158_ = ~new_n38156_ & ~new_n38157_;
  assign new_n38159_ = ~new_n24565_ & ~new_n38158_;
  assign new_n38160_ = new_n24576_ & new_n38159_;
  assign new_n38161_ = new_n23784_ & ~new_n24576_;
  assign new_n38162_ = ~new_n38160_ & ~new_n38161_;
  assign new_n38163_ = ~new_n37679_ & ~new_n38162_;
  assign new_n38164_ = ~new_n38153_ & ~new_n38163_;
  assign new_n38165_ = new_n13344_ & ~new_n38164_;
  assign new_n38166_ = new_n37686_ & ~new_n38164_;
  assign ys__n29100 = new_n38165_ | new_n38166_;
  assign new_n38168_ = ~new_n23807_ & new_n37679_;
  assign new_n38169_ = ys__n30066 & new_n38002_;
  assign new_n38170_ = ~new_n38004_ & ~new_n38169_;
  assign new_n38171_ = ~new_n24561_ & ~new_n38170_;
  assign new_n38172_ = ys__n30066 & new_n24561_;
  assign new_n38173_ = ~new_n38171_ & ~new_n38172_;
  assign new_n38174_ = ~new_n24565_ & ~new_n38173_;
  assign new_n38175_ = new_n24576_ & new_n38174_;
  assign new_n38176_ = new_n23799_ & ~new_n24576_;
  assign new_n38177_ = ~new_n38175_ & ~new_n38176_;
  assign new_n38178_ = ~new_n37679_ & ~new_n38177_;
  assign new_n38179_ = ~new_n38168_ & ~new_n38178_;
  assign new_n38180_ = new_n13344_ & ~new_n38179_;
  assign new_n38181_ = new_n37686_ & ~new_n38179_;
  assign ys__n29103 = new_n38180_ | new_n38181_;
  assign new_n38183_ = ~new_n23822_ & new_n37679_;
  assign new_n38184_ = ys__n30068 & new_n38002_;
  assign new_n38185_ = ~new_n38004_ & ~new_n38184_;
  assign new_n38186_ = ~new_n24561_ & ~new_n38185_;
  assign new_n38187_ = ys__n30068 & new_n24561_;
  assign new_n38188_ = ~new_n38186_ & ~new_n38187_;
  assign new_n38189_ = ~new_n24565_ & ~new_n38188_;
  assign new_n38190_ = new_n24576_ & new_n38189_;
  assign new_n38191_ = new_n23814_ & ~new_n24576_;
  assign new_n38192_ = ~new_n38190_ & ~new_n38191_;
  assign new_n38193_ = ~new_n37679_ & ~new_n38192_;
  assign new_n38194_ = ~new_n38183_ & ~new_n38193_;
  assign new_n38195_ = new_n13344_ & ~new_n38194_;
  assign new_n38196_ = new_n37686_ & ~new_n38194_;
  assign ys__n29106 = new_n38195_ | new_n38196_;
  assign new_n38198_ = ~new_n23837_ & new_n37679_;
  assign new_n38199_ = ys__n30070 & new_n38002_;
  assign new_n38200_ = ~new_n38004_ & ~new_n38199_;
  assign new_n38201_ = ~new_n24561_ & ~new_n38200_;
  assign new_n38202_ = ys__n30070 & new_n24561_;
  assign new_n38203_ = ~new_n38201_ & ~new_n38202_;
  assign new_n38204_ = ~new_n24565_ & ~new_n38203_;
  assign new_n38205_ = new_n24576_ & new_n38204_;
  assign new_n38206_ = new_n23829_ & ~new_n24576_;
  assign new_n38207_ = ~new_n38205_ & ~new_n38206_;
  assign new_n38208_ = ~new_n37679_ & ~new_n38207_;
  assign new_n38209_ = ~new_n38198_ & ~new_n38208_;
  assign new_n38210_ = new_n13344_ & ~new_n38209_;
  assign new_n38211_ = new_n37686_ & ~new_n38209_;
  assign ys__n29109 = new_n38210_ | new_n38211_;
  assign new_n38213_ = ~new_n23852_ & new_n37679_;
  assign new_n38214_ = ys__n30072 & new_n38002_;
  assign new_n38215_ = ~new_n38004_ & ~new_n38214_;
  assign new_n38216_ = ~new_n24561_ & ~new_n38215_;
  assign new_n38217_ = ys__n30072 & new_n24561_;
  assign new_n38218_ = ~new_n38216_ & ~new_n38217_;
  assign new_n38219_ = ~new_n24565_ & ~new_n38218_;
  assign new_n38220_ = new_n24576_ & new_n38219_;
  assign new_n38221_ = new_n23844_ & ~new_n24576_;
  assign new_n38222_ = ~new_n38220_ & ~new_n38221_;
  assign new_n38223_ = ~new_n37679_ & ~new_n38222_;
  assign new_n38224_ = ~new_n38213_ & ~new_n38223_;
  assign new_n38225_ = new_n13344_ & ~new_n38224_;
  assign new_n38226_ = new_n37686_ & ~new_n38224_;
  assign ys__n29112 = new_n38225_ | new_n38226_;
  assign new_n38228_ = ~new_n23867_ & new_n37679_;
  assign new_n38229_ = ys__n30074 & new_n38002_;
  assign new_n38230_ = ~new_n38004_ & ~new_n38229_;
  assign new_n38231_ = ~new_n24561_ & ~new_n38230_;
  assign new_n38232_ = ys__n30074 & new_n24561_;
  assign new_n38233_ = ~new_n38231_ & ~new_n38232_;
  assign new_n38234_ = ~new_n24565_ & ~new_n38233_;
  assign new_n38235_ = new_n24576_ & new_n38234_;
  assign new_n38236_ = new_n23859_ & ~new_n24576_;
  assign new_n38237_ = ~new_n38235_ & ~new_n38236_;
  assign new_n38238_ = ~new_n37679_ & ~new_n38237_;
  assign new_n38239_ = ~new_n38228_ & ~new_n38238_;
  assign new_n38240_ = new_n13344_ & ~new_n38239_;
  assign new_n38241_ = new_n37686_ & ~new_n38239_;
  assign ys__n29115 = new_n38240_ | new_n38241_;
  assign new_n38243_ = new_n22682_ & new_n22684_;
  assign new_n38244_ = new_n22668_ & new_n22672_;
  assign new_n38245_ = ~new_n38243_ & ~new_n38244_;
  assign new_n38246_ = ~new_n22689_ & new_n22695_;
  assign new_n38247_ = ~new_n38245_ & new_n38246_;
  assign new_n38248_ = ~new_n22695_ & new_n22721_;
  assign new_n38249_ = new_n22717_ & new_n38248_;
  assign new_n38250_ = ~new_n38247_ & ~new_n38249_;
  assign new_n38251_ = ~ys__n28243 & ~ys__n29117;
  assign ys__n29118 = ~new_n38250_ & new_n38251_;
  assign new_n38253_ = ys__n29119 & ~ys__n29121;
  assign new_n38254_ = ys__n29120 & ys__n29121;
  assign ys__n29122 = new_n38253_ | new_n38254_;
  assign new_n38256_ = ~ys__n29121 & ys__n29123;
  assign new_n38257_ = ys__n29121 & ys__n29124;
  assign ys__n29125 = new_n38256_ | new_n38257_;
  assign new_n38259_ = ~ys__n29121 & ys__n29126;
  assign new_n38260_ = ys__n29121 & ys__n29127;
  assign ys__n29128 = new_n38259_ | new_n38260_;
  assign new_n38262_ = ~ys__n29121 & ys__n29129;
  assign new_n38263_ = ys__n29121 & ys__n29130;
  assign ys__n29131 = new_n38262_ | new_n38263_;
  assign new_n38265_ = ~ys__n29121 & ys__n29132;
  assign new_n38266_ = ys__n29121 & ys__n29133;
  assign ys__n29134 = new_n38265_ | new_n38266_;
  assign new_n38268_ = ~ys__n29121 & ys__n29135;
  assign new_n38269_ = ys__n29121 & ys__n29136;
  assign ys__n29137 = new_n38268_ | new_n38269_;
  assign new_n38271_ = ~ys__n29121 & ys__n29138;
  assign new_n38272_ = ys__n29121 & ys__n29139;
  assign ys__n29140 = new_n38271_ | new_n38272_;
  assign new_n38274_ = ~ys__n29121 & ys__n29141;
  assign new_n38275_ = ys__n29121 & ys__n29142;
  assign ys__n29143 = new_n38274_ | new_n38275_;
  assign new_n38277_ = ~ys__n29121 & ys__n29144;
  assign new_n38278_ = ys__n29121 & ys__n29145;
  assign ys__n29146 = new_n38277_ | new_n38278_;
  assign new_n38280_ = ~ys__n29121 & ys__n29147;
  assign new_n38281_ = ys__n29121 & ys__n29148;
  assign ys__n29149 = new_n38280_ | new_n38281_;
  assign new_n38283_ = ~ys__n29121 & ys__n29150;
  assign new_n38284_ = ys__n29121 & ys__n29151;
  assign ys__n29152 = new_n38283_ | new_n38284_;
  assign new_n38286_ = ~ys__n29121 & ys__n29153;
  assign new_n38287_ = ys__n29121 & ys__n29154;
  assign ys__n29155 = new_n38286_ | new_n38287_;
  assign new_n38289_ = ~ys__n29121 & ys__n29156;
  assign new_n38290_ = ys__n29121 & ys__n29157;
  assign ys__n29158 = new_n38289_ | new_n38290_;
  assign new_n38292_ = ~ys__n29121 & ys__n29159;
  assign new_n38293_ = ys__n29121 & ys__n29160;
  assign ys__n29161 = new_n38292_ | new_n38293_;
  assign new_n38295_ = ~ys__n29121 & ys__n29162;
  assign new_n38296_ = ys__n29121 & ys__n29163;
  assign ys__n29164 = new_n38295_ | new_n38296_;
  assign new_n38298_ = ~ys__n29121 & ys__n29165;
  assign new_n38299_ = ys__n29121 & ys__n29166;
  assign ys__n29167 = new_n38298_ | new_n38299_;
  assign new_n38301_ = ~ys__n29121 & ys__n29168;
  assign new_n38302_ = ys__n29121 & ys__n29169;
  assign ys__n29170 = new_n38301_ | new_n38302_;
  assign new_n38304_ = ~ys__n29121 & ys__n29171;
  assign new_n38305_ = ys__n29121 & ys__n29172;
  assign ys__n29173 = new_n38304_ | new_n38305_;
  assign new_n38307_ = ~ys__n29121 & ys__n29174;
  assign new_n38308_ = ys__n29121 & ys__n29175;
  assign ys__n29176 = new_n38307_ | new_n38308_;
  assign new_n38310_ = ~ys__n29121 & ys__n29177;
  assign new_n38311_ = ys__n29121 & ys__n29178;
  assign ys__n29179 = new_n38310_ | new_n38311_;
  assign new_n38313_ = ~ys__n29121 & ys__n29180;
  assign new_n38314_ = ys__n29121 & ys__n29181;
  assign ys__n29182 = new_n38313_ | new_n38314_;
  assign new_n38316_ = ~ys__n29121 & ys__n29183;
  assign new_n38317_ = ys__n29121 & ys__n29184;
  assign ys__n29185 = new_n38316_ | new_n38317_;
  assign new_n38319_ = ~ys__n29121 & ys__n29186;
  assign new_n38320_ = ys__n29121 & ys__n29187;
  assign ys__n29188 = new_n38319_ | new_n38320_;
  assign new_n38322_ = ~ys__n29121 & ys__n29189;
  assign new_n38323_ = ys__n29121 & ys__n29190;
  assign ys__n29191 = new_n38322_ | new_n38323_;
  assign new_n38325_ = ~ys__n29121 & ys__n29192;
  assign new_n38326_ = ys__n29121 & ys__n29193;
  assign ys__n29194 = new_n38325_ | new_n38326_;
  assign new_n38328_ = ~ys__n29121 & ys__n29195;
  assign new_n38329_ = ys__n29121 & ys__n29196;
  assign ys__n29197 = new_n38328_ | new_n38329_;
  assign new_n38331_ = ~ys__n29121 & ys__n29198;
  assign new_n38332_ = ys__n29121 & ys__n29199;
  assign ys__n29200 = new_n38331_ | new_n38332_;
  assign new_n38334_ = ~ys__n29121 & ys__n29201;
  assign new_n38335_ = ys__n29121 & ys__n29202;
  assign ys__n29203 = new_n38334_ | new_n38335_;
  assign new_n38337_ = ~ys__n29121 & ys__n29204;
  assign new_n38338_ = ys__n29121 & ys__n29205;
  assign ys__n29206 = new_n38337_ | new_n38338_;
  assign new_n38340_ = ~ys__n29121 & ys__n29207;
  assign new_n38341_ = ys__n29121 & ys__n29208;
  assign ys__n29209 = new_n38340_ | new_n38341_;
  assign new_n38343_ = ~ys__n29121 & ys__n29210;
  assign new_n38344_ = ys__n29121 & ys__n29211;
  assign ys__n29212 = new_n38343_ | new_n38344_;
  assign new_n38346_ = ~ys__n29121 & ys__n29213;
  assign new_n38347_ = ys__n29121 & ys__n29214;
  assign ys__n29215 = new_n38346_ | new_n38347_;
  assign new_n38349_ = ~ys__n28243 & new_n22679_;
  assign new_n38350_ = new_n22695_ & new_n38349_;
  assign ys__n29217 = ~ys__n4566 & new_n38350_;
  assign ys__n29219 = ys__n29218 & ~ys__n4566;
  assign ys__n29221 = ys__n29220 & ~ys__n4566;
  assign new_n38354_ = new_n22676_ & new_n22695_;
  assign new_n38355_ = ~new_n22721_ & new_n22724_;
  assign new_n38356_ = ~new_n22695_ & new_n38355_;
  assign new_n38357_ = ~new_n38354_ & ~new_n38356_;
  assign new_n38358_ = ~ys__n28243 & ~ys__n4566;
  assign ys__n29223 = ~new_n38357_ & new_n38358_;
  assign ys__n29225 = ys__n29224 & ~ys__n4566;
  assign ys__n29226 = ys__n18114 & ~ys__n4566;
  assign ys__n29227 = ~ys__n28243 & ys__n23795;
  assign ys__n29228 = ~ys__n28243 & ys__n23798;
  assign ys__n29229 = ~ys__n28243 & ys__n23801;
  assign ys__n29230 = ~ys__n28243 & ys__n23804;
  assign ys__n29231 = ~ys__n28243 & ys__n23807;
  assign new_n38367_ = ~new_n38246_ & ~new_n38248_;
  assign ys__n29232 = ~ys__n28243 & ~new_n38367_;
  assign new_n38369_ = ~ys__n28243 & new_n22684_;
  assign new_n38370_ = new_n22695_ & new_n38369_;
  assign ys__n29233 = ~new_n22682_ & new_n38370_;
  assign new_n38372_ = new_n22672_ & new_n22695_;
  assign new_n38373_ = ~new_n22668_ & new_n38372_;
  assign new_n38374_ = ~new_n22717_ & new_n38248_;
  assign new_n38375_ = ~new_n38373_ & ~new_n38374_;
  assign ys__n29234 = ~ys__n28243 & ~new_n38375_;
  assign new_n38377_ = ~new_n22721_ & ~new_n38355_;
  assign new_n38378_ = ~ys__n28243 & ~new_n22695_;
  assign ys__n29235 = ~new_n38377_ & new_n38378_;
  assign new_n38380_ = ~ys__n4625 & ~ys__n38502;
  assign new_n38381_ = new_n13359_ & new_n38380_;
  assign new_n38382_ = ~new_n24254_ & new_n38381_;
  assign new_n38383_ = ~new_n23753_ & ~new_n37682_;
  assign new_n38384_ = ~new_n24250_ & ~new_n38383_;
  assign new_n38385_ = ~new_n38381_ & ~new_n38384_;
  assign new_n38386_ = ~new_n38382_ & ~new_n38385_;
  assign new_n38387_ = new_n13322_ & ~new_n38386_;
  assign new_n38388_ = ~ys__n740 & ~new_n13322_;
  assign new_n38389_ = ~new_n38386_ & new_n38388_;
  assign ys__n29336 = new_n38387_ | new_n38389_;
  assign new_n38391_ = ~new_n24273_ & new_n38381_;
  assign new_n38392_ = ~new_n23753_ & ~new_n37705_;
  assign new_n38393_ = ~new_n24269_ & ~new_n38392_;
  assign new_n38394_ = ~new_n38381_ & ~new_n38393_;
  assign new_n38395_ = ~new_n38391_ & ~new_n38394_;
  assign new_n38396_ = new_n13322_ & ~new_n38395_;
  assign new_n38397_ = new_n38388_ & ~new_n38395_;
  assign ys__n29339 = new_n38396_ | new_n38397_;
  assign new_n38399_ = ~new_n24292_ & new_n38381_;
  assign new_n38400_ = ~new_n23753_ & ~new_n37727_;
  assign new_n38401_ = ~new_n24288_ & ~new_n38400_;
  assign new_n38402_ = ~new_n38381_ & ~new_n38401_;
  assign new_n38403_ = ~new_n38399_ & ~new_n38402_;
  assign new_n38404_ = new_n13322_ & ~new_n38403_;
  assign new_n38405_ = new_n38388_ & ~new_n38403_;
  assign ys__n29342 = new_n38404_ | new_n38405_;
  assign new_n38407_ = ~new_n24311_ & new_n38381_;
  assign new_n38408_ = ~new_n23753_ & ~new_n37749_;
  assign new_n38409_ = ~new_n24307_ & ~new_n38408_;
  assign new_n38410_ = ~new_n38381_ & ~new_n38409_;
  assign new_n38411_ = ~new_n38407_ & ~new_n38410_;
  assign new_n38412_ = new_n13322_ & ~new_n38411_;
  assign new_n38413_ = new_n38388_ & ~new_n38411_;
  assign ys__n29345 = new_n38412_ | new_n38413_;
  assign new_n38415_ = ~new_n24330_ & new_n38381_;
  assign new_n38416_ = ~new_n23753_ & ~new_n37771_;
  assign new_n38417_ = ~new_n24326_ & ~new_n38416_;
  assign new_n38418_ = ~new_n38381_ & ~new_n38417_;
  assign new_n38419_ = ~new_n38415_ & ~new_n38418_;
  assign new_n38420_ = new_n13322_ & ~new_n38419_;
  assign new_n38421_ = new_n38388_ & ~new_n38419_;
  assign ys__n29348 = new_n38420_ | new_n38421_;
  assign new_n38423_ = ~new_n24349_ & new_n38381_;
  assign new_n38424_ = ~new_n23753_ & ~new_n37793_;
  assign new_n38425_ = ~new_n24345_ & ~new_n38424_;
  assign new_n38426_ = ~new_n38381_ & ~new_n38425_;
  assign new_n38427_ = ~new_n38423_ & ~new_n38426_;
  assign new_n38428_ = new_n13322_ & ~new_n38427_;
  assign new_n38429_ = new_n38388_ & ~new_n38427_;
  assign ys__n29351 = new_n38428_ | new_n38429_;
  assign new_n38431_ = ~new_n24368_ & new_n38381_;
  assign new_n38432_ = ~new_n23753_ & ~new_n37815_;
  assign new_n38433_ = ~new_n24364_ & ~new_n38432_;
  assign new_n38434_ = ~new_n38381_ & ~new_n38433_;
  assign new_n38435_ = ~new_n38431_ & ~new_n38434_;
  assign new_n38436_ = new_n13322_ & ~new_n38435_;
  assign new_n38437_ = new_n38388_ & ~new_n38435_;
  assign ys__n29354 = new_n38436_ | new_n38437_;
  assign new_n38439_ = ~new_n24387_ & new_n38381_;
  assign new_n38440_ = ~new_n23753_ & ~new_n37837_;
  assign new_n38441_ = ~new_n24383_ & ~new_n38440_;
  assign new_n38442_ = ~new_n38381_ & ~new_n38441_;
  assign new_n38443_ = ~new_n38439_ & ~new_n38442_;
  assign new_n38444_ = new_n13322_ & ~new_n38443_;
  assign new_n38445_ = new_n38388_ & ~new_n38443_;
  assign ys__n29357 = new_n38444_ | new_n38445_;
  assign new_n38447_ = ~new_n24068_ & new_n38381_;
  assign new_n38448_ = ~new_n23753_ & ~new_n37888_;
  assign new_n38449_ = ~new_n24064_ & ~new_n38448_;
  assign new_n38450_ = ~new_n38381_ & ~new_n38449_;
  assign new_n38451_ = ~new_n38447_ & ~new_n38450_;
  assign new_n38452_ = new_n13322_ & ~new_n38451_;
  assign new_n38453_ = new_n38388_ & ~new_n38451_;
  assign ys__n29360 = new_n38452_ | new_n38453_;
  assign new_n38455_ = ~new_n24086_ & new_n38381_;
  assign new_n38456_ = ~new_n23753_ & ~new_n37903_;
  assign new_n38457_ = ~new_n24082_ & ~new_n38456_;
  assign new_n38458_ = ~new_n38381_ & ~new_n38457_;
  assign new_n38459_ = ~new_n38455_ & ~new_n38458_;
  assign new_n38460_ = new_n13322_ & ~new_n38459_;
  assign new_n38461_ = new_n38388_ & ~new_n38459_;
  assign ys__n29363 = new_n38460_ | new_n38461_;
  assign new_n38463_ = ~new_n24104_ & new_n38381_;
  assign new_n38464_ = ~new_n23753_ & ~new_n37918_;
  assign new_n38465_ = ~new_n24100_ & ~new_n38464_;
  assign new_n38466_ = ~new_n38381_ & ~new_n38465_;
  assign new_n38467_ = ~new_n38463_ & ~new_n38466_;
  assign new_n38468_ = new_n13322_ & ~new_n38467_;
  assign new_n38469_ = new_n38388_ & ~new_n38467_;
  assign ys__n29366 = new_n38468_ | new_n38469_;
  assign new_n38471_ = ~new_n24122_ & new_n38381_;
  assign new_n38472_ = ~new_n23753_ & ~new_n37933_;
  assign new_n38473_ = ~new_n24118_ & ~new_n38472_;
  assign new_n38474_ = ~new_n38381_ & ~new_n38473_;
  assign new_n38475_ = ~new_n38471_ & ~new_n38474_;
  assign new_n38476_ = new_n13322_ & ~new_n38475_;
  assign new_n38477_ = new_n38388_ & ~new_n38475_;
  assign ys__n29369 = new_n38476_ | new_n38477_;
  assign new_n38479_ = ~new_n24140_ & new_n38381_;
  assign new_n38480_ = ~new_n23753_ & ~new_n37948_;
  assign new_n38481_ = ~new_n24136_ & ~new_n38480_;
  assign new_n38482_ = ~new_n38381_ & ~new_n38481_;
  assign new_n38483_ = ~new_n38479_ & ~new_n38482_;
  assign new_n38484_ = new_n13322_ & ~new_n38483_;
  assign new_n38485_ = new_n38388_ & ~new_n38483_;
  assign ys__n29372 = new_n38484_ | new_n38485_;
  assign new_n38487_ = ~new_n24158_ & new_n38381_;
  assign new_n38488_ = ~new_n23753_ & ~new_n37963_;
  assign new_n38489_ = ~new_n24154_ & ~new_n38488_;
  assign new_n38490_ = ~new_n38381_ & ~new_n38489_;
  assign new_n38491_ = ~new_n38487_ & ~new_n38490_;
  assign new_n38492_ = new_n13322_ & ~new_n38491_;
  assign new_n38493_ = new_n38388_ & ~new_n38491_;
  assign ys__n29375 = new_n38492_ | new_n38493_;
  assign new_n38495_ = ~new_n24176_ & new_n38381_;
  assign new_n38496_ = ~new_n23753_ & ~new_n37978_;
  assign new_n38497_ = ~new_n24172_ & ~new_n38496_;
  assign new_n38498_ = ~new_n38381_ & ~new_n38497_;
  assign new_n38499_ = ~new_n38495_ & ~new_n38498_;
  assign new_n38500_ = new_n13322_ & ~new_n38499_;
  assign new_n38501_ = new_n38388_ & ~new_n38499_;
  assign ys__n29378 = new_n38500_ | new_n38501_;
  assign new_n38503_ = ~new_n24194_ & new_n38381_;
  assign new_n38504_ = ~new_n23753_ & ~new_n37993_;
  assign new_n38505_ = ~new_n24190_ & ~new_n38504_;
  assign new_n38506_ = ~new_n38381_ & ~new_n38505_;
  assign new_n38507_ = ~new_n38503_ & ~new_n38506_;
  assign new_n38508_ = new_n13322_ & ~new_n38507_;
  assign new_n38509_ = new_n38388_ & ~new_n38507_;
  assign ys__n29381 = new_n38508_ | new_n38509_;
  assign new_n38511_ = ~new_n23908_ & new_n38381_;
  assign new_n38512_ = ~new_n23753_ & ~new_n38012_;
  assign new_n38513_ = ~new_n23904_ & ~new_n38512_;
  assign new_n38514_ = ~new_n38381_ & ~new_n38513_;
  assign new_n38515_ = ~new_n38511_ & ~new_n38514_;
  assign new_n38516_ = new_n13322_ & ~new_n38515_;
  assign new_n38517_ = new_n38388_ & ~new_n38515_;
  assign ys__n29384 = new_n38516_ | new_n38517_;
  assign new_n38519_ = ~new_n23923_ & new_n38381_;
  assign new_n38520_ = ~new_n23753_ & ~new_n38027_;
  assign new_n38521_ = ~new_n23919_ & ~new_n38520_;
  assign new_n38522_ = ~new_n38381_ & ~new_n38521_;
  assign new_n38523_ = ~new_n38519_ & ~new_n38522_;
  assign new_n38524_ = new_n13322_ & ~new_n38523_;
  assign new_n38525_ = new_n38388_ & ~new_n38523_;
  assign ys__n29387 = new_n38524_ | new_n38525_;
  assign new_n38527_ = ~new_n23938_ & new_n38381_;
  assign new_n38528_ = ~new_n23753_ & ~new_n38042_;
  assign new_n38529_ = ~new_n23934_ & ~new_n38528_;
  assign new_n38530_ = ~new_n38381_ & ~new_n38529_;
  assign new_n38531_ = ~new_n38527_ & ~new_n38530_;
  assign new_n38532_ = new_n13322_ & ~new_n38531_;
  assign new_n38533_ = new_n38388_ & ~new_n38531_;
  assign ys__n29390 = new_n38532_ | new_n38533_;
  assign new_n38535_ = ~new_n23953_ & new_n38381_;
  assign new_n38536_ = ~new_n23753_ & ~new_n38057_;
  assign new_n38537_ = ~new_n23949_ & ~new_n38536_;
  assign new_n38538_ = ~new_n38381_ & ~new_n38537_;
  assign new_n38539_ = ~new_n38535_ & ~new_n38538_;
  assign new_n38540_ = new_n13322_ & ~new_n38539_;
  assign new_n38541_ = new_n38388_ & ~new_n38539_;
  assign ys__n29393 = new_n38540_ | new_n38541_;
  assign new_n38543_ = ~new_n23968_ & new_n38381_;
  assign new_n38544_ = ~new_n23753_ & ~new_n38072_;
  assign new_n38545_ = ~new_n23964_ & ~new_n38544_;
  assign new_n38546_ = ~new_n38381_ & ~new_n38545_;
  assign new_n38547_ = ~new_n38543_ & ~new_n38546_;
  assign new_n38548_ = new_n13322_ & ~new_n38547_;
  assign new_n38549_ = new_n38388_ & ~new_n38547_;
  assign ys__n29396 = new_n38548_ | new_n38549_;
  assign new_n38551_ = ~new_n23983_ & new_n38381_;
  assign new_n38552_ = ~new_n23753_ & ~new_n38087_;
  assign new_n38553_ = ~new_n23979_ & ~new_n38552_;
  assign new_n38554_ = ~new_n38381_ & ~new_n38553_;
  assign new_n38555_ = ~new_n38551_ & ~new_n38554_;
  assign new_n38556_ = new_n13322_ & ~new_n38555_;
  assign new_n38557_ = new_n38388_ & ~new_n38555_;
  assign ys__n29399 = new_n38556_ | new_n38557_;
  assign new_n38559_ = ~new_n23998_ & new_n38381_;
  assign new_n38560_ = ~new_n23753_ & ~new_n38102_;
  assign new_n38561_ = ~new_n23994_ & ~new_n38560_;
  assign new_n38562_ = ~new_n38381_ & ~new_n38561_;
  assign new_n38563_ = ~new_n38559_ & ~new_n38562_;
  assign new_n38564_ = new_n13322_ & ~new_n38563_;
  assign new_n38565_ = new_n38388_ & ~new_n38563_;
  assign ys__n29402 = new_n38564_ | new_n38565_;
  assign new_n38567_ = ~new_n24013_ & new_n38381_;
  assign new_n38568_ = ~new_n23753_ & ~new_n38117_;
  assign new_n38569_ = ~new_n24009_ & ~new_n38568_;
  assign new_n38570_ = ~new_n38381_ & ~new_n38569_;
  assign new_n38571_ = ~new_n38567_ & ~new_n38570_;
  assign new_n38572_ = new_n13322_ & ~new_n38571_;
  assign new_n38573_ = new_n38388_ & ~new_n38571_;
  assign ys__n29405 = new_n38572_ | new_n38573_;
  assign new_n38575_ = ~new_n23760_ & new_n38381_;
  assign new_n38576_ = ~new_n23753_ & ~new_n38132_;
  assign new_n38577_ = ~new_n23754_ & ~new_n38576_;
  assign new_n38578_ = ~new_n38381_ & ~new_n38577_;
  assign new_n38579_ = ~new_n38575_ & ~new_n38578_;
  assign new_n38580_ = new_n13322_ & ~new_n38579_;
  assign new_n38581_ = new_n38388_ & ~new_n38579_;
  assign ys__n29408 = new_n38580_ | new_n38581_;
  assign new_n38583_ = ~new_n23775_ & new_n38381_;
  assign new_n38584_ = ~new_n23753_ & ~new_n38147_;
  assign new_n38585_ = ~new_n23771_ & ~new_n38584_;
  assign new_n38586_ = ~new_n38381_ & ~new_n38585_;
  assign new_n38587_ = ~new_n38583_ & ~new_n38586_;
  assign new_n38588_ = new_n13322_ & ~new_n38587_;
  assign new_n38589_ = new_n38388_ & ~new_n38587_;
  assign ys__n29411 = new_n38588_ | new_n38589_;
  assign new_n38591_ = ~new_n23790_ & new_n38381_;
  assign new_n38592_ = ~new_n23753_ & ~new_n38162_;
  assign new_n38593_ = ~new_n23786_ & ~new_n38592_;
  assign new_n38594_ = ~new_n38381_ & ~new_n38593_;
  assign new_n38595_ = ~new_n38591_ & ~new_n38594_;
  assign new_n38596_ = new_n13322_ & ~new_n38595_;
  assign new_n38597_ = new_n38388_ & ~new_n38595_;
  assign ys__n29414 = new_n38596_ | new_n38597_;
  assign new_n38599_ = ~new_n23805_ & new_n38381_;
  assign new_n38600_ = ~new_n23753_ & ~new_n38177_;
  assign new_n38601_ = ~new_n23801_ & ~new_n38600_;
  assign new_n38602_ = ~new_n38381_ & ~new_n38601_;
  assign new_n38603_ = ~new_n38599_ & ~new_n38602_;
  assign new_n38604_ = new_n13322_ & ~new_n38603_;
  assign new_n38605_ = new_n38388_ & ~new_n38603_;
  assign ys__n29417 = new_n38604_ | new_n38605_;
  assign new_n38607_ = ~new_n23820_ & new_n38381_;
  assign new_n38608_ = ~new_n23753_ & ~new_n38192_;
  assign new_n38609_ = ~new_n23816_ & ~new_n38608_;
  assign new_n38610_ = ~new_n38381_ & ~new_n38609_;
  assign new_n38611_ = ~new_n38607_ & ~new_n38610_;
  assign new_n38612_ = new_n13322_ & ~new_n38611_;
  assign new_n38613_ = new_n38388_ & ~new_n38611_;
  assign ys__n29420 = new_n38612_ | new_n38613_;
  assign new_n38615_ = ~new_n23835_ & new_n38381_;
  assign new_n38616_ = ~new_n23753_ & ~new_n38207_;
  assign new_n38617_ = ~new_n23831_ & ~new_n38616_;
  assign new_n38618_ = ~new_n38381_ & ~new_n38617_;
  assign new_n38619_ = ~new_n38615_ & ~new_n38618_;
  assign new_n38620_ = new_n13322_ & ~new_n38619_;
  assign new_n38621_ = new_n38388_ & ~new_n38619_;
  assign ys__n29423 = new_n38620_ | new_n38621_;
  assign new_n38623_ = ~new_n23850_ & new_n38381_;
  assign new_n38624_ = ~new_n23753_ & ~new_n38222_;
  assign new_n38625_ = ~new_n23846_ & ~new_n38624_;
  assign new_n38626_ = ~new_n38381_ & ~new_n38625_;
  assign new_n38627_ = ~new_n38623_ & ~new_n38626_;
  assign new_n38628_ = new_n13322_ & ~new_n38627_;
  assign new_n38629_ = new_n38388_ & ~new_n38627_;
  assign ys__n29426 = new_n38628_ | new_n38629_;
  assign new_n38631_ = ~new_n23865_ & new_n38381_;
  assign new_n38632_ = ~new_n23753_ & ~new_n38237_;
  assign new_n38633_ = ~new_n23861_ & ~new_n38632_;
  assign new_n38634_ = ~new_n38381_ & ~new_n38633_;
  assign new_n38635_ = ~new_n38631_ & ~new_n38634_;
  assign new_n38636_ = new_n13322_ & ~new_n38635_;
  assign new_n38637_ = new_n38388_ & ~new_n38635_;
  assign ys__n29429 = new_n38636_ | new_n38637_;
  assign new_n38639_ = new_n22829_ & new_n22831_;
  assign new_n38640_ = new_n22815_ & new_n22819_;
  assign new_n38641_ = ~new_n38639_ & ~new_n38640_;
  assign new_n38642_ = ~new_n22836_ & new_n22842_;
  assign new_n38643_ = ~new_n38641_ & new_n38642_;
  assign new_n38644_ = ~new_n22842_ & new_n22868_;
  assign new_n38645_ = new_n22864_ & new_n38644_;
  assign new_n38646_ = ~new_n38643_ & ~new_n38645_;
  assign ys__n29431 = new_n38251_ & ~new_n38646_;
  assign new_n38648_ = ys__n29432 & ~ys__n29434;
  assign new_n38649_ = ys__n29433 & ys__n29434;
  assign ys__n29435 = new_n38648_ | new_n38649_;
  assign new_n38651_ = ~ys__n29434 & ys__n29436;
  assign new_n38652_ = ys__n29434 & ys__n29437;
  assign ys__n29438 = new_n38651_ | new_n38652_;
  assign new_n38654_ = ~ys__n29434 & ys__n29439;
  assign new_n38655_ = ys__n29434 & ys__n29440;
  assign ys__n29441 = new_n38654_ | new_n38655_;
  assign new_n38657_ = ~ys__n29434 & ys__n29442;
  assign new_n38658_ = ys__n29434 & ys__n29443;
  assign ys__n29444 = new_n38657_ | new_n38658_;
  assign new_n38660_ = ~ys__n29434 & ys__n29445;
  assign new_n38661_ = ys__n29434 & ys__n29446;
  assign ys__n29447 = new_n38660_ | new_n38661_;
  assign new_n38663_ = ~ys__n29434 & ys__n29448;
  assign new_n38664_ = ys__n29434 & ys__n29449;
  assign ys__n29450 = new_n38663_ | new_n38664_;
  assign new_n38666_ = ~ys__n29434 & ys__n29451;
  assign new_n38667_ = ys__n29434 & ys__n29452;
  assign ys__n29453 = new_n38666_ | new_n38667_;
  assign new_n38669_ = ~ys__n29434 & ys__n29454;
  assign new_n38670_ = ys__n29434 & ys__n29455;
  assign ys__n29456 = new_n38669_ | new_n38670_;
  assign new_n38672_ = ~ys__n29434 & ys__n29457;
  assign new_n38673_ = ys__n29434 & ys__n29458;
  assign ys__n29459 = new_n38672_ | new_n38673_;
  assign new_n38675_ = ~ys__n29434 & ys__n29460;
  assign new_n38676_ = ys__n29434 & ys__n29461;
  assign ys__n29462 = new_n38675_ | new_n38676_;
  assign new_n38678_ = ~ys__n29434 & ys__n29463;
  assign new_n38679_ = ys__n29434 & ys__n29464;
  assign ys__n29465 = new_n38678_ | new_n38679_;
  assign new_n38681_ = ~ys__n29434 & ys__n29466;
  assign new_n38682_ = ys__n29434 & ys__n29467;
  assign ys__n29468 = new_n38681_ | new_n38682_;
  assign new_n38684_ = ~ys__n29434 & ys__n29469;
  assign new_n38685_ = ys__n29434 & ys__n29470;
  assign ys__n29471 = new_n38684_ | new_n38685_;
  assign new_n38687_ = ~ys__n29434 & ys__n29472;
  assign new_n38688_ = ys__n29434 & ys__n29473;
  assign ys__n29474 = new_n38687_ | new_n38688_;
  assign new_n38690_ = ~ys__n29434 & ys__n29475;
  assign new_n38691_ = ys__n29434 & ys__n29476;
  assign ys__n29477 = new_n38690_ | new_n38691_;
  assign new_n38693_ = ~ys__n29434 & ys__n29478;
  assign new_n38694_ = ys__n29434 & ys__n29479;
  assign ys__n29480 = new_n38693_ | new_n38694_;
  assign new_n38696_ = ~ys__n29434 & ys__n29481;
  assign new_n38697_ = ys__n29434 & ys__n29482;
  assign ys__n29483 = new_n38696_ | new_n38697_;
  assign new_n38699_ = ~ys__n29434 & ys__n29484;
  assign new_n38700_ = ys__n29434 & ys__n29485;
  assign ys__n29486 = new_n38699_ | new_n38700_;
  assign new_n38702_ = ~ys__n29434 & ys__n29487;
  assign new_n38703_ = ys__n29434 & ys__n29488;
  assign ys__n29489 = new_n38702_ | new_n38703_;
  assign new_n38705_ = ~ys__n29434 & ys__n29490;
  assign new_n38706_ = ys__n29434 & ys__n29491;
  assign ys__n29492 = new_n38705_ | new_n38706_;
  assign new_n38708_ = ~ys__n29434 & ys__n29493;
  assign new_n38709_ = ys__n29434 & ys__n29494;
  assign ys__n29495 = new_n38708_ | new_n38709_;
  assign new_n38711_ = ~ys__n29434 & ys__n29496;
  assign new_n38712_ = ys__n29434 & ys__n29497;
  assign ys__n29498 = new_n38711_ | new_n38712_;
  assign new_n38714_ = ~ys__n29434 & ys__n29499;
  assign new_n38715_ = ys__n29434 & ys__n29500;
  assign ys__n29501 = new_n38714_ | new_n38715_;
  assign new_n38717_ = ~ys__n29434 & ys__n29502;
  assign new_n38718_ = ys__n29434 & ys__n29503;
  assign ys__n29504 = new_n38717_ | new_n38718_;
  assign new_n38720_ = ~ys__n29434 & ys__n29505;
  assign new_n38721_ = ys__n29434 & ys__n29506;
  assign ys__n29507 = new_n38720_ | new_n38721_;
  assign new_n38723_ = ~ys__n29434 & ys__n29508;
  assign new_n38724_ = ys__n29434 & ys__n29509;
  assign ys__n29510 = new_n38723_ | new_n38724_;
  assign new_n38726_ = ~ys__n29434 & ys__n29511;
  assign new_n38727_ = ys__n29434 & ys__n29512;
  assign ys__n29513 = new_n38726_ | new_n38727_;
  assign new_n38729_ = ~ys__n29434 & ys__n29514;
  assign new_n38730_ = ys__n29434 & ys__n29515;
  assign ys__n29516 = new_n38729_ | new_n38730_;
  assign new_n38732_ = ~ys__n29434 & ys__n29517;
  assign new_n38733_ = ys__n29434 & ys__n29518;
  assign ys__n29519 = new_n38732_ | new_n38733_;
  assign new_n38735_ = ~ys__n29434 & ys__n29520;
  assign new_n38736_ = ys__n29434 & ys__n29521;
  assign ys__n29522 = new_n38735_ | new_n38736_;
  assign new_n38738_ = ~ys__n29434 & ys__n29523;
  assign new_n38739_ = ys__n29434 & ys__n29524;
  assign ys__n29525 = new_n38738_ | new_n38739_;
  assign new_n38741_ = ~ys__n29434 & ys__n29526;
  assign new_n38742_ = ys__n29434 & ys__n29527;
  assign ys__n29528 = new_n38741_ | new_n38742_;
  assign new_n38744_ = ~ys__n28243 & new_n22826_;
  assign new_n38745_ = new_n22842_ & new_n38744_;
  assign ys__n29530 = ~ys__n4566 & new_n38745_;
  assign ys__n29532 = ys__n29531 & ~ys__n4566;
  assign ys__n29534 = ys__n29533 & ~ys__n4566;
  assign new_n38749_ = new_n22823_ & new_n22842_;
  assign new_n38750_ = ~new_n22868_ & new_n22871_;
  assign new_n38751_ = ~new_n22842_ & new_n38750_;
  assign new_n38752_ = ~new_n38749_ & ~new_n38751_;
  assign ys__n29536 = new_n38358_ & ~new_n38752_;
  assign ys__n29538 = ys__n29537 & ~ys__n4566;
  assign ys__n29539 = ys__n18116 & ~ys__n4566;
  assign ys__n29540 = ~ys__n28243 & ys__n23865;
  assign ys__n29541 = ~ys__n28243 & ys__n23868;
  assign ys__n29542 = ~ys__n28243 & ys__n23871;
  assign ys__n29543 = ~ys__n28243 & ys__n23874;
  assign ys__n29544 = ~ys__n28243 & ys__n23877;
  assign new_n38761_ = ~new_n38642_ & ~new_n38644_;
  assign ys__n29545 = ~ys__n28243 & ~new_n38761_;
  assign new_n38763_ = ~ys__n28243 & new_n22831_;
  assign new_n38764_ = new_n22842_ & new_n38763_;
  assign ys__n29546 = ~new_n22829_ & new_n38764_;
  assign new_n38766_ = new_n22819_ & new_n22842_;
  assign new_n38767_ = ~new_n22815_ & new_n38766_;
  assign new_n38768_ = ~new_n22864_ & new_n38644_;
  assign new_n38769_ = ~new_n38767_ & ~new_n38768_;
  assign ys__n29547 = ~ys__n28243 & ~new_n38769_;
  assign new_n38771_ = ~new_n22868_ & ~new_n38750_;
  assign new_n38772_ = ~ys__n28243 & ~new_n22842_;
  assign ys__n29548 = ~new_n38771_ & new_n38772_;
  assign new_n38774_ = ~ys__n4625 & ~ys__n38513;
  assign new_n38775_ = new_n13359_ & new_n38774_;
  assign new_n38776_ = ys__n28462 & new_n38775_;
  assign new_n38777_ = ~new_n23755_ & ~new_n38384_;
  assign new_n38778_ = ~new_n24251_ & ~new_n38777_;
  assign new_n38779_ = ~new_n38775_ & ~new_n38778_;
  assign new_n38780_ = ~new_n38776_ & ~new_n38779_;
  assign new_n38781_ = new_n13311_ & ~new_n38780_;
  assign new_n38782_ = ~ys__n740 & ~new_n13311_;
  assign new_n38783_ = ~new_n38780_ & new_n38782_;
  assign ys__n29611 = new_n38781_ | new_n38783_;
  assign new_n38785_ = ys__n28464 & new_n38775_;
  assign new_n38786_ = ~new_n23755_ & ~new_n38393_;
  assign new_n38787_ = ~new_n24270_ & ~new_n38786_;
  assign new_n38788_ = ~new_n38775_ & ~new_n38787_;
  assign new_n38789_ = ~new_n38785_ & ~new_n38788_;
  assign new_n38790_ = new_n13311_ & ~new_n38789_;
  assign new_n38791_ = new_n38782_ & ~new_n38789_;
  assign ys__n29614 = new_n38790_ | new_n38791_;
  assign new_n38793_ = ys__n28466 & new_n38775_;
  assign new_n38794_ = ~new_n23755_ & ~new_n38401_;
  assign new_n38795_ = ~new_n24289_ & ~new_n38794_;
  assign new_n38796_ = ~new_n38775_ & ~new_n38795_;
  assign new_n38797_ = ~new_n38793_ & ~new_n38796_;
  assign new_n38798_ = new_n13311_ & ~new_n38797_;
  assign new_n38799_ = new_n38782_ & ~new_n38797_;
  assign ys__n29617 = new_n38798_ | new_n38799_;
  assign new_n38801_ = ys__n28468 & new_n38775_;
  assign new_n38802_ = ~new_n23755_ & ~new_n38409_;
  assign new_n38803_ = ~new_n24308_ & ~new_n38802_;
  assign new_n38804_ = ~new_n38775_ & ~new_n38803_;
  assign new_n38805_ = ~new_n38801_ & ~new_n38804_;
  assign new_n38806_ = new_n13311_ & ~new_n38805_;
  assign new_n38807_ = new_n38782_ & ~new_n38805_;
  assign ys__n29620 = new_n38806_ | new_n38807_;
  assign new_n38809_ = ys__n28470 & new_n38775_;
  assign new_n38810_ = ~new_n23755_ & ~new_n38417_;
  assign new_n38811_ = ~new_n24327_ & ~new_n38810_;
  assign new_n38812_ = ~new_n38775_ & ~new_n38811_;
  assign new_n38813_ = ~new_n38809_ & ~new_n38812_;
  assign new_n38814_ = new_n13311_ & ~new_n38813_;
  assign new_n38815_ = new_n38782_ & ~new_n38813_;
  assign ys__n29623 = new_n38814_ | new_n38815_;
  assign new_n38817_ = ys__n28472 & new_n38775_;
  assign new_n38818_ = ~new_n23755_ & ~new_n38425_;
  assign new_n38819_ = ~new_n24346_ & ~new_n38818_;
  assign new_n38820_ = ~new_n38775_ & ~new_n38819_;
  assign new_n38821_ = ~new_n38817_ & ~new_n38820_;
  assign new_n38822_ = new_n13311_ & ~new_n38821_;
  assign new_n38823_ = new_n38782_ & ~new_n38821_;
  assign ys__n29626 = new_n38822_ | new_n38823_;
  assign new_n38825_ = ys__n29558 & new_n38775_;
  assign new_n38826_ = ~new_n23755_ & ~new_n38433_;
  assign new_n38827_ = ~new_n24365_ & ~new_n38826_;
  assign new_n38828_ = ~new_n38775_ & ~new_n38827_;
  assign new_n38829_ = ~new_n38825_ & ~new_n38828_;
  assign new_n38830_ = new_n13311_ & ~new_n38829_;
  assign new_n38831_ = new_n38782_ & ~new_n38829_;
  assign ys__n29629 = new_n38830_ | new_n38831_;
  assign new_n38833_ = ys__n29560 & new_n38775_;
  assign new_n38834_ = ~new_n23755_ & ~new_n38441_;
  assign new_n38835_ = ~new_n24384_ & ~new_n38834_;
  assign new_n38836_ = ~new_n38775_ & ~new_n38835_;
  assign new_n38837_ = ~new_n38833_ & ~new_n38836_;
  assign new_n38838_ = new_n13311_ & ~new_n38837_;
  assign new_n38839_ = new_n38782_ & ~new_n38837_;
  assign ys__n29632 = new_n38838_ | new_n38839_;
  assign new_n38841_ = ys__n29562 & new_n38775_;
  assign new_n38842_ = ~new_n23755_ & ~new_n38449_;
  assign new_n38843_ = ~new_n24065_ & ~new_n38842_;
  assign new_n38844_ = ~new_n38775_ & ~new_n38843_;
  assign new_n38845_ = ~new_n38841_ & ~new_n38844_;
  assign new_n38846_ = new_n13311_ & ~new_n38845_;
  assign new_n38847_ = new_n38782_ & ~new_n38845_;
  assign ys__n29635 = new_n38846_ | new_n38847_;
  assign new_n38849_ = ys__n29564 & new_n38775_;
  assign new_n38850_ = ~new_n23755_ & ~new_n38457_;
  assign new_n38851_ = ~new_n24083_ & ~new_n38850_;
  assign new_n38852_ = ~new_n38775_ & ~new_n38851_;
  assign new_n38853_ = ~new_n38849_ & ~new_n38852_;
  assign new_n38854_ = new_n13311_ & ~new_n38853_;
  assign new_n38855_ = new_n38782_ & ~new_n38853_;
  assign ys__n29638 = new_n38854_ | new_n38855_;
  assign new_n38857_ = ys__n29566 & new_n38775_;
  assign new_n38858_ = ~new_n23755_ & ~new_n38465_;
  assign new_n38859_ = ~new_n24101_ & ~new_n38858_;
  assign new_n38860_ = ~new_n38775_ & ~new_n38859_;
  assign new_n38861_ = ~new_n38857_ & ~new_n38860_;
  assign new_n38862_ = new_n13311_ & ~new_n38861_;
  assign new_n38863_ = new_n38782_ & ~new_n38861_;
  assign ys__n29641 = new_n38862_ | new_n38863_;
  assign new_n38865_ = ys__n29568 & new_n38775_;
  assign new_n38866_ = ~new_n23755_ & ~new_n38473_;
  assign new_n38867_ = ~new_n24119_ & ~new_n38866_;
  assign new_n38868_ = ~new_n38775_ & ~new_n38867_;
  assign new_n38869_ = ~new_n38865_ & ~new_n38868_;
  assign new_n38870_ = new_n13311_ & ~new_n38869_;
  assign new_n38871_ = new_n38782_ & ~new_n38869_;
  assign ys__n29644 = new_n38870_ | new_n38871_;
  assign new_n38873_ = ys__n29570 & new_n38775_;
  assign new_n38874_ = ~new_n23755_ & ~new_n38481_;
  assign new_n38875_ = ~new_n24137_ & ~new_n38874_;
  assign new_n38876_ = ~new_n38775_ & ~new_n38875_;
  assign new_n38877_ = ~new_n38873_ & ~new_n38876_;
  assign new_n38878_ = new_n13311_ & ~new_n38877_;
  assign new_n38879_ = new_n38782_ & ~new_n38877_;
  assign ys__n29647 = new_n38878_ | new_n38879_;
  assign new_n38881_ = ys__n29572 & new_n38775_;
  assign new_n38882_ = ~new_n23755_ & ~new_n38489_;
  assign new_n38883_ = ~new_n24155_ & ~new_n38882_;
  assign new_n38884_ = ~new_n38775_ & ~new_n38883_;
  assign new_n38885_ = ~new_n38881_ & ~new_n38884_;
  assign new_n38886_ = new_n13311_ & ~new_n38885_;
  assign new_n38887_ = new_n38782_ & ~new_n38885_;
  assign ys__n29650 = new_n38886_ | new_n38887_;
  assign new_n38889_ = ys__n29574 & new_n38775_;
  assign new_n38890_ = ~new_n23755_ & ~new_n38497_;
  assign new_n38891_ = ~new_n24173_ & ~new_n38890_;
  assign new_n38892_ = ~new_n38775_ & ~new_n38891_;
  assign new_n38893_ = ~new_n38889_ & ~new_n38892_;
  assign new_n38894_ = new_n13311_ & ~new_n38893_;
  assign new_n38895_ = new_n38782_ & ~new_n38893_;
  assign ys__n29653 = new_n38894_ | new_n38895_;
  assign new_n38897_ = ys__n29576 & new_n38775_;
  assign new_n38898_ = ~new_n23755_ & ~new_n38505_;
  assign new_n38899_ = ~new_n24191_ & ~new_n38898_;
  assign new_n38900_ = ~new_n38775_ & ~new_n38899_;
  assign new_n38901_ = ~new_n38897_ & ~new_n38900_;
  assign new_n38902_ = new_n13311_ & ~new_n38901_;
  assign new_n38903_ = new_n38782_ & ~new_n38901_;
  assign ys__n29656 = new_n38902_ | new_n38903_;
  assign new_n38905_ = ys__n29578 & new_n38775_;
  assign new_n38906_ = ~new_n23755_ & ~new_n38513_;
  assign new_n38907_ = ~new_n23905_ & ~new_n38906_;
  assign new_n38908_ = ~new_n38775_ & ~new_n38907_;
  assign new_n38909_ = ~new_n38905_ & ~new_n38908_;
  assign new_n38910_ = new_n13311_ & ~new_n38909_;
  assign new_n38911_ = new_n38782_ & ~new_n38909_;
  assign ys__n29659 = new_n38910_ | new_n38911_;
  assign new_n38913_ = ys__n29580 & new_n38775_;
  assign new_n38914_ = ~new_n23755_ & ~new_n38521_;
  assign new_n38915_ = ~new_n23920_ & ~new_n38914_;
  assign new_n38916_ = ~new_n38775_ & ~new_n38915_;
  assign new_n38917_ = ~new_n38913_ & ~new_n38916_;
  assign new_n38918_ = new_n13311_ & ~new_n38917_;
  assign new_n38919_ = new_n38782_ & ~new_n38917_;
  assign ys__n29662 = new_n38918_ | new_n38919_;
  assign new_n38921_ = ys__n29582 & new_n38775_;
  assign new_n38922_ = ~new_n23755_ & ~new_n38529_;
  assign new_n38923_ = ~new_n23935_ & ~new_n38922_;
  assign new_n38924_ = ~new_n38775_ & ~new_n38923_;
  assign new_n38925_ = ~new_n38921_ & ~new_n38924_;
  assign new_n38926_ = new_n13311_ & ~new_n38925_;
  assign new_n38927_ = new_n38782_ & ~new_n38925_;
  assign ys__n29665 = new_n38926_ | new_n38927_;
  assign new_n38929_ = ys__n29584 & new_n38775_;
  assign new_n38930_ = ~new_n23755_ & ~new_n38537_;
  assign new_n38931_ = ~new_n23950_ & ~new_n38930_;
  assign new_n38932_ = ~new_n38775_ & ~new_n38931_;
  assign new_n38933_ = ~new_n38929_ & ~new_n38932_;
  assign new_n38934_ = new_n13311_ & ~new_n38933_;
  assign new_n38935_ = new_n38782_ & ~new_n38933_;
  assign ys__n29668 = new_n38934_ | new_n38935_;
  assign new_n38937_ = ys__n29586 & new_n38775_;
  assign new_n38938_ = ~new_n23755_ & ~new_n38545_;
  assign new_n38939_ = ~new_n23965_ & ~new_n38938_;
  assign new_n38940_ = ~new_n38775_ & ~new_n38939_;
  assign new_n38941_ = ~new_n38937_ & ~new_n38940_;
  assign new_n38942_ = new_n13311_ & ~new_n38941_;
  assign new_n38943_ = new_n38782_ & ~new_n38941_;
  assign ys__n29671 = new_n38942_ | new_n38943_;
  assign new_n38945_ = ys__n29588 & new_n38775_;
  assign new_n38946_ = ~new_n23755_ & ~new_n38553_;
  assign new_n38947_ = ~new_n23980_ & ~new_n38946_;
  assign new_n38948_ = ~new_n38775_ & ~new_n38947_;
  assign new_n38949_ = ~new_n38945_ & ~new_n38948_;
  assign new_n38950_ = new_n13311_ & ~new_n38949_;
  assign new_n38951_ = new_n38782_ & ~new_n38949_;
  assign ys__n29674 = new_n38950_ | new_n38951_;
  assign new_n38953_ = ys__n29590 & new_n38775_;
  assign new_n38954_ = ~new_n23755_ & ~new_n38561_;
  assign new_n38955_ = ~new_n23995_ & ~new_n38954_;
  assign new_n38956_ = ~new_n38775_ & ~new_n38955_;
  assign new_n38957_ = ~new_n38953_ & ~new_n38956_;
  assign new_n38958_ = new_n13311_ & ~new_n38957_;
  assign new_n38959_ = new_n38782_ & ~new_n38957_;
  assign ys__n29677 = new_n38958_ | new_n38959_;
  assign new_n38961_ = ys__n29592 & new_n38775_;
  assign new_n38962_ = ~new_n23755_ & ~new_n38569_;
  assign new_n38963_ = ~new_n24010_ & ~new_n38962_;
  assign new_n38964_ = ~new_n38775_ & ~new_n38963_;
  assign new_n38965_ = ~new_n38961_ & ~new_n38964_;
  assign new_n38966_ = new_n13311_ & ~new_n38965_;
  assign new_n38967_ = new_n38782_ & ~new_n38965_;
  assign ys__n29680 = new_n38966_ | new_n38967_;
  assign new_n38969_ = ys__n29594 & new_n38775_;
  assign new_n38970_ = ~new_n23755_ & ~new_n38577_;
  assign new_n38971_ = ~new_n23756_ & ~new_n38970_;
  assign new_n38972_ = ~new_n38775_ & ~new_n38971_;
  assign new_n38973_ = ~new_n38969_ & ~new_n38972_;
  assign new_n38974_ = new_n13311_ & ~new_n38973_;
  assign new_n38975_ = new_n38782_ & ~new_n38973_;
  assign ys__n29683 = new_n38974_ | new_n38975_;
  assign new_n38977_ = ys__n29596 & new_n38775_;
  assign new_n38978_ = ~new_n23755_ & ~new_n38585_;
  assign new_n38979_ = ~new_n23772_ & ~new_n38978_;
  assign new_n38980_ = ~new_n38775_ & ~new_n38979_;
  assign new_n38981_ = ~new_n38977_ & ~new_n38980_;
  assign new_n38982_ = new_n13311_ & ~new_n38981_;
  assign new_n38983_ = new_n38782_ & ~new_n38981_;
  assign ys__n29686 = new_n38982_ | new_n38983_;
  assign new_n38985_ = ys__n29598 & new_n38775_;
  assign new_n38986_ = ~new_n23755_ & ~new_n38593_;
  assign new_n38987_ = ~new_n23787_ & ~new_n38986_;
  assign new_n38988_ = ~new_n38775_ & ~new_n38987_;
  assign new_n38989_ = ~new_n38985_ & ~new_n38988_;
  assign new_n38990_ = new_n13311_ & ~new_n38989_;
  assign new_n38991_ = new_n38782_ & ~new_n38989_;
  assign ys__n29689 = new_n38990_ | new_n38991_;
  assign new_n38993_ = ys__n29600 & new_n38775_;
  assign new_n38994_ = ~new_n23755_ & ~new_n38601_;
  assign new_n38995_ = ~new_n23802_ & ~new_n38994_;
  assign new_n38996_ = ~new_n38775_ & ~new_n38995_;
  assign new_n38997_ = ~new_n38993_ & ~new_n38996_;
  assign new_n38998_ = new_n13311_ & ~new_n38997_;
  assign new_n38999_ = new_n38782_ & ~new_n38997_;
  assign ys__n29692 = new_n38998_ | new_n38999_;
  assign new_n39001_ = ys__n29602 & new_n38775_;
  assign new_n39002_ = ~new_n23755_ & ~new_n38609_;
  assign new_n39003_ = ~new_n23817_ & ~new_n39002_;
  assign new_n39004_ = ~new_n38775_ & ~new_n39003_;
  assign new_n39005_ = ~new_n39001_ & ~new_n39004_;
  assign new_n39006_ = new_n13311_ & ~new_n39005_;
  assign new_n39007_ = new_n38782_ & ~new_n39005_;
  assign ys__n29695 = new_n39006_ | new_n39007_;
  assign new_n39009_ = ys__n29604 & new_n38775_;
  assign new_n39010_ = ~new_n23755_ & ~new_n38617_;
  assign new_n39011_ = ~new_n23832_ & ~new_n39010_;
  assign new_n39012_ = ~new_n38775_ & ~new_n39011_;
  assign new_n39013_ = ~new_n39009_ & ~new_n39012_;
  assign new_n39014_ = new_n13311_ & ~new_n39013_;
  assign new_n39015_ = new_n38782_ & ~new_n39013_;
  assign ys__n29698 = new_n39014_ | new_n39015_;
  assign new_n39017_ = ys__n29606 & new_n38775_;
  assign new_n39018_ = ~new_n23755_ & ~new_n38625_;
  assign new_n39019_ = ~new_n23847_ & ~new_n39018_;
  assign new_n39020_ = ~new_n38775_ & ~new_n39019_;
  assign new_n39021_ = ~new_n39017_ & ~new_n39020_;
  assign new_n39022_ = new_n13311_ & ~new_n39021_;
  assign new_n39023_ = new_n38782_ & ~new_n39021_;
  assign ys__n29701 = new_n39022_ | new_n39023_;
  assign new_n39025_ = ys__n29608 & new_n38775_;
  assign new_n39026_ = ~new_n23755_ & ~new_n38633_;
  assign new_n39027_ = ~new_n23862_ & ~new_n39026_;
  assign new_n39028_ = ~new_n38775_ & ~new_n39027_;
  assign new_n39029_ = ~new_n39025_ & ~new_n39028_;
  assign new_n39030_ = new_n13311_ & ~new_n39029_;
  assign new_n39031_ = new_n38782_ & ~new_n39029_;
  assign ys__n29704 = new_n39030_ | new_n39031_;
  assign new_n39033_ = new_n22976_ & new_n22978_;
  assign new_n39034_ = new_n22962_ & new_n22966_;
  assign new_n39035_ = ~new_n39033_ & ~new_n39034_;
  assign new_n39036_ = ~new_n22983_ & new_n22989_;
  assign new_n39037_ = ~new_n39035_ & new_n39036_;
  assign new_n39038_ = ~new_n22989_ & new_n23015_;
  assign new_n39039_ = new_n23011_ & new_n39038_;
  assign new_n39040_ = ~new_n39037_ & ~new_n39039_;
  assign ys__n29706 = new_n38251_ & ~new_n39040_;
  assign new_n39042_ = ys__n29707 & ~ys__n29709;
  assign new_n39043_ = ys__n29708 & ys__n29709;
  assign ys__n29710 = new_n39042_ | new_n39043_;
  assign new_n39045_ = ~ys__n29709 & ys__n29711;
  assign new_n39046_ = ys__n29709 & ys__n29712;
  assign ys__n29713 = new_n39045_ | new_n39046_;
  assign new_n39048_ = ~ys__n29709 & ys__n29714;
  assign new_n39049_ = ys__n29709 & ys__n29715;
  assign ys__n29716 = new_n39048_ | new_n39049_;
  assign new_n39051_ = ~ys__n29709 & ys__n29717;
  assign new_n39052_ = ys__n29709 & ys__n29718;
  assign ys__n29719 = new_n39051_ | new_n39052_;
  assign new_n39054_ = ~ys__n29709 & ys__n29720;
  assign new_n39055_ = ys__n29709 & ys__n29721;
  assign ys__n29722 = new_n39054_ | new_n39055_;
  assign new_n39057_ = ~ys__n29709 & ys__n29723;
  assign new_n39058_ = ys__n29709 & ys__n29724;
  assign ys__n29725 = new_n39057_ | new_n39058_;
  assign new_n39060_ = ~ys__n29709 & ys__n29726;
  assign new_n39061_ = ys__n29709 & ys__n29727;
  assign ys__n29728 = new_n39060_ | new_n39061_;
  assign new_n39063_ = ~ys__n29709 & ys__n29729;
  assign new_n39064_ = ys__n29709 & ys__n29730;
  assign ys__n29731 = new_n39063_ | new_n39064_;
  assign new_n39066_ = ~ys__n29709 & ys__n29732;
  assign new_n39067_ = ys__n29709 & ys__n29733;
  assign ys__n29734 = new_n39066_ | new_n39067_;
  assign new_n39069_ = ~ys__n29709 & ys__n29735;
  assign new_n39070_ = ys__n29709 & ys__n29736;
  assign ys__n29737 = new_n39069_ | new_n39070_;
  assign new_n39072_ = ~ys__n29709 & ys__n29738;
  assign new_n39073_ = ys__n29709 & ys__n29739;
  assign ys__n29740 = new_n39072_ | new_n39073_;
  assign new_n39075_ = ~ys__n29709 & ys__n29741;
  assign new_n39076_ = ys__n29709 & ys__n29742;
  assign ys__n29743 = new_n39075_ | new_n39076_;
  assign new_n39078_ = ~ys__n29709 & ys__n29744;
  assign new_n39079_ = ys__n29709 & ys__n29745;
  assign ys__n29746 = new_n39078_ | new_n39079_;
  assign new_n39081_ = ~ys__n29709 & ys__n29747;
  assign new_n39082_ = ys__n29709 & ys__n29748;
  assign ys__n29749 = new_n39081_ | new_n39082_;
  assign new_n39084_ = ~ys__n29709 & ys__n29750;
  assign new_n39085_ = ys__n29709 & ys__n29751;
  assign ys__n29752 = new_n39084_ | new_n39085_;
  assign new_n39087_ = ~ys__n29709 & ys__n29753;
  assign new_n39088_ = ys__n29709 & ys__n29754;
  assign ys__n29755 = new_n39087_ | new_n39088_;
  assign new_n39090_ = ~ys__n29709 & ys__n29756;
  assign new_n39091_ = ys__n29709 & ys__n29757;
  assign ys__n29758 = new_n39090_ | new_n39091_;
  assign new_n39093_ = ~ys__n29709 & ys__n29759;
  assign new_n39094_ = ys__n29709 & ys__n29760;
  assign ys__n29761 = new_n39093_ | new_n39094_;
  assign new_n39096_ = ~ys__n29709 & ys__n29762;
  assign new_n39097_ = ys__n29709 & ys__n29763;
  assign ys__n29764 = new_n39096_ | new_n39097_;
  assign new_n39099_ = ~ys__n29709 & ys__n29765;
  assign new_n39100_ = ys__n29709 & ys__n29766;
  assign ys__n29767 = new_n39099_ | new_n39100_;
  assign new_n39102_ = ~ys__n29709 & ys__n29768;
  assign new_n39103_ = ys__n29709 & ys__n29769;
  assign ys__n29770 = new_n39102_ | new_n39103_;
  assign new_n39105_ = ~ys__n29709 & ys__n29771;
  assign new_n39106_ = ys__n29709 & ys__n29772;
  assign ys__n29773 = new_n39105_ | new_n39106_;
  assign new_n39108_ = ~ys__n29709 & ys__n29774;
  assign new_n39109_ = ys__n29709 & ys__n29775;
  assign ys__n29776 = new_n39108_ | new_n39109_;
  assign new_n39111_ = ~ys__n29709 & ys__n29777;
  assign new_n39112_ = ys__n29709 & ys__n29778;
  assign ys__n29779 = new_n39111_ | new_n39112_;
  assign new_n39114_ = ~ys__n29709 & ys__n29780;
  assign new_n39115_ = ys__n29709 & ys__n29781;
  assign ys__n29782 = new_n39114_ | new_n39115_;
  assign new_n39117_ = ~ys__n29709 & ys__n29783;
  assign new_n39118_ = ys__n29709 & ys__n29784;
  assign ys__n29785 = new_n39117_ | new_n39118_;
  assign new_n39120_ = ~ys__n29709 & ys__n29786;
  assign new_n39121_ = ys__n29709 & ys__n29787;
  assign ys__n29788 = new_n39120_ | new_n39121_;
  assign new_n39123_ = ~ys__n29709 & ys__n29789;
  assign new_n39124_ = ys__n29709 & ys__n29790;
  assign ys__n29791 = new_n39123_ | new_n39124_;
  assign new_n39126_ = ~ys__n29709 & ys__n29792;
  assign new_n39127_ = ys__n29709 & ys__n29793;
  assign ys__n29794 = new_n39126_ | new_n39127_;
  assign new_n39129_ = ~ys__n29709 & ys__n29795;
  assign new_n39130_ = ys__n29709 & ys__n29796;
  assign ys__n29797 = new_n39129_ | new_n39130_;
  assign new_n39132_ = ~ys__n29709 & ys__n29798;
  assign new_n39133_ = ys__n29709 & ys__n29799;
  assign ys__n29800 = new_n39132_ | new_n39133_;
  assign new_n39135_ = ~ys__n29709 & ys__n29801;
  assign new_n39136_ = ys__n29709 & ys__n29802;
  assign ys__n29803 = new_n39135_ | new_n39136_;
  assign new_n39138_ = ~ys__n28243 & new_n22973_;
  assign new_n39139_ = new_n22989_ & new_n39138_;
  assign ys__n29805 = ~ys__n4566 & new_n39139_;
  assign ys__n29807 = ys__n29806 & ~ys__n4566;
  assign ys__n29809 = ys__n29808 & ~ys__n4566;
  assign new_n39143_ = new_n22970_ & new_n22989_;
  assign new_n39144_ = ~new_n23015_ & new_n23018_;
  assign new_n39145_ = ~new_n22989_ & new_n39144_;
  assign new_n39146_ = ~new_n39143_ & ~new_n39145_;
  assign ys__n29811 = new_n38358_ & ~new_n39146_;
  assign ys__n29813 = ys__n29812 & ~ys__n4566;
  assign ys__n29814 = ys__n18118 & ~ys__n4566;
  assign ys__n29815 = ~ys__n28243 & ys__n23933;
  assign ys__n29816 = ~ys__n28243 & ys__n23936;
  assign ys__n29817 = ~ys__n28243 & ys__n23939;
  assign ys__n29818 = ~ys__n28243 & ys__n23942;
  assign ys__n29819 = ~ys__n28243 & ys__n23945;
  assign new_n39155_ = ~new_n39036_ & ~new_n39038_;
  assign ys__n29820 = ~ys__n28243 & ~new_n39155_;
  assign new_n39157_ = ~ys__n28243 & new_n22978_;
  assign new_n39158_ = new_n22989_ & new_n39157_;
  assign ys__n29821 = ~new_n22976_ & new_n39158_;
  assign new_n39160_ = new_n22966_ & new_n22989_;
  assign new_n39161_ = ~new_n22962_ & new_n39160_;
  assign new_n39162_ = ~new_n23011_ & new_n39038_;
  assign new_n39163_ = ~new_n39161_ & ~new_n39162_;
  assign ys__n29822 = ~ys__n28243 & ~new_n39163_;
  assign new_n39165_ = ~new_n23015_ & ~new_n39144_;
  assign new_n39166_ = ~ys__n28243 & ~new_n22989_;
  assign ys__n29823 = ~new_n39165_ & new_n39166_;
  assign new_n39168_ = ys__n29880 & ~new_n11737_;
  assign new_n39169_ = ys__n29881 & new_n11737_;
  assign ys__n29847 = new_n39168_ | new_n39169_;
  assign new_n39171_ = ys__n24389 & ~new_n13607_;
  assign new_n39172_ = new_n13607_ & ys__n24408;
  assign ys__n30010 = new_n39171_ | new_n39172_;
  assign new_n39174_ = ~new_n23747_ & ~new_n24579_;
  assign ys__n30080 = new_n24236_ | new_n39174_;
  assign new_n39176_ = ~new_n24277_ & ~new_n24576_;
  assign new_n39177_ = ~new_n37703_ & ~new_n39176_;
  assign ys__n30081 = ~new_n23747_ & ~new_n39177_;
  assign new_n39179_ = ~new_n24296_ & ~new_n24576_;
  assign new_n39180_ = ~new_n37725_ & ~new_n39179_;
  assign ys__n30082 = ~new_n23747_ & ~new_n39180_;
  assign new_n39182_ = ~new_n24315_ & ~new_n24576_;
  assign new_n39183_ = ~new_n37747_ & ~new_n39182_;
  assign ys__n30083 = ~new_n23747_ & ~new_n39183_;
  assign new_n39185_ = ~new_n24334_ & ~new_n24576_;
  assign new_n39186_ = ~new_n37769_ & ~new_n39185_;
  assign ys__n30084 = ~new_n23747_ & ~new_n39186_;
  assign new_n39188_ = ~new_n24353_ & ~new_n24576_;
  assign new_n39189_ = ~new_n37791_ & ~new_n39188_;
  assign ys__n30085 = ~new_n23747_ & ~new_n39189_;
  assign new_n39191_ = ~new_n24372_ & ~new_n24576_;
  assign new_n39192_ = ~new_n37813_ & ~new_n39191_;
  assign ys__n30086 = ~new_n23747_ & ~new_n39192_;
  assign new_n39194_ = ~new_n24391_ & ~new_n24576_;
  assign new_n39195_ = ~new_n37835_ & ~new_n39194_;
  assign ys__n30087 = ~new_n23747_ & ~new_n39195_;
  assign new_n39197_ = ~new_n24072_ & ~new_n24576_;
  assign new_n39198_ = ~new_n37886_ & ~new_n39197_;
  assign ys__n30089 = ~new_n23747_ & ~new_n39198_;
  assign new_n39200_ = ~new_n24090_ & ~new_n24576_;
  assign new_n39201_ = ~new_n37901_ & ~new_n39200_;
  assign ys__n30090 = ~new_n23747_ & ~new_n39201_;
  assign new_n39203_ = ~new_n24108_ & ~new_n24576_;
  assign new_n39204_ = ~new_n37916_ & ~new_n39203_;
  assign ys__n30091 = ~new_n23747_ & ~new_n39204_;
  assign new_n39206_ = ~new_n24126_ & ~new_n24576_;
  assign new_n39207_ = ~new_n37931_ & ~new_n39206_;
  assign ys__n30092 = ~new_n23747_ & ~new_n39207_;
  assign new_n39209_ = ~new_n24144_ & ~new_n24576_;
  assign new_n39210_ = ~new_n37946_ & ~new_n39209_;
  assign ys__n30093 = ~new_n23747_ & ~new_n39210_;
  assign new_n39212_ = ~new_n24162_ & ~new_n24576_;
  assign new_n39213_ = ~new_n37961_ & ~new_n39212_;
  assign ys__n30094 = ~new_n23747_ & ~new_n39213_;
  assign new_n39215_ = ~new_n24180_ & ~new_n24576_;
  assign new_n39216_ = ~new_n37976_ & ~new_n39215_;
  assign ys__n30095 = ~new_n23747_ & ~new_n39216_;
  assign new_n39218_ = ~new_n24198_ & ~new_n24576_;
  assign new_n39219_ = ~new_n37991_ & ~new_n39218_;
  assign ys__n30096 = ~new_n23747_ & ~new_n39219_;
  assign new_n39221_ = ~new_n23912_ & ~new_n24576_;
  assign new_n39222_ = ~new_n38010_ & ~new_n39221_;
  assign ys__n30098 = ~new_n23747_ & ~new_n39222_;
  assign new_n39224_ = ~new_n23927_ & ~new_n24576_;
  assign new_n39225_ = ~new_n38025_ & ~new_n39224_;
  assign ys__n30099 = ~new_n23747_ & ~new_n39225_;
  assign new_n39227_ = ~new_n23942_ & ~new_n24576_;
  assign new_n39228_ = ~new_n38040_ & ~new_n39227_;
  assign ys__n30100 = ~new_n23747_ & ~new_n39228_;
  assign new_n39230_ = ~new_n23957_ & ~new_n24576_;
  assign new_n39231_ = ~new_n38055_ & ~new_n39230_;
  assign ys__n30101 = ~new_n23747_ & ~new_n39231_;
  assign new_n39233_ = ~new_n23972_ & ~new_n24576_;
  assign new_n39234_ = ~new_n38070_ & ~new_n39233_;
  assign ys__n30102 = ~new_n23747_ & ~new_n39234_;
  assign new_n39236_ = ~new_n23987_ & ~new_n24576_;
  assign new_n39237_ = ~new_n38085_ & ~new_n39236_;
  assign ys__n30103 = ~new_n23747_ & ~new_n39237_;
  assign new_n39239_ = ~new_n24002_ & ~new_n24576_;
  assign new_n39240_ = ~new_n38100_ & ~new_n39239_;
  assign ys__n30104 = ~new_n23747_ & ~new_n39240_;
  assign new_n39242_ = ~new_n24017_ & ~new_n24576_;
  assign new_n39243_ = ~new_n38115_ & ~new_n39242_;
  assign ys__n30105 = ~new_n23747_ & ~new_n39243_;
  assign new_n39245_ = ~new_n23764_ & ~new_n24576_;
  assign new_n39246_ = ~new_n38130_ & ~new_n39245_;
  assign ys__n30106 = ~new_n23747_ & ~new_n39246_;
  assign new_n39248_ = ~new_n23779_ & ~new_n24576_;
  assign new_n39249_ = ~new_n38145_ & ~new_n39248_;
  assign ys__n30107 = ~new_n23747_ & ~new_n39249_;
  assign new_n39251_ = ~new_n23794_ & ~new_n24576_;
  assign new_n39252_ = ~new_n38160_ & ~new_n39251_;
  assign ys__n30108 = ~new_n23747_ & ~new_n39252_;
  assign new_n39254_ = ~new_n23809_ & ~new_n24576_;
  assign new_n39255_ = ~new_n38175_ & ~new_n39254_;
  assign ys__n30109 = ~new_n23747_ & ~new_n39255_;
  assign new_n39257_ = ~new_n23824_ & ~new_n24576_;
  assign new_n39258_ = ~new_n38190_ & ~new_n39257_;
  assign ys__n30110 = ~new_n23747_ & ~new_n39258_;
  assign new_n39260_ = ~new_n23839_ & ~new_n24576_;
  assign new_n39261_ = ~new_n38205_ & ~new_n39260_;
  assign ys__n30111 = ~new_n23747_ & ~new_n39261_;
  assign new_n39263_ = ~new_n23854_ & ~new_n24576_;
  assign new_n39264_ = ~new_n38220_ & ~new_n39263_;
  assign ys__n30112 = ~new_n23747_ & ~new_n39264_;
  assign new_n39266_ = ~new_n23869_ & ~new_n24576_;
  assign new_n39267_ = ~new_n38235_ & ~new_n39266_;
  assign ys__n30113 = ~new_n23747_ & ~new_n39267_;
  assign new_n39269_ = ~ys__n3039 & ys__n30080;
  assign new_n39270_ = ys__n3039 & ~new_n24246_;
  assign new_n39271_ = ~new_n39269_ & ~new_n39270_;
  assign new_n39272_ = ~ys__n740 & ~ys__n3039;
  assign new_n39273_ = ~new_n39271_ & new_n39272_;
  assign new_n39274_ = ys__n3039 & ~new_n39271_;
  assign ys__n30119 = new_n39273_ | new_n39274_;
  assign new_n39276_ = ~ys__n3039 & ys__n30081;
  assign new_n39277_ = ys__n3039 & ~new_n24266_;
  assign new_n39278_ = ~new_n39276_ & ~new_n39277_;
  assign new_n39279_ = new_n39272_ & ~new_n39278_;
  assign new_n39280_ = ys__n3039 & ~new_n39278_;
  assign ys__n30122 = new_n39279_ | new_n39280_;
  assign new_n39282_ = ~ys__n3039 & ys__n30082;
  assign new_n39283_ = ys__n3039 & ~new_n24285_;
  assign new_n39284_ = ~new_n39282_ & ~new_n39283_;
  assign new_n39285_ = new_n39272_ & ~new_n39284_;
  assign new_n39286_ = ys__n3039 & ~new_n39284_;
  assign ys__n30125 = new_n39285_ | new_n39286_;
  assign new_n39288_ = ~ys__n3039 & ys__n30083;
  assign new_n39289_ = ys__n3039 & ~new_n24304_;
  assign new_n39290_ = ~new_n39288_ & ~new_n39289_;
  assign new_n39291_ = new_n39272_ & ~new_n39290_;
  assign new_n39292_ = ys__n3039 & ~new_n39290_;
  assign ys__n30128 = new_n39291_ | new_n39292_;
  assign new_n39294_ = ~ys__n3039 & ys__n30084;
  assign new_n39295_ = ys__n3039 & ~new_n24323_;
  assign new_n39296_ = ~new_n39294_ & ~new_n39295_;
  assign new_n39297_ = new_n39272_ & ~new_n39296_;
  assign new_n39298_ = ys__n3039 & ~new_n39296_;
  assign ys__n30131 = new_n39297_ | new_n39298_;
  assign new_n39300_ = ~ys__n3039 & ys__n30085;
  assign new_n39301_ = ys__n3039 & ~new_n24342_;
  assign new_n39302_ = ~new_n39300_ & ~new_n39301_;
  assign new_n39303_ = new_n39272_ & ~new_n39302_;
  assign new_n39304_ = ys__n3039 & ~new_n39302_;
  assign ys__n30134 = new_n39303_ | new_n39304_;
  assign new_n39306_ = ~ys__n3039 & ys__n30086;
  assign new_n39307_ = ys__n3039 & ~new_n24361_;
  assign new_n39308_ = ~new_n39306_ & ~new_n39307_;
  assign new_n39309_ = new_n39272_ & ~new_n39308_;
  assign new_n39310_ = ys__n3039 & ~new_n39308_;
  assign ys__n30137 = new_n39309_ | new_n39310_;
  assign new_n39312_ = ~ys__n3039 & ys__n30087;
  assign new_n39313_ = ys__n3039 & ~new_n24380_;
  assign new_n39314_ = ~new_n39312_ & ~new_n39313_;
  assign new_n39315_ = new_n39272_ & ~new_n39314_;
  assign new_n39316_ = ys__n3039 & ~new_n39314_;
  assign ys__n30140 = new_n39315_ | new_n39316_;
  assign new_n39318_ = ~ys__n3039 & ys__n30089;
  assign new_n39319_ = ys__n3039 & ~new_n24061_;
  assign new_n39320_ = ~new_n39318_ & ~new_n39319_;
  assign new_n39321_ = new_n39272_ & ~new_n39320_;
  assign new_n39322_ = ys__n3039 & ~new_n39320_;
  assign ys__n30143 = new_n39321_ | new_n39322_;
  assign new_n39324_ = ~ys__n3039 & ys__n30090;
  assign new_n39325_ = ys__n3039 & ~new_n24079_;
  assign new_n39326_ = ~new_n39324_ & ~new_n39325_;
  assign new_n39327_ = new_n39272_ & ~new_n39326_;
  assign new_n39328_ = ys__n3039 & ~new_n39326_;
  assign ys__n30146 = new_n39327_ | new_n39328_;
  assign new_n39330_ = ~ys__n3039 & ys__n30091;
  assign new_n39331_ = ys__n3039 & ~new_n24097_;
  assign new_n39332_ = ~new_n39330_ & ~new_n39331_;
  assign new_n39333_ = new_n39272_ & ~new_n39332_;
  assign new_n39334_ = ys__n3039 & ~new_n39332_;
  assign ys__n30149 = new_n39333_ | new_n39334_;
  assign new_n39336_ = ~ys__n3039 & ys__n30092;
  assign new_n39337_ = ys__n3039 & ~new_n24115_;
  assign new_n39338_ = ~new_n39336_ & ~new_n39337_;
  assign new_n39339_ = new_n39272_ & ~new_n39338_;
  assign new_n39340_ = ys__n3039 & ~new_n39338_;
  assign ys__n30152 = new_n39339_ | new_n39340_;
  assign new_n39342_ = ~ys__n3039 & ys__n30093;
  assign new_n39343_ = ys__n3039 & ~new_n24133_;
  assign new_n39344_ = ~new_n39342_ & ~new_n39343_;
  assign new_n39345_ = new_n39272_ & ~new_n39344_;
  assign new_n39346_ = ys__n3039 & ~new_n39344_;
  assign ys__n30155 = new_n39345_ | new_n39346_;
  assign new_n39348_ = ~ys__n3039 & ys__n30094;
  assign new_n39349_ = ys__n3039 & ~new_n24151_;
  assign new_n39350_ = ~new_n39348_ & ~new_n39349_;
  assign new_n39351_ = new_n39272_ & ~new_n39350_;
  assign new_n39352_ = ys__n3039 & ~new_n39350_;
  assign ys__n30158 = new_n39351_ | new_n39352_;
  assign new_n39354_ = ~ys__n3039 & ys__n30095;
  assign new_n39355_ = ys__n3039 & ~new_n24169_;
  assign new_n39356_ = ~new_n39354_ & ~new_n39355_;
  assign new_n39357_ = new_n39272_ & ~new_n39356_;
  assign new_n39358_ = ys__n3039 & ~new_n39356_;
  assign ys__n30161 = new_n39357_ | new_n39358_;
  assign new_n39360_ = ~ys__n3039 & ys__n30096;
  assign new_n39361_ = ys__n3039 & ~new_n24187_;
  assign new_n39362_ = ~new_n39360_ & ~new_n39361_;
  assign new_n39363_ = new_n39272_ & ~new_n39362_;
  assign new_n39364_ = ys__n3039 & ~new_n39362_;
  assign ys__n30164 = new_n39363_ | new_n39364_;
  assign new_n39366_ = ~ys__n3039 & ys__n30098;
  assign new_n39367_ = ys__n3039 & ~new_n23901_;
  assign new_n39368_ = ~new_n39366_ & ~new_n39367_;
  assign new_n39369_ = new_n39272_ & ~new_n39368_;
  assign new_n39370_ = ys__n3039 & ~new_n39368_;
  assign ys__n30167 = new_n39369_ | new_n39370_;
  assign new_n39372_ = ~ys__n3039 & ys__n30099;
  assign new_n39373_ = ys__n3039 & ~new_n23916_;
  assign new_n39374_ = ~new_n39372_ & ~new_n39373_;
  assign new_n39375_ = new_n39272_ & ~new_n39374_;
  assign new_n39376_ = ys__n3039 & ~new_n39374_;
  assign ys__n30170 = new_n39375_ | new_n39376_;
  assign new_n39378_ = ~ys__n3039 & ys__n30100;
  assign new_n39379_ = ys__n3039 & ~new_n23931_;
  assign new_n39380_ = ~new_n39378_ & ~new_n39379_;
  assign new_n39381_ = new_n39272_ & ~new_n39380_;
  assign new_n39382_ = ys__n3039 & ~new_n39380_;
  assign ys__n30173 = new_n39381_ | new_n39382_;
  assign new_n39384_ = ~ys__n3039 & ys__n30101;
  assign new_n39385_ = ys__n3039 & ~new_n23946_;
  assign new_n39386_ = ~new_n39384_ & ~new_n39385_;
  assign new_n39387_ = new_n39272_ & ~new_n39386_;
  assign new_n39388_ = ys__n3039 & ~new_n39386_;
  assign ys__n30176 = new_n39387_ | new_n39388_;
  assign new_n39390_ = ~ys__n3039 & ys__n30102;
  assign new_n39391_ = ys__n3039 & ~new_n23961_;
  assign new_n39392_ = ~new_n39390_ & ~new_n39391_;
  assign new_n39393_ = new_n39272_ & ~new_n39392_;
  assign new_n39394_ = ys__n3039 & ~new_n39392_;
  assign ys__n30179 = new_n39393_ | new_n39394_;
  assign new_n39396_ = ~ys__n3039 & ys__n30103;
  assign new_n39397_ = ys__n3039 & ~new_n23976_;
  assign new_n39398_ = ~new_n39396_ & ~new_n39397_;
  assign new_n39399_ = new_n39272_ & ~new_n39398_;
  assign new_n39400_ = ys__n3039 & ~new_n39398_;
  assign ys__n30182 = new_n39399_ | new_n39400_;
  assign new_n39402_ = ~ys__n3039 & ys__n30104;
  assign new_n39403_ = ys__n3039 & ~new_n23991_;
  assign new_n39404_ = ~new_n39402_ & ~new_n39403_;
  assign new_n39405_ = new_n39272_ & ~new_n39404_;
  assign new_n39406_ = ys__n3039 & ~new_n39404_;
  assign ys__n30185 = new_n39405_ | new_n39406_;
  assign new_n39408_ = ~ys__n3039 & ys__n30105;
  assign new_n39409_ = ys__n3039 & ~new_n24006_;
  assign new_n39410_ = ~new_n39408_ & ~new_n39409_;
  assign new_n39411_ = new_n39272_ & ~new_n39410_;
  assign new_n39412_ = ys__n3039 & ~new_n39410_;
  assign ys__n30188 = new_n39411_ | new_n39412_;
  assign new_n39414_ = ~ys__n3039 & ys__n30106;
  assign new_n39415_ = ys__n3039 & ~new_n23742_;
  assign new_n39416_ = ~new_n39414_ & ~new_n39415_;
  assign new_n39417_ = new_n39272_ & ~new_n39416_;
  assign new_n39418_ = ys__n3039 & ~new_n39416_;
  assign ys__n30191 = new_n39417_ | new_n39418_;
  assign new_n39420_ = ~ys__n3039 & ys__n30107;
  assign new_n39421_ = ys__n3039 & ~new_n23768_;
  assign new_n39422_ = ~new_n39420_ & ~new_n39421_;
  assign new_n39423_ = new_n39272_ & ~new_n39422_;
  assign new_n39424_ = ys__n3039 & ~new_n39422_;
  assign ys__n30194 = new_n39423_ | new_n39424_;
  assign new_n39426_ = ~ys__n3039 & ys__n30108;
  assign new_n39427_ = ys__n3039 & ~new_n23783_;
  assign new_n39428_ = ~new_n39426_ & ~new_n39427_;
  assign new_n39429_ = new_n39272_ & ~new_n39428_;
  assign new_n39430_ = ys__n3039 & ~new_n39428_;
  assign ys__n30197 = new_n39429_ | new_n39430_;
  assign new_n39432_ = ~ys__n3039 & ys__n30109;
  assign new_n39433_ = ys__n3039 & ~new_n23798_;
  assign new_n39434_ = ~new_n39432_ & ~new_n39433_;
  assign new_n39435_ = new_n39272_ & ~new_n39434_;
  assign new_n39436_ = ys__n3039 & ~new_n39434_;
  assign ys__n30200 = new_n39435_ | new_n39436_;
  assign new_n39438_ = ~ys__n3039 & ys__n30110;
  assign new_n39439_ = ys__n3039 & ~new_n23813_;
  assign new_n39440_ = ~new_n39438_ & ~new_n39439_;
  assign new_n39441_ = new_n39272_ & ~new_n39440_;
  assign new_n39442_ = ys__n3039 & ~new_n39440_;
  assign ys__n30203 = new_n39441_ | new_n39442_;
  assign new_n39444_ = ~ys__n3039 & ys__n30111;
  assign new_n39445_ = ys__n3039 & ~new_n23828_;
  assign new_n39446_ = ~new_n39444_ & ~new_n39445_;
  assign new_n39447_ = new_n39272_ & ~new_n39446_;
  assign new_n39448_ = ys__n3039 & ~new_n39446_;
  assign ys__n30206 = new_n39447_ | new_n39448_;
  assign new_n39450_ = ~ys__n3039 & ys__n30112;
  assign new_n39451_ = ys__n3039 & ~new_n23843_;
  assign new_n39452_ = ~new_n39450_ & ~new_n39451_;
  assign new_n39453_ = new_n39272_ & ~new_n39452_;
  assign new_n39454_ = ys__n3039 & ~new_n39452_;
  assign ys__n30209 = new_n39453_ | new_n39454_;
  assign new_n39456_ = ~ys__n3039 & ys__n30113;
  assign new_n39457_ = ys__n3039 & ~new_n23858_;
  assign new_n39458_ = ~new_n39456_ & ~new_n39457_;
  assign new_n39459_ = new_n39272_ & ~new_n39458_;
  assign new_n39460_ = ys__n3039 & ~new_n39458_;
  assign ys__n30212 = new_n39459_ | new_n39460_;
  assign new_n39462_ = ys__n30220 & ~ys__n740;
  assign new_n39463_ = ~ys__n4566 & new_n39462_;
  assign new_n39464_ = ys__n30214 & ys__n740;
  assign ys__n30215 = new_n39463_ | new_n39464_;
  assign ys__n33414 = ~ys__n18120 & ~ys__n740;
  assign new_n39467_ = ys__n30225 & ys__n740;
  assign ys__n30226 = ys__n33414 | new_n39467_;
  assign new_n39469_ = ys__n352 & ys__n23335;
  assign new_n39470_ = new_n15136_ & new_n39469_;
  assign new_n39471_ = ~ys__n17867 & ~ys__n30334;
  assign new_n39472_ = ys__n17867 & ys__n30334;
  assign new_n39473_ = ~new_n39471_ & ~new_n39472_;
  assign new_n39474_ = ~ys__n17869 & ~ys__n30334;
  assign new_n39475_ = ys__n17869 & ys__n30334;
  assign new_n39476_ = ~new_n39474_ & ~new_n39475_;
  assign new_n39477_ = ~ys__n17803 & ~new_n39476_;
  assign new_n39478_ = ys__n17803 & new_n39476_;
  assign new_n39479_ = ~new_n39477_ & ~new_n39478_;
  assign new_n39480_ = ~new_n39473_ & new_n39479_;
  assign new_n39481_ = new_n39473_ & ~new_n39479_;
  assign new_n39482_ = ~new_n39480_ & ~new_n39481_;
  assign new_n39483_ = ~ys__n33581 & ~new_n39473_;
  assign new_n39484_ = ~ys__n17866 & ~ys__n30334;
  assign new_n39485_ = ys__n17866 & ys__n30334;
  assign new_n39486_ = ~new_n39484_ & ~new_n39485_;
  assign new_n39487_ = new_n39483_ & ~new_n39486_;
  assign new_n39488_ = new_n39473_ & new_n39486_;
  assign new_n39489_ = ys__n33581 & ~new_n39488_;
  assign new_n39490_ = ~new_n39487_ & ~new_n39489_;
  assign new_n39491_ = ~new_n39482_ & ~new_n39490_;
  assign new_n39492_ = new_n39482_ & ~new_n39490_;
  assign new_n39493_ = ~new_n39482_ & new_n39490_;
  assign new_n39494_ = ~new_n39492_ & ~new_n39493_;
  assign new_n39495_ = ys__n33581 & new_n39473_;
  assign new_n39496_ = ~new_n39483_ & ~new_n39495_;
  assign new_n39497_ = ~new_n39486_ & new_n39496_;
  assign new_n39498_ = new_n39486_ & ~new_n39496_;
  assign new_n39499_ = ~new_n39497_ & ~new_n39498_;
  assign new_n39500_ = ~ys__n33579 & ~new_n39486_;
  assign new_n39501_ = ~ys__n30334 & new_n39500_;
  assign new_n39502_ = ys__n30334 & new_n39486_;
  assign new_n39503_ = ys__n33579 & ~new_n39502_;
  assign new_n39504_ = ~new_n39501_ & ~new_n39503_;
  assign new_n39505_ = ~new_n39499_ & ~new_n39504_;
  assign new_n39506_ = ~new_n39494_ & new_n39505_;
  assign new_n39507_ = ~new_n39491_ & ~new_n39506_;
  assign new_n39508_ = ~ys__n17870 & ~ys__n30334;
  assign new_n39509_ = ys__n17870 & ys__n30334;
  assign new_n39510_ = ~new_n39508_ & ~new_n39509_;
  assign new_n39511_ = ~ys__n17872 & ~ys__n30334;
  assign new_n39512_ = ys__n17872 & ys__n30334;
  assign new_n39513_ = ~new_n39511_ & ~new_n39512_;
  assign new_n39514_ = ~ys__n17806 & ~new_n39513_;
  assign new_n39515_ = ys__n17806 & new_n39513_;
  assign new_n39516_ = ~new_n39514_ & ~new_n39515_;
  assign new_n39517_ = ~new_n39510_ & new_n39516_;
  assign new_n39518_ = new_n39510_ & ~new_n39516_;
  assign new_n39519_ = ~new_n39517_ & ~new_n39518_;
  assign new_n39520_ = ~ys__n17804 & ~new_n39510_;
  assign new_n39521_ = ~new_n39476_ & new_n39520_;
  assign new_n39522_ = new_n39476_ & new_n39510_;
  assign new_n39523_ = ys__n17804 & ~new_n39522_;
  assign new_n39524_ = ~new_n39521_ & ~new_n39523_;
  assign new_n39525_ = new_n39519_ & ~new_n39524_;
  assign new_n39526_ = ~new_n39519_ & new_n39524_;
  assign new_n39527_ = ~new_n39525_ & ~new_n39526_;
  assign new_n39528_ = ys__n17804 & new_n39510_;
  assign new_n39529_ = ~new_n39520_ & ~new_n39528_;
  assign new_n39530_ = ~new_n39476_ & new_n39529_;
  assign new_n39531_ = new_n39476_ & ~new_n39529_;
  assign new_n39532_ = ~new_n39530_ & ~new_n39531_;
  assign new_n39533_ = ~new_n39473_ & new_n39477_;
  assign new_n39534_ = new_n39473_ & new_n39476_;
  assign new_n39535_ = ys__n17803 & ~new_n39534_;
  assign new_n39536_ = ~new_n39533_ & ~new_n39535_;
  assign new_n39537_ = new_n39532_ & ~new_n39536_;
  assign new_n39538_ = ~new_n39532_ & new_n39536_;
  assign new_n39539_ = ~new_n39537_ & ~new_n39538_;
  assign new_n39540_ = ~new_n39527_ & ~new_n39539_;
  assign new_n39541_ = ~new_n39507_ & new_n39540_;
  assign new_n39542_ = ~new_n39519_ & ~new_n39524_;
  assign new_n39543_ = ~new_n39532_ & ~new_n39536_;
  assign new_n39544_ = ~new_n39527_ & new_n39543_;
  assign new_n39545_ = ~new_n39542_ & ~new_n39544_;
  assign new_n39546_ = ~new_n39541_ & new_n39545_;
  assign new_n39547_ = ~ys__n17876 & ~ys__n30334;
  assign new_n39548_ = ys__n17876 & ys__n30334;
  assign new_n39549_ = ~new_n39547_ & ~new_n39548_;
  assign new_n39550_ = ~ys__n17878 & ~ys__n30334;
  assign new_n39551_ = ys__n17878 & ys__n30334;
  assign new_n39552_ = ~new_n39550_ & ~new_n39551_;
  assign new_n39553_ = ~ys__n17812 & ~new_n39552_;
  assign new_n39554_ = ys__n17812 & new_n39552_;
  assign new_n39555_ = ~new_n39553_ & ~new_n39554_;
  assign new_n39556_ = ~new_n39549_ & new_n39555_;
  assign new_n39557_ = new_n39549_ & ~new_n39555_;
  assign new_n39558_ = ~new_n39556_ & ~new_n39557_;
  assign new_n39559_ = ~ys__n17810 & ~new_n39549_;
  assign new_n39560_ = ~ys__n17875 & ~ys__n30334;
  assign new_n39561_ = ys__n17875 & ys__n30334;
  assign new_n39562_ = ~new_n39560_ & ~new_n39561_;
  assign new_n39563_ = new_n39559_ & ~new_n39562_;
  assign new_n39564_ = new_n39549_ & new_n39562_;
  assign new_n39565_ = ys__n17810 & ~new_n39564_;
  assign new_n39566_ = ~new_n39563_ & ~new_n39565_;
  assign new_n39567_ = new_n39558_ & ~new_n39566_;
  assign new_n39568_ = ~new_n39558_ & new_n39566_;
  assign new_n39569_ = ~new_n39567_ & ~new_n39568_;
  assign new_n39570_ = ys__n17810 & new_n39549_;
  assign new_n39571_ = ~new_n39559_ & ~new_n39570_;
  assign new_n39572_ = ~new_n39562_ & new_n39571_;
  assign new_n39573_ = new_n39562_ & ~new_n39571_;
  assign new_n39574_ = ~new_n39572_ & ~new_n39573_;
  assign new_n39575_ = ~ys__n17809 & ~new_n39562_;
  assign new_n39576_ = ~ys__n17873 & ~ys__n30334;
  assign new_n39577_ = ys__n17873 & ys__n30334;
  assign new_n39578_ = ~new_n39576_ & ~new_n39577_;
  assign new_n39579_ = new_n39575_ & ~new_n39578_;
  assign new_n39580_ = new_n39562_ & new_n39578_;
  assign new_n39581_ = ys__n17809 & ~new_n39580_;
  assign new_n39582_ = ~new_n39579_ & ~new_n39581_;
  assign new_n39583_ = new_n39574_ & ~new_n39582_;
  assign new_n39584_ = ~new_n39574_ & new_n39582_;
  assign new_n39585_ = ~new_n39583_ & ~new_n39584_;
  assign new_n39586_ = ~new_n39569_ & ~new_n39585_;
  assign new_n39587_ = ys__n17809 & new_n39562_;
  assign new_n39588_ = ~new_n39575_ & ~new_n39587_;
  assign new_n39589_ = ~new_n39578_ & new_n39588_;
  assign new_n39590_ = new_n39578_ & ~new_n39588_;
  assign new_n39591_ = ~new_n39589_ & ~new_n39590_;
  assign new_n39592_ = ~ys__n17807 & ~new_n39578_;
  assign new_n39593_ = ~new_n39513_ & new_n39592_;
  assign new_n39594_ = new_n39513_ & new_n39578_;
  assign new_n39595_ = ys__n17807 & ~new_n39594_;
  assign new_n39596_ = ~new_n39593_ & ~new_n39595_;
  assign new_n39597_ = new_n39591_ & ~new_n39596_;
  assign new_n39598_ = ~new_n39591_ & new_n39596_;
  assign new_n39599_ = ~new_n39597_ & ~new_n39598_;
  assign new_n39600_ = ys__n17807 & new_n39578_;
  assign new_n39601_ = ~new_n39592_ & ~new_n39600_;
  assign new_n39602_ = ~new_n39513_ & new_n39601_;
  assign new_n39603_ = new_n39513_ & ~new_n39601_;
  assign new_n39604_ = ~new_n39602_ & ~new_n39603_;
  assign new_n39605_ = ~new_n39510_ & new_n39514_;
  assign new_n39606_ = new_n39510_ & new_n39513_;
  assign new_n39607_ = ys__n17806 & ~new_n39606_;
  assign new_n39608_ = ~new_n39605_ & ~new_n39607_;
  assign new_n39609_ = new_n39604_ & ~new_n39608_;
  assign new_n39610_ = ~new_n39604_ & new_n39608_;
  assign new_n39611_ = ~new_n39609_ & ~new_n39610_;
  assign new_n39612_ = ~new_n39599_ & ~new_n39611_;
  assign new_n39613_ = new_n39586_ & new_n39612_;
  assign new_n39614_ = ~new_n39546_ & new_n39613_;
  assign new_n39615_ = ~new_n39591_ & ~new_n39596_;
  assign new_n39616_ = ~new_n39604_ & ~new_n39608_;
  assign new_n39617_ = ~new_n39599_ & new_n39616_;
  assign new_n39618_ = ~new_n39615_ & ~new_n39617_;
  assign new_n39619_ = new_n39586_ & ~new_n39618_;
  assign new_n39620_ = ~new_n39558_ & ~new_n39566_;
  assign new_n39621_ = ~new_n39574_ & ~new_n39582_;
  assign new_n39622_ = ~new_n39569_ & new_n39621_;
  assign new_n39623_ = ~new_n39620_ & ~new_n39622_;
  assign new_n39624_ = ~new_n39619_ & new_n39623_;
  assign new_n39625_ = ~new_n39614_ & new_n39624_;
  assign new_n39626_ = ~ys__n17888 & ~ys__n30334;
  assign new_n39627_ = ys__n17888 & ys__n30334;
  assign new_n39628_ = ~new_n39626_ & ~new_n39627_;
  assign new_n39629_ = ~ys__n17890 & ~ys__n30334;
  assign new_n39630_ = ys__n17890 & ys__n30334;
  assign new_n39631_ = ~new_n39629_ & ~new_n39630_;
  assign new_n39632_ = ~ys__n17824 & ~new_n39631_;
  assign new_n39633_ = ys__n17824 & new_n39631_;
  assign new_n39634_ = ~new_n39632_ & ~new_n39633_;
  assign new_n39635_ = ~new_n39628_ & new_n39634_;
  assign new_n39636_ = new_n39628_ & ~new_n39634_;
  assign new_n39637_ = ~new_n39635_ & ~new_n39636_;
  assign new_n39638_ = ~ys__n17822 & ~new_n39628_;
  assign new_n39639_ = ~ys__n17887 & ~ys__n30334;
  assign new_n39640_ = ys__n17887 & ys__n30334;
  assign new_n39641_ = ~new_n39639_ & ~new_n39640_;
  assign new_n39642_ = new_n39638_ & ~new_n39641_;
  assign new_n39643_ = new_n39628_ & new_n39641_;
  assign new_n39644_ = ys__n17822 & ~new_n39643_;
  assign new_n39645_ = ~new_n39642_ & ~new_n39644_;
  assign new_n39646_ = new_n39637_ & ~new_n39645_;
  assign new_n39647_ = ~new_n39637_ & new_n39645_;
  assign new_n39648_ = ~new_n39646_ & ~new_n39647_;
  assign new_n39649_ = ys__n17822 & new_n39628_;
  assign new_n39650_ = ~new_n39638_ & ~new_n39649_;
  assign new_n39651_ = ~new_n39641_ & new_n39650_;
  assign new_n39652_ = new_n39641_ & ~new_n39650_;
  assign new_n39653_ = ~new_n39651_ & ~new_n39652_;
  assign new_n39654_ = ~ys__n17821 & ~new_n39641_;
  assign new_n39655_ = ~ys__n17885 & ~ys__n30334;
  assign new_n39656_ = ys__n17885 & ys__n30334;
  assign new_n39657_ = ~new_n39655_ & ~new_n39656_;
  assign new_n39658_ = new_n39654_ & ~new_n39657_;
  assign new_n39659_ = new_n39641_ & new_n39657_;
  assign new_n39660_ = ys__n17821 & ~new_n39659_;
  assign new_n39661_ = ~new_n39658_ & ~new_n39660_;
  assign new_n39662_ = new_n39653_ & ~new_n39661_;
  assign new_n39663_ = ~new_n39653_ & new_n39661_;
  assign new_n39664_ = ~new_n39662_ & ~new_n39663_;
  assign new_n39665_ = ~new_n39648_ & ~new_n39664_;
  assign new_n39666_ = ys__n17821 & new_n39641_;
  assign new_n39667_ = ~new_n39654_ & ~new_n39666_;
  assign new_n39668_ = ~new_n39657_ & new_n39667_;
  assign new_n39669_ = new_n39657_ & ~new_n39667_;
  assign new_n39670_ = ~new_n39668_ & ~new_n39669_;
  assign new_n39671_ = ~ys__n17819 & ~new_n39657_;
  assign new_n39672_ = ~ys__n17884 & ~ys__n30334;
  assign new_n39673_ = ys__n17884 & ys__n30334;
  assign new_n39674_ = ~new_n39672_ & ~new_n39673_;
  assign new_n39675_ = new_n39671_ & ~new_n39674_;
  assign new_n39676_ = new_n39657_ & new_n39674_;
  assign new_n39677_ = ys__n17819 & ~new_n39676_;
  assign new_n39678_ = ~new_n39675_ & ~new_n39677_;
  assign new_n39679_ = new_n39670_ & ~new_n39678_;
  assign new_n39680_ = ~new_n39670_ & new_n39678_;
  assign new_n39681_ = ~new_n39679_ & ~new_n39680_;
  assign new_n39682_ = ys__n17819 & new_n39657_;
  assign new_n39683_ = ~new_n39671_ & ~new_n39682_;
  assign new_n39684_ = ~new_n39674_ & new_n39683_;
  assign new_n39685_ = new_n39674_ & ~new_n39683_;
  assign new_n39686_ = ~new_n39684_ & ~new_n39685_;
  assign new_n39687_ = ~ys__n17818 & ~new_n39674_;
  assign new_n39688_ = ~ys__n17882 & ~ys__n30334;
  assign new_n39689_ = ys__n17882 & ys__n30334;
  assign new_n39690_ = ~new_n39688_ & ~new_n39689_;
  assign new_n39691_ = new_n39687_ & ~new_n39690_;
  assign new_n39692_ = new_n39674_ & new_n39690_;
  assign new_n39693_ = ys__n17818 & ~new_n39692_;
  assign new_n39694_ = ~new_n39691_ & ~new_n39693_;
  assign new_n39695_ = new_n39686_ & ~new_n39694_;
  assign new_n39696_ = ~new_n39686_ & new_n39694_;
  assign new_n39697_ = ~new_n39695_ & ~new_n39696_;
  assign new_n39698_ = ~new_n39681_ & ~new_n39697_;
  assign new_n39699_ = new_n39665_ & new_n39698_;
  assign new_n39700_ = ys__n17818 & new_n39674_;
  assign new_n39701_ = ~new_n39687_ & ~new_n39700_;
  assign new_n39702_ = ~new_n39690_ & new_n39701_;
  assign new_n39703_ = new_n39690_ & ~new_n39701_;
  assign new_n39704_ = ~new_n39702_ & ~new_n39703_;
  assign new_n39705_ = ~ys__n17816 & ~new_n39690_;
  assign new_n39706_ = ~ys__n17881 & ~ys__n30334;
  assign new_n39707_ = ys__n17881 & ys__n30334;
  assign new_n39708_ = ~new_n39706_ & ~new_n39707_;
  assign new_n39709_ = new_n39705_ & ~new_n39708_;
  assign new_n39710_ = new_n39690_ & new_n39708_;
  assign new_n39711_ = ys__n17816 & ~new_n39710_;
  assign new_n39712_ = ~new_n39709_ & ~new_n39711_;
  assign new_n39713_ = new_n39704_ & ~new_n39712_;
  assign new_n39714_ = ~new_n39704_ & new_n39712_;
  assign new_n39715_ = ~new_n39713_ & ~new_n39714_;
  assign new_n39716_ = ys__n17816 & new_n39690_;
  assign new_n39717_ = ~new_n39705_ & ~new_n39716_;
  assign new_n39718_ = ~new_n39708_ & new_n39717_;
  assign new_n39719_ = new_n39708_ & ~new_n39717_;
  assign new_n39720_ = ~new_n39718_ & ~new_n39719_;
  assign new_n39721_ = ~ys__n17815 & ~new_n39708_;
  assign new_n39722_ = ~ys__n17879 & ~ys__n30334;
  assign new_n39723_ = ys__n17879 & ys__n30334;
  assign new_n39724_ = ~new_n39722_ & ~new_n39723_;
  assign new_n39725_ = new_n39721_ & ~new_n39724_;
  assign new_n39726_ = new_n39708_ & new_n39724_;
  assign new_n39727_ = ys__n17815 & ~new_n39726_;
  assign new_n39728_ = ~new_n39725_ & ~new_n39727_;
  assign new_n39729_ = new_n39720_ & ~new_n39728_;
  assign new_n39730_ = ~new_n39720_ & new_n39728_;
  assign new_n39731_ = ~new_n39729_ & ~new_n39730_;
  assign new_n39732_ = ~new_n39715_ & ~new_n39731_;
  assign new_n39733_ = ys__n17815 & new_n39708_;
  assign new_n39734_ = ~new_n39721_ & ~new_n39733_;
  assign new_n39735_ = ~new_n39724_ & new_n39734_;
  assign new_n39736_ = new_n39724_ & ~new_n39734_;
  assign new_n39737_ = ~new_n39735_ & ~new_n39736_;
  assign new_n39738_ = ~ys__n17813 & ~new_n39724_;
  assign new_n39739_ = ~new_n39552_ & new_n39738_;
  assign new_n39740_ = new_n39552_ & new_n39724_;
  assign new_n39741_ = ys__n17813 & ~new_n39740_;
  assign new_n39742_ = ~new_n39739_ & ~new_n39741_;
  assign new_n39743_ = new_n39737_ & ~new_n39742_;
  assign new_n39744_ = ~new_n39737_ & new_n39742_;
  assign new_n39745_ = ~new_n39743_ & ~new_n39744_;
  assign new_n39746_ = ys__n17813 & new_n39724_;
  assign new_n39747_ = ~new_n39738_ & ~new_n39746_;
  assign new_n39748_ = ~new_n39552_ & new_n39747_;
  assign new_n39749_ = new_n39552_ & ~new_n39747_;
  assign new_n39750_ = ~new_n39748_ & ~new_n39749_;
  assign new_n39751_ = ~new_n39549_ & new_n39553_;
  assign new_n39752_ = new_n39549_ & new_n39552_;
  assign new_n39753_ = ys__n17812 & ~new_n39752_;
  assign new_n39754_ = ~new_n39751_ & ~new_n39753_;
  assign new_n39755_ = new_n39750_ & ~new_n39754_;
  assign new_n39756_ = ~new_n39750_ & new_n39754_;
  assign new_n39757_ = ~new_n39755_ & ~new_n39756_;
  assign new_n39758_ = ~new_n39745_ & ~new_n39757_;
  assign new_n39759_ = new_n39732_ & new_n39758_;
  assign new_n39760_ = new_n39699_ & new_n39759_;
  assign new_n39761_ = ~new_n39625_ & new_n39760_;
  assign new_n39762_ = ~new_n39737_ & ~new_n39742_;
  assign new_n39763_ = ~new_n39750_ & ~new_n39754_;
  assign new_n39764_ = ~new_n39745_ & new_n39763_;
  assign new_n39765_ = ~new_n39762_ & ~new_n39764_;
  assign new_n39766_ = new_n39732_ & ~new_n39765_;
  assign new_n39767_ = ~new_n39704_ & ~new_n39712_;
  assign new_n39768_ = ~new_n39720_ & ~new_n39728_;
  assign new_n39769_ = ~new_n39715_ & new_n39768_;
  assign new_n39770_ = ~new_n39767_ & ~new_n39769_;
  assign new_n39771_ = ~new_n39766_ & new_n39770_;
  assign new_n39772_ = new_n39699_ & ~new_n39771_;
  assign new_n39773_ = ~new_n39670_ & ~new_n39678_;
  assign new_n39774_ = ~new_n39686_ & ~new_n39694_;
  assign new_n39775_ = ~new_n39681_ & new_n39774_;
  assign new_n39776_ = ~new_n39773_ & ~new_n39775_;
  assign new_n39777_ = new_n39665_ & ~new_n39776_;
  assign new_n39778_ = ~new_n39637_ & ~new_n39645_;
  assign new_n39779_ = ~new_n39653_ & ~new_n39661_;
  assign new_n39780_ = ~new_n39648_ & new_n39779_;
  assign new_n39781_ = ~new_n39778_ & ~new_n39780_;
  assign new_n39782_ = ~new_n39777_ & new_n39781_;
  assign new_n39783_ = ~new_n39772_ & new_n39782_;
  assign new_n39784_ = ~new_n39761_ & new_n39783_;
  assign new_n39785_ = ~new_n39625_ & new_n39759_;
  assign new_n39786_ = new_n39771_ & ~new_n39785_;
  assign new_n39787_ = new_n39698_ & ~new_n39786_;
  assign new_n39788_ = new_n39776_ & ~new_n39787_;
  assign new_n39789_ = ~new_n39664_ & ~new_n39788_;
  assign new_n39790_ = ~new_n39779_ & ~new_n39789_;
  assign new_n39791_ = new_n39648_ & ~new_n39790_;
  assign new_n39792_ = ~new_n39648_ & new_n39790_;
  assign new_n39793_ = ~new_n39791_ & ~new_n39792_;
  assign new_n39794_ = ~new_n39625_ & new_n39758_;
  assign new_n39795_ = new_n39765_ & ~new_n39794_;
  assign new_n39796_ = ~new_n39731_ & ~new_n39795_;
  assign new_n39797_ = ~new_n39768_ & ~new_n39796_;
  assign new_n39798_ = new_n39715_ & ~new_n39797_;
  assign new_n39799_ = ~new_n39715_ & new_n39797_;
  assign new_n39800_ = ~new_n39798_ & ~new_n39799_;
  assign new_n39801_ = new_n39731_ & ~new_n39795_;
  assign new_n39802_ = ~new_n39731_ & new_n39795_;
  assign new_n39803_ = ~new_n39801_ & ~new_n39802_;
  assign new_n39804_ = ~new_n39625_ & ~new_n39757_;
  assign new_n39805_ = ~new_n39763_ & ~new_n39804_;
  assign new_n39806_ = new_n39745_ & ~new_n39805_;
  assign new_n39807_ = ~new_n39745_ & new_n39805_;
  assign new_n39808_ = ~new_n39806_ & ~new_n39807_;
  assign new_n39809_ = ~new_n39625_ & new_n39757_;
  assign new_n39810_ = new_n39625_ & ~new_n39757_;
  assign new_n39811_ = ~new_n39809_ & ~new_n39810_;
  assign new_n39812_ = ~new_n39808_ & ~new_n39811_;
  assign new_n39813_ = ~new_n39803_ & new_n39812_;
  assign new_n39814_ = ~new_n39800_ & new_n39813_;
  assign new_n39815_ = ~new_n39697_ & ~new_n39786_;
  assign new_n39816_ = ~new_n39774_ & ~new_n39815_;
  assign new_n39817_ = new_n39681_ & ~new_n39816_;
  assign new_n39818_ = ~new_n39681_ & new_n39816_;
  assign new_n39819_ = ~new_n39817_ & ~new_n39818_;
  assign new_n39820_ = new_n39697_ & ~new_n39786_;
  assign new_n39821_ = ~new_n39697_ & new_n39786_;
  assign new_n39822_ = ~new_n39820_ & ~new_n39821_;
  assign new_n39823_ = ~new_n39819_ & ~new_n39822_;
  assign new_n39824_ = new_n39664_ & ~new_n39788_;
  assign new_n39825_ = ~new_n39664_ & new_n39788_;
  assign new_n39826_ = ~new_n39824_ & ~new_n39825_;
  assign new_n39827_ = ~new_n39546_ & new_n39612_;
  assign new_n39828_ = new_n39618_ & ~new_n39827_;
  assign new_n39829_ = ~new_n39585_ & ~new_n39828_;
  assign new_n39830_ = ~new_n39621_ & ~new_n39829_;
  assign new_n39831_ = new_n39569_ & ~new_n39830_;
  assign new_n39832_ = ~new_n39569_ & new_n39830_;
  assign new_n39833_ = ~new_n39831_ & ~new_n39832_;
  assign new_n39834_ = ~new_n39546_ & ~new_n39611_;
  assign new_n39835_ = ~new_n39616_ & ~new_n39834_;
  assign new_n39836_ = new_n39599_ & ~new_n39835_;
  assign new_n39837_ = ~new_n39599_ & new_n39835_;
  assign new_n39838_ = ~new_n39836_ & ~new_n39837_;
  assign new_n39839_ = ~new_n39546_ & new_n39611_;
  assign new_n39840_ = new_n39546_ & ~new_n39611_;
  assign new_n39841_ = ~new_n39839_ & ~new_n39840_;
  assign new_n39842_ = ~new_n39838_ & ~new_n39841_;
  assign new_n39843_ = new_n39585_ & ~new_n39828_;
  assign new_n39844_ = ~new_n39585_ & new_n39828_;
  assign new_n39845_ = ~new_n39843_ & ~new_n39844_;
  assign new_n39846_ = ~new_n39507_ & ~new_n39539_;
  assign new_n39847_ = ~new_n39543_ & ~new_n39846_;
  assign new_n39848_ = new_n39527_ & ~new_n39847_;
  assign new_n39849_ = ~new_n39527_ & new_n39847_;
  assign new_n39850_ = ~new_n39848_ & ~new_n39849_;
  assign new_n39851_ = ~new_n39507_ & new_n39539_;
  assign new_n39852_ = new_n39507_ & ~new_n39539_;
  assign new_n39853_ = ~new_n39851_ & ~new_n39852_;
  assign new_n39854_ = new_n39494_ & new_n39505_;
  assign new_n39855_ = ~new_n39494_ & ~new_n39505_;
  assign new_n39856_ = ~new_n39854_ & ~new_n39855_;
  assign new_n39857_ = new_n39499_ & ~new_n39504_;
  assign new_n39858_ = ~new_n39499_ & new_n39504_;
  assign new_n39859_ = ~new_n39857_ & ~new_n39858_;
  assign new_n39860_ = ~ys__n30334 & ~new_n39859_;
  assign new_n39861_ = ~new_n39856_ & new_n39860_;
  assign new_n39862_ = ~new_n39853_ & new_n39861_;
  assign new_n39863_ = ~new_n39850_ & new_n39862_;
  assign new_n39864_ = ~new_n39845_ & new_n39863_;
  assign new_n39865_ = new_n39842_ & new_n39864_;
  assign new_n39866_ = ~new_n39833_ & new_n39865_;
  assign new_n39867_ = ~new_n39826_ & new_n39866_;
  assign new_n39868_ = new_n39823_ & new_n39867_;
  assign new_n39869_ = new_n39814_ & new_n39868_;
  assign new_n39870_ = ~new_n39793_ & new_n39869_;
  assign new_n39871_ = new_n39784_ & new_n39870_;
  assign new_n39872_ = ~new_n39784_ & ~new_n39870_;
  assign new_n39873_ = ~new_n39871_ & ~new_n39872_;
  assign new_n39874_ = ~ys__n17912 & ~ys__n30334;
  assign new_n39875_ = ys__n17912 & ys__n30334;
  assign new_n39876_ = ~new_n39874_ & ~new_n39875_;
  assign new_n39877_ = ~ys__n30333 & ~ys__n30334;
  assign new_n39878_ = ys__n30333 & ys__n30334;
  assign new_n39879_ = ~new_n39877_ & ~new_n39878_;
  assign new_n39880_ = ~ys__n17848 & ~new_n39879_;
  assign new_n39881_ = ys__n17848 & new_n39879_;
  assign new_n39882_ = ~new_n39880_ & ~new_n39881_;
  assign new_n39883_ = ~new_n39876_ & new_n39882_;
  assign new_n39884_ = new_n39876_ & ~new_n39882_;
  assign new_n39885_ = ~new_n39883_ & ~new_n39884_;
  assign new_n39886_ = ~ys__n17846 & ~new_n39876_;
  assign new_n39887_ = ~ys__n17911 & ~ys__n30334;
  assign new_n39888_ = ys__n17911 & ys__n30334;
  assign new_n39889_ = ~new_n39887_ & ~new_n39888_;
  assign new_n39890_ = new_n39886_ & ~new_n39889_;
  assign new_n39891_ = new_n39876_ & new_n39889_;
  assign new_n39892_ = ys__n17846 & ~new_n39891_;
  assign new_n39893_ = ~new_n39890_ & ~new_n39892_;
  assign new_n39894_ = new_n39885_ & ~new_n39893_;
  assign new_n39895_ = ~new_n39885_ & new_n39893_;
  assign new_n39896_ = ~new_n39894_ & ~new_n39895_;
  assign new_n39897_ = ys__n17846 & new_n39876_;
  assign new_n39898_ = ~new_n39886_ & ~new_n39897_;
  assign new_n39899_ = ~new_n39889_ & new_n39898_;
  assign new_n39900_ = new_n39889_ & ~new_n39898_;
  assign new_n39901_ = ~new_n39899_ & ~new_n39900_;
  assign new_n39902_ = ~ys__n17845 & ~new_n39889_;
  assign new_n39903_ = ~ys__n17909 & ~ys__n30334;
  assign new_n39904_ = ys__n17909 & ys__n30334;
  assign new_n39905_ = ~new_n39903_ & ~new_n39904_;
  assign new_n39906_ = new_n39902_ & ~new_n39905_;
  assign new_n39907_ = new_n39889_ & new_n39905_;
  assign new_n39908_ = ys__n17845 & ~new_n39907_;
  assign new_n39909_ = ~new_n39906_ & ~new_n39908_;
  assign new_n39910_ = ~new_n39901_ & ~new_n39909_;
  assign new_n39911_ = new_n39901_ & ~new_n39909_;
  assign new_n39912_ = ~new_n39901_ & new_n39909_;
  assign new_n39913_ = ~new_n39911_ & ~new_n39912_;
  assign new_n39914_ = ys__n17845 & new_n39889_;
  assign new_n39915_ = ~new_n39902_ & ~new_n39914_;
  assign new_n39916_ = ~new_n39905_ & new_n39915_;
  assign new_n39917_ = new_n39905_ & ~new_n39915_;
  assign new_n39918_ = ~new_n39916_ & ~new_n39917_;
  assign new_n39919_ = ~ys__n17843 & ~new_n39905_;
  assign new_n39920_ = ~ys__n17908 & ~ys__n30334;
  assign new_n39921_ = ys__n17908 & ys__n30334;
  assign new_n39922_ = ~new_n39920_ & ~new_n39921_;
  assign new_n39923_ = new_n39919_ & ~new_n39922_;
  assign new_n39924_ = new_n39905_ & new_n39922_;
  assign new_n39925_ = ys__n17843 & ~new_n39924_;
  assign new_n39926_ = ~new_n39923_ & ~new_n39925_;
  assign new_n39927_ = ~new_n39918_ & ~new_n39926_;
  assign new_n39928_ = new_n39918_ & ~new_n39926_;
  assign new_n39929_ = ~new_n39918_ & new_n39926_;
  assign new_n39930_ = ~new_n39928_ & ~new_n39929_;
  assign new_n39931_ = ys__n17843 & new_n39905_;
  assign new_n39932_ = ~new_n39919_ & ~new_n39931_;
  assign new_n39933_ = ~new_n39922_ & new_n39932_;
  assign new_n39934_ = new_n39922_ & ~new_n39932_;
  assign new_n39935_ = ~new_n39933_ & ~new_n39934_;
  assign new_n39936_ = ~ys__n17842 & ~new_n39922_;
  assign new_n39937_ = ~ys__n17906 & ~ys__n30334;
  assign new_n39938_ = ys__n17906 & ys__n30334;
  assign new_n39939_ = ~new_n39937_ & ~new_n39938_;
  assign new_n39940_ = new_n39936_ & ~new_n39939_;
  assign new_n39941_ = new_n39922_ & new_n39939_;
  assign new_n39942_ = ys__n17842 & ~new_n39941_;
  assign new_n39943_ = ~new_n39940_ & ~new_n39942_;
  assign new_n39944_ = ~new_n39935_ & ~new_n39943_;
  assign new_n39945_ = ~new_n39930_ & new_n39944_;
  assign new_n39946_ = ~new_n39927_ & ~new_n39945_;
  assign new_n39947_ = new_n39935_ & ~new_n39943_;
  assign new_n39948_ = ~new_n39935_ & new_n39943_;
  assign new_n39949_ = ~new_n39947_ & ~new_n39948_;
  assign new_n39950_ = ~new_n39930_ & ~new_n39949_;
  assign new_n39951_ = ys__n17842 & new_n39922_;
  assign new_n39952_ = ~new_n39936_ & ~new_n39951_;
  assign new_n39953_ = ~new_n39939_ & new_n39952_;
  assign new_n39954_ = new_n39939_ & ~new_n39952_;
  assign new_n39955_ = ~new_n39953_ & ~new_n39954_;
  assign new_n39956_ = ~ys__n17840 & ~new_n39939_;
  assign new_n39957_ = ~ys__n17905 & ~ys__n30334;
  assign new_n39958_ = ys__n17905 & ys__n30334;
  assign new_n39959_ = ~new_n39957_ & ~new_n39958_;
  assign new_n39960_ = new_n39956_ & ~new_n39959_;
  assign new_n39961_ = new_n39939_ & new_n39959_;
  assign new_n39962_ = ys__n17840 & ~new_n39961_;
  assign new_n39963_ = ~new_n39960_ & ~new_n39962_;
  assign new_n39964_ = new_n39955_ & ~new_n39963_;
  assign new_n39965_ = ~new_n39955_ & new_n39963_;
  assign new_n39966_ = ~new_n39964_ & ~new_n39965_;
  assign new_n39967_ = ys__n17840 & new_n39939_;
  assign new_n39968_ = ~new_n39956_ & ~new_n39967_;
  assign new_n39969_ = ~new_n39959_ & new_n39968_;
  assign new_n39970_ = new_n39959_ & ~new_n39968_;
  assign new_n39971_ = ~new_n39969_ & ~new_n39970_;
  assign new_n39972_ = ~ys__n17839 & ~new_n39959_;
  assign new_n39973_ = ~ys__n17903 & ~ys__n30334;
  assign new_n39974_ = ys__n17903 & ys__n30334;
  assign new_n39975_ = ~new_n39973_ & ~new_n39974_;
  assign new_n39976_ = new_n39972_ & ~new_n39975_;
  assign new_n39977_ = new_n39959_ & new_n39975_;
  assign new_n39978_ = ys__n17839 & ~new_n39977_;
  assign new_n39979_ = ~new_n39976_ & ~new_n39978_;
  assign new_n39980_ = new_n39971_ & ~new_n39979_;
  assign new_n39981_ = ~new_n39971_ & new_n39979_;
  assign new_n39982_ = ~new_n39980_ & ~new_n39981_;
  assign new_n39983_ = ~new_n39966_ & ~new_n39982_;
  assign new_n39984_ = ys__n17839 & new_n39959_;
  assign new_n39985_ = ~new_n39972_ & ~new_n39984_;
  assign new_n39986_ = ~new_n39975_ & new_n39985_;
  assign new_n39987_ = new_n39975_ & ~new_n39985_;
  assign new_n39988_ = ~new_n39986_ & ~new_n39987_;
  assign new_n39989_ = ~ys__n17837 & ~new_n39975_;
  assign new_n39990_ = ~ys__n17902 & ~ys__n30334;
  assign new_n39991_ = ys__n17902 & ys__n30334;
  assign new_n39992_ = ~new_n39990_ & ~new_n39991_;
  assign new_n39993_ = new_n39989_ & ~new_n39992_;
  assign new_n39994_ = new_n39975_ & new_n39992_;
  assign new_n39995_ = ys__n17837 & ~new_n39994_;
  assign new_n39996_ = ~new_n39993_ & ~new_n39995_;
  assign new_n39997_ = ~new_n39988_ & ~new_n39996_;
  assign new_n39998_ = new_n39988_ & ~new_n39996_;
  assign new_n39999_ = ~new_n39988_ & new_n39996_;
  assign new_n40000_ = ~new_n39998_ & ~new_n39999_;
  assign new_n40001_ = ys__n17837 & new_n39975_;
  assign new_n40002_ = ~new_n39989_ & ~new_n40001_;
  assign new_n40003_ = ~new_n39992_ & new_n40002_;
  assign new_n40004_ = new_n39992_ & ~new_n40002_;
  assign new_n40005_ = ~new_n40003_ & ~new_n40004_;
  assign new_n40006_ = ~ys__n17836 & ~new_n39992_;
  assign new_n40007_ = ~ys__n17900 & ~ys__n30334;
  assign new_n40008_ = ys__n17900 & ys__n30334;
  assign new_n40009_ = ~new_n40007_ & ~new_n40008_;
  assign new_n40010_ = new_n40006_ & ~new_n40009_;
  assign new_n40011_ = new_n39992_ & new_n40009_;
  assign new_n40012_ = ys__n17836 & ~new_n40011_;
  assign new_n40013_ = ~new_n40010_ & ~new_n40012_;
  assign new_n40014_ = ~new_n40005_ & ~new_n40013_;
  assign new_n40015_ = ~new_n40000_ & new_n40014_;
  assign new_n40016_ = ~new_n39997_ & ~new_n40015_;
  assign new_n40017_ = new_n39983_ & ~new_n40016_;
  assign new_n40018_ = ~new_n39955_ & ~new_n39963_;
  assign new_n40019_ = ~new_n39971_ & ~new_n39979_;
  assign new_n40020_ = ~new_n39966_ & new_n40019_;
  assign new_n40021_ = ~new_n40018_ & ~new_n40020_;
  assign new_n40022_ = ~new_n40017_ & new_n40021_;
  assign new_n40023_ = new_n40005_ & ~new_n40013_;
  assign new_n40024_ = ~new_n40005_ & new_n40013_;
  assign new_n40025_ = ~new_n40023_ & ~new_n40024_;
  assign new_n40026_ = ~new_n40000_ & ~new_n40025_;
  assign new_n40027_ = new_n39983_ & new_n40026_;
  assign new_n40028_ = ~ys__n17891 & ~ys__n30334;
  assign new_n40029_ = ys__n17891 & ys__n30334;
  assign new_n40030_ = ~new_n40028_ & ~new_n40029_;
  assign new_n40031_ = ~ys__n17893 & ~ys__n30334;
  assign new_n40032_ = ys__n17893 & ys__n30334;
  assign new_n40033_ = ~new_n40031_ & ~new_n40032_;
  assign new_n40034_ = ~ys__n17827 & ~new_n40033_;
  assign new_n40035_ = ys__n17827 & new_n40033_;
  assign new_n40036_ = ~new_n40034_ & ~new_n40035_;
  assign new_n40037_ = ~new_n40030_ & new_n40036_;
  assign new_n40038_ = new_n40030_ & ~new_n40036_;
  assign new_n40039_ = ~new_n40037_ & ~new_n40038_;
  assign new_n40040_ = ~ys__n17825 & ~new_n40030_;
  assign new_n40041_ = ~new_n39631_ & new_n40040_;
  assign new_n40042_ = new_n39631_ & new_n40030_;
  assign new_n40043_ = ys__n17825 & ~new_n40042_;
  assign new_n40044_ = ~new_n40041_ & ~new_n40043_;
  assign new_n40045_ = ~new_n40039_ & ~new_n40044_;
  assign new_n40046_ = new_n40039_ & ~new_n40044_;
  assign new_n40047_ = ~new_n40039_ & new_n40044_;
  assign new_n40048_ = ~new_n40046_ & ~new_n40047_;
  assign new_n40049_ = ys__n17825 & new_n40030_;
  assign new_n40050_ = ~new_n40040_ & ~new_n40049_;
  assign new_n40051_ = ~new_n39631_ & new_n40050_;
  assign new_n40052_ = new_n39631_ & ~new_n40050_;
  assign new_n40053_ = ~new_n40051_ & ~new_n40052_;
  assign new_n40054_ = ~new_n39628_ & new_n39632_;
  assign new_n40055_ = new_n39628_ & new_n39631_;
  assign new_n40056_ = ys__n17824 & ~new_n40055_;
  assign new_n40057_ = ~new_n40054_ & ~new_n40056_;
  assign new_n40058_ = ~new_n40053_ & ~new_n40057_;
  assign new_n40059_ = ~new_n40048_ & new_n40058_;
  assign new_n40060_ = ~new_n40045_ & ~new_n40059_;
  assign new_n40061_ = ~ys__n17894 & ~ys__n30334;
  assign new_n40062_ = ys__n17894 & ys__n30334;
  assign new_n40063_ = ~new_n40061_ & ~new_n40062_;
  assign new_n40064_ = ~ys__n17896 & ~ys__n30334;
  assign new_n40065_ = ys__n17896 & ys__n30334;
  assign new_n40066_ = ~new_n40064_ & ~new_n40065_;
  assign new_n40067_ = ~ys__n17830 & ~new_n40066_;
  assign new_n40068_ = ys__n17830 & new_n40066_;
  assign new_n40069_ = ~new_n40067_ & ~new_n40068_;
  assign new_n40070_ = ~new_n40063_ & new_n40069_;
  assign new_n40071_ = new_n40063_ & ~new_n40069_;
  assign new_n40072_ = ~new_n40070_ & ~new_n40071_;
  assign new_n40073_ = ~ys__n17828 & ~new_n40063_;
  assign new_n40074_ = ~new_n40033_ & new_n40073_;
  assign new_n40075_ = new_n40033_ & new_n40063_;
  assign new_n40076_ = ys__n17828 & ~new_n40075_;
  assign new_n40077_ = ~new_n40074_ & ~new_n40076_;
  assign new_n40078_ = new_n40072_ & ~new_n40077_;
  assign new_n40079_ = ~new_n40072_ & new_n40077_;
  assign new_n40080_ = ~new_n40078_ & ~new_n40079_;
  assign new_n40081_ = ys__n17828 & new_n40063_;
  assign new_n40082_ = ~new_n40073_ & ~new_n40081_;
  assign new_n40083_ = ~new_n40033_ & new_n40082_;
  assign new_n40084_ = new_n40033_ & ~new_n40082_;
  assign new_n40085_ = ~new_n40083_ & ~new_n40084_;
  assign new_n40086_ = ~new_n40030_ & new_n40034_;
  assign new_n40087_ = new_n40030_ & new_n40033_;
  assign new_n40088_ = ys__n17827 & ~new_n40087_;
  assign new_n40089_ = ~new_n40086_ & ~new_n40088_;
  assign new_n40090_ = new_n40085_ & ~new_n40089_;
  assign new_n40091_ = ~new_n40085_ & new_n40089_;
  assign new_n40092_ = ~new_n40090_ & ~new_n40091_;
  assign new_n40093_ = ~new_n40080_ & ~new_n40092_;
  assign new_n40094_ = ~new_n40060_ & new_n40093_;
  assign new_n40095_ = ~new_n40072_ & ~new_n40077_;
  assign new_n40096_ = ~new_n40085_ & ~new_n40089_;
  assign new_n40097_ = ~new_n40080_ & new_n40096_;
  assign new_n40098_ = ~new_n40095_ & ~new_n40097_;
  assign new_n40099_ = ~new_n40094_ & new_n40098_;
  assign new_n40100_ = ys__n17836 & new_n39992_;
  assign new_n40101_ = ~new_n40006_ & ~new_n40100_;
  assign new_n40102_ = ~new_n40009_ & new_n40101_;
  assign new_n40103_ = new_n40009_ & ~new_n40101_;
  assign new_n40104_ = ~new_n40102_ & ~new_n40103_;
  assign new_n40105_ = ~ys__n17834 & ~new_n40009_;
  assign new_n40106_ = ~ys__n17899 & ~ys__n30334;
  assign new_n40107_ = ys__n17899 & ys__n30334;
  assign new_n40108_ = ~new_n40106_ & ~new_n40107_;
  assign new_n40109_ = new_n40105_ & ~new_n40108_;
  assign new_n40110_ = new_n40009_ & new_n40108_;
  assign new_n40111_ = ys__n17834 & ~new_n40110_;
  assign new_n40112_ = ~new_n40109_ & ~new_n40111_;
  assign new_n40113_ = new_n40104_ & ~new_n40112_;
  assign new_n40114_ = ~new_n40104_ & new_n40112_;
  assign new_n40115_ = ~new_n40113_ & ~new_n40114_;
  assign new_n40116_ = ys__n17834 & new_n40009_;
  assign new_n40117_ = ~new_n40105_ & ~new_n40116_;
  assign new_n40118_ = ~new_n40108_ & new_n40117_;
  assign new_n40119_ = new_n40108_ & ~new_n40117_;
  assign new_n40120_ = ~new_n40118_ & ~new_n40119_;
  assign new_n40121_ = ~ys__n17833 & ~new_n40108_;
  assign new_n40122_ = ~ys__n17897 & ~ys__n30334;
  assign new_n40123_ = ys__n17897 & ys__n30334;
  assign new_n40124_ = ~new_n40122_ & ~new_n40123_;
  assign new_n40125_ = new_n40121_ & ~new_n40124_;
  assign new_n40126_ = new_n40108_ & new_n40124_;
  assign new_n40127_ = ys__n17833 & ~new_n40126_;
  assign new_n40128_ = ~new_n40125_ & ~new_n40127_;
  assign new_n40129_ = new_n40120_ & ~new_n40128_;
  assign new_n40130_ = ~new_n40120_ & new_n40128_;
  assign new_n40131_ = ~new_n40129_ & ~new_n40130_;
  assign new_n40132_ = ~new_n40115_ & ~new_n40131_;
  assign new_n40133_ = ys__n17833 & new_n40108_;
  assign new_n40134_ = ~new_n40121_ & ~new_n40133_;
  assign new_n40135_ = ~new_n40124_ & new_n40134_;
  assign new_n40136_ = new_n40124_ & ~new_n40134_;
  assign new_n40137_ = ~new_n40135_ & ~new_n40136_;
  assign new_n40138_ = ~ys__n17831 & ~new_n40124_;
  assign new_n40139_ = ~new_n40066_ & new_n40138_;
  assign new_n40140_ = new_n40066_ & new_n40124_;
  assign new_n40141_ = ys__n17831 & ~new_n40140_;
  assign new_n40142_ = ~new_n40139_ & ~new_n40141_;
  assign new_n40143_ = new_n40137_ & ~new_n40142_;
  assign new_n40144_ = ~new_n40137_ & new_n40142_;
  assign new_n40145_ = ~new_n40143_ & ~new_n40144_;
  assign new_n40146_ = ys__n17831 & new_n40124_;
  assign new_n40147_ = ~new_n40138_ & ~new_n40146_;
  assign new_n40148_ = ~new_n40066_ & new_n40147_;
  assign new_n40149_ = new_n40066_ & ~new_n40147_;
  assign new_n40150_ = ~new_n40148_ & ~new_n40149_;
  assign new_n40151_ = ~new_n40063_ & new_n40067_;
  assign new_n40152_ = new_n40063_ & new_n40066_;
  assign new_n40153_ = ys__n17830 & ~new_n40152_;
  assign new_n40154_ = ~new_n40151_ & ~new_n40153_;
  assign new_n40155_ = new_n40150_ & ~new_n40154_;
  assign new_n40156_ = ~new_n40150_ & new_n40154_;
  assign new_n40157_ = ~new_n40155_ & ~new_n40156_;
  assign new_n40158_ = ~new_n40145_ & ~new_n40157_;
  assign new_n40159_ = new_n40132_ & new_n40158_;
  assign new_n40160_ = ~new_n40099_ & new_n40159_;
  assign new_n40161_ = ~new_n40137_ & ~new_n40142_;
  assign new_n40162_ = ~new_n40150_ & ~new_n40154_;
  assign new_n40163_ = ~new_n40145_ & new_n40162_;
  assign new_n40164_ = ~new_n40161_ & ~new_n40163_;
  assign new_n40165_ = new_n40132_ & ~new_n40164_;
  assign new_n40166_ = ~new_n40104_ & ~new_n40112_;
  assign new_n40167_ = ~new_n40120_ & ~new_n40128_;
  assign new_n40168_ = ~new_n40115_ & new_n40167_;
  assign new_n40169_ = ~new_n40166_ & ~new_n40168_;
  assign new_n40170_ = ~new_n40165_ & new_n40169_;
  assign new_n40171_ = ~new_n40160_ & new_n40170_;
  assign new_n40172_ = new_n40027_ & ~new_n40171_;
  assign new_n40173_ = new_n40022_ & ~new_n40172_;
  assign new_n40174_ = new_n39950_ & ~new_n40173_;
  assign new_n40175_ = new_n39946_ & ~new_n40174_;
  assign new_n40176_ = ~new_n39913_ & ~new_n40175_;
  assign new_n40177_ = ~new_n39910_ & ~new_n40176_;
  assign new_n40178_ = new_n39896_ & ~new_n40177_;
  assign new_n40179_ = ~new_n39896_ & new_n40177_;
  assign new_n40180_ = ~new_n40178_ & ~new_n40179_;
  assign new_n40181_ = new_n39873_ & ~new_n40180_;
  assign new_n40182_ = new_n39913_ & ~new_n40175_;
  assign new_n40183_ = ~new_n39913_ & new_n40175_;
  assign new_n40184_ = ~new_n40182_ & ~new_n40183_;
  assign new_n40185_ = ~new_n39949_ & ~new_n40173_;
  assign new_n40186_ = ~new_n39944_ & ~new_n40185_;
  assign new_n40187_ = new_n39930_ & ~new_n40186_;
  assign new_n40188_ = ~new_n39930_ & new_n40186_;
  assign new_n40189_ = ~new_n40187_ & ~new_n40188_;
  assign new_n40190_ = new_n39949_ & ~new_n40173_;
  assign new_n40191_ = ~new_n39949_ & new_n40173_;
  assign new_n40192_ = ~new_n40190_ & ~new_n40191_;
  assign new_n40193_ = ~new_n40189_ & ~new_n40192_;
  assign new_n40194_ = new_n40026_ & ~new_n40171_;
  assign new_n40195_ = new_n40016_ & ~new_n40194_;
  assign new_n40196_ = ~new_n39982_ & ~new_n40195_;
  assign new_n40197_ = ~new_n40019_ & ~new_n40196_;
  assign new_n40198_ = new_n39966_ & ~new_n40197_;
  assign new_n40199_ = ~new_n39966_ & new_n40197_;
  assign new_n40200_ = ~new_n40198_ & ~new_n40199_;
  assign new_n40201_ = new_n39982_ & ~new_n40195_;
  assign new_n40202_ = ~new_n39982_ & new_n40195_;
  assign new_n40203_ = ~new_n40201_ & ~new_n40202_;
  assign new_n40204_ = ~new_n40025_ & ~new_n40171_;
  assign new_n40205_ = ~new_n40014_ & ~new_n40204_;
  assign new_n40206_ = new_n40000_ & ~new_n40205_;
  assign new_n40207_ = ~new_n40000_ & new_n40205_;
  assign new_n40208_ = ~new_n40206_ & ~new_n40207_;
  assign new_n40209_ = new_n40025_ & ~new_n40171_;
  assign new_n40210_ = ~new_n40025_ & new_n40171_;
  assign new_n40211_ = ~new_n40209_ & ~new_n40210_;
  assign new_n40212_ = ~new_n40208_ & ~new_n40211_;
  assign new_n40213_ = ~new_n40203_ & new_n40212_;
  assign new_n40214_ = ~new_n40200_ & new_n40213_;
  assign new_n40215_ = ~new_n40099_ & new_n40158_;
  assign new_n40216_ = new_n40164_ & ~new_n40215_;
  assign new_n40217_ = ~new_n40131_ & ~new_n40216_;
  assign new_n40218_ = ~new_n40167_ & ~new_n40217_;
  assign new_n40219_ = new_n40115_ & ~new_n40218_;
  assign new_n40220_ = ~new_n40115_ & new_n40218_;
  assign new_n40221_ = ~new_n40219_ & ~new_n40220_;
  assign new_n40222_ = ~new_n40099_ & ~new_n40157_;
  assign new_n40223_ = ~new_n40162_ & ~new_n40222_;
  assign new_n40224_ = new_n40145_ & ~new_n40223_;
  assign new_n40225_ = ~new_n40145_ & new_n40223_;
  assign new_n40226_ = ~new_n40224_ & ~new_n40225_;
  assign new_n40227_ = ~new_n40099_ & new_n40157_;
  assign new_n40228_ = new_n40099_ & ~new_n40157_;
  assign new_n40229_ = ~new_n40227_ & ~new_n40228_;
  assign new_n40230_ = ~new_n40226_ & ~new_n40229_;
  assign new_n40231_ = new_n40131_ & ~new_n40216_;
  assign new_n40232_ = ~new_n40131_ & new_n40216_;
  assign new_n40233_ = ~new_n40231_ & ~new_n40232_;
  assign new_n40234_ = ~new_n40060_ & ~new_n40092_;
  assign new_n40235_ = ~new_n40096_ & ~new_n40234_;
  assign new_n40236_ = new_n40080_ & ~new_n40235_;
  assign new_n40237_ = ~new_n40080_ & new_n40235_;
  assign new_n40238_ = ~new_n40236_ & ~new_n40237_;
  assign new_n40239_ = ~new_n40060_ & new_n40092_;
  assign new_n40240_ = new_n40060_ & ~new_n40092_;
  assign new_n40241_ = ~new_n40239_ & ~new_n40240_;
  assign new_n40242_ = new_n40048_ & new_n40058_;
  assign new_n40243_ = ~new_n40048_ & ~new_n40058_;
  assign new_n40244_ = ~new_n40242_ & ~new_n40243_;
  assign new_n40245_ = new_n40053_ & ~new_n40057_;
  assign new_n40246_ = ~new_n40053_ & new_n40057_;
  assign new_n40247_ = ~new_n40245_ & ~new_n40246_;
  assign new_n40248_ = ~new_n40244_ & ~new_n40247_;
  assign new_n40249_ = ~new_n40241_ & new_n40248_;
  assign new_n40250_ = ~new_n40238_ & new_n40249_;
  assign new_n40251_ = ~new_n40233_ & new_n40250_;
  assign new_n40252_ = new_n40230_ & new_n40251_;
  assign new_n40253_ = ~new_n40221_ & new_n40252_;
  assign new_n40254_ = new_n40214_ & new_n40253_;
  assign new_n40255_ = new_n40193_ & new_n40254_;
  assign new_n40256_ = ~new_n40184_ & new_n40255_;
  assign new_n40257_ = new_n40180_ & new_n40256_;
  assign new_n40258_ = ~new_n40180_ & ~new_n40256_;
  assign new_n40259_ = ~new_n40257_ & ~new_n40258_;
  assign new_n40260_ = ~new_n39873_ & ~new_n40259_;
  assign new_n40261_ = ~new_n40181_ & ~new_n40260_;
  assign new_n40262_ = ys__n18156 & ~new_n40261_;
  assign new_n40263_ = ~ys__n17849 & ~new_n39879_;
  assign new_n40264_ = ys__n17849 & new_n39879_;
  assign new_n40265_ = ~new_n40263_ & ~new_n40264_;
  assign new_n40266_ = ~new_n39879_ & new_n40265_;
  assign new_n40267_ = new_n39879_ & ~new_n40265_;
  assign new_n40268_ = ~new_n40266_ & ~new_n40267_;
  assign new_n40269_ = ~new_n39876_ & new_n39880_;
  assign new_n40270_ = new_n39876_ & new_n39879_;
  assign new_n40271_ = ys__n17848 & ~new_n40270_;
  assign new_n40272_ = ~new_n40269_ & ~new_n40271_;
  assign new_n40273_ = new_n40268_ & ~new_n40272_;
  assign new_n40274_ = ~new_n40268_ & new_n40272_;
  assign new_n40275_ = ~new_n40273_ & ~new_n40274_;
  assign new_n40276_ = ~new_n39896_ & ~new_n39913_;
  assign new_n40277_ = new_n39950_ & new_n40276_;
  assign new_n40278_ = new_n40027_ & new_n40277_;
  assign new_n40279_ = ~new_n40171_ & new_n40278_;
  assign new_n40280_ = ~new_n40022_ & new_n40277_;
  assign new_n40281_ = ~new_n39946_ & new_n40276_;
  assign new_n40282_ = ~new_n39885_ & ~new_n39893_;
  assign new_n40283_ = ~new_n39896_ & new_n39910_;
  assign new_n40284_ = ~new_n40282_ & ~new_n40283_;
  assign new_n40285_ = ~new_n40281_ & new_n40284_;
  assign new_n40286_ = ~new_n40280_ & new_n40285_;
  assign new_n40287_ = ~new_n40279_ & new_n40286_;
  assign new_n40288_ = new_n40275_ & ~new_n40287_;
  assign new_n40289_ = ~new_n40275_ & new_n40287_;
  assign new_n40290_ = ~new_n40288_ & ~new_n40289_;
  assign new_n40291_ = new_n39873_ & ~new_n40290_;
  assign new_n40292_ = ~new_n40184_ & new_n40253_;
  assign new_n40293_ = new_n40193_ & new_n40292_;
  assign new_n40294_ = new_n40214_ & new_n40293_;
  assign new_n40295_ = ~new_n40180_ & new_n40294_;
  assign new_n40296_ = new_n40290_ & new_n40295_;
  assign new_n40297_ = ~new_n40290_ & ~new_n40295_;
  assign new_n40298_ = ~new_n40296_ & ~new_n40297_;
  assign new_n40299_ = ~new_n39873_ & ~new_n40298_;
  assign new_n40300_ = ~new_n40291_ & ~new_n40299_;
  assign new_n40301_ = ~new_n40262_ & new_n40300_;
  assign new_n40302_ = ys__n33581 & ~new_n39486_;
  assign new_n40303_ = ~ys__n33581 & ~new_n39486_;
  assign new_n40304_ = ys__n33581 & new_n39486_;
  assign new_n40305_ = ~new_n40303_ & ~new_n40304_;
  assign new_n40306_ = ~ys__n30334 & ys__n33579;
  assign new_n40307_ = ~new_n40305_ & new_n40306_;
  assign new_n40308_ = ~new_n40302_ & ~new_n40307_;
  assign new_n40309_ = ~ys__n17804 & ~new_n39476_;
  assign new_n40310_ = ys__n17804 & new_n39476_;
  assign new_n40311_ = ~new_n40309_ & ~new_n40310_;
  assign new_n40312_ = ~ys__n17803 & ~new_n39473_;
  assign new_n40313_ = ys__n17803 & new_n39473_;
  assign new_n40314_ = ~new_n40312_ & ~new_n40313_;
  assign new_n40315_ = ~new_n40311_ & ~new_n40314_;
  assign new_n40316_ = ~new_n40308_ & new_n40315_;
  assign new_n40317_ = ys__n17804 & ~new_n39476_;
  assign new_n40318_ = ys__n17803 & ~new_n39473_;
  assign new_n40319_ = ~new_n40311_ & new_n40318_;
  assign new_n40320_ = ~new_n40317_ & ~new_n40319_;
  assign new_n40321_ = ~new_n40316_ & new_n40320_;
  assign new_n40322_ = ~ys__n17810 & ~new_n39562_;
  assign new_n40323_ = ys__n17810 & new_n39562_;
  assign new_n40324_ = ~new_n40322_ & ~new_n40323_;
  assign new_n40325_ = ~ys__n17809 & ~new_n39578_;
  assign new_n40326_ = ys__n17809 & new_n39578_;
  assign new_n40327_ = ~new_n40325_ & ~new_n40326_;
  assign new_n40328_ = ~new_n40324_ & ~new_n40327_;
  assign new_n40329_ = ~ys__n17807 & ~new_n39513_;
  assign new_n40330_ = ys__n17807 & new_n39513_;
  assign new_n40331_ = ~new_n40329_ & ~new_n40330_;
  assign new_n40332_ = ~ys__n17806 & ~new_n39510_;
  assign new_n40333_ = ys__n17806 & new_n39510_;
  assign new_n40334_ = ~new_n40332_ & ~new_n40333_;
  assign new_n40335_ = ~new_n40331_ & ~new_n40334_;
  assign new_n40336_ = new_n40328_ & new_n40335_;
  assign new_n40337_ = ~new_n40321_ & new_n40336_;
  assign new_n40338_ = ys__n17807 & ~new_n39513_;
  assign new_n40339_ = ys__n17806 & ~new_n39510_;
  assign new_n40340_ = ~new_n40331_ & new_n40339_;
  assign new_n40341_ = ~new_n40338_ & ~new_n40340_;
  assign new_n40342_ = new_n40328_ & ~new_n40341_;
  assign new_n40343_ = ys__n17810 & ~new_n39562_;
  assign new_n40344_ = ys__n17809 & ~new_n39578_;
  assign new_n40345_ = ~new_n40324_ & new_n40344_;
  assign new_n40346_ = ~new_n40343_ & ~new_n40345_;
  assign new_n40347_ = ~new_n40342_ & new_n40346_;
  assign new_n40348_ = ~new_n40337_ & new_n40347_;
  assign new_n40349_ = ~ys__n17822 & ~new_n39641_;
  assign new_n40350_ = ys__n17822 & new_n39641_;
  assign new_n40351_ = ~new_n40349_ & ~new_n40350_;
  assign new_n40352_ = ~ys__n17821 & ~new_n39657_;
  assign new_n40353_ = ys__n17821 & new_n39657_;
  assign new_n40354_ = ~new_n40352_ & ~new_n40353_;
  assign new_n40355_ = ~new_n40351_ & ~new_n40354_;
  assign new_n40356_ = ~ys__n17819 & ~new_n39674_;
  assign new_n40357_ = ys__n17819 & new_n39674_;
  assign new_n40358_ = ~new_n40356_ & ~new_n40357_;
  assign new_n40359_ = ~ys__n17818 & ~new_n39690_;
  assign new_n40360_ = ys__n17818 & new_n39690_;
  assign new_n40361_ = ~new_n40359_ & ~new_n40360_;
  assign new_n40362_ = ~new_n40358_ & ~new_n40361_;
  assign new_n40363_ = new_n40355_ & new_n40362_;
  assign new_n40364_ = ~ys__n17816 & ~new_n39708_;
  assign new_n40365_ = ys__n17816 & new_n39708_;
  assign new_n40366_ = ~new_n40364_ & ~new_n40365_;
  assign new_n40367_ = ~ys__n17815 & ~new_n39724_;
  assign new_n40368_ = ys__n17815 & new_n39724_;
  assign new_n40369_ = ~new_n40367_ & ~new_n40368_;
  assign new_n40370_ = ~new_n40366_ & ~new_n40369_;
  assign new_n40371_ = ~ys__n17813 & ~new_n39552_;
  assign new_n40372_ = ys__n17813 & new_n39552_;
  assign new_n40373_ = ~new_n40371_ & ~new_n40372_;
  assign new_n40374_ = ~ys__n17812 & ~new_n39549_;
  assign new_n40375_ = ys__n17812 & new_n39549_;
  assign new_n40376_ = ~new_n40374_ & ~new_n40375_;
  assign new_n40377_ = ~new_n40373_ & ~new_n40376_;
  assign new_n40378_ = new_n40370_ & new_n40377_;
  assign new_n40379_ = new_n40363_ & new_n40378_;
  assign new_n40380_ = ~new_n40348_ & new_n40379_;
  assign new_n40381_ = ys__n17813 & ~new_n39552_;
  assign new_n40382_ = ys__n17812 & ~new_n39549_;
  assign new_n40383_ = ~new_n40373_ & new_n40382_;
  assign new_n40384_ = ~new_n40381_ & ~new_n40383_;
  assign new_n40385_ = new_n40370_ & ~new_n40384_;
  assign new_n40386_ = ys__n17816 & ~new_n39708_;
  assign new_n40387_ = ys__n17815 & ~new_n39724_;
  assign new_n40388_ = ~new_n40366_ & new_n40387_;
  assign new_n40389_ = ~new_n40386_ & ~new_n40388_;
  assign new_n40390_ = ~new_n40385_ & new_n40389_;
  assign new_n40391_ = new_n40363_ & ~new_n40390_;
  assign new_n40392_ = ys__n17819 & ~new_n39674_;
  assign new_n40393_ = ys__n17818 & ~new_n39690_;
  assign new_n40394_ = ~new_n40358_ & new_n40393_;
  assign new_n40395_ = ~new_n40392_ & ~new_n40394_;
  assign new_n40396_ = new_n40355_ & ~new_n40395_;
  assign new_n40397_ = ys__n17822 & ~new_n39641_;
  assign new_n40398_ = ys__n17821 & ~new_n39657_;
  assign new_n40399_ = ~new_n40351_ & new_n40398_;
  assign new_n40400_ = ~new_n40397_ & ~new_n40399_;
  assign new_n40401_ = ~new_n40396_ & new_n40400_;
  assign new_n40402_ = ~new_n40391_ & new_n40401_;
  assign new_n40403_ = ~new_n40380_ & new_n40402_;
  assign new_n40404_ = ~new_n40348_ & new_n40378_;
  assign new_n40405_ = new_n40390_ & ~new_n40404_;
  assign new_n40406_ = new_n40362_ & ~new_n40405_;
  assign new_n40407_ = new_n40395_ & ~new_n40406_;
  assign new_n40408_ = ~new_n40354_ & ~new_n40407_;
  assign new_n40409_ = ~new_n40398_ & ~new_n40408_;
  assign new_n40410_ = new_n40351_ & ~new_n40409_;
  assign new_n40411_ = ~new_n40351_ & new_n40409_;
  assign new_n40412_ = ~new_n40410_ & ~new_n40411_;
  assign new_n40413_ = ~new_n40348_ & new_n40377_;
  assign new_n40414_ = new_n40384_ & ~new_n40413_;
  assign new_n40415_ = ~new_n40369_ & ~new_n40414_;
  assign new_n40416_ = ~new_n40387_ & ~new_n40415_;
  assign new_n40417_ = new_n40366_ & ~new_n40416_;
  assign new_n40418_ = ~new_n40366_ & new_n40416_;
  assign new_n40419_ = ~new_n40417_ & ~new_n40418_;
  assign new_n40420_ = new_n40369_ & ~new_n40414_;
  assign new_n40421_ = ~new_n40369_ & new_n40414_;
  assign new_n40422_ = ~new_n40420_ & ~new_n40421_;
  assign new_n40423_ = ~new_n40348_ & ~new_n40376_;
  assign new_n40424_ = ~new_n40382_ & ~new_n40423_;
  assign new_n40425_ = new_n40373_ & ~new_n40424_;
  assign new_n40426_ = ~new_n40373_ & new_n40424_;
  assign new_n40427_ = ~new_n40425_ & ~new_n40426_;
  assign new_n40428_ = ~new_n40348_ & new_n40376_;
  assign new_n40429_ = new_n40348_ & ~new_n40376_;
  assign new_n40430_ = ~new_n40428_ & ~new_n40429_;
  assign new_n40431_ = ~new_n40427_ & ~new_n40430_;
  assign new_n40432_ = ~new_n40422_ & new_n40431_;
  assign new_n40433_ = ~new_n40419_ & new_n40432_;
  assign new_n40434_ = ~new_n40361_ & ~new_n40405_;
  assign new_n40435_ = ~new_n40393_ & ~new_n40434_;
  assign new_n40436_ = new_n40358_ & ~new_n40435_;
  assign new_n40437_ = ~new_n40358_ & new_n40435_;
  assign new_n40438_ = ~new_n40436_ & ~new_n40437_;
  assign new_n40439_ = new_n40361_ & ~new_n40405_;
  assign new_n40440_ = ~new_n40361_ & new_n40405_;
  assign new_n40441_ = ~new_n40439_ & ~new_n40440_;
  assign new_n40442_ = ~new_n40438_ & ~new_n40441_;
  assign new_n40443_ = new_n40354_ & ~new_n40407_;
  assign new_n40444_ = ~new_n40354_ & new_n40407_;
  assign new_n40445_ = ~new_n40443_ & ~new_n40444_;
  assign new_n40446_ = ~new_n40321_ & new_n40335_;
  assign new_n40447_ = new_n40341_ & ~new_n40446_;
  assign new_n40448_ = ~new_n40327_ & ~new_n40447_;
  assign new_n40449_ = ~new_n40344_ & ~new_n40448_;
  assign new_n40450_ = new_n40324_ & ~new_n40449_;
  assign new_n40451_ = ~new_n40324_ & new_n40449_;
  assign new_n40452_ = ~new_n40450_ & ~new_n40451_;
  assign new_n40453_ = ~new_n40321_ & ~new_n40334_;
  assign new_n40454_ = ~new_n40339_ & ~new_n40453_;
  assign new_n40455_ = new_n40331_ & ~new_n40454_;
  assign new_n40456_ = ~new_n40331_ & new_n40454_;
  assign new_n40457_ = ~new_n40455_ & ~new_n40456_;
  assign new_n40458_ = ~new_n40321_ & new_n40334_;
  assign new_n40459_ = new_n40321_ & ~new_n40334_;
  assign new_n40460_ = ~new_n40458_ & ~new_n40459_;
  assign new_n40461_ = ~new_n40457_ & ~new_n40460_;
  assign new_n40462_ = new_n40327_ & ~new_n40447_;
  assign new_n40463_ = ~new_n40327_ & new_n40447_;
  assign new_n40464_ = ~new_n40462_ & ~new_n40463_;
  assign new_n40465_ = ~new_n40308_ & ~new_n40314_;
  assign new_n40466_ = ~new_n40318_ & ~new_n40465_;
  assign new_n40467_ = new_n40311_ & ~new_n40466_;
  assign new_n40468_ = ~new_n40311_ & new_n40466_;
  assign new_n40469_ = ~new_n40467_ & ~new_n40468_;
  assign new_n40470_ = ~new_n40308_ & new_n40314_;
  assign new_n40471_ = new_n40308_ & ~new_n40314_;
  assign new_n40472_ = ~new_n40470_ & ~new_n40471_;
  assign new_n40473_ = new_n40305_ & new_n40306_;
  assign new_n40474_ = ~new_n40305_ & ~new_n40306_;
  assign new_n40475_ = ~new_n40473_ & ~new_n40474_;
  assign new_n40476_ = ~ys__n30334 & ~ys__n33579;
  assign new_n40477_ = ys__n30334 & ys__n33579;
  assign new_n40478_ = ~new_n40476_ & ~new_n40477_;
  assign new_n40479_ = ~ys__n30334 & ~new_n40478_;
  assign new_n40480_ = ~new_n40475_ & new_n40479_;
  assign new_n40481_ = ~new_n40472_ & new_n40480_;
  assign new_n40482_ = ~new_n40469_ & new_n40481_;
  assign new_n40483_ = ~new_n40464_ & new_n40482_;
  assign new_n40484_ = new_n40461_ & new_n40483_;
  assign new_n40485_ = ~new_n40452_ & new_n40484_;
  assign new_n40486_ = ~new_n40445_ & new_n40485_;
  assign new_n40487_ = new_n40442_ & new_n40486_;
  assign new_n40488_ = new_n40433_ & new_n40487_;
  assign new_n40489_ = ~new_n40412_ & new_n40488_;
  assign new_n40490_ = new_n40403_ & new_n40489_;
  assign new_n40491_ = ~new_n40403_ & ~new_n40489_;
  assign new_n40492_ = ~new_n40490_ & ~new_n40491_;
  assign new_n40493_ = ~ys__n17848 & ~new_n39876_;
  assign new_n40494_ = ys__n17848 & new_n39876_;
  assign new_n40495_ = ~new_n40493_ & ~new_n40494_;
  assign new_n40496_ = ys__n17825 & ~new_n39631_;
  assign new_n40497_ = ~ys__n17825 & ~new_n39631_;
  assign new_n40498_ = ys__n17825 & new_n39631_;
  assign new_n40499_ = ~new_n40497_ & ~new_n40498_;
  assign new_n40500_ = ys__n17824 & ~new_n39628_;
  assign new_n40501_ = ~new_n40499_ & new_n40500_;
  assign new_n40502_ = ~new_n40496_ & ~new_n40501_;
  assign new_n40503_ = ~ys__n17828 & ~new_n40033_;
  assign new_n40504_ = ys__n17828 & new_n40033_;
  assign new_n40505_ = ~new_n40503_ & ~new_n40504_;
  assign new_n40506_ = ~ys__n17827 & ~new_n40030_;
  assign new_n40507_ = ys__n17827 & new_n40030_;
  assign new_n40508_ = ~new_n40506_ & ~new_n40507_;
  assign new_n40509_ = ~new_n40505_ & ~new_n40508_;
  assign new_n40510_ = ~new_n40502_ & new_n40509_;
  assign new_n40511_ = ys__n17828 & ~new_n40033_;
  assign new_n40512_ = ys__n17827 & ~new_n40030_;
  assign new_n40513_ = ~new_n40505_ & new_n40512_;
  assign new_n40514_ = ~new_n40511_ & ~new_n40513_;
  assign new_n40515_ = ~new_n40510_ & new_n40514_;
  assign new_n40516_ = ~ys__n17834 & ~new_n40108_;
  assign new_n40517_ = ys__n17834 & new_n40108_;
  assign new_n40518_ = ~new_n40516_ & ~new_n40517_;
  assign new_n40519_ = ~ys__n17833 & ~new_n40124_;
  assign new_n40520_ = ys__n17833 & new_n40124_;
  assign new_n40521_ = ~new_n40519_ & ~new_n40520_;
  assign new_n40522_ = ~new_n40518_ & ~new_n40521_;
  assign new_n40523_ = ~ys__n17831 & ~new_n40066_;
  assign new_n40524_ = ys__n17831 & new_n40066_;
  assign new_n40525_ = ~new_n40523_ & ~new_n40524_;
  assign new_n40526_ = ~ys__n17830 & ~new_n40063_;
  assign new_n40527_ = ys__n17830 & new_n40063_;
  assign new_n40528_ = ~new_n40526_ & ~new_n40527_;
  assign new_n40529_ = ~new_n40525_ & ~new_n40528_;
  assign new_n40530_ = new_n40522_ & new_n40529_;
  assign new_n40531_ = ~new_n40515_ & new_n40530_;
  assign new_n40532_ = ys__n17831 & ~new_n40066_;
  assign new_n40533_ = ys__n17830 & ~new_n40063_;
  assign new_n40534_ = ~new_n40525_ & new_n40533_;
  assign new_n40535_ = ~new_n40532_ & ~new_n40534_;
  assign new_n40536_ = new_n40522_ & ~new_n40535_;
  assign new_n40537_ = ys__n17834 & ~new_n40108_;
  assign new_n40538_ = ys__n17833 & ~new_n40124_;
  assign new_n40539_ = ~new_n40518_ & new_n40538_;
  assign new_n40540_ = ~new_n40537_ & ~new_n40539_;
  assign new_n40541_ = ~new_n40536_ & new_n40540_;
  assign new_n40542_ = ~new_n40531_ & new_n40541_;
  assign new_n40543_ = ~ys__n17846 & ~new_n39889_;
  assign new_n40544_ = ys__n17846 & new_n39889_;
  assign new_n40545_ = ~new_n40543_ & ~new_n40544_;
  assign new_n40546_ = ~ys__n17845 & ~new_n39905_;
  assign new_n40547_ = ys__n17845 & new_n39905_;
  assign new_n40548_ = ~new_n40546_ & ~new_n40547_;
  assign new_n40549_ = ~new_n40545_ & ~new_n40548_;
  assign new_n40550_ = ~ys__n17843 & ~new_n39922_;
  assign new_n40551_ = ys__n17843 & new_n39922_;
  assign new_n40552_ = ~new_n40550_ & ~new_n40551_;
  assign new_n40553_ = ~ys__n17842 & ~new_n39939_;
  assign new_n40554_ = ys__n17842 & new_n39939_;
  assign new_n40555_ = ~new_n40553_ & ~new_n40554_;
  assign new_n40556_ = ~new_n40552_ & ~new_n40555_;
  assign new_n40557_ = new_n40549_ & new_n40556_;
  assign new_n40558_ = ~ys__n17840 & ~new_n39959_;
  assign new_n40559_ = ys__n17840 & new_n39959_;
  assign new_n40560_ = ~new_n40558_ & ~new_n40559_;
  assign new_n40561_ = ~ys__n17839 & ~new_n39975_;
  assign new_n40562_ = ys__n17839 & new_n39975_;
  assign new_n40563_ = ~new_n40561_ & ~new_n40562_;
  assign new_n40564_ = ~new_n40560_ & ~new_n40563_;
  assign new_n40565_ = ~ys__n17837 & ~new_n39992_;
  assign new_n40566_ = ys__n17837 & new_n39992_;
  assign new_n40567_ = ~new_n40565_ & ~new_n40566_;
  assign new_n40568_ = ~ys__n17836 & ~new_n40009_;
  assign new_n40569_ = ys__n17836 & new_n40009_;
  assign new_n40570_ = ~new_n40568_ & ~new_n40569_;
  assign new_n40571_ = ~new_n40567_ & ~new_n40570_;
  assign new_n40572_ = new_n40564_ & new_n40571_;
  assign new_n40573_ = new_n40557_ & new_n40572_;
  assign new_n40574_ = ~new_n40542_ & new_n40573_;
  assign new_n40575_ = ys__n17837 & ~new_n39992_;
  assign new_n40576_ = ys__n17836 & ~new_n40009_;
  assign new_n40577_ = ~new_n40567_ & new_n40576_;
  assign new_n40578_ = ~new_n40575_ & ~new_n40577_;
  assign new_n40579_ = new_n40564_ & ~new_n40578_;
  assign new_n40580_ = ys__n17840 & ~new_n39959_;
  assign new_n40581_ = ys__n17839 & ~new_n39975_;
  assign new_n40582_ = ~new_n40560_ & new_n40581_;
  assign new_n40583_ = ~new_n40580_ & ~new_n40582_;
  assign new_n40584_ = ~new_n40579_ & new_n40583_;
  assign new_n40585_ = new_n40557_ & ~new_n40584_;
  assign new_n40586_ = ys__n17843 & ~new_n39922_;
  assign new_n40587_ = ys__n17842 & ~new_n39939_;
  assign new_n40588_ = ~new_n40552_ & new_n40587_;
  assign new_n40589_ = ~new_n40586_ & ~new_n40588_;
  assign new_n40590_ = new_n40549_ & ~new_n40589_;
  assign new_n40591_ = ys__n17846 & ~new_n39889_;
  assign new_n40592_ = ys__n17845 & ~new_n39905_;
  assign new_n40593_ = ~new_n40545_ & new_n40592_;
  assign new_n40594_ = ~new_n40591_ & ~new_n40593_;
  assign new_n40595_ = ~new_n40590_ & new_n40594_;
  assign new_n40596_ = ~new_n40585_ & new_n40595_;
  assign new_n40597_ = ~new_n40574_ & new_n40596_;
  assign new_n40598_ = new_n40495_ & ~new_n40597_;
  assign new_n40599_ = ~new_n40495_ & new_n40597_;
  assign new_n40600_ = ~new_n40598_ & ~new_n40599_;
  assign new_n40601_ = new_n40492_ & ~new_n40600_;
  assign new_n40602_ = ~new_n40542_ & new_n40572_;
  assign new_n40603_ = new_n40584_ & ~new_n40602_;
  assign new_n40604_ = new_n40556_ & ~new_n40603_;
  assign new_n40605_ = new_n40589_ & ~new_n40604_;
  assign new_n40606_ = ~new_n40548_ & ~new_n40605_;
  assign new_n40607_ = ~new_n40592_ & ~new_n40606_;
  assign new_n40608_ = new_n40545_ & ~new_n40607_;
  assign new_n40609_ = ~new_n40545_ & new_n40607_;
  assign new_n40610_ = ~new_n40608_ & ~new_n40609_;
  assign new_n40611_ = ~new_n40542_ & new_n40571_;
  assign new_n40612_ = new_n40578_ & ~new_n40611_;
  assign new_n40613_ = ~new_n40563_ & ~new_n40612_;
  assign new_n40614_ = ~new_n40581_ & ~new_n40613_;
  assign new_n40615_ = new_n40560_ & ~new_n40614_;
  assign new_n40616_ = ~new_n40560_ & new_n40614_;
  assign new_n40617_ = ~new_n40615_ & ~new_n40616_;
  assign new_n40618_ = new_n40563_ & ~new_n40612_;
  assign new_n40619_ = ~new_n40563_ & new_n40612_;
  assign new_n40620_ = ~new_n40618_ & ~new_n40619_;
  assign new_n40621_ = ~new_n40542_ & ~new_n40570_;
  assign new_n40622_ = ~new_n40576_ & ~new_n40621_;
  assign new_n40623_ = new_n40567_ & ~new_n40622_;
  assign new_n40624_ = ~new_n40567_ & new_n40622_;
  assign new_n40625_ = ~new_n40623_ & ~new_n40624_;
  assign new_n40626_ = ~new_n40542_ & new_n40570_;
  assign new_n40627_ = new_n40542_ & ~new_n40570_;
  assign new_n40628_ = ~new_n40626_ & ~new_n40627_;
  assign new_n40629_ = ~new_n40625_ & ~new_n40628_;
  assign new_n40630_ = ~new_n40620_ & new_n40629_;
  assign new_n40631_ = ~new_n40617_ & new_n40630_;
  assign new_n40632_ = ~new_n40555_ & ~new_n40603_;
  assign new_n40633_ = ~new_n40587_ & ~new_n40632_;
  assign new_n40634_ = new_n40552_ & ~new_n40633_;
  assign new_n40635_ = ~new_n40552_ & new_n40633_;
  assign new_n40636_ = ~new_n40634_ & ~new_n40635_;
  assign new_n40637_ = new_n40555_ & ~new_n40603_;
  assign new_n40638_ = ~new_n40555_ & new_n40603_;
  assign new_n40639_ = ~new_n40637_ & ~new_n40638_;
  assign new_n40640_ = ~new_n40636_ & ~new_n40639_;
  assign new_n40641_ = new_n40548_ & ~new_n40605_;
  assign new_n40642_ = ~new_n40548_ & new_n40605_;
  assign new_n40643_ = ~new_n40641_ & ~new_n40642_;
  assign new_n40644_ = ~new_n40515_ & new_n40529_;
  assign new_n40645_ = new_n40535_ & ~new_n40644_;
  assign new_n40646_ = ~new_n40521_ & ~new_n40645_;
  assign new_n40647_ = ~new_n40538_ & ~new_n40646_;
  assign new_n40648_ = new_n40518_ & ~new_n40647_;
  assign new_n40649_ = ~new_n40518_ & new_n40647_;
  assign new_n40650_ = ~new_n40648_ & ~new_n40649_;
  assign new_n40651_ = ~new_n40515_ & ~new_n40528_;
  assign new_n40652_ = ~new_n40533_ & ~new_n40651_;
  assign new_n40653_ = new_n40525_ & ~new_n40652_;
  assign new_n40654_ = ~new_n40525_ & new_n40652_;
  assign new_n40655_ = ~new_n40653_ & ~new_n40654_;
  assign new_n40656_ = ~new_n40515_ & new_n40528_;
  assign new_n40657_ = new_n40515_ & ~new_n40528_;
  assign new_n40658_ = ~new_n40656_ & ~new_n40657_;
  assign new_n40659_ = ~new_n40655_ & ~new_n40658_;
  assign new_n40660_ = new_n40521_ & ~new_n40645_;
  assign new_n40661_ = ~new_n40521_ & new_n40645_;
  assign new_n40662_ = ~new_n40660_ & ~new_n40661_;
  assign new_n40663_ = ~new_n40502_ & ~new_n40508_;
  assign new_n40664_ = ~new_n40512_ & ~new_n40663_;
  assign new_n40665_ = new_n40505_ & ~new_n40664_;
  assign new_n40666_ = ~new_n40505_ & new_n40664_;
  assign new_n40667_ = ~new_n40665_ & ~new_n40666_;
  assign new_n40668_ = ~new_n40502_ & new_n40508_;
  assign new_n40669_ = new_n40502_ & ~new_n40508_;
  assign new_n40670_ = ~new_n40668_ & ~new_n40669_;
  assign new_n40671_ = new_n40499_ & new_n40500_;
  assign new_n40672_ = ~new_n40499_ & ~new_n40500_;
  assign new_n40673_ = ~new_n40671_ & ~new_n40672_;
  assign new_n40674_ = ~ys__n17824 & ~new_n39628_;
  assign new_n40675_ = ys__n17824 & new_n39628_;
  assign new_n40676_ = ~new_n40674_ & ~new_n40675_;
  assign new_n40677_ = ~new_n40673_ & ~new_n40676_;
  assign new_n40678_ = ~new_n40670_ & new_n40677_;
  assign new_n40679_ = ~new_n40667_ & new_n40678_;
  assign new_n40680_ = ~new_n40662_ & new_n40679_;
  assign new_n40681_ = new_n40659_ & new_n40680_;
  assign new_n40682_ = ~new_n40650_ & new_n40681_;
  assign new_n40683_ = ~new_n40643_ & new_n40682_;
  assign new_n40684_ = new_n40640_ & new_n40683_;
  assign new_n40685_ = new_n40631_ & new_n40684_;
  assign new_n40686_ = ~new_n40610_ & new_n40685_;
  assign new_n40687_ = new_n40600_ & new_n40686_;
  assign new_n40688_ = ~new_n40600_ & ~new_n40686_;
  assign new_n40689_ = ~new_n40687_ & ~new_n40688_;
  assign new_n40690_ = ~new_n40492_ & ~new_n40689_;
  assign new_n40691_ = ~new_n40601_ & ~new_n40690_;
  assign new_n40692_ = ys__n18156 & ~new_n40691_;
  assign new_n40693_ = ys__n17848 & ~new_n39876_;
  assign new_n40694_ = ~new_n40495_ & ~new_n40597_;
  assign new_n40695_ = ~new_n40693_ & ~new_n40694_;
  assign new_n40696_ = new_n40265_ & ~new_n40695_;
  assign new_n40697_ = ~new_n40265_ & new_n40695_;
  assign new_n40698_ = ~new_n40696_ & ~new_n40697_;
  assign new_n40699_ = new_n40492_ & ~new_n40698_;
  assign new_n40700_ = ~new_n40600_ & new_n40686_;
  assign new_n40701_ = new_n40698_ & new_n40700_;
  assign new_n40702_ = ~new_n40698_ & ~new_n40700_;
  assign new_n40703_ = ~new_n40701_ & ~new_n40702_;
  assign new_n40704_ = ~new_n40492_ & ~new_n40703_;
  assign new_n40705_ = ~new_n40699_ & ~new_n40704_;
  assign new_n40706_ = ~new_n40692_ & new_n40705_;
  assign new_n40707_ = ~new_n40301_ & ~new_n40706_;
  assign new_n40708_ = ys__n33581 & ~new_n39473_;
  assign new_n40709_ = ys__n33579 & ~new_n39486_;
  assign new_n40710_ = ~new_n39496_ & new_n40709_;
  assign new_n40711_ = ~new_n40708_ & ~new_n40710_;
  assign new_n40712_ = ~new_n39479_ & ~new_n39529_;
  assign new_n40713_ = ~new_n40711_ & new_n40712_;
  assign new_n40714_ = ys__n17804 & ~new_n39510_;
  assign new_n40715_ = ys__n17803 & ~new_n39476_;
  assign new_n40716_ = ~new_n39529_ & new_n40715_;
  assign new_n40717_ = ~new_n40714_ & ~new_n40716_;
  assign new_n40718_ = ~new_n40713_ & new_n40717_;
  assign new_n40719_ = ~new_n39571_ & ~new_n39588_;
  assign new_n40720_ = ~new_n39516_ & ~new_n39601_;
  assign new_n40721_ = new_n40719_ & new_n40720_;
  assign new_n40722_ = ~new_n40718_ & new_n40721_;
  assign new_n40723_ = ys__n17807 & ~new_n39578_;
  assign new_n40724_ = ys__n17806 & ~new_n39513_;
  assign new_n40725_ = ~new_n39601_ & new_n40724_;
  assign new_n40726_ = ~new_n40723_ & ~new_n40725_;
  assign new_n40727_ = new_n40719_ & ~new_n40726_;
  assign new_n40728_ = ys__n17810 & ~new_n39549_;
  assign new_n40729_ = ys__n17809 & ~new_n39562_;
  assign new_n40730_ = ~new_n39571_ & new_n40729_;
  assign new_n40731_ = ~new_n40728_ & ~new_n40730_;
  assign new_n40732_ = ~new_n40727_ & new_n40731_;
  assign new_n40733_ = ~new_n40722_ & new_n40732_;
  assign new_n40734_ = ~new_n39650_ & ~new_n39667_;
  assign new_n40735_ = ~new_n39683_ & ~new_n39701_;
  assign new_n40736_ = new_n40734_ & new_n40735_;
  assign new_n40737_ = ~new_n39717_ & ~new_n39734_;
  assign new_n40738_ = ~new_n39555_ & ~new_n39747_;
  assign new_n40739_ = new_n40737_ & new_n40738_;
  assign new_n40740_ = new_n40736_ & new_n40739_;
  assign new_n40741_ = ~new_n40733_ & new_n40740_;
  assign new_n40742_ = ys__n17813 & ~new_n39724_;
  assign new_n40743_ = ys__n17812 & ~new_n39552_;
  assign new_n40744_ = ~new_n39747_ & new_n40743_;
  assign new_n40745_ = ~new_n40742_ & ~new_n40744_;
  assign new_n40746_ = new_n40737_ & ~new_n40745_;
  assign new_n40747_ = ys__n17816 & ~new_n39690_;
  assign new_n40748_ = ys__n17815 & ~new_n39708_;
  assign new_n40749_ = ~new_n39717_ & new_n40748_;
  assign new_n40750_ = ~new_n40747_ & ~new_n40749_;
  assign new_n40751_ = ~new_n40746_ & new_n40750_;
  assign new_n40752_ = new_n40736_ & ~new_n40751_;
  assign new_n40753_ = ys__n17819 & ~new_n39657_;
  assign new_n40754_ = ys__n17818 & ~new_n39674_;
  assign new_n40755_ = ~new_n39683_ & new_n40754_;
  assign new_n40756_ = ~new_n40753_ & ~new_n40755_;
  assign new_n40757_ = new_n40734_ & ~new_n40756_;
  assign new_n40758_ = ys__n17822 & ~new_n39628_;
  assign new_n40759_ = ys__n17821 & ~new_n39641_;
  assign new_n40760_ = ~new_n39650_ & new_n40759_;
  assign new_n40761_ = ~new_n40758_ & ~new_n40760_;
  assign new_n40762_ = ~new_n40757_ & new_n40761_;
  assign new_n40763_ = ~new_n40752_ & new_n40762_;
  assign new_n40764_ = ~new_n40741_ & new_n40763_;
  assign new_n40765_ = ~new_n40733_ & new_n40739_;
  assign new_n40766_ = new_n40751_ & ~new_n40765_;
  assign new_n40767_ = new_n40735_ & ~new_n40766_;
  assign new_n40768_ = new_n40756_ & ~new_n40767_;
  assign new_n40769_ = ~new_n39667_ & ~new_n40768_;
  assign new_n40770_ = ~new_n40759_ & ~new_n40769_;
  assign new_n40771_ = new_n39650_ & ~new_n40770_;
  assign new_n40772_ = ~new_n39650_ & new_n40770_;
  assign new_n40773_ = ~new_n40771_ & ~new_n40772_;
  assign new_n40774_ = ~new_n40733_ & new_n40738_;
  assign new_n40775_ = new_n40745_ & ~new_n40774_;
  assign new_n40776_ = ~new_n39734_ & ~new_n40775_;
  assign new_n40777_ = ~new_n40748_ & ~new_n40776_;
  assign new_n40778_ = new_n39717_ & ~new_n40777_;
  assign new_n40779_ = ~new_n39717_ & new_n40777_;
  assign new_n40780_ = ~new_n40778_ & ~new_n40779_;
  assign new_n40781_ = new_n39734_ & ~new_n40775_;
  assign new_n40782_ = ~new_n39734_ & new_n40775_;
  assign new_n40783_ = ~new_n40781_ & ~new_n40782_;
  assign new_n40784_ = ~new_n39555_ & ~new_n40733_;
  assign new_n40785_ = ~new_n40743_ & ~new_n40784_;
  assign new_n40786_ = new_n39747_ & ~new_n40785_;
  assign new_n40787_ = ~new_n39747_ & new_n40785_;
  assign new_n40788_ = ~new_n40786_ & ~new_n40787_;
  assign new_n40789_ = new_n39555_ & ~new_n40733_;
  assign new_n40790_ = ~new_n39555_ & new_n40733_;
  assign new_n40791_ = ~new_n40789_ & ~new_n40790_;
  assign new_n40792_ = ~new_n40788_ & ~new_n40791_;
  assign new_n40793_ = ~new_n40783_ & new_n40792_;
  assign new_n40794_ = ~new_n40780_ & new_n40793_;
  assign new_n40795_ = ~new_n39701_ & ~new_n40766_;
  assign new_n40796_ = ~new_n40754_ & ~new_n40795_;
  assign new_n40797_ = new_n39683_ & ~new_n40796_;
  assign new_n40798_ = ~new_n39683_ & new_n40796_;
  assign new_n40799_ = ~new_n40797_ & ~new_n40798_;
  assign new_n40800_ = new_n39701_ & ~new_n40766_;
  assign new_n40801_ = ~new_n39701_ & new_n40766_;
  assign new_n40802_ = ~new_n40800_ & ~new_n40801_;
  assign new_n40803_ = ~new_n40799_ & ~new_n40802_;
  assign new_n40804_ = new_n39667_ & ~new_n40768_;
  assign new_n40805_ = ~new_n39667_ & new_n40768_;
  assign new_n40806_ = ~new_n40804_ & ~new_n40805_;
  assign new_n40807_ = ~new_n40718_ & new_n40720_;
  assign new_n40808_ = new_n40726_ & ~new_n40807_;
  assign new_n40809_ = ~new_n39588_ & ~new_n40808_;
  assign new_n40810_ = ~new_n40729_ & ~new_n40809_;
  assign new_n40811_ = new_n39571_ & ~new_n40810_;
  assign new_n40812_ = ~new_n39571_ & new_n40810_;
  assign new_n40813_ = ~new_n40811_ & ~new_n40812_;
  assign new_n40814_ = ~new_n39516_ & ~new_n40718_;
  assign new_n40815_ = ~new_n40724_ & ~new_n40814_;
  assign new_n40816_ = new_n39601_ & ~new_n40815_;
  assign new_n40817_ = ~new_n39601_ & new_n40815_;
  assign new_n40818_ = ~new_n40816_ & ~new_n40817_;
  assign new_n40819_ = new_n39516_ & ~new_n40718_;
  assign new_n40820_ = ~new_n39516_ & new_n40718_;
  assign new_n40821_ = ~new_n40819_ & ~new_n40820_;
  assign new_n40822_ = ~new_n40818_ & ~new_n40821_;
  assign new_n40823_ = new_n39588_ & ~new_n40808_;
  assign new_n40824_ = ~new_n39588_ & new_n40808_;
  assign new_n40825_ = ~new_n40823_ & ~new_n40824_;
  assign new_n40826_ = ~new_n39479_ & ~new_n40711_;
  assign new_n40827_ = ~new_n40715_ & ~new_n40826_;
  assign new_n40828_ = new_n39529_ & ~new_n40827_;
  assign new_n40829_ = ~new_n39529_ & new_n40827_;
  assign new_n40830_ = ~new_n40828_ & ~new_n40829_;
  assign new_n40831_ = new_n39479_ & ~new_n40711_;
  assign new_n40832_ = ~new_n39479_ & new_n40711_;
  assign new_n40833_ = ~new_n40831_ & ~new_n40832_;
  assign new_n40834_ = new_n39496_ & new_n40709_;
  assign new_n40835_ = ~new_n39496_ & ~new_n40709_;
  assign new_n40836_ = ~new_n40834_ & ~new_n40835_;
  assign new_n40837_ = ys__n33579 & new_n39486_;
  assign new_n40838_ = ~new_n39500_ & ~new_n40837_;
  assign new_n40839_ = ~ys__n402 & ~ys__n30334;
  assign new_n40840_ = ~ys__n402 & ~new_n40839_;
  assign new_n40841_ = ~new_n40838_ & ~new_n40840_;
  assign new_n40842_ = ~new_n40836_ & new_n40841_;
  assign new_n40843_ = ~new_n40833_ & new_n40842_;
  assign new_n40844_ = ~new_n40830_ & new_n40843_;
  assign new_n40845_ = ~new_n40825_ & new_n40844_;
  assign new_n40846_ = new_n40822_ & new_n40845_;
  assign new_n40847_ = ~new_n40813_ & new_n40846_;
  assign new_n40848_ = ~new_n40806_ & new_n40847_;
  assign new_n40849_ = new_n40803_ & new_n40848_;
  assign new_n40850_ = new_n40794_ & new_n40849_;
  assign new_n40851_ = ~new_n40773_ & new_n40850_;
  assign new_n40852_ = new_n40764_ & new_n40851_;
  assign new_n40853_ = ~new_n40764_ & ~new_n40851_;
  assign new_n40854_ = ~new_n40852_ & ~new_n40853_;
  assign new_n40855_ = ys__n17825 & ~new_n40030_;
  assign new_n40856_ = ys__n17824 & ~new_n39631_;
  assign new_n40857_ = ~new_n40050_ & new_n40856_;
  assign new_n40858_ = ~new_n40855_ & ~new_n40857_;
  assign new_n40859_ = ~new_n40036_ & ~new_n40082_;
  assign new_n40860_ = ~new_n40858_ & new_n40859_;
  assign new_n40861_ = ys__n17828 & ~new_n40063_;
  assign new_n40862_ = ys__n17827 & ~new_n40033_;
  assign new_n40863_ = ~new_n40082_ & new_n40862_;
  assign new_n40864_ = ~new_n40861_ & ~new_n40863_;
  assign new_n40865_ = ~new_n40860_ & new_n40864_;
  assign new_n40866_ = ~new_n40117_ & ~new_n40134_;
  assign new_n40867_ = ~new_n40069_ & ~new_n40147_;
  assign new_n40868_ = new_n40866_ & new_n40867_;
  assign new_n40869_ = ~new_n40865_ & new_n40868_;
  assign new_n40870_ = ys__n17831 & ~new_n40124_;
  assign new_n40871_ = ys__n17830 & ~new_n40066_;
  assign new_n40872_ = ~new_n40147_ & new_n40871_;
  assign new_n40873_ = ~new_n40870_ & ~new_n40872_;
  assign new_n40874_ = new_n40866_ & ~new_n40873_;
  assign new_n40875_ = ys__n17834 & ~new_n40009_;
  assign new_n40876_ = ys__n17833 & ~new_n40108_;
  assign new_n40877_ = ~new_n40117_ & new_n40876_;
  assign new_n40878_ = ~new_n40875_ & ~new_n40877_;
  assign new_n40879_ = ~new_n40874_ & new_n40878_;
  assign new_n40880_ = ~new_n40869_ & new_n40879_;
  assign new_n40881_ = ~new_n39898_ & ~new_n39915_;
  assign new_n40882_ = ~new_n39932_ & ~new_n39952_;
  assign new_n40883_ = new_n40881_ & new_n40882_;
  assign new_n40884_ = ~new_n39968_ & ~new_n39985_;
  assign new_n40885_ = ~new_n40002_ & ~new_n40101_;
  assign new_n40886_ = new_n40884_ & new_n40885_;
  assign new_n40887_ = new_n40883_ & new_n40886_;
  assign new_n40888_ = ~new_n40880_ & new_n40887_;
  assign new_n40889_ = ys__n17837 & ~new_n39975_;
  assign new_n40890_ = ys__n17836 & ~new_n39992_;
  assign new_n40891_ = ~new_n40002_ & new_n40890_;
  assign new_n40892_ = ~new_n40889_ & ~new_n40891_;
  assign new_n40893_ = new_n40884_ & ~new_n40892_;
  assign new_n40894_ = ys__n17840 & ~new_n39939_;
  assign new_n40895_ = ys__n17839 & ~new_n39959_;
  assign new_n40896_ = ~new_n39968_ & new_n40895_;
  assign new_n40897_ = ~new_n40894_ & ~new_n40896_;
  assign new_n40898_ = ~new_n40893_ & new_n40897_;
  assign new_n40899_ = new_n40883_ & ~new_n40898_;
  assign new_n40900_ = ys__n17843 & ~new_n39905_;
  assign new_n40901_ = ys__n17842 & ~new_n39922_;
  assign new_n40902_ = ~new_n39932_ & new_n40901_;
  assign new_n40903_ = ~new_n40900_ & ~new_n40902_;
  assign new_n40904_ = new_n40881_ & ~new_n40903_;
  assign new_n40905_ = ys__n17846 & ~new_n39876_;
  assign new_n40906_ = ys__n17845 & ~new_n39889_;
  assign new_n40907_ = ~new_n39898_ & new_n40906_;
  assign new_n40908_ = ~new_n40905_ & ~new_n40907_;
  assign new_n40909_ = ~new_n40904_ & new_n40908_;
  assign new_n40910_ = ~new_n40899_ & new_n40909_;
  assign new_n40911_ = ~new_n40888_ & new_n40910_;
  assign new_n40912_ = new_n39882_ & ~new_n40911_;
  assign new_n40913_ = ~new_n39882_ & new_n40911_;
  assign new_n40914_ = ~new_n40912_ & ~new_n40913_;
  assign new_n40915_ = new_n40854_ & ~new_n40914_;
  assign new_n40916_ = ~new_n40880_ & new_n40886_;
  assign new_n40917_ = new_n40898_ & ~new_n40916_;
  assign new_n40918_ = new_n40882_ & ~new_n40917_;
  assign new_n40919_ = new_n40903_ & ~new_n40918_;
  assign new_n40920_ = ~new_n39915_ & ~new_n40919_;
  assign new_n40921_ = ~new_n40906_ & ~new_n40920_;
  assign new_n40922_ = new_n39898_ & ~new_n40921_;
  assign new_n40923_ = ~new_n39898_ & new_n40921_;
  assign new_n40924_ = ~new_n40922_ & ~new_n40923_;
  assign new_n40925_ = ~new_n40880_ & new_n40885_;
  assign new_n40926_ = new_n40892_ & ~new_n40925_;
  assign new_n40927_ = ~new_n39985_ & ~new_n40926_;
  assign new_n40928_ = ~new_n40895_ & ~new_n40927_;
  assign new_n40929_ = new_n39968_ & ~new_n40928_;
  assign new_n40930_ = ~new_n39968_ & new_n40928_;
  assign new_n40931_ = ~new_n40929_ & ~new_n40930_;
  assign new_n40932_ = new_n39985_ & ~new_n40926_;
  assign new_n40933_ = ~new_n39985_ & new_n40926_;
  assign new_n40934_ = ~new_n40932_ & ~new_n40933_;
  assign new_n40935_ = ~new_n40101_ & ~new_n40880_;
  assign new_n40936_ = ~new_n40890_ & ~new_n40935_;
  assign new_n40937_ = new_n40002_ & ~new_n40936_;
  assign new_n40938_ = ~new_n40002_ & new_n40936_;
  assign new_n40939_ = ~new_n40937_ & ~new_n40938_;
  assign new_n40940_ = new_n40101_ & ~new_n40880_;
  assign new_n40941_ = ~new_n40101_ & new_n40880_;
  assign new_n40942_ = ~new_n40940_ & ~new_n40941_;
  assign new_n40943_ = ~new_n40939_ & ~new_n40942_;
  assign new_n40944_ = ~new_n40934_ & new_n40943_;
  assign new_n40945_ = ~new_n40931_ & new_n40944_;
  assign new_n40946_ = ~new_n39952_ & ~new_n40917_;
  assign new_n40947_ = ~new_n40901_ & ~new_n40946_;
  assign new_n40948_ = new_n39932_ & ~new_n40947_;
  assign new_n40949_ = ~new_n39932_ & new_n40947_;
  assign new_n40950_ = ~new_n40948_ & ~new_n40949_;
  assign new_n40951_ = new_n39952_ & ~new_n40917_;
  assign new_n40952_ = ~new_n39952_ & new_n40917_;
  assign new_n40953_ = ~new_n40951_ & ~new_n40952_;
  assign new_n40954_ = ~new_n40950_ & ~new_n40953_;
  assign new_n40955_ = new_n39915_ & ~new_n40919_;
  assign new_n40956_ = ~new_n39915_ & new_n40919_;
  assign new_n40957_ = ~new_n40955_ & ~new_n40956_;
  assign new_n40958_ = ~new_n40865_ & new_n40867_;
  assign new_n40959_ = new_n40873_ & ~new_n40958_;
  assign new_n40960_ = ~new_n40134_ & ~new_n40959_;
  assign new_n40961_ = ~new_n40876_ & ~new_n40960_;
  assign new_n40962_ = new_n40117_ & ~new_n40961_;
  assign new_n40963_ = ~new_n40117_ & new_n40961_;
  assign new_n40964_ = ~new_n40962_ & ~new_n40963_;
  assign new_n40965_ = ~new_n40069_ & ~new_n40865_;
  assign new_n40966_ = ~new_n40871_ & ~new_n40965_;
  assign new_n40967_ = new_n40147_ & ~new_n40966_;
  assign new_n40968_ = ~new_n40147_ & new_n40966_;
  assign new_n40969_ = ~new_n40967_ & ~new_n40968_;
  assign new_n40970_ = new_n40069_ & ~new_n40865_;
  assign new_n40971_ = ~new_n40069_ & new_n40865_;
  assign new_n40972_ = ~new_n40970_ & ~new_n40971_;
  assign new_n40973_ = ~new_n40969_ & ~new_n40972_;
  assign new_n40974_ = new_n40134_ & ~new_n40959_;
  assign new_n40975_ = ~new_n40134_ & new_n40959_;
  assign new_n40976_ = ~new_n40974_ & ~new_n40975_;
  assign new_n40977_ = ~new_n40036_ & ~new_n40858_;
  assign new_n40978_ = ~new_n40862_ & ~new_n40977_;
  assign new_n40979_ = new_n40082_ & ~new_n40978_;
  assign new_n40980_ = ~new_n40082_ & new_n40978_;
  assign new_n40981_ = ~new_n40979_ & ~new_n40980_;
  assign new_n40982_ = new_n40036_ & ~new_n40858_;
  assign new_n40983_ = ~new_n40036_ & new_n40858_;
  assign new_n40984_ = ~new_n40982_ & ~new_n40983_;
  assign new_n40985_ = new_n40050_ & new_n40856_;
  assign new_n40986_ = ~new_n40050_ & ~new_n40856_;
  assign new_n40987_ = ~new_n40985_ & ~new_n40986_;
  assign new_n40988_ = ~new_n39634_ & ~new_n40987_;
  assign new_n40989_ = ~new_n40984_ & new_n40988_;
  assign new_n40990_ = ~new_n40981_ & new_n40989_;
  assign new_n40991_ = ~new_n40976_ & new_n40990_;
  assign new_n40992_ = new_n40973_ & new_n40991_;
  assign new_n40993_ = ~new_n40964_ & new_n40992_;
  assign new_n40994_ = ~new_n40957_ & new_n40993_;
  assign new_n40995_ = new_n40954_ & new_n40994_;
  assign new_n40996_ = new_n40945_ & new_n40995_;
  assign new_n40997_ = ~new_n40924_ & new_n40996_;
  assign new_n40998_ = new_n40914_ & new_n40997_;
  assign new_n40999_ = ~new_n40914_ & ~new_n40997_;
  assign new_n41000_ = ~new_n40998_ & ~new_n40999_;
  assign new_n41001_ = ~new_n40854_ & ~new_n41000_;
  assign new_n41002_ = ~new_n40915_ & ~new_n41001_;
  assign new_n41003_ = ys__n18156 & ~new_n41002_;
  assign new_n41004_ = ys__n17848 & ~new_n39879_;
  assign new_n41005_ = ~new_n39882_ & ~new_n40911_;
  assign new_n41006_ = ~new_n41004_ & ~new_n41005_;
  assign new_n41007_ = new_n40265_ & ~new_n41006_;
  assign new_n41008_ = ~new_n40265_ & new_n41006_;
  assign new_n41009_ = ~new_n41007_ & ~new_n41008_;
  assign new_n41010_ = new_n40854_ & ~new_n41009_;
  assign new_n41011_ = ~new_n40914_ & new_n40997_;
  assign new_n41012_ = new_n41009_ & new_n41011_;
  assign new_n41013_ = ~new_n41009_ & ~new_n41011_;
  assign new_n41014_ = ~new_n41012_ & ~new_n41013_;
  assign new_n41015_ = ~new_n40854_ & ~new_n41014_;
  assign new_n41016_ = ~new_n41010_ & ~new_n41015_;
  assign new_n41017_ = ~new_n41003_ & new_n41016_;
  assign new_n41018_ = ys__n408 & ~new_n41017_;
  assign new_n41019_ = new_n40707_ & new_n41018_;
  assign new_n41020_ = ys__n33579 & new_n41019_;
  assign new_n41021_ = ~ys__n30334 & new_n40838_;
  assign new_n41022_ = ys__n30334 & ~new_n40838_;
  assign new_n41023_ = ~new_n41021_ & ~new_n41022_;
  assign new_n41024_ = ys__n408 & new_n40301_;
  assign new_n41025_ = ~new_n41023_ & new_n41024_;
  assign new_n41026_ = ys__n402 & ys__n404;
  assign new_n41027_ = ys__n402 & ~new_n41026_;
  assign new_n41028_ = ~ys__n408 & ys__n17803;
  assign new_n41029_ = new_n41026_ & new_n41028_;
  assign new_n41030_ = ~new_n41027_ & new_n41029_;
  assign new_n41031_ = ~new_n41025_ & ~new_n41030_;
  assign new_n41032_ = ~new_n41020_ & new_n41031_;
  assign new_n41033_ = new_n40838_ & ~new_n40840_;
  assign new_n41034_ = ~new_n40838_ & new_n40840_;
  assign new_n41035_ = ~new_n41033_ & ~new_n41034_;
  assign new_n41036_ = ys__n408 & new_n41017_;
  assign new_n41037_ = new_n40707_ & new_n41036_;
  assign new_n41038_ = ~new_n41035_ & new_n41037_;
  assign new_n41039_ = ~ys__n30334 & new_n40478_;
  assign new_n41040_ = ys__n30334 & ~new_n40478_;
  assign new_n41041_ = ~new_n41039_ & ~new_n41040_;
  assign new_n41042_ = ~new_n40301_ & new_n40706_;
  assign new_n41043_ = ys__n408 & new_n41042_;
  assign new_n41044_ = ~new_n41041_ & new_n41043_;
  assign new_n41045_ = ~new_n41038_ & ~new_n41044_;
  assign new_n41046_ = new_n41032_ & new_n41045_;
  assign new_n41047_ = ys__n408 & ~new_n41024_;
  assign new_n41048_ = ~new_n41019_ & new_n41047_;
  assign new_n41049_ = ~new_n41037_ & ~new_n41043_;
  assign new_n41050_ = new_n41048_ & new_n41049_;
  assign new_n41051_ = ~new_n15136_ & ~new_n41050_;
  assign new_n41052_ = ~new_n41046_ & new_n41051_;
  assign ys__n30235 = new_n39470_ | new_n41052_;
  assign new_n41054_ = ys__n352 & ys__n23272;
  assign new_n41055_ = new_n15136_ & new_n41054_;
  assign new_n41056_ = ys__n33581 & new_n41019_;
  assign new_n41057_ = ~ys__n30334 & new_n39859_;
  assign new_n41058_ = ys__n30334 & ~new_n39859_;
  assign new_n41059_ = ~new_n41057_ & ~new_n41058_;
  assign new_n41060_ = new_n41024_ & ~new_n41059_;
  assign new_n41061_ = ~ys__n17803 & ys__n17804;
  assign new_n41062_ = ys__n17803 & ~ys__n17804;
  assign new_n41063_ = ~new_n41061_ & ~new_n41062_;
  assign new_n41064_ = ~ys__n408 & new_n41026_;
  assign new_n41065_ = ~new_n41063_ & new_n41064_;
  assign new_n41066_ = ~new_n41027_ & new_n41065_;
  assign new_n41067_ = ~new_n41060_ & ~new_n41066_;
  assign new_n41068_ = ~new_n41056_ & new_n41067_;
  assign new_n41069_ = new_n40836_ & new_n40841_;
  assign new_n41070_ = ~new_n40836_ & ~new_n40841_;
  assign new_n41071_ = ~new_n41069_ & ~new_n41070_;
  assign new_n41072_ = new_n41037_ & ~new_n41071_;
  assign new_n41073_ = new_n40475_ & new_n40479_;
  assign new_n41074_ = ~new_n40475_ & ~new_n40479_;
  assign new_n41075_ = ~new_n41073_ & ~new_n41074_;
  assign new_n41076_ = new_n41043_ & ~new_n41075_;
  assign new_n41077_ = ~new_n41072_ & ~new_n41076_;
  assign new_n41078_ = new_n41068_ & new_n41077_;
  assign new_n41079_ = new_n41051_ & ~new_n41078_;
  assign ys__n30238 = new_n41055_ | new_n41079_;
  assign new_n41081_ = ys__n352 & ys__n23274;
  assign new_n41082_ = new_n15136_ & new_n41081_;
  assign new_n41083_ = ys__n17803 & new_n41019_;
  assign new_n41084_ = new_n39856_ & new_n39860_;
  assign new_n41085_ = ~new_n39856_ & ~new_n39860_;
  assign new_n41086_ = ~new_n41084_ & ~new_n41085_;
  assign new_n41087_ = new_n41024_ & ~new_n41086_;
  assign new_n41088_ = ys__n17806 & new_n17806_;
  assign new_n41089_ = ~ys__n17806 & ~new_n17806_;
  assign new_n41090_ = ~new_n41088_ & ~new_n41089_;
  assign new_n41091_ = ~new_n41027_ & new_n41064_;
  assign new_n41092_ = ~new_n41090_ & new_n41091_;
  assign new_n41093_ = ~new_n41087_ & ~new_n41092_;
  assign new_n41094_ = ~new_n41083_ & new_n41093_;
  assign new_n41095_ = new_n40833_ & new_n40842_;
  assign new_n41096_ = ~new_n40833_ & ~new_n40842_;
  assign new_n41097_ = ~new_n41095_ & ~new_n41096_;
  assign new_n41098_ = new_n41037_ & ~new_n41097_;
  assign new_n41099_ = new_n40472_ & new_n40480_;
  assign new_n41100_ = ~new_n40472_ & ~new_n40480_;
  assign new_n41101_ = ~new_n41099_ & ~new_n41100_;
  assign new_n41102_ = new_n41043_ & ~new_n41101_;
  assign new_n41103_ = ~new_n41098_ & ~new_n41102_;
  assign new_n41104_ = new_n41094_ & new_n41103_;
  assign new_n41105_ = new_n41051_ & ~new_n41104_;
  assign ys__n30241 = new_n41082_ | new_n41105_;
  assign new_n41107_ = ys__n352 & ys__n23276;
  assign new_n41108_ = new_n15136_ & new_n41107_;
  assign new_n41109_ = ys__n17804 & new_n41019_;
  assign new_n41110_ = new_n39853_ & new_n39861_;
  assign new_n41111_ = ~new_n39853_ & ~new_n39861_;
  assign new_n41112_ = ~new_n41110_ & ~new_n41111_;
  assign new_n41113_ = new_n41024_ & ~new_n41112_;
  assign new_n41114_ = ~ys__n17806 & new_n17806_;
  assign new_n41115_ = ys__n17807 & new_n41114_;
  assign new_n41116_ = ~ys__n17807 & ~new_n41114_;
  assign new_n41117_ = ~new_n41115_ & ~new_n41116_;
  assign new_n41118_ = new_n41091_ & ~new_n41117_;
  assign new_n41119_ = ~new_n41113_ & ~new_n41118_;
  assign new_n41120_ = ~new_n41109_ & new_n41119_;
  assign new_n41121_ = new_n40830_ & new_n40843_;
  assign new_n41122_ = ~new_n40830_ & ~new_n40843_;
  assign new_n41123_ = ~new_n41121_ & ~new_n41122_;
  assign new_n41124_ = new_n41037_ & ~new_n41123_;
  assign new_n41125_ = new_n40469_ & new_n40481_;
  assign new_n41126_ = ~new_n40469_ & ~new_n40481_;
  assign new_n41127_ = ~new_n41125_ & ~new_n41126_;
  assign new_n41128_ = new_n41043_ & ~new_n41127_;
  assign new_n41129_ = ~new_n41124_ & ~new_n41128_;
  assign new_n41130_ = new_n41120_ & new_n41129_;
  assign new_n41131_ = new_n41051_ & ~new_n41130_;
  assign ys__n30244 = new_n41108_ | new_n41131_;
  assign new_n41133_ = ys__n352 & ys__n23278;
  assign new_n41134_ = new_n15136_ & new_n41133_;
  assign new_n41135_ = ys__n17806 & new_n41019_;
  assign new_n41136_ = new_n39850_ & new_n39862_;
  assign new_n41137_ = ~new_n39850_ & ~new_n39862_;
  assign new_n41138_ = ~new_n41136_ & ~new_n41137_;
  assign new_n41139_ = new_n41024_ & ~new_n41138_;
  assign new_n41140_ = ys__n17809 & new_n17808_;
  assign new_n41141_ = ~ys__n17809 & ~new_n17808_;
  assign new_n41142_ = ~new_n41140_ & ~new_n41141_;
  assign new_n41143_ = new_n41091_ & ~new_n41142_;
  assign new_n41144_ = ~new_n41139_ & ~new_n41143_;
  assign new_n41145_ = ~new_n41135_ & new_n41144_;
  assign new_n41146_ = new_n40821_ & new_n40844_;
  assign new_n41147_ = ~new_n40821_ & ~new_n40844_;
  assign new_n41148_ = ~new_n41146_ & ~new_n41147_;
  assign new_n41149_ = new_n41037_ & ~new_n41148_;
  assign new_n41150_ = new_n40460_ & new_n40482_;
  assign new_n41151_ = ~new_n40460_ & ~new_n40482_;
  assign new_n41152_ = ~new_n41150_ & ~new_n41151_;
  assign new_n41153_ = new_n41043_ & ~new_n41152_;
  assign new_n41154_ = ~new_n41149_ & ~new_n41153_;
  assign new_n41155_ = new_n41145_ & new_n41154_;
  assign new_n41156_ = new_n41051_ & ~new_n41155_;
  assign ys__n30247 = new_n41134_ | new_n41156_;
  assign new_n41158_ = ys__n352 & ys__n23280;
  assign new_n41159_ = new_n15136_ & new_n41158_;
  assign new_n41160_ = ys__n17807 & new_n41019_;
  assign new_n41161_ = new_n39841_ & new_n39863_;
  assign new_n41162_ = ~new_n39841_ & ~new_n39863_;
  assign new_n41163_ = ~new_n41161_ & ~new_n41162_;
  assign new_n41164_ = new_n41024_ & ~new_n41163_;
  assign new_n41165_ = ~ys__n17809 & new_n17808_;
  assign new_n41166_ = ys__n17810 & new_n41165_;
  assign new_n41167_ = ~ys__n17810 & ~new_n41165_;
  assign new_n41168_ = ~new_n41166_ & ~new_n41167_;
  assign new_n41169_ = new_n41091_ & ~new_n41168_;
  assign new_n41170_ = ~new_n41164_ & ~new_n41169_;
  assign new_n41171_ = ~new_n41160_ & new_n41170_;
  assign new_n41172_ = ~new_n40821_ & new_n40844_;
  assign new_n41173_ = new_n40818_ & new_n41172_;
  assign new_n41174_ = ~new_n40818_ & ~new_n41172_;
  assign new_n41175_ = ~new_n41173_ & ~new_n41174_;
  assign new_n41176_ = new_n41037_ & ~new_n41175_;
  assign new_n41177_ = ~new_n40460_ & new_n40482_;
  assign new_n41178_ = new_n40457_ & new_n41177_;
  assign new_n41179_ = ~new_n40457_ & ~new_n41177_;
  assign new_n41180_ = ~new_n41178_ & ~new_n41179_;
  assign new_n41181_ = new_n41043_ & ~new_n41180_;
  assign new_n41182_ = ~new_n41176_ & ~new_n41181_;
  assign new_n41183_ = new_n41171_ & new_n41182_;
  assign new_n41184_ = new_n41051_ & ~new_n41183_;
  assign ys__n30250 = new_n41159_ | new_n41184_;
  assign new_n41186_ = ys__n352 & ys__n23282;
  assign new_n41187_ = new_n15136_ & new_n41186_;
  assign new_n41188_ = ys__n17809 & new_n41019_;
  assign new_n41189_ = ~new_n39841_ & new_n39863_;
  assign new_n41190_ = new_n39838_ & new_n41189_;
  assign new_n41191_ = ~new_n39838_ & ~new_n41189_;
  assign new_n41192_ = ~new_n41190_ & ~new_n41191_;
  assign new_n41193_ = new_n41024_ & ~new_n41192_;
  assign new_n41194_ = new_n17808_ & new_n17809_;
  assign new_n41195_ = ys__n17812 & new_n41194_;
  assign new_n41196_ = ~ys__n17812 & ~new_n41194_;
  assign new_n41197_ = ~new_n41195_ & ~new_n41196_;
  assign new_n41198_ = new_n41091_ & ~new_n41197_;
  assign new_n41199_ = ~new_n41193_ & ~new_n41198_;
  assign new_n41200_ = ~new_n41188_ & new_n41199_;
  assign new_n41201_ = new_n40822_ & new_n40844_;
  assign new_n41202_ = new_n40825_ & new_n41201_;
  assign new_n41203_ = ~new_n40825_ & ~new_n41201_;
  assign new_n41204_ = ~new_n41202_ & ~new_n41203_;
  assign new_n41205_ = new_n41037_ & ~new_n41204_;
  assign new_n41206_ = new_n40461_ & new_n40482_;
  assign new_n41207_ = new_n40464_ & new_n41206_;
  assign new_n41208_ = ~new_n40464_ & ~new_n41206_;
  assign new_n41209_ = ~new_n41207_ & ~new_n41208_;
  assign new_n41210_ = new_n41043_ & ~new_n41209_;
  assign new_n41211_ = ~new_n41205_ & ~new_n41210_;
  assign new_n41212_ = new_n41200_ & new_n41211_;
  assign new_n41213_ = new_n41051_ & ~new_n41212_;
  assign ys__n30253 = new_n41187_ | new_n41213_;
  assign new_n41215_ = ys__n352 & ys__n23284;
  assign new_n41216_ = new_n15136_ & new_n41215_;
  assign new_n41217_ = ys__n17810 & new_n41019_;
  assign new_n41218_ = new_n39842_ & new_n39863_;
  assign new_n41219_ = new_n39845_ & new_n41218_;
  assign new_n41220_ = ~new_n39845_ & ~new_n41218_;
  assign new_n41221_ = ~new_n41219_ & ~new_n41220_;
  assign new_n41222_ = new_n41024_ & ~new_n41221_;
  assign new_n41223_ = ~ys__n17812 & new_n41194_;
  assign new_n41224_ = ys__n17813 & new_n41223_;
  assign new_n41225_ = ~ys__n17813 & ~new_n41223_;
  assign new_n41226_ = ~new_n41224_ & ~new_n41225_;
  assign new_n41227_ = new_n41091_ & ~new_n41226_;
  assign new_n41228_ = ~new_n41222_ & ~new_n41227_;
  assign new_n41229_ = ~new_n41217_ & new_n41228_;
  assign new_n41230_ = ~new_n40825_ & new_n41201_;
  assign new_n41231_ = new_n40813_ & new_n41230_;
  assign new_n41232_ = ~new_n40813_ & ~new_n41230_;
  assign new_n41233_ = ~new_n41231_ & ~new_n41232_;
  assign new_n41234_ = new_n41037_ & ~new_n41233_;
  assign new_n41235_ = ~new_n40464_ & new_n41206_;
  assign new_n41236_ = new_n40452_ & new_n41235_;
  assign new_n41237_ = ~new_n40452_ & ~new_n41235_;
  assign new_n41238_ = ~new_n41236_ & ~new_n41237_;
  assign new_n41239_ = new_n41043_ & ~new_n41238_;
  assign new_n41240_ = ~new_n41234_ & ~new_n41239_;
  assign new_n41241_ = new_n41229_ & new_n41240_;
  assign new_n41242_ = new_n41051_ & ~new_n41241_;
  assign ys__n30256 = new_n41216_ | new_n41242_;
  assign new_n41244_ = ys__n352 & ys__n23286;
  assign new_n41245_ = new_n15136_ & new_n41244_;
  assign new_n41246_ = ys__n17812 & new_n41019_;
  assign new_n41247_ = ~new_n39845_ & new_n41218_;
  assign new_n41248_ = new_n39833_ & new_n41247_;
  assign new_n41249_ = ~new_n39833_ & ~new_n41247_;
  assign new_n41250_ = ~new_n41248_ & ~new_n41249_;
  assign new_n41251_ = new_n41024_ & ~new_n41250_;
  assign new_n41252_ = ys__n17815 & new_n17812_;
  assign new_n41253_ = ~ys__n17815 & ~new_n17812_;
  assign new_n41254_ = ~new_n41252_ & ~new_n41253_;
  assign new_n41255_ = new_n41091_ & ~new_n41254_;
  assign new_n41256_ = ~new_n41251_ & ~new_n41255_;
  assign new_n41257_ = ~new_n41246_ & new_n41256_;
  assign new_n41258_ = new_n40791_ & new_n40847_;
  assign new_n41259_ = ~new_n40791_ & ~new_n40847_;
  assign new_n41260_ = ~new_n41258_ & ~new_n41259_;
  assign new_n41261_ = new_n41037_ & ~new_n41260_;
  assign new_n41262_ = new_n40430_ & new_n40485_;
  assign new_n41263_ = ~new_n40430_ & ~new_n40485_;
  assign new_n41264_ = ~new_n41262_ & ~new_n41263_;
  assign new_n41265_ = new_n41043_ & ~new_n41264_;
  assign new_n41266_ = ~new_n41261_ & ~new_n41265_;
  assign new_n41267_ = new_n41257_ & new_n41266_;
  assign new_n41268_ = new_n41051_ & ~new_n41267_;
  assign ys__n30259 = new_n41245_ | new_n41268_;
  assign new_n41270_ = ys__n352 & ys__n23288;
  assign new_n41271_ = new_n15136_ & new_n41270_;
  assign new_n41272_ = ys__n17813 & new_n41019_;
  assign new_n41273_ = new_n39811_ & new_n39866_;
  assign new_n41274_ = ~new_n39811_ & ~new_n39866_;
  assign new_n41275_ = ~new_n41273_ & ~new_n41274_;
  assign new_n41276_ = new_n41024_ & ~new_n41275_;
  assign new_n41277_ = ~ys__n17815 & new_n17812_;
  assign new_n41278_ = ys__n17816 & new_n41277_;
  assign new_n41279_ = ~ys__n17816 & ~new_n41277_;
  assign new_n41280_ = ~new_n41278_ & ~new_n41279_;
  assign new_n41281_ = new_n41091_ & ~new_n41280_;
  assign new_n41282_ = ~new_n41276_ & ~new_n41281_;
  assign new_n41283_ = ~new_n41272_ & new_n41282_;
  assign new_n41284_ = ~new_n40791_ & new_n40847_;
  assign new_n41285_ = new_n40788_ & new_n41284_;
  assign new_n41286_ = ~new_n40788_ & ~new_n41284_;
  assign new_n41287_ = ~new_n41285_ & ~new_n41286_;
  assign new_n41288_ = new_n41037_ & ~new_n41287_;
  assign new_n41289_ = ~new_n40430_ & new_n40485_;
  assign new_n41290_ = new_n40427_ & new_n41289_;
  assign new_n41291_ = ~new_n40427_ & ~new_n41289_;
  assign new_n41292_ = ~new_n41290_ & ~new_n41291_;
  assign new_n41293_ = new_n41043_ & ~new_n41292_;
  assign new_n41294_ = ~new_n41288_ & ~new_n41293_;
  assign new_n41295_ = new_n41283_ & new_n41294_;
  assign new_n41296_ = new_n41051_ & ~new_n41295_;
  assign ys__n30262 = new_n41271_ | new_n41296_;
  assign new_n41298_ = ys__n352 & ys__n23290;
  assign new_n41299_ = new_n15136_ & new_n41298_;
  assign new_n41300_ = ys__n17815 & new_n41019_;
  assign new_n41301_ = ~new_n39811_ & new_n39866_;
  assign new_n41302_ = new_n39808_ & new_n41301_;
  assign new_n41303_ = ~new_n39808_ & ~new_n41301_;
  assign new_n41304_ = ~new_n41302_ & ~new_n41303_;
  assign new_n41305_ = new_n41024_ & ~new_n41304_;
  assign new_n41306_ = new_n17812_ & new_n17813_;
  assign new_n41307_ = ys__n17818 & new_n41306_;
  assign new_n41308_ = ~ys__n17818 & ~new_n41306_;
  assign new_n41309_ = ~new_n41307_ & ~new_n41308_;
  assign new_n41310_ = new_n41091_ & ~new_n41309_;
  assign new_n41311_ = ~new_n41305_ & ~new_n41310_;
  assign new_n41312_ = ~new_n41300_ & new_n41311_;
  assign new_n41313_ = new_n40792_ & new_n40847_;
  assign new_n41314_ = new_n40783_ & new_n41313_;
  assign new_n41315_ = ~new_n40783_ & ~new_n41313_;
  assign new_n41316_ = ~new_n41314_ & ~new_n41315_;
  assign new_n41317_ = new_n41037_ & ~new_n41316_;
  assign new_n41318_ = new_n40431_ & new_n40485_;
  assign new_n41319_ = new_n40422_ & new_n41318_;
  assign new_n41320_ = ~new_n40422_ & ~new_n41318_;
  assign new_n41321_ = ~new_n41319_ & ~new_n41320_;
  assign new_n41322_ = new_n41043_ & ~new_n41321_;
  assign new_n41323_ = ~new_n41317_ & ~new_n41322_;
  assign new_n41324_ = new_n41312_ & new_n41323_;
  assign new_n41325_ = new_n41051_ & ~new_n41324_;
  assign ys__n30265 = new_n41299_ | new_n41325_;
  assign new_n41327_ = ys__n352 & ys__n23292;
  assign new_n41328_ = new_n15136_ & new_n41327_;
  assign new_n41329_ = ys__n17816 & new_n41019_;
  assign new_n41330_ = new_n39812_ & new_n39866_;
  assign new_n41331_ = new_n39803_ & new_n41330_;
  assign new_n41332_ = ~new_n39803_ & ~new_n41330_;
  assign new_n41333_ = ~new_n41331_ & ~new_n41332_;
  assign new_n41334_ = new_n41024_ & ~new_n41333_;
  assign new_n41335_ = ~ys__n17818 & new_n41306_;
  assign new_n41336_ = ys__n17819 & new_n41335_;
  assign new_n41337_ = ~ys__n17819 & ~new_n41335_;
  assign new_n41338_ = ~new_n41336_ & ~new_n41337_;
  assign new_n41339_ = new_n41091_ & ~new_n41338_;
  assign new_n41340_ = ~new_n41334_ & ~new_n41339_;
  assign new_n41341_ = ~new_n41329_ & new_n41340_;
  assign new_n41342_ = ~new_n40783_ & new_n41313_;
  assign new_n41343_ = new_n40780_ & new_n41342_;
  assign new_n41344_ = ~new_n40780_ & ~new_n41342_;
  assign new_n41345_ = ~new_n41343_ & ~new_n41344_;
  assign new_n41346_ = new_n41037_ & ~new_n41345_;
  assign new_n41347_ = ~new_n40422_ & new_n41318_;
  assign new_n41348_ = new_n40419_ & new_n41347_;
  assign new_n41349_ = ~new_n40419_ & ~new_n41347_;
  assign new_n41350_ = ~new_n41348_ & ~new_n41349_;
  assign new_n41351_ = new_n41043_ & ~new_n41350_;
  assign new_n41352_ = ~new_n41346_ & ~new_n41351_;
  assign new_n41353_ = new_n41341_ & new_n41352_;
  assign new_n41354_ = new_n41051_ & ~new_n41353_;
  assign ys__n30268 = new_n41328_ | new_n41354_;
  assign new_n41356_ = ys__n352 & ys__n23294;
  assign new_n41357_ = new_n15136_ & new_n41356_;
  assign new_n41358_ = ys__n17818 & new_n41019_;
  assign new_n41359_ = ~new_n39803_ & new_n41330_;
  assign new_n41360_ = new_n39800_ & new_n41359_;
  assign new_n41361_ = ~new_n39800_ & ~new_n41359_;
  assign new_n41362_ = ~new_n41360_ & ~new_n41361_;
  assign new_n41363_ = new_n41024_ & ~new_n41362_;
  assign new_n41364_ = new_n17812_ & new_n17815_;
  assign new_n41365_ = ys__n17821 & new_n41364_;
  assign new_n41366_ = ~ys__n17821 & ~new_n41364_;
  assign new_n41367_ = ~new_n41365_ & ~new_n41366_;
  assign new_n41368_ = new_n41091_ & ~new_n41367_;
  assign new_n41369_ = ~new_n41363_ & ~new_n41368_;
  assign new_n41370_ = ~new_n41358_ & new_n41369_;
  assign new_n41371_ = new_n40794_ & new_n40847_;
  assign new_n41372_ = new_n40802_ & new_n41371_;
  assign new_n41373_ = ~new_n40802_ & ~new_n41371_;
  assign new_n41374_ = ~new_n41372_ & ~new_n41373_;
  assign new_n41375_ = new_n41037_ & ~new_n41374_;
  assign new_n41376_ = new_n40433_ & new_n40485_;
  assign new_n41377_ = new_n40441_ & new_n41376_;
  assign new_n41378_ = ~new_n40441_ & ~new_n41376_;
  assign new_n41379_ = ~new_n41377_ & ~new_n41378_;
  assign new_n41380_ = new_n41043_ & ~new_n41379_;
  assign new_n41381_ = ~new_n41375_ & ~new_n41380_;
  assign new_n41382_ = new_n41370_ & new_n41381_;
  assign new_n41383_ = new_n41051_ & ~new_n41382_;
  assign ys__n30271 = new_n41357_ | new_n41383_;
  assign new_n41385_ = ys__n352 & ys__n23296;
  assign new_n41386_ = new_n15136_ & new_n41385_;
  assign new_n41387_ = ys__n17819 & new_n41019_;
  assign new_n41388_ = new_n39814_ & new_n39866_;
  assign new_n41389_ = new_n39822_ & new_n41388_;
  assign new_n41390_ = ~new_n39822_ & ~new_n41388_;
  assign new_n41391_ = ~new_n41389_ & ~new_n41390_;
  assign new_n41392_ = new_n41024_ & ~new_n41391_;
  assign new_n41393_ = ~ys__n17821 & new_n41364_;
  assign new_n41394_ = ys__n17822 & new_n41393_;
  assign new_n41395_ = ~ys__n17822 & ~new_n41393_;
  assign new_n41396_ = ~new_n41394_ & ~new_n41395_;
  assign new_n41397_ = new_n41091_ & ~new_n41396_;
  assign new_n41398_ = ~new_n41392_ & ~new_n41397_;
  assign new_n41399_ = ~new_n41387_ & new_n41398_;
  assign new_n41400_ = ~new_n40802_ & new_n41371_;
  assign new_n41401_ = new_n40799_ & new_n41400_;
  assign new_n41402_ = ~new_n40799_ & ~new_n41400_;
  assign new_n41403_ = ~new_n41401_ & ~new_n41402_;
  assign new_n41404_ = new_n41037_ & ~new_n41403_;
  assign new_n41405_ = ~new_n40441_ & new_n41376_;
  assign new_n41406_ = new_n40438_ & new_n41405_;
  assign new_n41407_ = ~new_n40438_ & ~new_n41405_;
  assign new_n41408_ = ~new_n41406_ & ~new_n41407_;
  assign new_n41409_ = new_n41043_ & ~new_n41408_;
  assign new_n41410_ = ~new_n41404_ & ~new_n41409_;
  assign new_n41411_ = new_n41399_ & new_n41410_;
  assign new_n41412_ = new_n41051_ & ~new_n41411_;
  assign ys__n30274 = new_n41386_ | new_n41412_;
  assign new_n41414_ = ys__n352 & ys__n23298;
  assign new_n41415_ = new_n15136_ & new_n41414_;
  assign new_n41416_ = ys__n17821 & new_n41019_;
  assign new_n41417_ = ~new_n39822_ & new_n41388_;
  assign new_n41418_ = new_n39819_ & new_n41417_;
  assign new_n41419_ = ~new_n39819_ & ~new_n41417_;
  assign new_n41420_ = ~new_n41418_ & ~new_n41419_;
  assign new_n41421_ = new_n41024_ & ~new_n41420_;
  assign new_n41422_ = new_n17816_ & new_n41364_;
  assign new_n41423_ = ys__n17824 & new_n41422_;
  assign new_n41424_ = ~ys__n17824 & ~new_n41422_;
  assign new_n41425_ = ~new_n41423_ & ~new_n41424_;
  assign new_n41426_ = new_n41091_ & ~new_n41425_;
  assign new_n41427_ = ~new_n41421_ & ~new_n41426_;
  assign new_n41428_ = ~new_n41416_ & new_n41427_;
  assign new_n41429_ = new_n40803_ & new_n41371_;
  assign new_n41430_ = new_n40806_ & new_n41429_;
  assign new_n41431_ = ~new_n40806_ & ~new_n41429_;
  assign new_n41432_ = ~new_n41430_ & ~new_n41431_;
  assign new_n41433_ = new_n41037_ & ~new_n41432_;
  assign new_n41434_ = new_n40442_ & new_n41376_;
  assign new_n41435_ = new_n40445_ & new_n41434_;
  assign new_n41436_ = ~new_n40445_ & ~new_n41434_;
  assign new_n41437_ = ~new_n41435_ & ~new_n41436_;
  assign new_n41438_ = new_n41043_ & ~new_n41437_;
  assign new_n41439_ = ~new_n41433_ & ~new_n41438_;
  assign new_n41440_ = new_n41428_ & new_n41439_;
  assign new_n41441_ = new_n41051_ & ~new_n41440_;
  assign ys__n30277 = new_n41415_ | new_n41441_;
  assign new_n41443_ = ys__n352 & ys__n23300;
  assign new_n41444_ = new_n15136_ & new_n41443_;
  assign new_n41445_ = ys__n17822 & new_n41019_;
  assign new_n41446_ = new_n39823_ & new_n41388_;
  assign new_n41447_ = new_n39826_ & new_n41446_;
  assign new_n41448_ = ~new_n39826_ & ~new_n41446_;
  assign new_n41449_ = ~new_n41447_ & ~new_n41448_;
  assign new_n41450_ = new_n41024_ & ~new_n41449_;
  assign new_n41451_ = ~ys__n17824 & new_n41422_;
  assign new_n41452_ = ys__n17825 & new_n41451_;
  assign new_n41453_ = ~ys__n17825 & ~new_n41451_;
  assign new_n41454_ = ~new_n41452_ & ~new_n41453_;
  assign new_n41455_ = new_n41091_ & ~new_n41454_;
  assign new_n41456_ = ~new_n41450_ & ~new_n41455_;
  assign new_n41457_ = ~new_n41445_ & new_n41456_;
  assign new_n41458_ = ~new_n40806_ & new_n41429_;
  assign new_n41459_ = new_n40773_ & new_n41458_;
  assign new_n41460_ = ~new_n40773_ & ~new_n41458_;
  assign new_n41461_ = ~new_n41459_ & ~new_n41460_;
  assign new_n41462_ = new_n41037_ & ~new_n41461_;
  assign new_n41463_ = ~new_n40445_ & new_n41434_;
  assign new_n41464_ = new_n40412_ & new_n41463_;
  assign new_n41465_ = ~new_n40412_ & ~new_n41463_;
  assign new_n41466_ = ~new_n41464_ & ~new_n41465_;
  assign new_n41467_ = new_n41043_ & ~new_n41466_;
  assign new_n41468_ = ~new_n41462_ & ~new_n41467_;
  assign new_n41469_ = new_n41457_ & new_n41468_;
  assign new_n41470_ = new_n41051_ & ~new_n41469_;
  assign ys__n30280 = new_n41444_ | new_n41470_;
  assign new_n41472_ = ys__n352 & ys__n23302;
  assign new_n41473_ = new_n15136_ & new_n41472_;
  assign new_n41474_ = ys__n17824 & new_n41019_;
  assign new_n41475_ = ~new_n39826_ & new_n41446_;
  assign new_n41476_ = new_n39793_ & new_n41475_;
  assign new_n41477_ = ~new_n39793_ & ~new_n41475_;
  assign new_n41478_ = ~new_n41476_ & ~new_n41477_;
  assign new_n41479_ = new_n41024_ & ~new_n41478_;
  assign new_n41480_ = ys__n17827 & new_n17820_;
  assign new_n41481_ = ~ys__n17827 & ~new_n17820_;
  assign new_n41482_ = ~new_n41480_ & ~new_n41481_;
  assign new_n41483_ = new_n41091_ & ~new_n41482_;
  assign new_n41484_ = ~new_n41479_ & ~new_n41483_;
  assign new_n41485_ = ~new_n41474_ & new_n41484_;
  assign new_n41486_ = ~new_n39634_ & new_n40854_;
  assign new_n41487_ = new_n39634_ & ~new_n40854_;
  assign new_n41488_ = ~new_n41486_ & ~new_n41487_;
  assign new_n41489_ = new_n41037_ & ~new_n41488_;
  assign new_n41490_ = new_n40492_ & ~new_n40676_;
  assign new_n41491_ = ~new_n40492_ & new_n40676_;
  assign new_n41492_ = ~new_n41490_ & ~new_n41491_;
  assign new_n41493_ = new_n41043_ & ~new_n41492_;
  assign new_n41494_ = ~new_n41489_ & ~new_n41493_;
  assign new_n41495_ = new_n41485_ & new_n41494_;
  assign new_n41496_ = new_n41051_ & ~new_n41495_;
  assign ys__n30283 = new_n41473_ | new_n41496_;
  assign new_n41498_ = ys__n352 & ys__n23304;
  assign new_n41499_ = new_n15136_ & new_n41498_;
  assign new_n41500_ = ys__n17825 & new_n41019_;
  assign new_n41501_ = new_n39873_ & ~new_n40247_;
  assign new_n41502_ = ~new_n39873_ & new_n40247_;
  assign new_n41503_ = ~new_n41501_ & ~new_n41502_;
  assign new_n41504_ = new_n41024_ & ~new_n41503_;
  assign new_n41505_ = ~ys__n17827 & new_n17820_;
  assign new_n41506_ = ys__n17828 & new_n41505_;
  assign new_n41507_ = ~ys__n17828 & ~new_n41505_;
  assign new_n41508_ = ~new_n41506_ & ~new_n41507_;
  assign new_n41509_ = new_n41091_ & ~new_n41508_;
  assign new_n41510_ = ~new_n41504_ & ~new_n41509_;
  assign new_n41511_ = ~new_n41500_ & new_n41510_;
  assign new_n41512_ = new_n40854_ & ~new_n40987_;
  assign new_n41513_ = ~new_n39634_ & new_n40987_;
  assign new_n41514_ = new_n39634_ & ~new_n40987_;
  assign new_n41515_ = ~new_n41513_ & ~new_n41514_;
  assign new_n41516_ = ~new_n40854_ & ~new_n41515_;
  assign new_n41517_ = ~new_n41512_ & ~new_n41516_;
  assign new_n41518_ = new_n41037_ & ~new_n41517_;
  assign new_n41519_ = new_n40492_ & ~new_n40673_;
  assign new_n41520_ = new_n40673_ & ~new_n40676_;
  assign new_n41521_ = ~new_n40673_ & new_n40676_;
  assign new_n41522_ = ~new_n41520_ & ~new_n41521_;
  assign new_n41523_ = ~new_n40492_ & ~new_n41522_;
  assign new_n41524_ = ~new_n41519_ & ~new_n41523_;
  assign new_n41525_ = new_n41043_ & ~new_n41524_;
  assign new_n41526_ = ~new_n41518_ & ~new_n41525_;
  assign new_n41527_ = new_n41511_ & new_n41526_;
  assign new_n41528_ = new_n41051_ & ~new_n41527_;
  assign ys__n30286 = new_n41499_ | new_n41528_;
  assign new_n41530_ = ys__n352 & ys__n23306;
  assign new_n41531_ = new_n15136_ & new_n41530_;
  assign new_n41532_ = ys__n17827 & new_n41019_;
  assign new_n41533_ = new_n39873_ & ~new_n40244_;
  assign new_n41534_ = new_n40244_ & ~new_n40247_;
  assign new_n41535_ = ~new_n40244_ & new_n40247_;
  assign new_n41536_ = ~new_n41534_ & ~new_n41535_;
  assign new_n41537_ = ~new_n39873_ & ~new_n41536_;
  assign new_n41538_ = ~new_n41533_ & ~new_n41537_;
  assign new_n41539_ = new_n41024_ & ~new_n41538_;
  assign new_n41540_ = new_n17790_ & new_n17820_;
  assign new_n41541_ = ys__n17830 & new_n41540_;
  assign new_n41542_ = ~ys__n17830 & ~new_n41540_;
  assign new_n41543_ = ~new_n41541_ & ~new_n41542_;
  assign new_n41544_ = new_n41091_ & ~new_n41543_;
  assign new_n41545_ = ~new_n41539_ & ~new_n41544_;
  assign new_n41546_ = ~new_n41532_ & new_n41545_;
  assign new_n41547_ = new_n40854_ & ~new_n40984_;
  assign new_n41548_ = new_n40984_ & new_n40988_;
  assign new_n41549_ = ~new_n40984_ & ~new_n40988_;
  assign new_n41550_ = ~new_n41548_ & ~new_n41549_;
  assign new_n41551_ = ~new_n40854_ & ~new_n41550_;
  assign new_n41552_ = ~new_n41547_ & ~new_n41551_;
  assign new_n41553_ = new_n41037_ & ~new_n41552_;
  assign new_n41554_ = new_n40492_ & ~new_n40670_;
  assign new_n41555_ = new_n40670_ & new_n40677_;
  assign new_n41556_ = ~new_n40670_ & ~new_n40677_;
  assign new_n41557_ = ~new_n41555_ & ~new_n41556_;
  assign new_n41558_ = ~new_n40492_ & ~new_n41557_;
  assign new_n41559_ = ~new_n41554_ & ~new_n41558_;
  assign new_n41560_ = new_n41043_ & ~new_n41559_;
  assign new_n41561_ = ~new_n41553_ & ~new_n41560_;
  assign new_n41562_ = new_n41546_ & new_n41561_;
  assign new_n41563_ = new_n41051_ & ~new_n41562_;
  assign ys__n30289 = new_n41531_ | new_n41563_;
  assign new_n41565_ = ys__n352 & ys__n23308;
  assign new_n41566_ = new_n15136_ & new_n41565_;
  assign new_n41567_ = ys__n17828 & new_n41019_;
  assign new_n41568_ = new_n39873_ & ~new_n40241_;
  assign new_n41569_ = new_n40241_ & new_n40248_;
  assign new_n41570_ = ~new_n40241_ & ~new_n40248_;
  assign new_n41571_ = ~new_n41569_ & ~new_n41570_;
  assign new_n41572_ = ~new_n39873_ & ~new_n41571_;
  assign new_n41573_ = ~new_n41568_ & ~new_n41572_;
  assign new_n41574_ = new_n41024_ & ~new_n41573_;
  assign new_n41575_ = ~ys__n17830 & new_n41540_;
  assign new_n41576_ = ys__n17831 & new_n41575_;
  assign new_n41577_ = ~ys__n17831 & ~new_n41575_;
  assign new_n41578_ = ~new_n41576_ & ~new_n41577_;
  assign new_n41579_ = new_n41091_ & ~new_n41578_;
  assign new_n41580_ = ~new_n41574_ & ~new_n41579_;
  assign new_n41581_ = ~new_n41567_ & new_n41580_;
  assign new_n41582_ = new_n40854_ & ~new_n40981_;
  assign new_n41583_ = new_n40981_ & new_n40989_;
  assign new_n41584_ = ~new_n40981_ & ~new_n40989_;
  assign new_n41585_ = ~new_n41583_ & ~new_n41584_;
  assign new_n41586_ = ~new_n40854_ & ~new_n41585_;
  assign new_n41587_ = ~new_n41582_ & ~new_n41586_;
  assign new_n41588_ = new_n41037_ & ~new_n41587_;
  assign new_n41589_ = new_n40492_ & ~new_n40667_;
  assign new_n41590_ = new_n40667_ & new_n40678_;
  assign new_n41591_ = ~new_n40667_ & ~new_n40678_;
  assign new_n41592_ = ~new_n41590_ & ~new_n41591_;
  assign new_n41593_ = ~new_n40492_ & ~new_n41592_;
  assign new_n41594_ = ~new_n41589_ & ~new_n41593_;
  assign new_n41595_ = new_n41043_ & ~new_n41594_;
  assign new_n41596_ = ~new_n41588_ & ~new_n41595_;
  assign new_n41597_ = new_n41581_ & new_n41596_;
  assign new_n41598_ = new_n41051_ & ~new_n41597_;
  assign ys__n30292 = new_n41566_ | new_n41598_;
  assign new_n41600_ = ys__n352 & ys__n23310;
  assign new_n41601_ = new_n15136_ & new_n41600_;
  assign new_n41602_ = ys__n17830 & new_n41019_;
  assign new_n41603_ = new_n39873_ & ~new_n40238_;
  assign new_n41604_ = new_n40238_ & new_n40249_;
  assign new_n41605_ = ~new_n40238_ & ~new_n40249_;
  assign new_n41606_ = ~new_n41604_ & ~new_n41605_;
  assign new_n41607_ = ~new_n39873_ & ~new_n41606_;
  assign new_n41608_ = ~new_n41603_ & ~new_n41607_;
  assign new_n41609_ = new_n41024_ & ~new_n41608_;
  assign new_n41610_ = new_n17792_ & new_n17820_;
  assign new_n41611_ = ys__n17833 & new_n41610_;
  assign new_n41612_ = ~ys__n17833 & ~new_n41610_;
  assign new_n41613_ = ~new_n41611_ & ~new_n41612_;
  assign new_n41614_ = new_n41091_ & ~new_n41613_;
  assign new_n41615_ = ~new_n41609_ & ~new_n41614_;
  assign new_n41616_ = ~new_n41602_ & new_n41615_;
  assign new_n41617_ = new_n40854_ & ~new_n40972_;
  assign new_n41618_ = new_n40972_ & new_n40990_;
  assign new_n41619_ = ~new_n40972_ & ~new_n40990_;
  assign new_n41620_ = ~new_n41618_ & ~new_n41619_;
  assign new_n41621_ = ~new_n40854_ & ~new_n41620_;
  assign new_n41622_ = ~new_n41617_ & ~new_n41621_;
  assign new_n41623_ = new_n41037_ & ~new_n41622_;
  assign new_n41624_ = new_n40492_ & ~new_n40658_;
  assign new_n41625_ = new_n40658_ & new_n40679_;
  assign new_n41626_ = ~new_n40658_ & ~new_n40679_;
  assign new_n41627_ = ~new_n41625_ & ~new_n41626_;
  assign new_n41628_ = ~new_n40492_ & ~new_n41627_;
  assign new_n41629_ = ~new_n41624_ & ~new_n41628_;
  assign new_n41630_ = new_n41043_ & ~new_n41629_;
  assign new_n41631_ = ~new_n41623_ & ~new_n41630_;
  assign new_n41632_ = new_n41616_ & new_n41631_;
  assign new_n41633_ = new_n41051_ & ~new_n41632_;
  assign ys__n30295 = new_n41601_ | new_n41633_;
  assign new_n41635_ = ys__n352 & ys__n23312;
  assign new_n41636_ = new_n15136_ & new_n41635_;
  assign new_n41637_ = ys__n17831 & new_n41019_;
  assign new_n41638_ = new_n39873_ & ~new_n40229_;
  assign new_n41639_ = new_n40229_ & new_n40250_;
  assign new_n41640_ = ~new_n40229_ & ~new_n40250_;
  assign new_n41641_ = ~new_n41639_ & ~new_n41640_;
  assign new_n41642_ = ~new_n39873_ & ~new_n41641_;
  assign new_n41643_ = ~new_n41638_ & ~new_n41642_;
  assign new_n41644_ = new_n41024_ & ~new_n41643_;
  assign new_n41645_ = ~ys__n17833 & new_n41610_;
  assign new_n41646_ = ys__n17834 & new_n41645_;
  assign new_n41647_ = ~ys__n17834 & ~new_n41645_;
  assign new_n41648_ = ~new_n41646_ & ~new_n41647_;
  assign new_n41649_ = new_n41091_ & ~new_n41648_;
  assign new_n41650_ = ~new_n41644_ & ~new_n41649_;
  assign new_n41651_ = ~new_n41637_ & new_n41650_;
  assign new_n41652_ = new_n40854_ & ~new_n40969_;
  assign new_n41653_ = ~new_n40972_ & new_n40990_;
  assign new_n41654_ = new_n40969_ & new_n41653_;
  assign new_n41655_ = ~new_n40969_ & ~new_n41653_;
  assign new_n41656_ = ~new_n41654_ & ~new_n41655_;
  assign new_n41657_ = ~new_n40854_ & ~new_n41656_;
  assign new_n41658_ = ~new_n41652_ & ~new_n41657_;
  assign new_n41659_ = new_n41037_ & ~new_n41658_;
  assign new_n41660_ = new_n40492_ & ~new_n40655_;
  assign new_n41661_ = ~new_n40658_ & new_n40679_;
  assign new_n41662_ = new_n40655_ & new_n41661_;
  assign new_n41663_ = ~new_n40655_ & ~new_n41661_;
  assign new_n41664_ = ~new_n41662_ & ~new_n41663_;
  assign new_n41665_ = ~new_n40492_ & ~new_n41664_;
  assign new_n41666_ = ~new_n41660_ & ~new_n41665_;
  assign new_n41667_ = new_n41043_ & ~new_n41666_;
  assign new_n41668_ = ~new_n41659_ & ~new_n41667_;
  assign new_n41669_ = new_n41651_ & new_n41668_;
  assign new_n41670_ = new_n41051_ & ~new_n41669_;
  assign ys__n30298 = new_n41636_ | new_n41670_;
  assign new_n41672_ = ys__n352 & ys__n23314;
  assign new_n41673_ = new_n15136_ & new_n41672_;
  assign new_n41674_ = ys__n17833 & new_n41019_;
  assign new_n41675_ = new_n39873_ & ~new_n40226_;
  assign new_n41676_ = ~new_n40229_ & new_n40250_;
  assign new_n41677_ = new_n40226_ & new_n41676_;
  assign new_n41678_ = ~new_n40226_ & ~new_n41676_;
  assign new_n41679_ = ~new_n41677_ & ~new_n41678_;
  assign new_n41680_ = ~new_n39873_ & ~new_n41679_;
  assign new_n41681_ = ~new_n41675_ & ~new_n41680_;
  assign new_n41682_ = new_n41024_ & ~new_n41681_;
  assign new_n41683_ = new_n17793_ & new_n41610_;
  assign new_n41684_ = ys__n17836 & new_n41683_;
  assign new_n41685_ = ~ys__n17836 & ~new_n41683_;
  assign new_n41686_ = ~new_n41684_ & ~new_n41685_;
  assign new_n41687_ = new_n41091_ & ~new_n41686_;
  assign new_n41688_ = ~new_n41682_ & ~new_n41687_;
  assign new_n41689_ = ~new_n41674_ & new_n41688_;
  assign new_n41690_ = new_n40854_ & ~new_n40976_;
  assign new_n41691_ = new_n40973_ & new_n40990_;
  assign new_n41692_ = new_n40976_ & new_n41691_;
  assign new_n41693_ = ~new_n40976_ & ~new_n41691_;
  assign new_n41694_ = ~new_n41692_ & ~new_n41693_;
  assign new_n41695_ = ~new_n40854_ & ~new_n41694_;
  assign new_n41696_ = ~new_n41690_ & ~new_n41695_;
  assign new_n41697_ = new_n41037_ & ~new_n41696_;
  assign new_n41698_ = new_n40492_ & ~new_n40662_;
  assign new_n41699_ = new_n40659_ & new_n40679_;
  assign new_n41700_ = new_n40662_ & new_n41699_;
  assign new_n41701_ = ~new_n40662_ & ~new_n41699_;
  assign new_n41702_ = ~new_n41700_ & ~new_n41701_;
  assign new_n41703_ = ~new_n40492_ & ~new_n41702_;
  assign new_n41704_ = ~new_n41698_ & ~new_n41703_;
  assign new_n41705_ = new_n41043_ & ~new_n41704_;
  assign new_n41706_ = ~new_n41697_ & ~new_n41705_;
  assign new_n41707_ = new_n41689_ & new_n41706_;
  assign new_n41708_ = new_n41051_ & ~new_n41707_;
  assign ys__n30301 = new_n41673_ | new_n41708_;
  assign new_n41710_ = ys__n352 & ys__n23316;
  assign new_n41711_ = new_n15136_ & new_n41710_;
  assign new_n41712_ = ys__n17834 & new_n41019_;
  assign new_n41713_ = new_n39873_ & ~new_n40233_;
  assign new_n41714_ = new_n40230_ & new_n40250_;
  assign new_n41715_ = new_n40233_ & new_n41714_;
  assign new_n41716_ = ~new_n40233_ & ~new_n41714_;
  assign new_n41717_ = ~new_n41715_ & ~new_n41716_;
  assign new_n41718_ = ~new_n39873_ & ~new_n41717_;
  assign new_n41719_ = ~new_n41713_ & ~new_n41718_;
  assign new_n41720_ = new_n41024_ & ~new_n41719_;
  assign new_n41721_ = ~ys__n17836 & new_n41683_;
  assign new_n41722_ = ys__n17837 & new_n41721_;
  assign new_n41723_ = ~ys__n17837 & ~new_n41721_;
  assign new_n41724_ = ~new_n41722_ & ~new_n41723_;
  assign new_n41725_ = new_n41091_ & ~new_n41724_;
  assign new_n41726_ = ~new_n41720_ & ~new_n41725_;
  assign new_n41727_ = ~new_n41712_ & new_n41726_;
  assign new_n41728_ = new_n40854_ & ~new_n40964_;
  assign new_n41729_ = ~new_n40976_ & new_n41691_;
  assign new_n41730_ = new_n40964_ & new_n41729_;
  assign new_n41731_ = ~new_n40964_ & ~new_n41729_;
  assign new_n41732_ = ~new_n41730_ & ~new_n41731_;
  assign new_n41733_ = ~new_n40854_ & ~new_n41732_;
  assign new_n41734_ = ~new_n41728_ & ~new_n41733_;
  assign new_n41735_ = new_n41037_ & ~new_n41734_;
  assign new_n41736_ = new_n40492_ & ~new_n40650_;
  assign new_n41737_ = ~new_n40662_ & new_n41699_;
  assign new_n41738_ = new_n40650_ & new_n41737_;
  assign new_n41739_ = ~new_n40650_ & ~new_n41737_;
  assign new_n41740_ = ~new_n41738_ & ~new_n41739_;
  assign new_n41741_ = ~new_n40492_ & ~new_n41740_;
  assign new_n41742_ = ~new_n41736_ & ~new_n41741_;
  assign new_n41743_ = new_n41043_ & ~new_n41742_;
  assign new_n41744_ = ~new_n41735_ & ~new_n41743_;
  assign new_n41745_ = new_n41727_ & new_n41744_;
  assign new_n41746_ = new_n41051_ & ~new_n41745_;
  assign ys__n30304 = new_n41711_ | new_n41746_;
  assign new_n41748_ = ys__n352 & ys__n23318;
  assign new_n41749_ = new_n15136_ & new_n41748_;
  assign new_n41750_ = ys__n17836 & new_n41019_;
  assign new_n41751_ = new_n39873_ & ~new_n40221_;
  assign new_n41752_ = ~new_n40233_ & new_n41714_;
  assign new_n41753_ = new_n40221_ & new_n41752_;
  assign new_n41754_ = ~new_n40221_ & ~new_n41752_;
  assign new_n41755_ = ~new_n41753_ & ~new_n41754_;
  assign new_n41756_ = ~new_n39873_ & ~new_n41755_;
  assign new_n41757_ = ~new_n41751_ & ~new_n41756_;
  assign new_n41758_ = new_n41024_ & ~new_n41757_;
  assign new_n41759_ = new_n17796_ & new_n17820_;
  assign new_n41760_ = ys__n17839 & new_n41759_;
  assign new_n41761_ = ~ys__n17839 & ~new_n41759_;
  assign new_n41762_ = ~new_n41760_ & ~new_n41761_;
  assign new_n41763_ = new_n41091_ & ~new_n41762_;
  assign new_n41764_ = ~new_n41758_ & ~new_n41763_;
  assign new_n41765_ = ~new_n41750_ & new_n41764_;
  assign new_n41766_ = new_n40854_ & ~new_n40942_;
  assign new_n41767_ = new_n40942_ & new_n40993_;
  assign new_n41768_ = ~new_n40942_ & ~new_n40993_;
  assign new_n41769_ = ~new_n41767_ & ~new_n41768_;
  assign new_n41770_ = ~new_n40854_ & ~new_n41769_;
  assign new_n41771_ = ~new_n41766_ & ~new_n41770_;
  assign new_n41772_ = new_n41037_ & ~new_n41771_;
  assign new_n41773_ = new_n40492_ & ~new_n40628_;
  assign new_n41774_ = new_n40628_ & new_n40682_;
  assign new_n41775_ = ~new_n40628_ & ~new_n40682_;
  assign new_n41776_ = ~new_n41774_ & ~new_n41775_;
  assign new_n41777_ = ~new_n40492_ & ~new_n41776_;
  assign new_n41778_ = ~new_n41773_ & ~new_n41777_;
  assign new_n41779_ = new_n41043_ & ~new_n41778_;
  assign new_n41780_ = ~new_n41772_ & ~new_n41779_;
  assign new_n41781_ = new_n41765_ & new_n41780_;
  assign new_n41782_ = new_n41051_ & ~new_n41781_;
  assign ys__n30307 = new_n41749_ | new_n41782_;
  assign new_n41784_ = ys__n352 & ys__n23320;
  assign new_n41785_ = new_n15136_ & new_n41784_;
  assign new_n41786_ = ys__n17837 & new_n41019_;
  assign new_n41787_ = new_n39873_ & ~new_n40211_;
  assign new_n41788_ = new_n40211_ & new_n40253_;
  assign new_n41789_ = ~new_n40211_ & ~new_n40253_;
  assign new_n41790_ = ~new_n41788_ & ~new_n41789_;
  assign new_n41791_ = ~new_n39873_ & ~new_n41790_;
  assign new_n41792_ = ~new_n41787_ & ~new_n41791_;
  assign new_n41793_ = new_n41024_ & ~new_n41792_;
  assign new_n41794_ = ~ys__n17839 & new_n41759_;
  assign new_n41795_ = ys__n17840 & new_n41794_;
  assign new_n41796_ = ~ys__n17840 & ~new_n41794_;
  assign new_n41797_ = ~new_n41795_ & ~new_n41796_;
  assign new_n41798_ = new_n41091_ & ~new_n41797_;
  assign new_n41799_ = ~new_n41793_ & ~new_n41798_;
  assign new_n41800_ = ~new_n41786_ & new_n41799_;
  assign new_n41801_ = new_n40854_ & ~new_n40939_;
  assign new_n41802_ = ~new_n40942_ & new_n40993_;
  assign new_n41803_ = new_n40939_ & new_n41802_;
  assign new_n41804_ = ~new_n40939_ & ~new_n41802_;
  assign new_n41805_ = ~new_n41803_ & ~new_n41804_;
  assign new_n41806_ = ~new_n40854_ & ~new_n41805_;
  assign new_n41807_ = ~new_n41801_ & ~new_n41806_;
  assign new_n41808_ = new_n41037_ & ~new_n41807_;
  assign new_n41809_ = new_n40492_ & ~new_n40625_;
  assign new_n41810_ = ~new_n40628_ & new_n40682_;
  assign new_n41811_ = new_n40625_ & new_n41810_;
  assign new_n41812_ = ~new_n40625_ & ~new_n41810_;
  assign new_n41813_ = ~new_n41811_ & ~new_n41812_;
  assign new_n41814_ = ~new_n40492_ & ~new_n41813_;
  assign new_n41815_ = ~new_n41809_ & ~new_n41814_;
  assign new_n41816_ = new_n41043_ & ~new_n41815_;
  assign new_n41817_ = ~new_n41808_ & ~new_n41816_;
  assign new_n41818_ = new_n41800_ & new_n41817_;
  assign new_n41819_ = new_n41051_ & ~new_n41818_;
  assign ys__n30310 = new_n41785_ | new_n41819_;
  assign new_n41821_ = ys__n352 & ys__n23322;
  assign new_n41822_ = new_n15136_ & new_n41821_;
  assign new_n41823_ = ys__n17839 & new_n41019_;
  assign new_n41824_ = new_n39873_ & ~new_n40208_;
  assign new_n41825_ = ~new_n40211_ & new_n40253_;
  assign new_n41826_ = new_n40208_ & new_n41825_;
  assign new_n41827_ = ~new_n40208_ & ~new_n41825_;
  assign new_n41828_ = ~new_n41826_ & ~new_n41827_;
  assign new_n41829_ = ~new_n39873_ & ~new_n41828_;
  assign new_n41830_ = ~new_n41824_ & ~new_n41829_;
  assign new_n41831_ = new_n41024_ & ~new_n41830_;
  assign new_n41832_ = new_n17828_ & new_n41759_;
  assign new_n41833_ = ys__n17842 & new_n41832_;
  assign new_n41834_ = ~ys__n17842 & ~new_n41832_;
  assign new_n41835_ = ~new_n41833_ & ~new_n41834_;
  assign new_n41836_ = new_n41091_ & ~new_n41835_;
  assign new_n41837_ = ~new_n41831_ & ~new_n41836_;
  assign new_n41838_ = ~new_n41823_ & new_n41837_;
  assign new_n41839_ = new_n40854_ & ~new_n40934_;
  assign new_n41840_ = new_n40943_ & new_n40993_;
  assign new_n41841_ = new_n40934_ & new_n41840_;
  assign new_n41842_ = ~new_n40934_ & ~new_n41840_;
  assign new_n41843_ = ~new_n41841_ & ~new_n41842_;
  assign new_n41844_ = ~new_n40854_ & ~new_n41843_;
  assign new_n41845_ = ~new_n41839_ & ~new_n41844_;
  assign new_n41846_ = new_n41037_ & ~new_n41845_;
  assign new_n41847_ = new_n40492_ & ~new_n40620_;
  assign new_n41848_ = new_n40629_ & new_n40682_;
  assign new_n41849_ = new_n40620_ & new_n41848_;
  assign new_n41850_ = ~new_n40620_ & ~new_n41848_;
  assign new_n41851_ = ~new_n41849_ & ~new_n41850_;
  assign new_n41852_ = ~new_n40492_ & ~new_n41851_;
  assign new_n41853_ = ~new_n41847_ & ~new_n41852_;
  assign new_n41854_ = new_n41043_ & ~new_n41853_;
  assign new_n41855_ = ~new_n41846_ & ~new_n41854_;
  assign new_n41856_ = new_n41838_ & new_n41855_;
  assign new_n41857_ = new_n41051_ & ~new_n41856_;
  assign ys__n30313 = new_n41822_ | new_n41857_;
  assign new_n41859_ = ys__n352 & ys__n23324;
  assign new_n41860_ = new_n15136_ & new_n41859_;
  assign new_n41861_ = ys__n17840 & new_n41019_;
  assign new_n41862_ = new_n39873_ & ~new_n40203_;
  assign new_n41863_ = new_n40212_ & new_n40253_;
  assign new_n41864_ = new_n40203_ & new_n41863_;
  assign new_n41865_ = ~new_n40203_ & ~new_n41863_;
  assign new_n41866_ = ~new_n41864_ & ~new_n41865_;
  assign new_n41867_ = ~new_n39873_ & ~new_n41866_;
  assign new_n41868_ = ~new_n41862_ & ~new_n41867_;
  assign new_n41869_ = new_n41024_ & ~new_n41868_;
  assign new_n41870_ = ~ys__n17842 & new_n41832_;
  assign new_n41871_ = ys__n17843 & new_n41870_;
  assign new_n41872_ = ~ys__n17843 & ~new_n41870_;
  assign new_n41873_ = ~new_n41871_ & ~new_n41872_;
  assign new_n41874_ = new_n41091_ & ~new_n41873_;
  assign new_n41875_ = ~new_n41869_ & ~new_n41874_;
  assign new_n41876_ = ~new_n41861_ & new_n41875_;
  assign new_n41877_ = new_n40854_ & ~new_n40931_;
  assign new_n41878_ = ~new_n40934_ & new_n41840_;
  assign new_n41879_ = new_n40931_ & new_n41878_;
  assign new_n41880_ = ~new_n40931_ & ~new_n41878_;
  assign new_n41881_ = ~new_n41879_ & ~new_n41880_;
  assign new_n41882_ = ~new_n40854_ & ~new_n41881_;
  assign new_n41883_ = ~new_n41877_ & ~new_n41882_;
  assign new_n41884_ = new_n41037_ & ~new_n41883_;
  assign new_n41885_ = new_n40492_ & ~new_n40617_;
  assign new_n41886_ = ~new_n40620_ & new_n41848_;
  assign new_n41887_ = new_n40617_ & new_n41886_;
  assign new_n41888_ = ~new_n40617_ & ~new_n41886_;
  assign new_n41889_ = ~new_n41887_ & ~new_n41888_;
  assign new_n41890_ = ~new_n40492_ & ~new_n41889_;
  assign new_n41891_ = ~new_n41885_ & ~new_n41890_;
  assign new_n41892_ = new_n41043_ & ~new_n41891_;
  assign new_n41893_ = ~new_n41884_ & ~new_n41892_;
  assign new_n41894_ = new_n41876_ & new_n41893_;
  assign new_n41895_ = new_n41051_ & ~new_n41894_;
  assign ys__n30316 = new_n41860_ | new_n41895_;
  assign new_n41897_ = ys__n352 & ys__n23326;
  assign new_n41898_ = new_n15136_ & new_n41897_;
  assign new_n41899_ = ys__n17842 & new_n41019_;
  assign new_n41900_ = new_n39873_ & ~new_n40200_;
  assign new_n41901_ = ~new_n40203_ & new_n41863_;
  assign new_n41902_ = new_n40200_ & new_n41901_;
  assign new_n41903_ = ~new_n40200_ & ~new_n41901_;
  assign new_n41904_ = ~new_n41902_ & ~new_n41903_;
  assign new_n41905_ = ~new_n39873_ & ~new_n41904_;
  assign new_n41906_ = ~new_n41900_ & ~new_n41905_;
  assign new_n41907_ = new_n41024_ & ~new_n41906_;
  assign new_n41908_ = new_n17830_ & new_n41759_;
  assign new_n41909_ = ys__n17845 & new_n41908_;
  assign new_n41910_ = ~ys__n17845 & ~new_n41908_;
  assign new_n41911_ = ~new_n41909_ & ~new_n41910_;
  assign new_n41912_ = new_n41091_ & ~new_n41911_;
  assign new_n41913_ = ~new_n41907_ & ~new_n41912_;
  assign new_n41914_ = ~new_n41899_ & new_n41913_;
  assign new_n41915_ = new_n40854_ & ~new_n40953_;
  assign new_n41916_ = new_n40945_ & new_n40993_;
  assign new_n41917_ = new_n40953_ & new_n41916_;
  assign new_n41918_ = ~new_n40953_ & ~new_n41916_;
  assign new_n41919_ = ~new_n41917_ & ~new_n41918_;
  assign new_n41920_ = ~new_n40854_ & ~new_n41919_;
  assign new_n41921_ = ~new_n41915_ & ~new_n41920_;
  assign new_n41922_ = new_n41037_ & ~new_n41921_;
  assign new_n41923_ = new_n40492_ & ~new_n40639_;
  assign new_n41924_ = new_n40631_ & new_n40682_;
  assign new_n41925_ = new_n40639_ & new_n41924_;
  assign new_n41926_ = ~new_n40639_ & ~new_n41924_;
  assign new_n41927_ = ~new_n41925_ & ~new_n41926_;
  assign new_n41928_ = ~new_n40492_ & ~new_n41927_;
  assign new_n41929_ = ~new_n41923_ & ~new_n41928_;
  assign new_n41930_ = new_n41043_ & ~new_n41929_;
  assign new_n41931_ = ~new_n41922_ & ~new_n41930_;
  assign new_n41932_ = new_n41914_ & new_n41931_;
  assign new_n41933_ = new_n41051_ & ~new_n41932_;
  assign ys__n30319 = new_n41898_ | new_n41933_;
  assign new_n41935_ = ys__n352 & ys__n23328;
  assign new_n41936_ = new_n15136_ & new_n41935_;
  assign new_n41937_ = ys__n17843 & new_n41019_;
  assign new_n41938_ = new_n39873_ & ~new_n40192_;
  assign new_n41939_ = new_n40192_ & new_n40254_;
  assign new_n41940_ = ~new_n40192_ & ~new_n40254_;
  assign new_n41941_ = ~new_n41939_ & ~new_n41940_;
  assign new_n41942_ = ~new_n39873_ & ~new_n41941_;
  assign new_n41943_ = ~new_n41938_ & ~new_n41942_;
  assign new_n41944_ = new_n41024_ & ~new_n41943_;
  assign new_n41945_ = ~ys__n17845 & new_n41908_;
  assign new_n41946_ = ys__n17846 & new_n41945_;
  assign new_n41947_ = ~ys__n17846 & ~new_n41945_;
  assign new_n41948_ = ~new_n41946_ & ~new_n41947_;
  assign new_n41949_ = new_n41091_ & ~new_n41948_;
  assign new_n41950_ = ~new_n41944_ & ~new_n41949_;
  assign new_n41951_ = ~new_n41937_ & new_n41950_;
  assign new_n41952_ = new_n40854_ & ~new_n40950_;
  assign new_n41953_ = ~new_n40953_ & new_n41916_;
  assign new_n41954_ = new_n40950_ & new_n41953_;
  assign new_n41955_ = ~new_n40950_ & ~new_n41953_;
  assign new_n41956_ = ~new_n41954_ & ~new_n41955_;
  assign new_n41957_ = ~new_n40854_ & ~new_n41956_;
  assign new_n41958_ = ~new_n41952_ & ~new_n41957_;
  assign new_n41959_ = new_n41037_ & ~new_n41958_;
  assign new_n41960_ = new_n40492_ & ~new_n40636_;
  assign new_n41961_ = ~new_n40639_ & new_n41924_;
  assign new_n41962_ = new_n40636_ & new_n41961_;
  assign new_n41963_ = ~new_n40636_ & ~new_n41961_;
  assign new_n41964_ = ~new_n41962_ & ~new_n41963_;
  assign new_n41965_ = ~new_n40492_ & ~new_n41964_;
  assign new_n41966_ = ~new_n41960_ & ~new_n41965_;
  assign new_n41967_ = new_n41043_ & ~new_n41966_;
  assign new_n41968_ = ~new_n41959_ & ~new_n41967_;
  assign new_n41969_ = new_n41951_ & new_n41968_;
  assign new_n41970_ = new_n41051_ & ~new_n41969_;
  assign ys__n30322 = new_n41936_ | new_n41970_;
  assign new_n41972_ = ys__n352 & ys__n23330;
  assign new_n41973_ = new_n15136_ & new_n41972_;
  assign new_n41974_ = ys__n17845 & new_n41019_;
  assign new_n41975_ = new_n39873_ & ~new_n40189_;
  assign new_n41976_ = ~new_n40192_ & new_n40254_;
  assign new_n41977_ = new_n40189_ & new_n41976_;
  assign new_n41978_ = ~new_n40189_ & ~new_n41976_;
  assign new_n41979_ = ~new_n41977_ & ~new_n41978_;
  assign new_n41980_ = ~new_n39873_ & ~new_n41979_;
  assign new_n41981_ = ~new_n41975_ & ~new_n41980_;
  assign new_n41982_ = new_n41024_ & ~new_n41981_;
  assign new_n41983_ = new_n17800_ & new_n41908_;
  assign new_n41984_ = ys__n17848 & new_n41983_;
  assign new_n41985_ = ~ys__n17848 & ~new_n41983_;
  assign new_n41986_ = ~new_n41984_ & ~new_n41985_;
  assign new_n41987_ = new_n41091_ & ~new_n41986_;
  assign new_n41988_ = ~new_n41982_ & ~new_n41987_;
  assign new_n41989_ = ~new_n41974_ & new_n41988_;
  assign new_n41990_ = new_n40854_ & ~new_n40957_;
  assign new_n41991_ = new_n40954_ & new_n41916_;
  assign new_n41992_ = new_n40957_ & new_n41991_;
  assign new_n41993_ = ~new_n40957_ & ~new_n41991_;
  assign new_n41994_ = ~new_n41992_ & ~new_n41993_;
  assign new_n41995_ = ~new_n40854_ & ~new_n41994_;
  assign new_n41996_ = ~new_n41990_ & ~new_n41995_;
  assign new_n41997_ = new_n41037_ & ~new_n41996_;
  assign new_n41998_ = new_n40492_ & ~new_n40643_;
  assign new_n41999_ = new_n40640_ & new_n41924_;
  assign new_n42000_ = new_n40643_ & new_n41999_;
  assign new_n42001_ = ~new_n40643_ & ~new_n41999_;
  assign new_n42002_ = ~new_n42000_ & ~new_n42001_;
  assign new_n42003_ = ~new_n40492_ & ~new_n42002_;
  assign new_n42004_ = ~new_n41998_ & ~new_n42003_;
  assign new_n42005_ = new_n41043_ & ~new_n42004_;
  assign new_n42006_ = ~new_n41997_ & ~new_n42005_;
  assign new_n42007_ = new_n41989_ & new_n42006_;
  assign new_n42008_ = new_n41051_ & ~new_n42007_;
  assign ys__n30325 = new_n41973_ | new_n42008_;
  assign new_n42010_ = ys__n352 & ys__n23332;
  assign new_n42011_ = new_n15136_ & new_n42010_;
  assign new_n42012_ = ys__n17846 & new_n41019_;
  assign new_n42013_ = new_n39873_ & ~new_n40184_;
  assign new_n42014_ = new_n40184_ & new_n40255_;
  assign new_n42015_ = ~new_n40184_ & ~new_n40255_;
  assign new_n42016_ = ~new_n42014_ & ~new_n42015_;
  assign new_n42017_ = ~new_n39873_ & ~new_n42016_;
  assign new_n42018_ = ~new_n42013_ & ~new_n42017_;
  assign new_n42019_ = new_n41024_ & ~new_n42018_;
  assign new_n42020_ = ~ys__n17848 & new_n41983_;
  assign new_n42021_ = ys__n17849 & new_n42020_;
  assign new_n42022_ = ~ys__n17849 & ~new_n42020_;
  assign new_n42023_ = ~new_n42021_ & ~new_n42022_;
  assign new_n42024_ = new_n41091_ & ~new_n42023_;
  assign new_n42025_ = ~new_n42019_ & ~new_n42024_;
  assign new_n42026_ = ~new_n42012_ & new_n42025_;
  assign new_n42027_ = new_n40854_ & ~new_n40924_;
  assign new_n42028_ = ~new_n40957_ & new_n41991_;
  assign new_n42029_ = new_n40924_ & new_n42028_;
  assign new_n42030_ = ~new_n40924_ & ~new_n42028_;
  assign new_n42031_ = ~new_n42029_ & ~new_n42030_;
  assign new_n42032_ = ~new_n40854_ & ~new_n42031_;
  assign new_n42033_ = ~new_n42027_ & ~new_n42032_;
  assign new_n42034_ = new_n41037_ & ~new_n42033_;
  assign new_n42035_ = new_n40492_ & ~new_n40610_;
  assign new_n42036_ = ~new_n40643_ & new_n41999_;
  assign new_n42037_ = new_n40610_ & new_n42036_;
  assign new_n42038_ = ~new_n40610_ & ~new_n42036_;
  assign new_n42039_ = ~new_n42037_ & ~new_n42038_;
  assign new_n42040_ = ~new_n40492_ & ~new_n42039_;
  assign new_n42041_ = ~new_n42035_ & ~new_n42040_;
  assign new_n42042_ = new_n41043_ & ~new_n42041_;
  assign new_n42043_ = ~new_n42034_ & ~new_n42042_;
  assign new_n42044_ = new_n42026_ & new_n42043_;
  assign new_n42045_ = new_n41051_ & ~new_n42044_;
  assign ys__n30328 = new_n42011_ | new_n42045_;
  assign ys__n30331 = ys__n2652 & ys__n30330;
  assign new_n42048_ = ys__n174 & ~ys__n196;
  assign new_n42049_ = ys__n2830 & new_n42048_;
  assign new_n42050_ = new_n41443_ & new_n42049_;
  assign new_n42051_ = ys__n174 & ys__n196;
  assign new_n42052_ = ys__n24786 & new_n42051_;
  assign new_n42053_ = ~ys__n2830 & new_n42048_;
  assign new_n42054_ = new_n41443_ & new_n42053_;
  assign new_n42055_ = ~new_n42052_ & ~new_n42054_;
  assign new_n42056_ = ~new_n42050_ & new_n42055_;
  assign new_n42057_ = ~ys__n174 & ys__n196;
  assign new_n42058_ = ~new_n42051_ & ~new_n42057_;
  assign new_n42059_ = ~new_n42053_ & new_n42058_;
  assign new_n42060_ = ~ys__n196 & ys__n2830;
  assign new_n42061_ = ~ys__n174 & new_n42060_;
  assign new_n42062_ = ~ys__n174 & ~ys__n196;
  assign new_n42063_ = ~ys__n2830 & new_n42062_;
  assign new_n42064_ = ~new_n42049_ & ~new_n42063_;
  assign new_n42065_ = ~new_n42061_ & new_n42064_;
  assign new_n42066_ = new_n42059_ & new_n42065_;
  assign ys__n33095 = ~new_n42056_ & ~new_n42066_;
  assign new_n42068_ = ys__n24789 & new_n42051_;
  assign new_n42069_ = new_n41472_ & new_n42053_;
  assign new_n42070_ = ~new_n42068_ & ~new_n42069_;
  assign new_n42071_ = new_n39469_ & new_n42061_;
  assign new_n42072_ = new_n39469_ & new_n42063_;
  assign new_n42073_ = new_n41472_ & new_n42049_;
  assign new_n42074_ = ~new_n42072_ & ~new_n42073_;
  assign new_n42075_ = ~new_n42071_ & new_n42074_;
  assign new_n42076_ = new_n42070_ & new_n42075_;
  assign ys__n33096 = ~new_n42066_ & ~new_n42076_;
  assign new_n42078_ = ~ys__n33095 & ys__n33096;
  assign new_n42079_ = ys__n33095 & ~ys__n33096;
  assign new_n42080_ = ~new_n42078_ & ~new_n42079_;
  assign new_n42081_ = new_n41081_ & new_n42049_;
  assign new_n42082_ = ys__n24747 & new_n42051_;
  assign new_n42083_ = new_n41081_ & new_n42053_;
  assign new_n42084_ = ~new_n42082_ & ~new_n42083_;
  assign new_n42085_ = ~new_n42081_ & new_n42084_;
  assign ys__n33082 = ~new_n42066_ & ~new_n42085_;
  assign new_n42087_ = new_n41054_ & new_n42049_;
  assign new_n42088_ = ys__n24744 & new_n42051_;
  assign new_n42089_ = new_n41054_ & new_n42053_;
  assign new_n42090_ = ~new_n42088_ & ~new_n42089_;
  assign new_n42091_ = ~new_n42087_ & new_n42090_;
  assign ys__n33081 = ~new_n42066_ & ~new_n42091_;
  assign new_n42093_ = ~ys__n33082 & ys__n33081;
  assign new_n42094_ = ys__n33082 & ~ys__n33081;
  assign new_n42095_ = ~new_n42093_ & ~new_n42094_;
  assign new_n42096_ = new_n41107_ & new_n42049_;
  assign new_n42097_ = ys__n24750 & new_n42051_;
  assign new_n42098_ = new_n41107_ & new_n42053_;
  assign new_n42099_ = ~new_n42097_ & ~new_n42098_;
  assign new_n42100_ = ~new_n42096_ & new_n42099_;
  assign ys__n33083 = ~new_n42066_ & ~new_n42100_;
  assign new_n42102_ = ys__n33082 & ~ys__n33083;
  assign new_n42103_ = ~ys__n33082 & ys__n33083;
  assign new_n42104_ = ~new_n42102_ & ~new_n42103_;
  assign new_n42105_ = new_n39469_ & new_n42049_;
  assign new_n42106_ = ys__n24741 & new_n42051_;
  assign new_n42107_ = new_n39469_ & new_n42053_;
  assign new_n42108_ = ~new_n42106_ & ~new_n42107_;
  assign new_n42109_ = ~new_n42105_ & new_n42108_;
  assign ys__n33080 = ~new_n42066_ & ~new_n42109_;
  assign new_n42111_ = ys__n33081 & ys__n33080;
  assign new_n42112_ = ~new_n42104_ & new_n42111_;
  assign new_n42113_ = ~new_n42095_ & new_n42112_;
  assign new_n42114_ = ys__n33082 & ys__n33083;
  assign new_n42115_ = ys__n33082 & ys__n33081;
  assign new_n42116_ = ~new_n42104_ & new_n42115_;
  assign new_n42117_ = ~new_n42114_ & ~new_n42116_;
  assign new_n42118_ = ~new_n42113_ & new_n42117_;
  assign new_n42119_ = new_n41215_ & new_n42049_;
  assign new_n42120_ = ys__n24762 & new_n42051_;
  assign new_n42121_ = new_n41215_ & new_n42053_;
  assign new_n42122_ = ~new_n42120_ & ~new_n42121_;
  assign new_n42123_ = ~new_n42119_ & new_n42122_;
  assign ys__n33087 = ~new_n42066_ & ~new_n42123_;
  assign new_n42125_ = new_n41186_ & new_n42049_;
  assign new_n42126_ = ys__n24759 & new_n42051_;
  assign new_n42127_ = new_n41186_ & new_n42053_;
  assign new_n42128_ = ~new_n42126_ & ~new_n42127_;
  assign new_n42129_ = ~new_n42125_ & new_n42128_;
  assign ys__n33086 = ~new_n42066_ & ~new_n42129_;
  assign new_n42131_ = ~ys__n33087 & ys__n33086;
  assign new_n42132_ = ys__n33087 & ~ys__n33086;
  assign new_n42133_ = ~new_n42131_ & ~new_n42132_;
  assign new_n42134_ = new_n41158_ & new_n42049_;
  assign new_n42135_ = ys__n24756 & new_n42051_;
  assign new_n42136_ = new_n41158_ & new_n42053_;
  assign new_n42137_ = ~new_n42135_ & ~new_n42136_;
  assign new_n42138_ = ~new_n42134_ & new_n42137_;
  assign ys__n33085 = ~new_n42066_ & ~new_n42138_;
  assign new_n42140_ = ~ys__n33086 & ys__n33085;
  assign new_n42141_ = ys__n33086 & ~ys__n33085;
  assign new_n42142_ = ~new_n42140_ & ~new_n42141_;
  assign new_n42143_ = ~new_n42133_ & ~new_n42142_;
  assign new_n42144_ = new_n41133_ & new_n42049_;
  assign new_n42145_ = ys__n24753 & new_n42051_;
  assign new_n42146_ = new_n41133_ & new_n42053_;
  assign new_n42147_ = ~new_n42145_ & ~new_n42146_;
  assign new_n42148_ = ~new_n42144_ & new_n42147_;
  assign ys__n33084 = ~new_n42066_ & ~new_n42148_;
  assign new_n42150_ = ~ys__n33085 & ys__n33084;
  assign new_n42151_ = ys__n33085 & ~ys__n33084;
  assign new_n42152_ = ~new_n42150_ & ~new_n42151_;
  assign new_n42153_ = ys__n33083 & ~ys__n33084;
  assign new_n42154_ = ~ys__n33083 & ys__n33084;
  assign new_n42155_ = ~new_n42153_ & ~new_n42154_;
  assign new_n42156_ = ~new_n42152_ & ~new_n42155_;
  assign new_n42157_ = new_n42143_ & new_n42156_;
  assign new_n42158_ = ~new_n42118_ & new_n42157_;
  assign new_n42159_ = ys__n33085 & ys__n33084;
  assign new_n42160_ = ys__n33083 & ys__n33084;
  assign new_n42161_ = ~new_n42152_ & new_n42160_;
  assign new_n42162_ = ~new_n42159_ & ~new_n42161_;
  assign new_n42163_ = new_n42143_ & ~new_n42162_;
  assign new_n42164_ = ys__n33087 & ys__n33086;
  assign new_n42165_ = ys__n33086 & ys__n33085;
  assign new_n42166_ = ~new_n42133_ & new_n42165_;
  assign new_n42167_ = ~new_n42164_ & ~new_n42166_;
  assign new_n42168_ = ~new_n42163_ & new_n42167_;
  assign new_n42169_ = ~new_n42158_ & new_n42168_;
  assign new_n42170_ = new_n41414_ & new_n42049_;
  assign new_n42171_ = ys__n24783 & new_n42051_;
  assign new_n42172_ = new_n41414_ & new_n42053_;
  assign new_n42173_ = ~new_n42171_ & ~new_n42172_;
  assign new_n42174_ = ~new_n42170_ & new_n42173_;
  assign ys__n33094 = ~new_n42066_ & ~new_n42174_;
  assign new_n42176_ = ~ys__n33095 & ys__n33094;
  assign new_n42177_ = ys__n33095 & ~ys__n33094;
  assign new_n42178_ = ~new_n42176_ & ~new_n42177_;
  assign new_n42179_ = new_n41385_ & new_n42049_;
  assign new_n42180_ = ys__n24780 & new_n42051_;
  assign new_n42181_ = new_n41385_ & new_n42053_;
  assign new_n42182_ = ~new_n42180_ & ~new_n42181_;
  assign new_n42183_ = ~new_n42179_ & new_n42182_;
  assign ys__n33093 = ~new_n42066_ & ~new_n42183_;
  assign new_n42185_ = ~ys__n33094 & ys__n33093;
  assign new_n42186_ = ys__n33094 & ~ys__n33093;
  assign new_n42187_ = ~new_n42185_ & ~new_n42186_;
  assign new_n42188_ = ~new_n42178_ & ~new_n42187_;
  assign new_n42189_ = new_n41356_ & new_n42049_;
  assign new_n42190_ = ys__n24777 & new_n42051_;
  assign new_n42191_ = new_n41356_ & new_n42053_;
  assign new_n42192_ = ~new_n42190_ & ~new_n42191_;
  assign new_n42193_ = ~new_n42189_ & new_n42192_;
  assign ys__n33092 = ~new_n42066_ & ~new_n42193_;
  assign new_n42195_ = ~ys__n33093 & ys__n33092;
  assign new_n42196_ = ys__n33093 & ~ys__n33092;
  assign new_n42197_ = ~new_n42195_ & ~new_n42196_;
  assign new_n42198_ = new_n41327_ & new_n42049_;
  assign new_n42199_ = ys__n24774 & new_n42051_;
  assign new_n42200_ = new_n41327_ & new_n42053_;
  assign new_n42201_ = ~new_n42199_ & ~new_n42200_;
  assign new_n42202_ = ~new_n42198_ & new_n42201_;
  assign ys__n33091 = ~new_n42066_ & ~new_n42202_;
  assign new_n42204_ = ~ys__n33092 & ys__n33091;
  assign new_n42205_ = ys__n33092 & ~ys__n33091;
  assign new_n42206_ = ~new_n42204_ & ~new_n42205_;
  assign new_n42207_ = ~new_n42197_ & ~new_n42206_;
  assign new_n42208_ = new_n42188_ & new_n42207_;
  assign new_n42209_ = new_n41298_ & new_n42049_;
  assign new_n42210_ = ys__n24771 & new_n42051_;
  assign new_n42211_ = new_n41298_ & new_n42053_;
  assign new_n42212_ = ~new_n42210_ & ~new_n42211_;
  assign new_n42213_ = ~new_n42209_ & new_n42212_;
  assign ys__n33090 = ~new_n42066_ & ~new_n42213_;
  assign new_n42215_ = ~ys__n33091 & ys__n33090;
  assign new_n42216_ = ys__n33091 & ~ys__n33090;
  assign new_n42217_ = ~new_n42215_ & ~new_n42216_;
  assign new_n42218_ = new_n41270_ & new_n42049_;
  assign new_n42219_ = ys__n24768 & new_n42051_;
  assign new_n42220_ = new_n41270_ & new_n42053_;
  assign new_n42221_ = ~new_n42219_ & ~new_n42220_;
  assign new_n42222_ = ~new_n42218_ & new_n42221_;
  assign ys__n33089 = ~new_n42066_ & ~new_n42222_;
  assign new_n42224_ = ~ys__n33090 & ys__n33089;
  assign new_n42225_ = ys__n33090 & ~ys__n33089;
  assign new_n42226_ = ~new_n42224_ & ~new_n42225_;
  assign new_n42227_ = ~new_n42217_ & ~new_n42226_;
  assign new_n42228_ = new_n41244_ & new_n42049_;
  assign new_n42229_ = ys__n24765 & new_n42051_;
  assign new_n42230_ = new_n41244_ & new_n42053_;
  assign new_n42231_ = ~new_n42229_ & ~new_n42230_;
  assign new_n42232_ = ~new_n42228_ & new_n42231_;
  assign ys__n33088 = ~new_n42066_ & ~new_n42232_;
  assign new_n42234_ = ~ys__n33089 & ys__n33088;
  assign new_n42235_ = ys__n33089 & ~ys__n33088;
  assign new_n42236_ = ~new_n42234_ & ~new_n42235_;
  assign new_n42237_ = ys__n33087 & ~ys__n33088;
  assign new_n42238_ = ~ys__n33087 & ys__n33088;
  assign new_n42239_ = ~new_n42237_ & ~new_n42238_;
  assign new_n42240_ = ~new_n42236_ & ~new_n42239_;
  assign new_n42241_ = new_n42227_ & new_n42240_;
  assign new_n42242_ = new_n42208_ & new_n42241_;
  assign new_n42243_ = ~new_n42169_ & new_n42242_;
  assign new_n42244_ = ys__n33089 & ys__n33088;
  assign new_n42245_ = ys__n33087 & ys__n33088;
  assign new_n42246_ = ~new_n42236_ & new_n42245_;
  assign new_n42247_ = ~new_n42244_ & ~new_n42246_;
  assign new_n42248_ = new_n42227_ & ~new_n42247_;
  assign new_n42249_ = ys__n33091 & ys__n33090;
  assign new_n42250_ = ys__n33090 & ys__n33089;
  assign new_n42251_ = ~new_n42217_ & new_n42250_;
  assign new_n42252_ = ~new_n42249_ & ~new_n42251_;
  assign new_n42253_ = ~new_n42248_ & new_n42252_;
  assign new_n42254_ = new_n42208_ & ~new_n42253_;
  assign new_n42255_ = ys__n33093 & ys__n33092;
  assign new_n42256_ = ys__n33092 & ys__n33091;
  assign new_n42257_ = ~new_n42197_ & new_n42256_;
  assign new_n42258_ = ~new_n42255_ & ~new_n42257_;
  assign new_n42259_ = new_n42188_ & ~new_n42258_;
  assign new_n42260_ = ys__n33095 & ys__n33094;
  assign new_n42261_ = ys__n33094 & ys__n33093;
  assign new_n42262_ = ~new_n42178_ & new_n42261_;
  assign new_n42263_ = ~new_n42260_ & ~new_n42262_;
  assign new_n42264_ = ~new_n42259_ & new_n42263_;
  assign new_n42265_ = ~new_n42254_ & new_n42264_;
  assign new_n42266_ = ~new_n42243_ & new_n42265_;
  assign new_n42267_ = ~new_n42080_ & new_n42266_;
  assign new_n42268_ = new_n42080_ & ~new_n42266_;
  assign ys__n30616 = new_n42267_ | new_n42268_;
  assign new_n42270_ = ys__n24792 & new_n42051_;
  assign new_n42271_ = new_n41498_ & new_n42053_;
  assign new_n42272_ = ~new_n42270_ & ~new_n42271_;
  assign new_n42273_ = new_n41054_ & new_n42061_;
  assign new_n42274_ = new_n41054_ & new_n42063_;
  assign new_n42275_ = new_n41498_ & new_n42049_;
  assign new_n42276_ = ~new_n42274_ & ~new_n42275_;
  assign new_n42277_ = ~new_n42273_ & new_n42276_;
  assign new_n42278_ = new_n42272_ & new_n42277_;
  assign ys__n33097 = ~new_n42066_ & ~new_n42278_;
  assign new_n42280_ = ~ys__n33096 & ys__n33097;
  assign new_n42281_ = ys__n33096 & ~ys__n33097;
  assign new_n42282_ = ~new_n42280_ & ~new_n42281_;
  assign new_n42283_ = ys__n33095 & ys__n33096;
  assign new_n42284_ = new_n42282_ & new_n42283_;
  assign new_n42285_ = ~new_n42282_ & ~new_n42283_;
  assign new_n42286_ = ~new_n42284_ & ~new_n42285_;
  assign new_n42287_ = new_n42266_ & ~new_n42286_;
  assign new_n42288_ = ~new_n42080_ & new_n42286_;
  assign new_n42289_ = new_n42080_ & ~new_n42286_;
  assign new_n42290_ = ~new_n42288_ & ~new_n42289_;
  assign new_n42291_ = ~new_n42266_ & ~new_n42290_;
  assign ys__n30619 = new_n42287_ | new_n42291_;
  assign new_n42293_ = ys__n24795 & new_n42051_;
  assign new_n42294_ = new_n41530_ & new_n42053_;
  assign new_n42295_ = ~new_n42293_ & ~new_n42294_;
  assign new_n42296_ = new_n41081_ & new_n42061_;
  assign new_n42297_ = new_n41081_ & new_n42063_;
  assign new_n42298_ = new_n41530_ & new_n42049_;
  assign new_n42299_ = ~new_n42297_ & ~new_n42298_;
  assign new_n42300_ = ~new_n42296_ & new_n42299_;
  assign new_n42301_ = new_n42295_ & new_n42300_;
  assign ys__n33098 = ~new_n42066_ & ~new_n42301_;
  assign new_n42303_ = ~ys__n33097 & ys__n33098;
  assign new_n42304_ = ys__n33097 & ~ys__n33098;
  assign new_n42305_ = ~new_n42303_ & ~new_n42304_;
  assign new_n42306_ = ys__n33096 & ys__n33097;
  assign new_n42307_ = ~new_n42282_ & new_n42283_;
  assign new_n42308_ = ~new_n42306_ & ~new_n42307_;
  assign new_n42309_ = new_n42305_ & ~new_n42308_;
  assign new_n42310_ = ~new_n42305_ & new_n42308_;
  assign new_n42311_ = ~new_n42309_ & ~new_n42310_;
  assign new_n42312_ = new_n42266_ & ~new_n42311_;
  assign new_n42313_ = ~new_n42080_ & ~new_n42286_;
  assign new_n42314_ = new_n42311_ & new_n42313_;
  assign new_n42315_ = ~new_n42311_ & ~new_n42313_;
  assign new_n42316_ = ~new_n42314_ & ~new_n42315_;
  assign new_n42317_ = ~new_n42266_ & ~new_n42316_;
  assign ys__n30622 = new_n42312_ | new_n42317_;
  assign new_n42319_ = ys__n24798 & new_n42051_;
  assign new_n42320_ = new_n41565_ & new_n42053_;
  assign new_n42321_ = ~new_n42319_ & ~new_n42320_;
  assign new_n42322_ = new_n41107_ & new_n42061_;
  assign new_n42323_ = new_n41107_ & new_n42063_;
  assign new_n42324_ = new_n41565_ & new_n42049_;
  assign new_n42325_ = ~new_n42323_ & ~new_n42324_;
  assign new_n42326_ = ~new_n42322_ & new_n42325_;
  assign new_n42327_ = new_n42321_ & new_n42326_;
  assign ys__n33099 = ~new_n42066_ & ~new_n42327_;
  assign new_n42329_ = ~ys__n33098 & ys__n33099;
  assign new_n42330_ = ys__n33098 & ~ys__n33099;
  assign new_n42331_ = ~new_n42329_ & ~new_n42330_;
  assign new_n42332_ = ys__n33097 & ys__n33098;
  assign new_n42333_ = ~new_n42305_ & ~new_n42308_;
  assign new_n42334_ = ~new_n42332_ & ~new_n42333_;
  assign new_n42335_ = new_n42331_ & ~new_n42334_;
  assign new_n42336_ = ~new_n42331_ & new_n42334_;
  assign new_n42337_ = ~new_n42335_ & ~new_n42336_;
  assign new_n42338_ = new_n42266_ & ~new_n42337_;
  assign new_n42339_ = ~new_n42311_ & new_n42313_;
  assign new_n42340_ = new_n42337_ & new_n42339_;
  assign new_n42341_ = ~new_n42337_ & ~new_n42339_;
  assign new_n42342_ = ~new_n42340_ & ~new_n42341_;
  assign new_n42343_ = ~new_n42266_ & ~new_n42342_;
  assign ys__n30625 = new_n42338_ | new_n42343_;
  assign new_n42345_ = ys__n24801 & new_n42051_;
  assign new_n42346_ = new_n41600_ & new_n42053_;
  assign new_n42347_ = ~new_n42345_ & ~new_n42346_;
  assign new_n42348_ = new_n41133_ & new_n42061_;
  assign new_n42349_ = new_n41133_ & new_n42063_;
  assign new_n42350_ = new_n41600_ & new_n42049_;
  assign new_n42351_ = ~new_n42349_ & ~new_n42350_;
  assign new_n42352_ = ~new_n42348_ & new_n42351_;
  assign new_n42353_ = new_n42347_ & new_n42352_;
  assign ys__n33100 = ~new_n42066_ & ~new_n42353_;
  assign new_n42355_ = ~ys__n33099 & ys__n33100;
  assign new_n42356_ = ys__n33099 & ~ys__n33100;
  assign new_n42357_ = ~new_n42355_ & ~new_n42356_;
  assign new_n42358_ = ~new_n42305_ & ~new_n42331_;
  assign new_n42359_ = ~new_n42308_ & new_n42358_;
  assign new_n42360_ = ys__n33098 & ys__n33099;
  assign new_n42361_ = ~new_n42331_ & new_n42332_;
  assign new_n42362_ = ~new_n42360_ & ~new_n42361_;
  assign new_n42363_ = ~new_n42359_ & new_n42362_;
  assign new_n42364_ = new_n42357_ & ~new_n42363_;
  assign new_n42365_ = ~new_n42357_ & new_n42363_;
  assign new_n42366_ = ~new_n42364_ & ~new_n42365_;
  assign new_n42367_ = new_n42266_ & ~new_n42366_;
  assign new_n42368_ = ~new_n42337_ & new_n42339_;
  assign new_n42369_ = new_n42366_ & new_n42368_;
  assign new_n42370_ = ~new_n42366_ & ~new_n42368_;
  assign new_n42371_ = ~new_n42369_ & ~new_n42370_;
  assign new_n42372_ = ~new_n42266_ & ~new_n42371_;
  assign ys__n30628 = new_n42367_ | new_n42372_;
  assign new_n42374_ = ys__n24804 & new_n42051_;
  assign new_n42375_ = new_n41635_ & new_n42053_;
  assign new_n42376_ = ~new_n42374_ & ~new_n42375_;
  assign new_n42377_ = new_n41158_ & new_n42061_;
  assign new_n42378_ = new_n41158_ & new_n42063_;
  assign new_n42379_ = new_n41635_ & new_n42049_;
  assign new_n42380_ = ~new_n42378_ & ~new_n42379_;
  assign new_n42381_ = ~new_n42377_ & new_n42380_;
  assign new_n42382_ = new_n42376_ & new_n42381_;
  assign ys__n33101 = ~new_n42066_ & ~new_n42382_;
  assign new_n42384_ = ~ys__n33100 & ys__n33101;
  assign new_n42385_ = ys__n33100 & ~ys__n33101;
  assign new_n42386_ = ~new_n42384_ & ~new_n42385_;
  assign new_n42387_ = ys__n33099 & ys__n33100;
  assign new_n42388_ = ~new_n42357_ & ~new_n42363_;
  assign new_n42389_ = ~new_n42387_ & ~new_n42388_;
  assign new_n42390_ = new_n42386_ & ~new_n42389_;
  assign new_n42391_ = ~new_n42386_ & new_n42389_;
  assign new_n42392_ = ~new_n42390_ & ~new_n42391_;
  assign new_n42393_ = new_n42266_ & ~new_n42392_;
  assign new_n42394_ = ~new_n42366_ & new_n42368_;
  assign new_n42395_ = new_n42392_ & new_n42394_;
  assign new_n42396_ = ~new_n42392_ & ~new_n42394_;
  assign new_n42397_ = ~new_n42395_ & ~new_n42396_;
  assign new_n42398_ = ~new_n42266_ & ~new_n42397_;
  assign ys__n30631 = new_n42393_ | new_n42398_;
  assign new_n42400_ = ys__n24807 & new_n42051_;
  assign new_n42401_ = new_n41672_ & new_n42053_;
  assign new_n42402_ = ~new_n42400_ & ~new_n42401_;
  assign new_n42403_ = new_n41186_ & new_n42061_;
  assign new_n42404_ = new_n41186_ & new_n42063_;
  assign new_n42405_ = new_n41672_ & new_n42049_;
  assign new_n42406_ = ~new_n42404_ & ~new_n42405_;
  assign new_n42407_ = ~new_n42403_ & new_n42406_;
  assign new_n42408_ = new_n42402_ & new_n42407_;
  assign ys__n33102 = ~new_n42066_ & ~new_n42408_;
  assign new_n42410_ = ~ys__n33101 & ys__n33102;
  assign new_n42411_ = ys__n33101 & ~ys__n33102;
  assign new_n42412_ = ~new_n42410_ & ~new_n42411_;
  assign new_n42413_ = ys__n33100 & ys__n33101;
  assign new_n42414_ = ~new_n42386_ & new_n42387_;
  assign new_n42415_ = ~new_n42413_ & ~new_n42414_;
  assign new_n42416_ = ~new_n42357_ & ~new_n42386_;
  assign new_n42417_ = ~new_n42363_ & new_n42416_;
  assign new_n42418_ = new_n42415_ & ~new_n42417_;
  assign new_n42419_ = new_n42412_ & ~new_n42418_;
  assign new_n42420_ = ~new_n42412_ & new_n42418_;
  assign new_n42421_ = ~new_n42419_ & ~new_n42420_;
  assign new_n42422_ = new_n42266_ & ~new_n42421_;
  assign new_n42423_ = ~new_n42366_ & ~new_n42392_;
  assign new_n42424_ = new_n42368_ & new_n42423_;
  assign new_n42425_ = new_n42421_ & new_n42424_;
  assign new_n42426_ = ~new_n42421_ & ~new_n42424_;
  assign new_n42427_ = ~new_n42425_ & ~new_n42426_;
  assign new_n42428_ = ~new_n42266_ & ~new_n42427_;
  assign ys__n30634 = new_n42422_ | new_n42428_;
  assign new_n42430_ = ys__n24810 & new_n42051_;
  assign new_n42431_ = new_n41710_ & new_n42053_;
  assign new_n42432_ = ~new_n42430_ & ~new_n42431_;
  assign new_n42433_ = new_n41215_ & new_n42061_;
  assign new_n42434_ = new_n41215_ & new_n42063_;
  assign new_n42435_ = new_n41710_ & new_n42049_;
  assign new_n42436_ = ~new_n42434_ & ~new_n42435_;
  assign new_n42437_ = ~new_n42433_ & new_n42436_;
  assign new_n42438_ = new_n42432_ & new_n42437_;
  assign ys__n33103 = ~new_n42066_ & ~new_n42438_;
  assign new_n42440_ = ~ys__n33102 & ys__n33103;
  assign new_n42441_ = ys__n33102 & ~ys__n33103;
  assign new_n42442_ = ~new_n42440_ & ~new_n42441_;
  assign new_n42443_ = ys__n33101 & ys__n33102;
  assign new_n42444_ = ~new_n42412_ & ~new_n42418_;
  assign new_n42445_ = ~new_n42443_ & ~new_n42444_;
  assign new_n42446_ = new_n42442_ & ~new_n42445_;
  assign new_n42447_ = ~new_n42442_ & new_n42445_;
  assign new_n42448_ = ~new_n42446_ & ~new_n42447_;
  assign new_n42449_ = new_n42266_ & ~new_n42448_;
  assign new_n42450_ = ~new_n42421_ & new_n42424_;
  assign new_n42451_ = new_n42448_ & new_n42450_;
  assign new_n42452_ = ~new_n42448_ & ~new_n42450_;
  assign new_n42453_ = ~new_n42451_ & ~new_n42452_;
  assign new_n42454_ = ~new_n42266_ & ~new_n42453_;
  assign ys__n30637 = new_n42449_ | new_n42454_;
  assign new_n42456_ = ys__n24813 & new_n42051_;
  assign new_n42457_ = new_n41748_ & new_n42053_;
  assign new_n42458_ = ~new_n42456_ & ~new_n42457_;
  assign new_n42459_ = new_n41244_ & new_n42061_;
  assign new_n42460_ = new_n41244_ & new_n42063_;
  assign new_n42461_ = new_n41748_ & new_n42049_;
  assign new_n42462_ = ~new_n42460_ & ~new_n42461_;
  assign new_n42463_ = ~new_n42459_ & new_n42462_;
  assign new_n42464_ = new_n42458_ & new_n42463_;
  assign ys__n33104 = ~new_n42066_ & ~new_n42464_;
  assign new_n42466_ = ~ys__n33103 & ys__n33104;
  assign new_n42467_ = ys__n33103 & ~ys__n33104;
  assign new_n42468_ = ~new_n42466_ & ~new_n42467_;
  assign new_n42469_ = ~new_n42412_ & ~new_n42442_;
  assign new_n42470_ = new_n42416_ & new_n42469_;
  assign new_n42471_ = ~new_n42363_ & new_n42470_;
  assign new_n42472_ = ~new_n42415_ & new_n42469_;
  assign new_n42473_ = ys__n33102 & ys__n33103;
  assign new_n42474_ = ~new_n42442_ & new_n42443_;
  assign new_n42475_ = ~new_n42473_ & ~new_n42474_;
  assign new_n42476_ = ~new_n42472_ & new_n42475_;
  assign new_n42477_ = ~new_n42471_ & new_n42476_;
  assign new_n42478_ = new_n42468_ & ~new_n42477_;
  assign new_n42479_ = ~new_n42468_ & new_n42477_;
  assign new_n42480_ = ~new_n42478_ & ~new_n42479_;
  assign new_n42481_ = new_n42266_ & ~new_n42480_;
  assign new_n42482_ = new_n42368_ & ~new_n42421_;
  assign new_n42483_ = new_n42423_ & new_n42482_;
  assign new_n42484_ = ~new_n42448_ & new_n42483_;
  assign new_n42485_ = new_n42480_ & new_n42484_;
  assign new_n42486_ = ~new_n42480_ & ~new_n42484_;
  assign new_n42487_ = ~new_n42485_ & ~new_n42486_;
  assign new_n42488_ = ~new_n42266_ & ~new_n42487_;
  assign ys__n30640 = new_n42481_ | new_n42488_;
  assign new_n42490_ = ys__n24816 & new_n42051_;
  assign new_n42491_ = new_n41784_ & new_n42053_;
  assign new_n42492_ = ~new_n42490_ & ~new_n42491_;
  assign new_n42493_ = new_n41270_ & new_n42061_;
  assign new_n42494_ = new_n41270_ & new_n42063_;
  assign new_n42495_ = new_n41784_ & new_n42049_;
  assign new_n42496_ = ~new_n42494_ & ~new_n42495_;
  assign new_n42497_ = ~new_n42493_ & new_n42496_;
  assign new_n42498_ = new_n42492_ & new_n42497_;
  assign ys__n33105 = ~new_n42066_ & ~new_n42498_;
  assign new_n42500_ = ~ys__n33104 & ys__n33105;
  assign new_n42501_ = ys__n33104 & ~ys__n33105;
  assign new_n42502_ = ~new_n42500_ & ~new_n42501_;
  assign new_n42503_ = ys__n33103 & ys__n33104;
  assign new_n42504_ = ~new_n42468_ & ~new_n42477_;
  assign new_n42505_ = ~new_n42503_ & ~new_n42504_;
  assign new_n42506_ = new_n42502_ & ~new_n42505_;
  assign new_n42507_ = ~new_n42502_ & new_n42505_;
  assign new_n42508_ = ~new_n42506_ & ~new_n42507_;
  assign new_n42509_ = new_n42266_ & ~new_n42508_;
  assign new_n42510_ = ~new_n42480_ & new_n42484_;
  assign new_n42511_ = new_n42508_ & new_n42510_;
  assign new_n42512_ = ~new_n42508_ & ~new_n42510_;
  assign new_n42513_ = ~new_n42511_ & ~new_n42512_;
  assign new_n42514_ = ~new_n42266_ & ~new_n42513_;
  assign ys__n30643 = new_n42509_ | new_n42514_;
  assign new_n42516_ = ys__n24819 & new_n42051_;
  assign new_n42517_ = new_n41821_ & new_n42053_;
  assign new_n42518_ = ~new_n42516_ & ~new_n42517_;
  assign new_n42519_ = new_n41298_ & new_n42061_;
  assign new_n42520_ = new_n41298_ & new_n42063_;
  assign new_n42521_ = new_n41821_ & new_n42049_;
  assign new_n42522_ = ~new_n42520_ & ~new_n42521_;
  assign new_n42523_ = ~new_n42519_ & new_n42522_;
  assign new_n42524_ = new_n42518_ & new_n42523_;
  assign ys__n33106 = ~new_n42066_ & ~new_n42524_;
  assign new_n42526_ = ~ys__n33105 & ys__n33106;
  assign new_n42527_ = ys__n33105 & ~ys__n33106;
  assign new_n42528_ = ~new_n42526_ & ~new_n42527_;
  assign new_n42529_ = ys__n33104 & ys__n33105;
  assign new_n42530_ = ~new_n42502_ & new_n42503_;
  assign new_n42531_ = ~new_n42529_ & ~new_n42530_;
  assign new_n42532_ = ~new_n42468_ & ~new_n42502_;
  assign new_n42533_ = ~new_n42477_ & new_n42532_;
  assign new_n42534_ = new_n42531_ & ~new_n42533_;
  assign new_n42535_ = new_n42528_ & ~new_n42534_;
  assign new_n42536_ = ~new_n42528_ & new_n42534_;
  assign new_n42537_ = ~new_n42535_ & ~new_n42536_;
  assign new_n42538_ = new_n42266_ & ~new_n42537_;
  assign new_n42539_ = ~new_n42480_ & ~new_n42508_;
  assign new_n42540_ = new_n42484_ & new_n42539_;
  assign new_n42541_ = new_n42537_ & new_n42540_;
  assign new_n42542_ = ~new_n42537_ & ~new_n42540_;
  assign new_n42543_ = ~new_n42541_ & ~new_n42542_;
  assign new_n42544_ = ~new_n42266_ & ~new_n42543_;
  assign ys__n30646 = new_n42538_ | new_n42544_;
  assign new_n42546_ = ys__n24822 & new_n42051_;
  assign new_n42547_ = new_n41859_ & new_n42053_;
  assign new_n42548_ = ~new_n42546_ & ~new_n42547_;
  assign new_n42549_ = new_n41327_ & new_n42061_;
  assign new_n42550_ = new_n41327_ & new_n42063_;
  assign new_n42551_ = new_n41859_ & new_n42049_;
  assign new_n42552_ = ~new_n42550_ & ~new_n42551_;
  assign new_n42553_ = ~new_n42549_ & new_n42552_;
  assign new_n42554_ = new_n42548_ & new_n42553_;
  assign ys__n33107 = ~new_n42066_ & ~new_n42554_;
  assign new_n42556_ = ~ys__n33106 & ys__n33107;
  assign new_n42557_ = ys__n33106 & ~ys__n33107;
  assign new_n42558_ = ~new_n42556_ & ~new_n42557_;
  assign new_n42559_ = ys__n33105 & ys__n33106;
  assign new_n42560_ = ~new_n42528_ & ~new_n42534_;
  assign new_n42561_ = ~new_n42559_ & ~new_n42560_;
  assign new_n42562_ = new_n42558_ & ~new_n42561_;
  assign new_n42563_ = ~new_n42558_ & new_n42561_;
  assign new_n42564_ = ~new_n42562_ & ~new_n42563_;
  assign new_n42565_ = new_n42266_ & ~new_n42564_;
  assign new_n42566_ = ~new_n42537_ & new_n42540_;
  assign new_n42567_ = new_n42564_ & new_n42566_;
  assign new_n42568_ = ~new_n42564_ & ~new_n42566_;
  assign new_n42569_ = ~new_n42567_ & ~new_n42568_;
  assign new_n42570_ = ~new_n42266_ & ~new_n42569_;
  assign ys__n30649 = new_n42565_ | new_n42570_;
  assign new_n42572_ = ys__n24825 & new_n42051_;
  assign new_n42573_ = new_n41897_ & new_n42053_;
  assign new_n42574_ = ~new_n42572_ & ~new_n42573_;
  assign new_n42575_ = new_n41356_ & new_n42061_;
  assign new_n42576_ = new_n41356_ & new_n42063_;
  assign new_n42577_ = new_n41897_ & new_n42049_;
  assign new_n42578_ = ~new_n42576_ & ~new_n42577_;
  assign new_n42579_ = ~new_n42575_ & new_n42578_;
  assign new_n42580_ = new_n42574_ & new_n42579_;
  assign ys__n33108 = ~new_n42066_ & ~new_n42580_;
  assign new_n42582_ = ~ys__n33107 & ys__n33108;
  assign new_n42583_ = ys__n33107 & ~ys__n33108;
  assign new_n42584_ = ~new_n42582_ & ~new_n42583_;
  assign new_n42585_ = ~new_n42528_ & ~new_n42558_;
  assign new_n42586_ = ~new_n42531_ & new_n42585_;
  assign new_n42587_ = ys__n33106 & ys__n33107;
  assign new_n42588_ = ~new_n42558_ & new_n42559_;
  assign new_n42589_ = ~new_n42587_ & ~new_n42588_;
  assign new_n42590_ = ~new_n42586_ & new_n42589_;
  assign new_n42591_ = new_n42532_ & new_n42585_;
  assign new_n42592_ = ~new_n42477_ & new_n42591_;
  assign new_n42593_ = new_n42590_ & ~new_n42592_;
  assign new_n42594_ = new_n42584_ & ~new_n42593_;
  assign new_n42595_ = ~new_n42584_ & new_n42593_;
  assign new_n42596_ = ~new_n42594_ & ~new_n42595_;
  assign new_n42597_ = new_n42266_ & ~new_n42596_;
  assign new_n42598_ = ~new_n42537_ & new_n42539_;
  assign new_n42599_ = ~new_n42564_ & new_n42598_;
  assign new_n42600_ = new_n42484_ & new_n42599_;
  assign new_n42601_ = new_n42596_ & new_n42600_;
  assign new_n42602_ = ~new_n42596_ & ~new_n42600_;
  assign new_n42603_ = ~new_n42601_ & ~new_n42602_;
  assign new_n42604_ = ~new_n42266_ & ~new_n42603_;
  assign ys__n30652 = new_n42597_ | new_n42604_;
  assign new_n42606_ = ys__n24828 & new_n42051_;
  assign new_n42607_ = new_n41935_ & new_n42053_;
  assign new_n42608_ = ~new_n42606_ & ~new_n42607_;
  assign new_n42609_ = new_n41385_ & new_n42061_;
  assign new_n42610_ = new_n41385_ & new_n42063_;
  assign new_n42611_ = new_n41935_ & new_n42049_;
  assign new_n42612_ = ~new_n42610_ & ~new_n42611_;
  assign new_n42613_ = ~new_n42609_ & new_n42612_;
  assign new_n42614_ = new_n42608_ & new_n42613_;
  assign ys__n33109 = ~new_n42066_ & ~new_n42614_;
  assign new_n42616_ = ~ys__n33108 & ys__n33109;
  assign new_n42617_ = ys__n33108 & ~ys__n33109;
  assign new_n42618_ = ~new_n42616_ & ~new_n42617_;
  assign new_n42619_ = ys__n33107 & ys__n33108;
  assign new_n42620_ = ~new_n42584_ & ~new_n42593_;
  assign new_n42621_ = ~new_n42619_ & ~new_n42620_;
  assign new_n42622_ = new_n42618_ & ~new_n42621_;
  assign new_n42623_ = ~new_n42618_ & new_n42621_;
  assign new_n42624_ = ~new_n42622_ & ~new_n42623_;
  assign new_n42625_ = new_n42266_ & ~new_n42624_;
  assign new_n42626_ = ~new_n42596_ & new_n42600_;
  assign new_n42627_ = new_n42624_ & new_n42626_;
  assign new_n42628_ = ~new_n42624_ & ~new_n42626_;
  assign new_n42629_ = ~new_n42627_ & ~new_n42628_;
  assign new_n42630_ = ~new_n42266_ & ~new_n42629_;
  assign ys__n30655 = new_n42625_ | new_n42630_;
  assign new_n42632_ = ys__n24831 & new_n42051_;
  assign new_n42633_ = new_n41972_ & new_n42053_;
  assign new_n42634_ = ~new_n42632_ & ~new_n42633_;
  assign new_n42635_ = new_n41414_ & new_n42061_;
  assign new_n42636_ = new_n41414_ & new_n42063_;
  assign new_n42637_ = new_n41972_ & new_n42049_;
  assign new_n42638_ = ~new_n42636_ & ~new_n42637_;
  assign new_n42639_ = ~new_n42635_ & new_n42638_;
  assign new_n42640_ = new_n42634_ & new_n42639_;
  assign ys__n33110 = ~new_n42066_ & ~new_n42640_;
  assign new_n42642_ = ~ys__n33109 & ys__n33110;
  assign new_n42643_ = ys__n33109 & ~ys__n33110;
  assign new_n42644_ = ~new_n42642_ & ~new_n42643_;
  assign new_n42645_ = ys__n33108 & ys__n33109;
  assign new_n42646_ = ~new_n42618_ & new_n42619_;
  assign new_n42647_ = ~new_n42645_ & ~new_n42646_;
  assign new_n42648_ = ~new_n42584_ & ~new_n42618_;
  assign new_n42649_ = ~new_n42593_ & new_n42648_;
  assign new_n42650_ = new_n42647_ & ~new_n42649_;
  assign new_n42651_ = new_n42644_ & ~new_n42650_;
  assign new_n42652_ = ~new_n42644_ & new_n42650_;
  assign new_n42653_ = ~new_n42651_ & ~new_n42652_;
  assign new_n42654_ = new_n42266_ & ~new_n42653_;
  assign new_n42655_ = ~new_n42596_ & ~new_n42624_;
  assign new_n42656_ = new_n42600_ & new_n42655_;
  assign new_n42657_ = new_n42653_ & new_n42656_;
  assign new_n42658_ = ~new_n42653_ & ~new_n42656_;
  assign new_n42659_ = ~new_n42657_ & ~new_n42658_;
  assign new_n42660_ = ~new_n42266_ & ~new_n42659_;
  assign ys__n30658 = new_n42654_ | new_n42660_;
  assign new_n42662_ = new_n42010_ & new_n42053_;
  assign new_n42663_ = new_n41443_ & new_n42063_;
  assign new_n42664_ = ~new_n42662_ & ~new_n42663_;
  assign new_n42665_ = new_n41443_ & new_n42061_;
  assign new_n42666_ = ys__n24834 & new_n42051_;
  assign new_n42667_ = new_n42010_ & new_n42049_;
  assign new_n42668_ = ~new_n42666_ & ~new_n42667_;
  assign new_n42669_ = ~new_n42665_ & new_n42668_;
  assign new_n42670_ = new_n42664_ & new_n42669_;
  assign ys__n33111 = ~new_n42066_ & ~new_n42670_;
  assign new_n42672_ = ~ys__n33110 & ys__n33111;
  assign new_n42673_ = ys__n33110 & ~ys__n33111;
  assign new_n42674_ = ~new_n42672_ & ~new_n42673_;
  assign new_n42675_ = ys__n33109 & ys__n33110;
  assign new_n42676_ = ~new_n42644_ & ~new_n42650_;
  assign new_n42677_ = ~new_n42675_ & ~new_n42676_;
  assign new_n42678_ = new_n42674_ & ~new_n42677_;
  assign new_n42679_ = ~new_n42674_ & new_n42677_;
  assign new_n42680_ = ~new_n42678_ & ~new_n42679_;
  assign new_n42681_ = new_n42266_ & ~new_n42680_;
  assign new_n42682_ = ~new_n42653_ & new_n42656_;
  assign new_n42683_ = new_n42680_ & new_n42682_;
  assign new_n42684_ = ~new_n42680_ & ~new_n42682_;
  assign new_n42685_ = ~new_n42683_ & ~new_n42684_;
  assign new_n42686_ = ~new_n42266_ & ~new_n42685_;
  assign ys__n30661 = new_n42681_ | new_n42686_;
  assign new_n42688_ = ys__n39518 & new_n42051_;
  assign new_n42689_ = new_n42664_ & ~new_n42688_;
  assign ys__n30668 = ~new_n42066_ & ~new_n42689_;
  assign new_n42691_ = ~ys__n33111 & ys__n30668;
  assign new_n42692_ = ys__n33111 & ~ys__n30668;
  assign new_n42693_ = ~new_n42691_ & ~new_n42692_;
  assign new_n42694_ = ~new_n42644_ & ~new_n42674_;
  assign new_n42695_ = new_n42648_ & new_n42694_;
  assign new_n42696_ = new_n42591_ & new_n42695_;
  assign new_n42697_ = ~new_n42477_ & new_n42696_;
  assign new_n42698_ = ~new_n42590_ & new_n42695_;
  assign new_n42699_ = ~new_n42647_ & new_n42694_;
  assign new_n42700_ = ys__n33110 & ys__n33111;
  assign new_n42701_ = ~new_n42674_ & new_n42675_;
  assign new_n42702_ = ~new_n42700_ & ~new_n42701_;
  assign new_n42703_ = ~new_n42699_ & new_n42702_;
  assign new_n42704_ = ~new_n42698_ & new_n42703_;
  assign new_n42705_ = ~new_n42697_ & new_n42704_;
  assign new_n42706_ = new_n42693_ & ~new_n42705_;
  assign new_n42707_ = ~new_n42693_ & new_n42705_;
  assign new_n42708_ = ~new_n42706_ & ~new_n42707_;
  assign new_n42709_ = new_n42266_ & ~new_n42708_;
  assign new_n42710_ = new_n42484_ & ~new_n42653_;
  assign new_n42711_ = new_n42599_ & new_n42710_;
  assign new_n42712_ = new_n42655_ & new_n42711_;
  assign new_n42713_ = ~new_n42680_ & new_n42712_;
  assign new_n42714_ = new_n42708_ & new_n42713_;
  assign new_n42715_ = ~new_n42708_ & ~new_n42713_;
  assign new_n42716_ = ~new_n42714_ & ~new_n42715_;
  assign new_n42717_ = ~new_n42266_ & ~new_n42716_;
  assign ys__n30664 = new_n42709_ | new_n42717_;
  assign new_n42719_ = ys__n33111 & ys__n30668;
  assign new_n42720_ = ~new_n42693_ & ~new_n42705_;
  assign new_n42721_ = ~new_n42719_ & ~new_n42720_;
  assign new_n42722_ = new_n42266_ & ~new_n42721_;
  assign new_n42723_ = ~new_n42708_ & new_n42713_;
  assign new_n42724_ = new_n42721_ & new_n42723_;
  assign new_n42725_ = ~new_n42721_ & ~new_n42723_;
  assign new_n42726_ = ~new_n42724_ & ~new_n42725_;
  assign new_n42727_ = ~new_n42266_ & ~new_n42726_;
  assign ys__n30667 = new_n42722_ | new_n42727_;
  assign new_n42729_ = new_n42266_ & ys__n30668;
  assign new_n42730_ = ~new_n42708_ & ~new_n42721_;
  assign new_n42731_ = new_n42713_ & new_n42730_;
  assign new_n42732_ = ~ys__n30668 & new_n42731_;
  assign new_n42733_ = ys__n30668 & ~new_n42731_;
  assign new_n42734_ = ~new_n42732_ & ~new_n42733_;
  assign new_n42735_ = ~new_n42266_ & ~new_n42734_;
  assign ys__n30670 = new_n42729_ | new_n42735_;
  assign new_n42737_ = ~ys__n2535 & ~new_n25368_;
  assign new_n42738_ = ys__n2535 & ~new_n26642_;
  assign ys__n30797 = new_n42737_ | new_n42738_;
  assign new_n42740_ = ~ys__n2535 & ~new_n25446_;
  assign new_n42741_ = ys__n2535 & ~new_n26667_;
  assign ys__n30798 = new_n42740_ | new_n42741_;
  assign new_n42743_ = ~ys__n2535 & ~new_n25518_;
  assign new_n42744_ = ys__n2535 & ~new_n26694_;
  assign ys__n30799 = new_n42743_ | new_n42744_;
  assign new_n42746_ = ~ys__n2535 & ~new_n25593_;
  assign new_n42747_ = ys__n2535 & ~new_n26721_;
  assign ys__n30800 = new_n42746_ | new_n42747_;
  assign new_n42749_ = ~ys__n2535 & ~new_n25670_;
  assign new_n42750_ = ys__n2535 & ~new_n26751_;
  assign ys__n30801 = new_n42749_ | new_n42750_;
  assign new_n42752_ = ~ys__n2535 & ~new_n25745_;
  assign new_n42753_ = ys__n2535 & ~new_n26778_;
  assign ys__n30802 = new_n42752_ | new_n42753_;
  assign new_n42755_ = ~ys__n2535 & ~new_n25825_;
  assign new_n42756_ = ys__n2535 & ~new_n26808_;
  assign ys__n30803 = new_n42755_ | new_n42756_;
  assign new_n42758_ = ~ys__n2535 & ~new_n25901_;
  assign new_n42759_ = ys__n2535 & ~new_n26835_;
  assign ys__n30804 = new_n42758_ | new_n42759_;
  assign new_n42761_ = ~ys__n2535 & ~new_n25983_;
  assign new_n42762_ = ys__n2535 & ~new_n26868_;
  assign ys__n30805 = new_n42761_ | new_n42762_;
  assign new_n42764_ = ~ys__n2535 & ~new_n26058_;
  assign new_n42765_ = ys__n2535 & ~new_n26895_;
  assign ys__n30806 = new_n42764_ | new_n42765_;
  assign new_n42767_ = ~ys__n2535 & ~new_n26138_;
  assign new_n42768_ = ys__n2535 & ~new_n26925_;
  assign ys__n30807 = new_n42767_ | new_n42768_;
  assign new_n42770_ = ~ys__n2535 & ~new_n26214_;
  assign new_n42771_ = ys__n2535 & ~new_n26952_;
  assign ys__n30808 = new_n42770_ | new_n42771_;
  assign new_n42773_ = ~ys__n2535 & ~new_n26298_;
  assign new_n42774_ = ys__n2535 & ~new_n26985_;
  assign ys__n30809 = new_n42773_ | new_n42774_;
  assign new_n42776_ = ~ys__n2535 & ~new_n26374_;
  assign new_n42777_ = ys__n2535 & ~new_n27012_;
  assign ys__n30810 = new_n42776_ | new_n42777_;
  assign new_n42779_ = ~ys__n2535 & ~new_n26454_;
  assign new_n42780_ = ys__n2535 & ~new_n27042_;
  assign ys__n30811 = new_n42779_ | new_n42780_;
  assign new_n42782_ = ~ys__n2535 & ~new_n26528_;
  assign new_n42783_ = ys__n2535 & ~new_n27069_;
  assign ys__n30812 = new_n42782_ | new_n42783_;
  assign new_n42785_ = ~ys__n2535 & ~new_n25394_;
  assign new_n42786_ = ys__n2535 & new_n27095_;
  assign ys__n30813 = new_n42785_ | new_n42786_;
  assign new_n42788_ = ~ys__n152 & ys__n158;
  assign new_n42789_ = ~ys__n150 & ~ys__n156;
  assign new_n42790_ = new_n42788_ & new_n42789_;
  assign new_n42791_ = ys__n148 & new_n42790_;
  assign new_n42792_ = ys__n152 & ys__n158;
  assign new_n42793_ = ys__n148 & new_n42789_;
  assign new_n42794_ = new_n42792_ & new_n42793_;
  assign new_n42795_ = ~new_n42791_ & ~new_n42794_;
  assign new_n42796_ = ~ys__n150 & ys__n156;
  assign new_n42797_ = ~ys__n152 & ~ys__n158;
  assign new_n42798_ = ys__n148 & new_n42797_;
  assign new_n42799_ = new_n42796_ & new_n42798_;
  assign new_n42800_ = ys__n148 & new_n42788_;
  assign new_n42801_ = new_n42796_ & new_n42800_;
  assign new_n42802_ = ~new_n42799_ & ~new_n42801_;
  assign new_n42803_ = new_n42795_ & new_n42802_;
  assign new_n42804_ = ~ys__n30837 & ~new_n42803_;
  assign new_n42805_ = ys__n948 & new_n42804_;
  assign new_n42806_ = new_n13729_ & new_n13739_;
  assign new_n42807_ = ys__n352 & new_n13728_;
  assign new_n42808_ = new_n42806_ & new_n42807_;
  assign new_n42809_ = new_n13734_ & new_n13739_;
  assign new_n42810_ = new_n42807_ & new_n42809_;
  assign new_n42811_ = ~new_n42808_ & ~new_n42810_;
  assign new_n42812_ = new_n13738_ & new_n42811_;
  assign new_n42813_ = new_n13478_ & new_n13739_;
  assign new_n42814_ = new_n13741_ & new_n42813_;
  assign new_n42815_ = ~new_n13742_ & ~new_n42814_;
  assign new_n42816_ = new_n13476_ & new_n42809_;
  assign new_n42817_ = new_n13476_ & new_n13740_;
  assign new_n42818_ = ~new_n42816_ & ~new_n42817_;
  assign new_n42819_ = ys__n352 & new_n13470_;
  assign new_n42820_ = new_n13729_ & new_n42819_;
  assign new_n42821_ = new_n13475_ & new_n42820_;
  assign new_n42822_ = new_n13734_ & new_n42819_;
  assign new_n42823_ = new_n13475_ & new_n42822_;
  assign new_n42824_ = ~new_n42821_ & ~new_n42823_;
  assign new_n42825_ = new_n42818_ & new_n42824_;
  assign new_n42826_ = new_n42815_ & new_n42825_;
  assign new_n42827_ = new_n42812_ & new_n42826_;
  assign new_n42828_ = ys__n30832 & ~new_n42827_;
  assign ys__n30833 = new_n42805_ | new_n42828_;
  assign new_n42830_ = ~ys__n30837 & new_n42801_;
  assign new_n42831_ = ~ys__n4566 & new_n42830_;
  assign new_n42832_ = ~ys__n30832 & new_n42831_;
  assign new_n42833_ = ~new_n13737_ & ~new_n42823_;
  assign new_n42834_ = ~new_n42810_ & new_n42833_;
  assign new_n42835_ = ys__n30832 & ~new_n42834_;
  assign ys__n30835 = new_n42832_ | new_n42835_;
  assign new_n42837_ = ys__n30861 & ~ys__n30863;
  assign new_n42838_ = ys__n30862 & ys__n30863;
  assign ys__n30864 = new_n42837_ | new_n42838_;
  assign new_n42840_ = ys__n30865 & ~new_n15093_;
  assign new_n42841_ = new_n15096_ & new_n42840_;
  assign new_n42842_ = new_n15093_ & ys__n25842;
  assign ys__n30873 = new_n42841_ | new_n42842_;
  assign new_n42844_ = ys__n30867 & ~new_n15093_;
  assign new_n42845_ = new_n15096_ & new_n42844_;
  assign new_n42846_ = new_n15093_ & ys__n25844;
  assign ys__n30874 = new_n42845_ | new_n42846_;
  assign new_n42848_ = ys__n30869 & ~new_n15093_;
  assign new_n42849_ = new_n15096_ & new_n42848_;
  assign new_n42850_ = new_n15093_ & ys__n25846;
  assign ys__n30875 = new_n42849_ | new_n42850_;
  assign new_n42852_ = ys__n30871 & ~new_n15093_;
  assign new_n42853_ = new_n15096_ & new_n42852_;
  assign new_n42854_ = new_n15093_ & ys__n25852;
  assign ys__n30876 = new_n42853_ | new_n42854_;
  assign ys__n30942 = ys__n26425 & ~ys__n30941;
  assign ys__n30943 = ys__n26440 & ~ys__n30941;
  assign ys__n30944 = ys__n26446 & ~ys__n30941;
  assign new_n42859_ = ys__n26449 & ~ys__n30941;
  assign ys__n30945 = ys__n30941 | new_n42859_;
  assign ys__n30946 = ys__n26452 & ~ys__n30941;
  assign ys__n30947 = ys__n26466 & ~ys__n30941;
  assign ys__n30948 = ys__n26469 & ~ys__n30941;
  assign ys__n30949 = ys__n26472 & ~ys__n30941;
  assign new_n42865_ = ys__n26475 & ~ys__n30941;
  assign ys__n30950 = ys__n30941 | new_n42865_;
  assign new_n42867_ = ys__n26478 & ~ys__n30941;
  assign ys__n30951 = ys__n30941 | new_n42867_;
  assign ys__n30952 = ys__n26484 & ~ys__n30941;
  assign ys__n30953 = ys__n26496 & ~ys__n30941;
  assign ys__n30954 = ys__n26499 & ~ys__n30941;
  assign ys__n30955 = ys__n26502 & ~ys__n30941;
  assign ys__n30956 = ys__n26517 & ~ys__n30941;
  assign new_n42874_ = ~ys__n536 & ys__n538;
  assign new_n42875_ = new_n36479_ & new_n42874_;
  assign new_n42876_ = ys__n536 & ys__n538;
  assign new_n42877_ = new_n36477_ & new_n42876_;
  assign new_n42878_ = ~new_n42875_ & ~new_n42877_;
  assign new_n42879_ = new_n36479_ & new_n42876_;
  assign new_n42880_ = ys__n182 & ~ys__n536;
  assign new_n42881_ = ys__n538 & new_n42880_;
  assign new_n42882_ = ys__n182 & ys__n536;
  assign new_n42883_ = ys__n538 & new_n42882_;
  assign new_n42884_ = ~new_n42881_ & ~new_n42883_;
  assign new_n42885_ = ~new_n42879_ & new_n42884_;
  assign new_n42886_ = new_n36477_ & new_n42874_;
  assign new_n42887_ = ys__n538 & ~new_n42886_;
  assign new_n42888_ = new_n42878_ & new_n42887_;
  assign new_n42889_ = new_n42885_ & new_n42888_;
  assign new_n42890_ = ~new_n42878_ & ~new_n42889_;
  assign new_n42891_ = ~ys__n1386 & new_n13763_;
  assign new_n42892_ = new_n42890_ & new_n42891_;
  assign new_n42893_ = ys__n564 & new_n36477_;
  assign new_n42894_ = ys__n564 & ~new_n42893_;
  assign new_n42895_ = ys__n564 & new_n36479_;
  assign new_n42896_ = ys__n564 & ~new_n42895_;
  assign new_n42897_ = ys__n182 & ys__n564;
  assign new_n42898_ = ~new_n42893_ & ~new_n42897_;
  assign new_n42899_ = new_n42896_ & new_n42898_;
  assign new_n42900_ = ~new_n42894_ & ~new_n42899_;
  assign new_n42901_ = ys__n1386 & new_n42900_;
  assign new_n42902_ = ~new_n42892_ & ~new_n42901_;
  assign new_n42903_ = ~ys__n1386 & ~new_n42891_;
  assign ys__n31202 = ~new_n42902_ & ~new_n42903_;
  assign new_n42905_ = new_n42879_ & ~new_n42889_;
  assign new_n42906_ = new_n42891_ & new_n42905_;
  assign new_n42907_ = ~new_n42896_ & ~new_n42899_;
  assign new_n42908_ = ys__n1386 & new_n42907_;
  assign new_n42909_ = ~new_n42906_ & ~new_n42908_;
  assign ys__n31203 = ~new_n42903_ & ~new_n42909_;
  assign new_n42911_ = new_n40707_ & new_n41017_;
  assign new_n42912_ = ~new_n40301_ & ~new_n42911_;
  assign new_n42913_ = new_n40707_ & ~new_n41017_;
  assign new_n42914_ = ~new_n40301_ & ~new_n41042_;
  assign new_n42915_ = ~new_n42911_ & new_n42914_;
  assign new_n42916_ = ~new_n42913_ & new_n42915_;
  assign new_n42917_ = ~new_n42912_ & ~new_n42916_;
  assign new_n42918_ = ~ys__n30553 & ys__n30330;
  assign new_n42919_ = ys__n30553 & ~ys__n30330;
  assign new_n42920_ = ~new_n42918_ & ~new_n42919_;
  assign new_n42921_ = ~new_n42917_ & ~new_n42920_;
  assign new_n42922_ = new_n42917_ & new_n42920_;
  assign new_n42923_ = ~new_n42921_ & ~new_n42922_;
  assign new_n42924_ = ys__n39167 & ~new_n42923_;
  assign new_n42925_ = ys__n562 & ys__n47010;
  assign new_n42926_ = ys__n398 & ~ys__n33614;
  assign new_n42927_ = new_n42925_ & new_n42926_;
  assign new_n42928_ = ys__n2652 & ys__n17803;
  assign new_n42929_ = ys__n398 & ys__n33614;
  assign new_n42930_ = ~new_n42925_ & new_n42929_;
  assign new_n42931_ = ~new_n42928_ & ~new_n42930_;
  assign new_n42932_ = ~new_n42927_ & new_n42931_;
  assign new_n42933_ = ~new_n42924_ & new_n42932_;
  assign new_n42934_ = new_n13353_ & ~new_n42933_;
  assign new_n42935_ = ys__n30820 & ~new_n24611_;
  assign new_n42936_ = ys__n30819 & ~new_n24611_;
  assign new_n42937_ = ~new_n42935_ & ~new_n42936_;
  assign new_n42938_ = ys__n314 & new_n42937_;
  assign new_n42939_ = ~new_n25394_ & ~new_n42937_;
  assign new_n42940_ = ~new_n42938_ & ~new_n42939_;
  assign new_n42941_ = ~new_n13350_ & ~new_n42940_;
  assign new_n42942_ = ys__n314 & new_n13350_;
  assign new_n42943_ = ~new_n42941_ & ~new_n42942_;
  assign new_n42944_ = new_n13352_ & ~new_n42943_;
  assign new_n42945_ = ~new_n42934_ & ~new_n42944_;
  assign ys__n31207 = ys__n888 & ~new_n42945_;
  assign new_n42947_ = ~new_n42914_ & ~new_n42916_;
  assign new_n42948_ = ~new_n42920_ & ~new_n42947_;
  assign new_n42949_ = new_n42920_ & new_n42947_;
  assign new_n42950_ = ~new_n42948_ & ~new_n42949_;
  assign new_n42951_ = ys__n39167 & ~new_n42950_;
  assign new_n42952_ = ys__n562 & ys__n47011;
  assign new_n42953_ = new_n42925_ & ~new_n42952_;
  assign new_n42954_ = ~new_n42925_ & new_n42952_;
  assign new_n42955_ = ~new_n42953_ & ~new_n42954_;
  assign new_n42956_ = new_n42929_ & ~new_n42955_;
  assign new_n42957_ = ys__n2652 & ys__n17804;
  assign new_n42958_ = new_n42926_ & new_n42952_;
  assign new_n42959_ = ~new_n42957_ & ~new_n42958_;
  assign new_n42960_ = ~new_n42956_ & new_n42959_;
  assign new_n42961_ = ~new_n42951_ & new_n42960_;
  assign new_n42962_ = new_n13353_ & ~new_n42961_;
  assign new_n42963_ = ys__n170 & new_n42937_;
  assign new_n42964_ = ~new_n25463_ & ~new_n42937_;
  assign new_n42965_ = ~new_n42963_ & ~new_n42964_;
  assign new_n42966_ = ~new_n13350_ & ~new_n42965_;
  assign new_n42967_ = ys__n170 & new_n13350_;
  assign new_n42968_ = ~new_n42966_ & ~new_n42967_;
  assign new_n42969_ = new_n13352_ & ~new_n42968_;
  assign new_n42970_ = ~new_n42962_ & ~new_n42969_;
  assign ys__n31208 = ys__n888 & ~new_n42970_;
  assign new_n42972_ = ys__n562 & ys__n47012;
  assign new_n42973_ = new_n42925_ & new_n42952_;
  assign new_n42974_ = ~new_n42972_ & new_n42973_;
  assign new_n42975_ = new_n42972_ & ~new_n42973_;
  assign new_n42976_ = ~new_n42974_ & ~new_n42975_;
  assign new_n42977_ = new_n42929_ & ~new_n42976_;
  assign new_n42978_ = new_n42926_ & new_n42972_;
  assign new_n42979_ = ys__n2652 & ys__n17806;
  assign new_n42980_ = ys__n39167 & new_n42925_;
  assign new_n42981_ = ~new_n42979_ & ~new_n42980_;
  assign new_n42982_ = ~new_n42978_ & new_n42981_;
  assign new_n42983_ = ~new_n42977_ & new_n42982_;
  assign new_n42984_ = new_n13353_ & ~new_n42983_;
  assign new_n42985_ = ys__n380 & new_n42937_;
  assign new_n42986_ = ~new_n25535_ & ~new_n42937_;
  assign new_n42987_ = ~new_n42985_ & ~new_n42986_;
  assign new_n42988_ = ~new_n13350_ & ~new_n42987_;
  assign new_n42989_ = ys__n380 & new_n13350_;
  assign new_n42990_ = ~new_n42988_ & ~new_n42989_;
  assign new_n42991_ = new_n13352_ & ~new_n42990_;
  assign new_n42992_ = ~new_n42984_ & ~new_n42991_;
  assign ys__n31209 = ys__n888 & ~new_n42992_;
  assign new_n42994_ = ys__n562 & ys__n47013;
  assign new_n42995_ = new_n42972_ & new_n42973_;
  assign new_n42996_ = ~new_n42994_ & new_n42995_;
  assign new_n42997_ = new_n42994_ & ~new_n42995_;
  assign new_n42998_ = ~new_n42996_ & ~new_n42997_;
  assign new_n42999_ = new_n42929_ & ~new_n42998_;
  assign new_n43000_ = new_n42926_ & new_n42994_;
  assign new_n43001_ = ys__n2652 & ys__n17807;
  assign new_n43002_ = ys__n39167 & new_n42952_;
  assign new_n43003_ = ~new_n43001_ & ~new_n43002_;
  assign new_n43004_ = ~new_n43000_ & new_n43003_;
  assign new_n43005_ = ~new_n42999_ & new_n43004_;
  assign new_n43006_ = new_n13353_ & ~new_n43005_;
  assign new_n43007_ = ys__n378 & new_n42937_;
  assign new_n43008_ = ~new_n25610_ & ~new_n42937_;
  assign new_n43009_ = ~new_n43007_ & ~new_n43008_;
  assign new_n43010_ = ~new_n13350_ & ~new_n43009_;
  assign new_n43011_ = ys__n378 & new_n13350_;
  assign new_n43012_ = ~new_n43010_ & ~new_n43011_;
  assign new_n43013_ = new_n13352_ & ~new_n43012_;
  assign new_n43014_ = ~new_n43006_ & ~new_n43013_;
  assign ys__n31210 = ys__n888 & ~new_n43014_;
  assign new_n43016_ = ys__n562 & ys__n47014;
  assign new_n43017_ = new_n42972_ & new_n42994_;
  assign new_n43018_ = new_n42973_ & new_n43017_;
  assign new_n43019_ = ~new_n43016_ & new_n43018_;
  assign new_n43020_ = new_n43016_ & ~new_n43018_;
  assign new_n43021_ = ~new_n43019_ & ~new_n43020_;
  assign new_n43022_ = new_n42929_ & ~new_n43021_;
  assign new_n43023_ = new_n42926_ & new_n43016_;
  assign new_n43024_ = ys__n2652 & ys__n17809;
  assign new_n43025_ = ys__n39167 & new_n42972_;
  assign new_n43026_ = ~new_n43024_ & ~new_n43025_;
  assign new_n43027_ = ~new_n43023_ & new_n43026_;
  assign new_n43028_ = ~new_n43022_ & new_n43027_;
  assign new_n43029_ = new_n13353_ & ~new_n43028_;
  assign new_n43030_ = ys__n382 & new_n42937_;
  assign new_n43031_ = ~new_n25687_ & ~new_n42937_;
  assign new_n43032_ = ~new_n43030_ & ~new_n43031_;
  assign new_n43033_ = ~new_n13350_ & ~new_n43032_;
  assign new_n43034_ = ys__n382 & new_n13350_;
  assign new_n43035_ = ~new_n43033_ & ~new_n43034_;
  assign new_n43036_ = new_n13352_ & ~new_n43035_;
  assign new_n43037_ = ~new_n43029_ & ~new_n43036_;
  assign ys__n31211 = ys__n888 & ~new_n43037_;
  assign new_n43039_ = ys__n562 & ys__n47015;
  assign new_n43040_ = new_n43016_ & new_n43018_;
  assign new_n43041_ = ~new_n43039_ & new_n43040_;
  assign new_n43042_ = new_n43039_ & ~new_n43040_;
  assign new_n43043_ = ~new_n43041_ & ~new_n43042_;
  assign new_n43044_ = new_n42929_ & ~new_n43043_;
  assign new_n43045_ = new_n42926_ & new_n43039_;
  assign new_n43046_ = ys__n2652 & ys__n17810;
  assign new_n43047_ = ys__n39167 & new_n42994_;
  assign new_n43048_ = ~new_n43046_ & ~new_n43047_;
  assign new_n43049_ = ~new_n43045_ & new_n43048_;
  assign new_n43050_ = ~new_n43044_ & new_n43049_;
  assign new_n43051_ = new_n13353_ & ~new_n43050_;
  assign new_n43052_ = ys__n374 & new_n42937_;
  assign new_n43053_ = ~new_n25763_ & ~new_n42937_;
  assign new_n43054_ = ~new_n43052_ & ~new_n43053_;
  assign new_n43055_ = ~new_n13350_ & ~new_n43054_;
  assign new_n43056_ = ys__n374 & new_n13350_;
  assign new_n43057_ = ~new_n43055_ & ~new_n43056_;
  assign new_n43058_ = new_n13352_ & ~new_n43057_;
  assign new_n43059_ = ~new_n43051_ & ~new_n43058_;
  assign ys__n31212 = ys__n888 & ~new_n43059_;
  assign new_n43061_ = ys__n562 & ys__n47016;
  assign new_n43062_ = new_n43016_ & new_n43039_;
  assign new_n43063_ = new_n43018_ & new_n43062_;
  assign new_n43064_ = ~new_n43061_ & new_n43063_;
  assign new_n43065_ = new_n43061_ & ~new_n43063_;
  assign new_n43066_ = ~new_n43064_ & ~new_n43065_;
  assign new_n43067_ = new_n42929_ & ~new_n43066_;
  assign new_n43068_ = new_n42926_ & new_n43061_;
  assign new_n43069_ = ys__n2652 & ys__n17812;
  assign new_n43070_ = ys__n39167 & new_n43016_;
  assign new_n43071_ = ~new_n43069_ & ~new_n43070_;
  assign new_n43072_ = ~new_n43068_ & new_n43071_;
  assign new_n43073_ = ~new_n43067_ & new_n43072_;
  assign new_n43074_ = new_n13353_ & ~new_n43073_;
  assign new_n43075_ = ys__n376 & new_n42937_;
  assign new_n43076_ = ~new_n25843_ & ~new_n42937_;
  assign new_n43077_ = ~new_n43075_ & ~new_n43076_;
  assign new_n43078_ = ~new_n13350_ & ~new_n43077_;
  assign new_n43079_ = ys__n376 & new_n13350_;
  assign new_n43080_ = ~new_n43078_ & ~new_n43079_;
  assign new_n43081_ = new_n13352_ & ~new_n43080_;
  assign new_n43082_ = ~new_n43074_ & ~new_n43081_;
  assign ys__n31213 = ys__n888 & ~new_n43082_;
  assign new_n43084_ = ys__n562 & ys__n47017;
  assign new_n43085_ = new_n43061_ & new_n43063_;
  assign new_n43086_ = ~new_n43084_ & new_n43085_;
  assign new_n43087_ = new_n43084_ & ~new_n43085_;
  assign new_n43088_ = ~new_n43086_ & ~new_n43087_;
  assign new_n43089_ = new_n42929_ & ~new_n43088_;
  assign new_n43090_ = new_n42926_ & new_n43084_;
  assign new_n43091_ = ys__n2652 & ys__n17813;
  assign new_n43092_ = ys__n39167 & new_n43039_;
  assign new_n43093_ = ~new_n43091_ & ~new_n43092_;
  assign new_n43094_ = ~new_n43090_ & new_n43093_;
  assign new_n43095_ = ~new_n43089_ & new_n43094_;
  assign new_n43096_ = new_n13353_ & ~new_n43095_;
  assign new_n43097_ = ys__n372 & new_n42937_;
  assign new_n43098_ = ~new_n25919_ & ~new_n42937_;
  assign new_n43099_ = ~new_n43097_ & ~new_n43098_;
  assign new_n43100_ = ~new_n13350_ & ~new_n43099_;
  assign new_n43101_ = ys__n372 & new_n13350_;
  assign new_n43102_ = ~new_n43100_ & ~new_n43101_;
  assign new_n43103_ = new_n13352_ & ~new_n43102_;
  assign new_n43104_ = ~new_n43096_ & ~new_n43103_;
  assign ys__n31214 = ys__n888 & ~new_n43104_;
  assign new_n43106_ = ys__n562 & ys__n47018;
  assign new_n43107_ = new_n43061_ & new_n43084_;
  assign new_n43108_ = new_n43062_ & new_n43107_;
  assign new_n43109_ = new_n43018_ & new_n43108_;
  assign new_n43110_ = ~new_n43106_ & new_n43109_;
  assign new_n43111_ = new_n43106_ & ~new_n43109_;
  assign new_n43112_ = ~new_n43110_ & ~new_n43111_;
  assign new_n43113_ = new_n42929_ & ~new_n43112_;
  assign new_n43114_ = new_n42926_ & new_n43106_;
  assign new_n43115_ = ys__n2652 & ys__n17815;
  assign new_n43116_ = ys__n39167 & new_n43061_;
  assign new_n43117_ = ~new_n43115_ & ~new_n43116_;
  assign new_n43118_ = ~new_n43114_ & new_n43117_;
  assign new_n43119_ = ~new_n43113_ & new_n43118_;
  assign new_n43120_ = new_n13353_ & ~new_n43119_;
  assign new_n43121_ = ys__n384 & new_n42937_;
  assign new_n43122_ = ~new_n26000_ & ~new_n42937_;
  assign new_n43123_ = ~new_n43121_ & ~new_n43122_;
  assign new_n43124_ = ~new_n13350_ & ~new_n43123_;
  assign new_n43125_ = ys__n384 & new_n13350_;
  assign new_n43126_ = ~new_n43124_ & ~new_n43125_;
  assign new_n43127_ = new_n13352_ & ~new_n43126_;
  assign new_n43128_ = ~new_n43120_ & ~new_n43127_;
  assign ys__n31215 = ys__n888 & ~new_n43128_;
  assign new_n43130_ = ys__n562 & ys__n47019;
  assign new_n43131_ = new_n43106_ & new_n43109_;
  assign new_n43132_ = ~new_n43130_ & new_n43131_;
  assign new_n43133_ = new_n43130_ & ~new_n43131_;
  assign new_n43134_ = ~new_n43132_ & ~new_n43133_;
  assign new_n43135_ = new_n42929_ & ~new_n43134_;
  assign new_n43136_ = new_n42926_ & new_n43130_;
  assign new_n43137_ = ys__n2652 & ys__n17816;
  assign new_n43138_ = ys__n39167 & new_n43084_;
  assign new_n43139_ = ~new_n43137_ & ~new_n43138_;
  assign new_n43140_ = ~new_n43136_ & new_n43139_;
  assign new_n43141_ = ~new_n43135_ & new_n43140_;
  assign new_n43142_ = new_n13353_ & ~new_n43141_;
  assign new_n43143_ = ys__n366 & new_n42937_;
  assign new_n43144_ = ~new_n26076_ & ~new_n42937_;
  assign new_n43145_ = ~new_n43143_ & ~new_n43144_;
  assign new_n43146_ = ~new_n13350_ & ~new_n43145_;
  assign new_n43147_ = ys__n366 & new_n13350_;
  assign new_n43148_ = ~new_n43146_ & ~new_n43147_;
  assign new_n43149_ = new_n13352_ & ~new_n43148_;
  assign new_n43150_ = ~new_n43142_ & ~new_n43149_;
  assign ys__n31216 = ys__n888 & ~new_n43150_;
  assign new_n43152_ = ys__n562 & ys__n47020;
  assign new_n43153_ = new_n43106_ & new_n43130_;
  assign new_n43154_ = new_n43109_ & new_n43153_;
  assign new_n43155_ = ~new_n43152_ & new_n43154_;
  assign new_n43156_ = new_n43152_ & ~new_n43154_;
  assign new_n43157_ = ~new_n43155_ & ~new_n43156_;
  assign new_n43158_ = new_n42929_ & ~new_n43157_;
  assign new_n43159_ = new_n42926_ & new_n43152_;
  assign new_n43160_ = ys__n2652 & ys__n17818;
  assign new_n43161_ = ys__n39167 & new_n43106_;
  assign new_n43162_ = ~new_n43160_ & ~new_n43161_;
  assign new_n43163_ = ~new_n43159_ & new_n43162_;
  assign new_n43164_ = ~new_n43158_ & new_n43163_;
  assign new_n43165_ = new_n13353_ & ~new_n43164_;
  assign new_n43166_ = ys__n368 & new_n42937_;
  assign new_n43167_ = ~new_n26156_ & ~new_n42937_;
  assign new_n43168_ = ~new_n43166_ & ~new_n43167_;
  assign new_n43169_ = ~new_n13350_ & ~new_n43168_;
  assign new_n43170_ = ys__n368 & new_n13350_;
  assign new_n43171_ = ~new_n43169_ & ~new_n43170_;
  assign new_n43172_ = new_n13352_ & ~new_n43171_;
  assign new_n43173_ = ~new_n43165_ & ~new_n43172_;
  assign ys__n31217 = ys__n888 & ~new_n43173_;
  assign new_n43175_ = ys__n562 & ys__n47021;
  assign new_n43176_ = new_n43152_ & new_n43154_;
  assign new_n43177_ = ~new_n43175_ & new_n43176_;
  assign new_n43178_ = new_n43175_ & ~new_n43176_;
  assign new_n43179_ = ~new_n43177_ & ~new_n43178_;
  assign new_n43180_ = new_n42929_ & ~new_n43179_;
  assign new_n43181_ = new_n42926_ & new_n43175_;
  assign new_n43182_ = ys__n2652 & ys__n17819;
  assign new_n43183_ = ys__n39167 & new_n43130_;
  assign new_n43184_ = ~new_n43182_ & ~new_n43183_;
  assign new_n43185_ = ~new_n43181_ & new_n43184_;
  assign new_n43186_ = ~new_n43180_ & new_n43185_;
  assign new_n43187_ = new_n13353_ & ~new_n43186_;
  assign new_n43188_ = ys__n364 & new_n42937_;
  assign new_n43189_ = ~new_n26232_ & ~new_n42937_;
  assign new_n43190_ = ~new_n43188_ & ~new_n43189_;
  assign new_n43191_ = ~new_n13350_ & ~new_n43190_;
  assign new_n43192_ = ys__n364 & new_n13350_;
  assign new_n43193_ = ~new_n43191_ & ~new_n43192_;
  assign new_n43194_ = new_n13352_ & ~new_n43193_;
  assign new_n43195_ = ~new_n43187_ & ~new_n43194_;
  assign ys__n31218 = ys__n888 & ~new_n43195_;
  assign new_n43197_ = ys__n562 & ys__n47022;
  assign new_n43198_ = new_n43152_ & new_n43175_;
  assign new_n43199_ = new_n43153_ & new_n43198_;
  assign new_n43200_ = new_n43109_ & new_n43199_;
  assign new_n43201_ = ~new_n43197_ & new_n43200_;
  assign new_n43202_ = new_n43197_ & ~new_n43200_;
  assign new_n43203_ = ~new_n43201_ & ~new_n43202_;
  assign new_n43204_ = new_n42929_ & ~new_n43203_;
  assign new_n43205_ = new_n42926_ & new_n43197_;
  assign new_n43206_ = ys__n2652 & ys__n17821;
  assign new_n43207_ = ys__n39167 & new_n43152_;
  assign new_n43208_ = ~new_n43206_ & ~new_n43207_;
  assign new_n43209_ = ~new_n43205_ & new_n43208_;
  assign new_n43210_ = ~new_n43204_ & new_n43209_;
  assign new_n43211_ = new_n13353_ & ~new_n43210_;
  assign new_n43212_ = ys__n370 & new_n42937_;
  assign new_n43213_ = ~new_n26316_ & ~new_n42937_;
  assign new_n43214_ = ~new_n43212_ & ~new_n43213_;
  assign new_n43215_ = ~new_n13350_ & ~new_n43214_;
  assign new_n43216_ = ys__n370 & new_n13350_;
  assign new_n43217_ = ~new_n43215_ & ~new_n43216_;
  assign new_n43218_ = new_n13352_ & ~new_n43217_;
  assign new_n43219_ = ~new_n43211_ & ~new_n43218_;
  assign ys__n31219 = ys__n888 & ~new_n43219_;
  assign new_n43221_ = ys__n562 & ys__n47023;
  assign new_n43222_ = new_n43197_ & new_n43200_;
  assign new_n43223_ = ~new_n43221_ & new_n43222_;
  assign new_n43224_ = new_n43221_ & ~new_n43222_;
  assign new_n43225_ = ~new_n43223_ & ~new_n43224_;
  assign new_n43226_ = new_n42929_ & ~new_n43225_;
  assign new_n43227_ = new_n42926_ & new_n43221_;
  assign new_n43228_ = ys__n2652 & ys__n17822;
  assign new_n43229_ = ys__n39167 & new_n43175_;
  assign new_n43230_ = ~new_n43228_ & ~new_n43229_;
  assign new_n43231_ = ~new_n43227_ & new_n43230_;
  assign new_n43232_ = ~new_n43226_ & new_n43231_;
  assign new_n43233_ = new_n13353_ & ~new_n43232_;
  assign new_n43234_ = ys__n360 & new_n42937_;
  assign new_n43235_ = ~new_n26392_ & ~new_n42937_;
  assign new_n43236_ = ~new_n43234_ & ~new_n43235_;
  assign new_n43237_ = ~new_n13350_ & ~new_n43236_;
  assign new_n43238_ = ys__n360 & new_n13350_;
  assign new_n43239_ = ~new_n43237_ & ~new_n43238_;
  assign new_n43240_ = new_n13352_ & ~new_n43239_;
  assign new_n43241_ = ~new_n43233_ & ~new_n43240_;
  assign ys__n31220 = ys__n888 & ~new_n43241_;
  assign new_n43243_ = ys__n562 & ys__n47024;
  assign new_n43244_ = new_n43197_ & new_n43221_;
  assign new_n43245_ = new_n43200_ & new_n43244_;
  assign new_n43246_ = ~new_n43243_ & new_n43245_;
  assign new_n43247_ = new_n43243_ & ~new_n43245_;
  assign new_n43248_ = ~new_n43246_ & ~new_n43247_;
  assign new_n43249_ = new_n42929_ & ~new_n43248_;
  assign new_n43250_ = new_n42926_ & new_n43243_;
  assign new_n43251_ = ys__n2652 & ys__n17824;
  assign new_n43252_ = ys__n39167 & new_n43197_;
  assign new_n43253_ = ~new_n43251_ & ~new_n43252_;
  assign new_n43254_ = ~new_n43250_ & new_n43253_;
  assign new_n43255_ = ~new_n43249_ & new_n43254_;
  assign new_n43256_ = new_n13353_ & ~new_n43255_;
  assign new_n43257_ = ys__n362 & new_n42937_;
  assign new_n43258_ = ~new_n26472_ & ~new_n42937_;
  assign new_n43259_ = ~new_n43257_ & ~new_n43258_;
  assign new_n43260_ = ~new_n13350_ & ~new_n43259_;
  assign new_n43261_ = ys__n362 & new_n13350_;
  assign new_n43262_ = ~new_n43260_ & ~new_n43261_;
  assign new_n43263_ = new_n13352_ & ~new_n43262_;
  assign new_n43264_ = ~new_n43256_ & ~new_n43263_;
  assign ys__n31221 = ys__n888 & ~new_n43264_;
  assign new_n43266_ = ys__n562 & ys__n47025;
  assign new_n43267_ = new_n43243_ & new_n43245_;
  assign new_n43268_ = ~new_n43266_ & new_n43267_;
  assign new_n43269_ = new_n43266_ & ~new_n43267_;
  assign new_n43270_ = ~new_n43268_ & ~new_n43269_;
  assign new_n43271_ = new_n42929_ & ~new_n43270_;
  assign new_n43272_ = new_n42926_ & new_n43266_;
  assign new_n43273_ = ys__n2652 & ys__n17825;
  assign new_n43274_ = ys__n39167 & new_n43221_;
  assign new_n43275_ = ~new_n43273_ & ~new_n43274_;
  assign new_n43276_ = ~new_n43272_ & new_n43275_;
  assign new_n43277_ = ~new_n43271_ & new_n43276_;
  assign new_n43278_ = new_n13353_ & ~new_n43277_;
  assign new_n43279_ = ys__n358 & new_n42937_;
  assign new_n43280_ = ~new_n26546_ & ~new_n42937_;
  assign new_n43281_ = ~new_n43279_ & ~new_n43280_;
  assign new_n43282_ = ~new_n13350_ & ~new_n43281_;
  assign new_n43283_ = ys__n358 & new_n13350_;
  assign new_n43284_ = ~new_n43282_ & ~new_n43283_;
  assign new_n43285_ = new_n13352_ & ~new_n43284_;
  assign new_n43286_ = ~new_n43278_ & ~new_n43285_;
  assign ys__n31222 = ys__n888 & ~new_n43286_;
  assign new_n43288_ = ys__n562 & ys__n47026;
  assign new_n43289_ = new_n43243_ & new_n43266_;
  assign new_n43290_ = new_n43244_ & new_n43289_;
  assign new_n43291_ = new_n43199_ & new_n43290_;
  assign new_n43292_ = new_n43109_ & new_n43291_;
  assign new_n43293_ = ~new_n43288_ & new_n43292_;
  assign new_n43294_ = new_n43288_ & ~new_n43292_;
  assign new_n43295_ = ~new_n43293_ & ~new_n43294_;
  assign new_n43296_ = new_n42929_ & ~new_n43295_;
  assign new_n43297_ = new_n42926_ & new_n43288_;
  assign new_n43298_ = ys__n2652 & ys__n17827;
  assign new_n43299_ = ys__n39167 & new_n43243_;
  assign new_n43300_ = ~new_n43298_ & ~new_n43299_;
  assign new_n43301_ = ~new_n43297_ & new_n43300_;
  assign new_n43302_ = ~new_n43296_ & new_n43301_;
  assign new_n43303_ = new_n13353_ & ~new_n43302_;
  assign new_n43304_ = ~new_n25368_ & new_n42937_;
  assign new_n43305_ = ~new_n25361_ & ~new_n42937_;
  assign new_n43306_ = ~new_n43304_ & ~new_n43305_;
  assign new_n43307_ = ~new_n13350_ & ~new_n43306_;
  assign new_n43308_ = new_n13350_ & ~new_n25368_;
  assign new_n43309_ = ~new_n43307_ & ~new_n43308_;
  assign new_n43310_ = new_n13352_ & ~new_n43309_;
  assign new_n43311_ = ~new_n43303_ & ~new_n43310_;
  assign ys__n31223 = ys__n888 & ~new_n43311_;
  assign new_n43313_ = ys__n562 & ys__n47027;
  assign new_n43314_ = new_n43288_ & new_n43292_;
  assign new_n43315_ = ~new_n43313_ & new_n43314_;
  assign new_n43316_ = new_n43313_ & ~new_n43314_;
  assign new_n43317_ = ~new_n43315_ & ~new_n43316_;
  assign new_n43318_ = new_n42929_ & ~new_n43317_;
  assign new_n43319_ = new_n42926_ & new_n43313_;
  assign new_n43320_ = ys__n2652 & ys__n17828;
  assign new_n43321_ = ys__n39167 & new_n43266_;
  assign new_n43322_ = ~new_n43320_ & ~new_n43321_;
  assign new_n43323_ = ~new_n43319_ & new_n43322_;
  assign new_n43324_ = ~new_n43318_ & new_n43323_;
  assign new_n43325_ = new_n13353_ & ~new_n43324_;
  assign new_n43326_ = ~new_n25446_ & new_n42937_;
  assign new_n43327_ = ~new_n25440_ & ~new_n42937_;
  assign new_n43328_ = ~new_n43326_ & ~new_n43327_;
  assign new_n43329_ = ~new_n13350_ & ~new_n43328_;
  assign new_n43330_ = new_n13350_ & ~new_n25446_;
  assign new_n43331_ = ~new_n43329_ & ~new_n43330_;
  assign new_n43332_ = new_n13352_ & ~new_n43331_;
  assign new_n43333_ = ~new_n43325_ & ~new_n43332_;
  assign ys__n31224 = ys__n888 & ~new_n43333_;
  assign new_n43335_ = ys__n562 & ys__n47028;
  assign new_n43336_ = new_n43288_ & new_n43313_;
  assign new_n43337_ = new_n43292_ & new_n43336_;
  assign new_n43338_ = ~new_n43335_ & new_n43337_;
  assign new_n43339_ = new_n43335_ & ~new_n43337_;
  assign new_n43340_ = ~new_n43338_ & ~new_n43339_;
  assign new_n43341_ = new_n42929_ & ~new_n43340_;
  assign new_n43342_ = new_n42926_ & new_n43335_;
  assign new_n43343_ = ys__n2652 & ys__n17830;
  assign new_n43344_ = ys__n39167 & new_n43288_;
  assign new_n43345_ = ~new_n43343_ & ~new_n43344_;
  assign new_n43346_ = ~new_n43342_ & new_n43345_;
  assign new_n43347_ = ~new_n43341_ & new_n43346_;
  assign new_n43348_ = new_n13353_ & ~new_n43347_;
  assign new_n43349_ = ~new_n25518_ & new_n42937_;
  assign new_n43350_ = ~new_n25512_ & ~new_n42937_;
  assign new_n43351_ = ~new_n43349_ & ~new_n43350_;
  assign new_n43352_ = ~new_n13350_ & ~new_n43351_;
  assign new_n43353_ = new_n13350_ & ~new_n25518_;
  assign new_n43354_ = ~new_n43352_ & ~new_n43353_;
  assign new_n43355_ = new_n13352_ & ~new_n43354_;
  assign new_n43356_ = ~new_n43348_ & ~new_n43355_;
  assign ys__n31225 = ys__n888 & ~new_n43356_;
  assign new_n43358_ = ys__n562 & ys__n47029;
  assign new_n43359_ = new_n43335_ & new_n43337_;
  assign new_n43360_ = ~new_n43358_ & new_n43359_;
  assign new_n43361_ = new_n43358_ & ~new_n43359_;
  assign new_n43362_ = ~new_n43360_ & ~new_n43361_;
  assign new_n43363_ = new_n42929_ & ~new_n43362_;
  assign new_n43364_ = new_n42926_ & new_n43358_;
  assign new_n43365_ = ys__n2652 & ys__n17831;
  assign new_n43366_ = ys__n39167 & new_n43313_;
  assign new_n43367_ = ~new_n43365_ & ~new_n43366_;
  assign new_n43368_ = ~new_n43364_ & new_n43367_;
  assign new_n43369_ = ~new_n43363_ & new_n43368_;
  assign new_n43370_ = new_n13353_ & ~new_n43369_;
  assign new_n43371_ = ~new_n25593_ & new_n42937_;
  assign new_n43372_ = ~new_n25585_ & ~new_n42937_;
  assign new_n43373_ = ~new_n43371_ & ~new_n43372_;
  assign new_n43374_ = ~new_n13350_ & ~new_n43373_;
  assign new_n43375_ = new_n13350_ & ~new_n25593_;
  assign new_n43376_ = ~new_n43374_ & ~new_n43375_;
  assign new_n43377_ = new_n13352_ & ~new_n43376_;
  assign new_n43378_ = ~new_n43370_ & ~new_n43377_;
  assign ys__n31226 = ys__n888 & ~new_n43378_;
  assign new_n43380_ = ys__n562 & ys__n47030;
  assign new_n43381_ = new_n43335_ & new_n43358_;
  assign new_n43382_ = new_n43336_ & new_n43381_;
  assign new_n43383_ = new_n43292_ & new_n43382_;
  assign new_n43384_ = ~new_n43380_ & new_n43383_;
  assign new_n43385_ = new_n43380_ & ~new_n43383_;
  assign new_n43386_ = ~new_n43384_ & ~new_n43385_;
  assign new_n43387_ = new_n42929_ & ~new_n43386_;
  assign new_n43388_ = new_n42926_ & new_n43380_;
  assign new_n43389_ = ys__n2652 & ys__n17833;
  assign new_n43390_ = ys__n39167 & new_n43335_;
  assign new_n43391_ = ~new_n43389_ & ~new_n43390_;
  assign new_n43392_ = ~new_n43388_ & new_n43391_;
  assign new_n43393_ = ~new_n43387_ & new_n43392_;
  assign new_n43394_ = new_n13353_ & ~new_n43393_;
  assign new_n43395_ = ~new_n25670_ & new_n42937_;
  assign new_n43396_ = ~new_n25664_ & ~new_n42937_;
  assign new_n43397_ = ~new_n43395_ & ~new_n43396_;
  assign new_n43398_ = ~new_n13350_ & ~new_n43397_;
  assign new_n43399_ = new_n13350_ & ~new_n25670_;
  assign new_n43400_ = ~new_n43398_ & ~new_n43399_;
  assign new_n43401_ = new_n13352_ & ~new_n43400_;
  assign new_n43402_ = ~new_n43394_ & ~new_n43401_;
  assign ys__n31227 = ys__n888 & ~new_n43402_;
  assign new_n43404_ = ys__n562 & ys__n47031;
  assign new_n43405_ = new_n43380_ & new_n43383_;
  assign new_n43406_ = ~new_n43404_ & new_n43405_;
  assign new_n43407_ = new_n43404_ & ~new_n43405_;
  assign new_n43408_ = ~new_n43406_ & ~new_n43407_;
  assign new_n43409_ = new_n42929_ & ~new_n43408_;
  assign new_n43410_ = new_n42926_ & new_n43404_;
  assign new_n43411_ = ys__n2652 & ys__n17834;
  assign new_n43412_ = ys__n39167 & new_n43358_;
  assign new_n43413_ = ~new_n43411_ & ~new_n43412_;
  assign new_n43414_ = ~new_n43410_ & new_n43413_;
  assign new_n43415_ = ~new_n43409_ & new_n43414_;
  assign new_n43416_ = new_n13353_ & ~new_n43415_;
  assign new_n43417_ = ~new_n25745_ & new_n42937_;
  assign new_n43418_ = ~new_n25737_ & ~new_n42937_;
  assign new_n43419_ = ~new_n43417_ & ~new_n43418_;
  assign new_n43420_ = ~new_n13350_ & ~new_n43419_;
  assign new_n43421_ = new_n13350_ & ~new_n25745_;
  assign new_n43422_ = ~new_n43420_ & ~new_n43421_;
  assign new_n43423_ = new_n13352_ & ~new_n43422_;
  assign new_n43424_ = ~new_n43416_ & ~new_n43423_;
  assign ys__n31228 = ys__n888 & ~new_n43424_;
  assign new_n43426_ = ys__n562 & ys__n47032;
  assign new_n43427_ = new_n43380_ & new_n43404_;
  assign new_n43428_ = new_n43383_ & new_n43427_;
  assign new_n43429_ = ~new_n43426_ & new_n43428_;
  assign new_n43430_ = new_n43426_ & ~new_n43428_;
  assign new_n43431_ = ~new_n43429_ & ~new_n43430_;
  assign new_n43432_ = new_n42929_ & ~new_n43431_;
  assign new_n43433_ = new_n42926_ & new_n43426_;
  assign new_n43434_ = ys__n2652 & ys__n17836;
  assign new_n43435_ = ys__n39167 & new_n43380_;
  assign new_n43436_ = ~new_n43434_ & ~new_n43435_;
  assign new_n43437_ = ~new_n43433_ & new_n43436_;
  assign new_n43438_ = ~new_n43432_ & new_n43437_;
  assign new_n43439_ = new_n13353_ & ~new_n43438_;
  assign new_n43440_ = ~new_n25825_ & new_n42937_;
  assign new_n43441_ = ~new_n25817_ & ~new_n42937_;
  assign new_n43442_ = ~new_n43440_ & ~new_n43441_;
  assign new_n43443_ = ~new_n13350_ & ~new_n43442_;
  assign new_n43444_ = new_n13350_ & ~new_n25825_;
  assign new_n43445_ = ~new_n43443_ & ~new_n43444_;
  assign new_n43446_ = new_n13352_ & ~new_n43445_;
  assign new_n43447_ = ~new_n43439_ & ~new_n43446_;
  assign ys__n31229 = ys__n888 & ~new_n43447_;
  assign new_n43449_ = ys__n562 & ys__n47033;
  assign new_n43450_ = new_n43426_ & new_n43428_;
  assign new_n43451_ = ~new_n43449_ & new_n43450_;
  assign new_n43452_ = new_n43449_ & ~new_n43450_;
  assign new_n43453_ = ~new_n43451_ & ~new_n43452_;
  assign new_n43454_ = new_n42929_ & ~new_n43453_;
  assign new_n43455_ = new_n42926_ & new_n43449_;
  assign new_n43456_ = ys__n2652 & ys__n17837;
  assign new_n43457_ = ys__n39167 & new_n43404_;
  assign new_n43458_ = ~new_n43456_ & ~new_n43457_;
  assign new_n43459_ = ~new_n43455_ & new_n43458_;
  assign new_n43460_ = ~new_n43454_ & new_n43459_;
  assign new_n43461_ = new_n13353_ & ~new_n43460_;
  assign new_n43462_ = ~new_n25901_ & new_n42937_;
  assign new_n43463_ = ~new_n25893_ & ~new_n42937_;
  assign new_n43464_ = ~new_n43462_ & ~new_n43463_;
  assign new_n43465_ = ~new_n13350_ & ~new_n43464_;
  assign new_n43466_ = new_n13350_ & ~new_n25901_;
  assign new_n43467_ = ~new_n43465_ & ~new_n43466_;
  assign new_n43468_ = new_n13352_ & ~new_n43467_;
  assign new_n43469_ = ~new_n43461_ & ~new_n43468_;
  assign ys__n31230 = ys__n888 & ~new_n43469_;
  assign new_n43471_ = ys__n562 & ys__n47034;
  assign new_n43472_ = new_n43426_ & new_n43449_;
  assign new_n43473_ = new_n43427_ & new_n43472_;
  assign new_n43474_ = new_n43382_ & new_n43473_;
  assign new_n43475_ = new_n43292_ & new_n43474_;
  assign new_n43476_ = ~new_n43471_ & new_n43475_;
  assign new_n43477_ = new_n43471_ & ~new_n43475_;
  assign new_n43478_ = ~new_n43476_ & ~new_n43477_;
  assign new_n43479_ = new_n42929_ & ~new_n43478_;
  assign new_n43480_ = new_n42926_ & new_n43471_;
  assign new_n43481_ = ys__n2652 & ys__n17839;
  assign new_n43482_ = ys__n39167 & new_n43426_;
  assign new_n43483_ = ~new_n43481_ & ~new_n43482_;
  assign new_n43484_ = ~new_n43480_ & new_n43483_;
  assign new_n43485_ = ~new_n43479_ & new_n43484_;
  assign new_n43486_ = new_n13353_ & ~new_n43485_;
  assign new_n43487_ = ~new_n25983_ & new_n42937_;
  assign new_n43488_ = ~new_n25977_ & ~new_n42937_;
  assign new_n43489_ = ~new_n43487_ & ~new_n43488_;
  assign new_n43490_ = ~new_n13350_ & ~new_n43489_;
  assign new_n43491_ = new_n13350_ & ~new_n25983_;
  assign new_n43492_ = ~new_n43490_ & ~new_n43491_;
  assign new_n43493_ = new_n13352_ & ~new_n43492_;
  assign new_n43494_ = ~new_n43486_ & ~new_n43493_;
  assign ys__n31231 = ys__n888 & ~new_n43494_;
  assign new_n43496_ = ys__n562 & ys__n47035;
  assign new_n43497_ = new_n43471_ & new_n43475_;
  assign new_n43498_ = ~new_n43496_ & new_n43497_;
  assign new_n43499_ = new_n43496_ & ~new_n43497_;
  assign new_n43500_ = ~new_n43498_ & ~new_n43499_;
  assign new_n43501_ = new_n42929_ & ~new_n43500_;
  assign new_n43502_ = new_n42926_ & new_n43496_;
  assign new_n43503_ = ys__n2652 & ys__n17840;
  assign new_n43504_ = ys__n39167 & new_n43449_;
  assign new_n43505_ = ~new_n43503_ & ~new_n43504_;
  assign new_n43506_ = ~new_n43502_ & new_n43505_;
  assign new_n43507_ = ~new_n43501_ & new_n43506_;
  assign new_n43508_ = new_n13353_ & ~new_n43507_;
  assign new_n43509_ = ~new_n26058_ & new_n42937_;
  assign new_n43510_ = ~new_n26050_ & ~new_n42937_;
  assign new_n43511_ = ~new_n43509_ & ~new_n43510_;
  assign new_n43512_ = ~new_n13350_ & ~new_n43511_;
  assign new_n43513_ = new_n13350_ & ~new_n26058_;
  assign new_n43514_ = ~new_n43512_ & ~new_n43513_;
  assign new_n43515_ = new_n13352_ & ~new_n43514_;
  assign new_n43516_ = ~new_n43508_ & ~new_n43515_;
  assign ys__n31232 = ys__n888 & ~new_n43516_;
  assign new_n43518_ = ys__n562 & ys__n47036;
  assign new_n43519_ = new_n43471_ & new_n43496_;
  assign new_n43520_ = new_n43475_ & new_n43519_;
  assign new_n43521_ = ~new_n43518_ & new_n43520_;
  assign new_n43522_ = new_n43518_ & ~new_n43520_;
  assign new_n43523_ = ~new_n43521_ & ~new_n43522_;
  assign new_n43524_ = new_n42929_ & ~new_n43523_;
  assign new_n43525_ = new_n42926_ & new_n43518_;
  assign new_n43526_ = ys__n2652 & ys__n17842;
  assign new_n43527_ = ys__n39167 & new_n43471_;
  assign new_n43528_ = ~new_n43526_ & ~new_n43527_;
  assign new_n43529_ = ~new_n43525_ & new_n43528_;
  assign new_n43530_ = ~new_n43524_ & new_n43529_;
  assign new_n43531_ = new_n13353_ & ~new_n43530_;
  assign new_n43532_ = ~new_n26138_ & new_n42937_;
  assign new_n43533_ = ~new_n26130_ & ~new_n42937_;
  assign new_n43534_ = ~new_n43532_ & ~new_n43533_;
  assign new_n43535_ = ~new_n13350_ & ~new_n43534_;
  assign new_n43536_ = new_n13350_ & ~new_n26138_;
  assign new_n43537_ = ~new_n43535_ & ~new_n43536_;
  assign new_n43538_ = new_n13352_ & ~new_n43537_;
  assign new_n43539_ = ~new_n43531_ & ~new_n43538_;
  assign ys__n31233 = ys__n888 & ~new_n43539_;
  assign new_n43541_ = ys__n562 & ys__n47037;
  assign new_n43542_ = new_n43518_ & new_n43520_;
  assign new_n43543_ = ~new_n43541_ & new_n43542_;
  assign new_n43544_ = new_n43541_ & ~new_n43542_;
  assign new_n43545_ = ~new_n43543_ & ~new_n43544_;
  assign new_n43546_ = new_n42929_ & ~new_n43545_;
  assign new_n43547_ = new_n42926_ & new_n43541_;
  assign new_n43548_ = ys__n2652 & ys__n17843;
  assign new_n43549_ = ys__n39167 & new_n43496_;
  assign new_n43550_ = ~new_n43548_ & ~new_n43549_;
  assign new_n43551_ = ~new_n43547_ & new_n43550_;
  assign new_n43552_ = ~new_n43546_ & new_n43551_;
  assign new_n43553_ = new_n13353_ & ~new_n43552_;
  assign new_n43554_ = ~new_n26214_ & new_n42937_;
  assign new_n43555_ = ~new_n26206_ & ~new_n42937_;
  assign new_n43556_ = ~new_n43554_ & ~new_n43555_;
  assign new_n43557_ = ~new_n13350_ & ~new_n43556_;
  assign new_n43558_ = new_n13350_ & ~new_n26214_;
  assign new_n43559_ = ~new_n43557_ & ~new_n43558_;
  assign new_n43560_ = new_n13352_ & ~new_n43559_;
  assign new_n43561_ = ~new_n43553_ & ~new_n43560_;
  assign ys__n31234 = ys__n888 & ~new_n43561_;
  assign new_n43563_ = ys__n562 & ys__n47038;
  assign new_n43564_ = new_n43518_ & new_n43541_;
  assign new_n43565_ = new_n43519_ & new_n43564_;
  assign new_n43566_ = new_n43475_ & new_n43565_;
  assign new_n43567_ = ~new_n43563_ & new_n43566_;
  assign new_n43568_ = new_n43563_ & ~new_n43566_;
  assign new_n43569_ = ~new_n43567_ & ~new_n43568_;
  assign new_n43570_ = new_n42929_ & ~new_n43569_;
  assign new_n43571_ = new_n42926_ & new_n43563_;
  assign new_n43572_ = ys__n2652 & ys__n17845;
  assign new_n43573_ = ys__n39167 & new_n43518_;
  assign new_n43574_ = ~new_n43572_ & ~new_n43573_;
  assign new_n43575_ = ~new_n43571_ & new_n43574_;
  assign new_n43576_ = ~new_n43570_ & new_n43575_;
  assign new_n43577_ = new_n13353_ & ~new_n43576_;
  assign new_n43578_ = ~new_n26298_ & new_n42937_;
  assign new_n43579_ = ~new_n26290_ & ~new_n42937_;
  assign new_n43580_ = ~new_n43578_ & ~new_n43579_;
  assign new_n43581_ = ~new_n13350_ & ~new_n43580_;
  assign new_n43582_ = new_n13350_ & ~new_n26298_;
  assign new_n43583_ = ~new_n43581_ & ~new_n43582_;
  assign new_n43584_ = new_n13352_ & ~new_n43583_;
  assign new_n43585_ = ~new_n43577_ & ~new_n43584_;
  assign ys__n31235 = ys__n888 & ~new_n43585_;
  assign new_n43587_ = ys__n562 & ys__n47039;
  assign new_n43588_ = new_n43563_ & new_n43566_;
  assign new_n43589_ = ~new_n43587_ & new_n43588_;
  assign new_n43590_ = new_n43587_ & ~new_n43588_;
  assign new_n43591_ = ~new_n43589_ & ~new_n43590_;
  assign new_n43592_ = new_n42929_ & ~new_n43591_;
  assign new_n43593_ = new_n42926_ & new_n43587_;
  assign new_n43594_ = ys__n2652 & ys__n17846;
  assign new_n43595_ = ys__n39167 & new_n43541_;
  assign new_n43596_ = ~new_n43594_ & ~new_n43595_;
  assign new_n43597_ = ~new_n43593_ & new_n43596_;
  assign new_n43598_ = ~new_n43592_ & new_n43597_;
  assign new_n43599_ = new_n13353_ & ~new_n43598_;
  assign new_n43600_ = ~new_n26374_ & new_n42937_;
  assign new_n43601_ = ~new_n26366_ & ~new_n42937_;
  assign new_n43602_ = ~new_n43600_ & ~new_n43601_;
  assign new_n43603_ = ~new_n13350_ & ~new_n43602_;
  assign new_n43604_ = new_n13350_ & ~new_n26374_;
  assign new_n43605_ = ~new_n43603_ & ~new_n43604_;
  assign new_n43606_ = new_n13352_ & ~new_n43605_;
  assign new_n43607_ = ~new_n43599_ & ~new_n43606_;
  assign ys__n31236 = ys__n888 & ~new_n43607_;
  assign new_n43609_ = ys__n562 & ys__n47040;
  assign new_n43610_ = new_n43563_ & new_n43587_;
  assign new_n43611_ = new_n43566_ & new_n43610_;
  assign new_n43612_ = ~new_n43609_ & new_n43611_;
  assign new_n43613_ = new_n43609_ & ~new_n43611_;
  assign new_n43614_ = ~new_n43612_ & ~new_n43613_;
  assign new_n43615_ = new_n42929_ & ~new_n43614_;
  assign new_n43616_ = new_n42926_ & new_n43609_;
  assign new_n43617_ = ys__n2652 & ys__n17848;
  assign new_n43618_ = ys__n39167 & new_n43563_;
  assign new_n43619_ = ~new_n43617_ & ~new_n43618_;
  assign new_n43620_ = ~new_n43616_ & new_n43619_;
  assign ys__n39392 = new_n43615_ | ~new_n43620_;
  assign new_n43622_ = new_n13353_ & ys__n39392;
  assign new_n43623_ = ~new_n26454_ & new_n42937_;
  assign new_n43624_ = ~new_n26446_ & ~new_n42937_;
  assign new_n43625_ = ~new_n43623_ & ~new_n43624_;
  assign new_n43626_ = ~new_n13350_ & ~new_n43625_;
  assign new_n43627_ = new_n13350_ & ~new_n26454_;
  assign new_n43628_ = ~new_n43626_ & ~new_n43627_;
  assign new_n43629_ = new_n13352_ & ~new_n43628_;
  assign new_n43630_ = ~new_n43622_ & ~new_n43629_;
  assign ys__n31237 = ys__n888 & ~new_n43630_;
  assign new_n43632_ = ys__n562 & ys__n47041;
  assign new_n43633_ = new_n43609_ & new_n43611_;
  assign new_n43634_ = ~new_n43632_ & new_n43633_;
  assign new_n43635_ = new_n43632_ & ~new_n43633_;
  assign new_n43636_ = ~new_n43634_ & ~new_n43635_;
  assign new_n43637_ = new_n42929_ & ~new_n43636_;
  assign new_n43638_ = new_n42926_ & new_n43632_;
  assign new_n43639_ = ys__n2652 & ys__n17849;
  assign new_n43640_ = ys__n39167 & new_n43587_;
  assign new_n43641_ = ~new_n43639_ & ~new_n43640_;
  assign new_n43642_ = ~new_n43638_ & new_n43641_;
  assign ys__n39393 = new_n43637_ | ~new_n43642_;
  assign new_n43644_ = new_n13353_ & ys__n39393;
  assign new_n43645_ = ~new_n26528_ & new_n42937_;
  assign new_n43646_ = ~new_n26520_ & ~new_n42937_;
  assign new_n43647_ = ~new_n43645_ & ~new_n43646_;
  assign new_n43648_ = ~new_n13350_ & ~new_n43647_;
  assign new_n43649_ = new_n13350_ & ~new_n26528_;
  assign new_n43650_ = ~new_n43648_ & ~new_n43649_;
  assign new_n43651_ = new_n13352_ & ~new_n43650_;
  assign new_n43652_ = ~new_n43644_ & ~new_n43651_;
  assign ys__n31238 = ys__n888 & ~new_n43652_;
  assign new_n43654_ = ys__n842 & new_n13240_;
  assign new_n43655_ = ys__n47234 & new_n43654_;
  assign new_n43656_ = ~ys__n844 & ~new_n13240_;
  assign new_n43657_ = ~ys__n842 & new_n13240_;
  assign new_n43658_ = ~new_n43656_ & ~new_n43657_;
  assign new_n43659_ = ys__n47202 & ~new_n43658_;
  assign new_n43660_ = ~new_n43655_ & ~new_n43659_;
  assign new_n43661_ = ~new_n43654_ & new_n43658_;
  assign ys__n31326 = ~new_n43660_ & ~new_n43661_;
  assign new_n43663_ = ys__n47235 & new_n43654_;
  assign new_n43664_ = ys__n47203 & ~new_n43658_;
  assign new_n43665_ = ~new_n43663_ & ~new_n43664_;
  assign ys__n31327 = ~new_n43661_ & ~new_n43665_;
  assign new_n43667_ = ys__n47236 & new_n43654_;
  assign new_n43668_ = ys__n47204 & ~new_n43658_;
  assign new_n43669_ = ~new_n43667_ & ~new_n43668_;
  assign ys__n31328 = ~new_n43661_ & ~new_n43669_;
  assign new_n43671_ = ys__n47237 & new_n43654_;
  assign new_n43672_ = ys__n47205 & ~new_n43658_;
  assign new_n43673_ = ~new_n43671_ & ~new_n43672_;
  assign ys__n31329 = ~new_n43661_ & ~new_n43673_;
  assign new_n43675_ = ys__n47238 & new_n43654_;
  assign new_n43676_ = ys__n47206 & ~new_n43658_;
  assign new_n43677_ = ~new_n43675_ & ~new_n43676_;
  assign ys__n31330 = ~new_n43661_ & ~new_n43677_;
  assign new_n43679_ = ys__n47239 & new_n43654_;
  assign new_n43680_ = ys__n47207 & ~new_n43658_;
  assign new_n43681_ = ~new_n43679_ & ~new_n43680_;
  assign ys__n31331 = ~new_n43661_ & ~new_n43681_;
  assign new_n43683_ = ys__n47240 & new_n43654_;
  assign new_n43684_ = ys__n47208 & ~new_n43658_;
  assign new_n43685_ = ~new_n43683_ & ~new_n43684_;
  assign ys__n31332 = ~new_n43661_ & ~new_n43685_;
  assign new_n43687_ = ys__n47241 & new_n43654_;
  assign new_n43688_ = ys__n47209 & ~new_n43658_;
  assign new_n43689_ = ~new_n43687_ & ~new_n43688_;
  assign ys__n31333 = ~new_n43661_ & ~new_n43689_;
  assign new_n43691_ = ys__n47242 & new_n43654_;
  assign new_n43692_ = ys__n47210 & ~new_n43658_;
  assign new_n43693_ = ~new_n43691_ & ~new_n43692_;
  assign ys__n31334 = ~new_n43661_ & ~new_n43693_;
  assign new_n43695_ = ys__n47243 & new_n43654_;
  assign new_n43696_ = ys__n47211 & ~new_n43658_;
  assign new_n43697_ = ~new_n43695_ & ~new_n43696_;
  assign ys__n31335 = ~new_n43661_ & ~new_n43697_;
  assign new_n43699_ = ys__n47244 & new_n43654_;
  assign new_n43700_ = ys__n47212 & ~new_n43658_;
  assign new_n43701_ = ~new_n43699_ & ~new_n43700_;
  assign ys__n31336 = ~new_n43661_ & ~new_n43701_;
  assign new_n43703_ = ys__n47245 & new_n43654_;
  assign new_n43704_ = ys__n47213 & ~new_n43658_;
  assign new_n43705_ = ~new_n43703_ & ~new_n43704_;
  assign ys__n31337 = ~new_n43661_ & ~new_n43705_;
  assign new_n43707_ = ys__n47246 & new_n43654_;
  assign new_n43708_ = ys__n47214 & ~new_n43658_;
  assign new_n43709_ = ~new_n43707_ & ~new_n43708_;
  assign ys__n31338 = ~new_n43661_ & ~new_n43709_;
  assign new_n43711_ = ys__n47247 & new_n43654_;
  assign new_n43712_ = ys__n47215 & ~new_n43658_;
  assign new_n43713_ = ~new_n43711_ & ~new_n43712_;
  assign ys__n31339 = ~new_n43661_ & ~new_n43713_;
  assign new_n43715_ = ys__n47248 & new_n43654_;
  assign new_n43716_ = ys__n47216 & ~new_n43658_;
  assign new_n43717_ = ~new_n43715_ & ~new_n43716_;
  assign ys__n31340 = ~new_n43661_ & ~new_n43717_;
  assign new_n43719_ = ys__n47249 & new_n43654_;
  assign new_n43720_ = ys__n47217 & ~new_n43658_;
  assign new_n43721_ = ~new_n43719_ & ~new_n43720_;
  assign ys__n31341 = ~new_n43661_ & ~new_n43721_;
  assign new_n43723_ = ys__n47250 & new_n43654_;
  assign new_n43724_ = ys__n47218 & ~new_n43658_;
  assign new_n43725_ = ~new_n43723_ & ~new_n43724_;
  assign ys__n31342 = ~new_n43661_ & ~new_n43725_;
  assign new_n43727_ = ys__n47251 & new_n43654_;
  assign new_n43728_ = ys__n47219 & ~new_n43658_;
  assign new_n43729_ = ~new_n43727_ & ~new_n43728_;
  assign ys__n31343 = ~new_n43661_ & ~new_n43729_;
  assign new_n43731_ = ys__n47252 & new_n43654_;
  assign new_n43732_ = ys__n47220 & ~new_n43658_;
  assign new_n43733_ = ~new_n43731_ & ~new_n43732_;
  assign ys__n31344 = ~new_n43661_ & ~new_n43733_;
  assign new_n43735_ = ys__n47253 & new_n43654_;
  assign new_n43736_ = ys__n47221 & ~new_n43658_;
  assign new_n43737_ = ~new_n43735_ & ~new_n43736_;
  assign ys__n31345 = ~new_n43661_ & ~new_n43737_;
  assign new_n43739_ = ys__n47254 & new_n43654_;
  assign new_n43740_ = ys__n47222 & ~new_n43658_;
  assign new_n43741_ = ~new_n43739_ & ~new_n43740_;
  assign ys__n31346 = ~new_n43661_ & ~new_n43741_;
  assign new_n43743_ = ys__n47255 & new_n43654_;
  assign new_n43744_ = ys__n47223 & ~new_n43658_;
  assign new_n43745_ = ~new_n43743_ & ~new_n43744_;
  assign ys__n31347 = ~new_n43661_ & ~new_n43745_;
  assign new_n43747_ = ys__n47256 & new_n43654_;
  assign new_n43748_ = ys__n47224 & ~new_n43658_;
  assign new_n43749_ = ~new_n43747_ & ~new_n43748_;
  assign ys__n31348 = ~new_n43661_ & ~new_n43749_;
  assign new_n43751_ = ys__n47257 & new_n43654_;
  assign new_n43752_ = ys__n47225 & ~new_n43658_;
  assign new_n43753_ = ~new_n43751_ & ~new_n43752_;
  assign ys__n31349 = ~new_n43661_ & ~new_n43753_;
  assign new_n43755_ = ys__n47258 & new_n43654_;
  assign new_n43756_ = ys__n47226 & ~new_n43658_;
  assign new_n43757_ = ~new_n43755_ & ~new_n43756_;
  assign ys__n31350 = ~new_n43661_ & ~new_n43757_;
  assign new_n43759_ = ys__n47259 & new_n43654_;
  assign new_n43760_ = ys__n47227 & ~new_n43658_;
  assign new_n43761_ = ~new_n43759_ & ~new_n43760_;
  assign ys__n31351 = ~new_n43661_ & ~new_n43761_;
  assign new_n43763_ = ys__n47260 & new_n43654_;
  assign new_n43764_ = ys__n47228 & ~new_n43658_;
  assign new_n43765_ = ~new_n43763_ & ~new_n43764_;
  assign ys__n31352 = ~new_n43661_ & ~new_n43765_;
  assign new_n43767_ = ys__n47261 & new_n43654_;
  assign new_n43768_ = ys__n47229 & ~new_n43658_;
  assign new_n43769_ = ~new_n43767_ & ~new_n43768_;
  assign ys__n31353 = ~new_n43661_ & ~new_n43769_;
  assign new_n43771_ = ys__n47262 & new_n43654_;
  assign new_n43772_ = ys__n47230 & ~new_n43658_;
  assign new_n43773_ = ~new_n43771_ & ~new_n43772_;
  assign ys__n31354 = ~new_n43661_ & ~new_n43773_;
  assign new_n43775_ = ys__n47263 & new_n43654_;
  assign new_n43776_ = ys__n47231 & ~new_n43658_;
  assign new_n43777_ = ~new_n43775_ & ~new_n43776_;
  assign ys__n31355 = ~new_n43661_ & ~new_n43777_;
  assign new_n43779_ = ys__n47264 & new_n43654_;
  assign new_n43780_ = ys__n47232 & ~new_n43658_;
  assign new_n43781_ = ~new_n43779_ & ~new_n43780_;
  assign ys__n31356 = ~new_n43661_ & ~new_n43781_;
  assign new_n43783_ = ys__n47265 & new_n43654_;
  assign new_n43784_ = ys__n47233 & ~new_n43658_;
  assign new_n43785_ = ~new_n43783_ & ~new_n43784_;
  assign ys__n31357 = ~new_n43661_ & ~new_n43785_;
  assign new_n43787_ = ys__n47266 & new_n43654_;
  assign new_n43788_ = ys__n18762 & ~new_n43658_;
  assign new_n43789_ = ~new_n43787_ & ~new_n43788_;
  assign ys__n31358 = ~new_n43661_ & ~new_n43789_;
  assign new_n43791_ = ys__n47267 & new_n43654_;
  assign new_n43792_ = ys__n18750 & ~new_n43658_;
  assign new_n43793_ = ~new_n43791_ & ~new_n43792_;
  assign ys__n31359 = ~new_n43661_ & ~new_n43793_;
  assign new_n43795_ = ys__n47268 & new_n43654_;
  assign new_n43796_ = ys__n18753 & ~new_n43658_;
  assign new_n43797_ = ~new_n43795_ & ~new_n43796_;
  assign ys__n31360 = ~new_n43661_ & ~new_n43797_;
  assign new_n43799_ = ys__n840 & new_n13240_;
  assign new_n43800_ = ys__n47269 & new_n43799_;
  assign new_n43801_ = ~ys__n842 & ~new_n13240_;
  assign new_n43802_ = ~ys__n840 & new_n13240_;
  assign new_n43803_ = ~new_n43801_ & ~new_n43802_;
  assign new_n43804_ = ys__n47202 & ~new_n43803_;
  assign new_n43805_ = ~new_n43800_ & ~new_n43804_;
  assign new_n43806_ = ~new_n43799_ & new_n43803_;
  assign ys__n31361 = ~new_n43805_ & ~new_n43806_;
  assign new_n43808_ = ys__n47270 & new_n43799_;
  assign new_n43809_ = ys__n47203 & ~new_n43803_;
  assign new_n43810_ = ~new_n43808_ & ~new_n43809_;
  assign ys__n31362 = ~new_n43806_ & ~new_n43810_;
  assign new_n43812_ = ys__n47271 & new_n43799_;
  assign new_n43813_ = ys__n47204 & ~new_n43803_;
  assign new_n43814_ = ~new_n43812_ & ~new_n43813_;
  assign ys__n31363 = ~new_n43806_ & ~new_n43814_;
  assign new_n43816_ = ys__n47272 & new_n43799_;
  assign new_n43817_ = ys__n47205 & ~new_n43803_;
  assign new_n43818_ = ~new_n43816_ & ~new_n43817_;
  assign ys__n31364 = ~new_n43806_ & ~new_n43818_;
  assign new_n43820_ = ys__n47273 & new_n43799_;
  assign new_n43821_ = ys__n47206 & ~new_n43803_;
  assign new_n43822_ = ~new_n43820_ & ~new_n43821_;
  assign ys__n31365 = ~new_n43806_ & ~new_n43822_;
  assign new_n43824_ = ys__n47274 & new_n43799_;
  assign new_n43825_ = ys__n47207 & ~new_n43803_;
  assign new_n43826_ = ~new_n43824_ & ~new_n43825_;
  assign ys__n31366 = ~new_n43806_ & ~new_n43826_;
  assign new_n43828_ = ys__n47275 & new_n43799_;
  assign new_n43829_ = ys__n47208 & ~new_n43803_;
  assign new_n43830_ = ~new_n43828_ & ~new_n43829_;
  assign ys__n31367 = ~new_n43806_ & ~new_n43830_;
  assign new_n43832_ = ys__n47276 & new_n43799_;
  assign new_n43833_ = ys__n47209 & ~new_n43803_;
  assign new_n43834_ = ~new_n43832_ & ~new_n43833_;
  assign ys__n31368 = ~new_n43806_ & ~new_n43834_;
  assign new_n43836_ = ys__n47277 & new_n43799_;
  assign new_n43837_ = ys__n47210 & ~new_n43803_;
  assign new_n43838_ = ~new_n43836_ & ~new_n43837_;
  assign ys__n31369 = ~new_n43806_ & ~new_n43838_;
  assign new_n43840_ = ys__n47278 & new_n43799_;
  assign new_n43841_ = ys__n47211 & ~new_n43803_;
  assign new_n43842_ = ~new_n43840_ & ~new_n43841_;
  assign ys__n31370 = ~new_n43806_ & ~new_n43842_;
  assign new_n43844_ = ys__n47279 & new_n43799_;
  assign new_n43845_ = ys__n47212 & ~new_n43803_;
  assign new_n43846_ = ~new_n43844_ & ~new_n43845_;
  assign ys__n31371 = ~new_n43806_ & ~new_n43846_;
  assign new_n43848_ = ys__n47280 & new_n43799_;
  assign new_n43849_ = ys__n47213 & ~new_n43803_;
  assign new_n43850_ = ~new_n43848_ & ~new_n43849_;
  assign ys__n31372 = ~new_n43806_ & ~new_n43850_;
  assign new_n43852_ = ys__n47281 & new_n43799_;
  assign new_n43853_ = ys__n47214 & ~new_n43803_;
  assign new_n43854_ = ~new_n43852_ & ~new_n43853_;
  assign ys__n31373 = ~new_n43806_ & ~new_n43854_;
  assign new_n43856_ = ys__n47282 & new_n43799_;
  assign new_n43857_ = ys__n47215 & ~new_n43803_;
  assign new_n43858_ = ~new_n43856_ & ~new_n43857_;
  assign ys__n31374 = ~new_n43806_ & ~new_n43858_;
  assign new_n43860_ = ys__n47283 & new_n43799_;
  assign new_n43861_ = ys__n47216 & ~new_n43803_;
  assign new_n43862_ = ~new_n43860_ & ~new_n43861_;
  assign ys__n31375 = ~new_n43806_ & ~new_n43862_;
  assign new_n43864_ = ys__n47284 & new_n43799_;
  assign new_n43865_ = ys__n47217 & ~new_n43803_;
  assign new_n43866_ = ~new_n43864_ & ~new_n43865_;
  assign ys__n31376 = ~new_n43806_ & ~new_n43866_;
  assign new_n43868_ = ys__n47285 & new_n43799_;
  assign new_n43869_ = ys__n47218 & ~new_n43803_;
  assign new_n43870_ = ~new_n43868_ & ~new_n43869_;
  assign ys__n31377 = ~new_n43806_ & ~new_n43870_;
  assign new_n43872_ = ys__n47286 & new_n43799_;
  assign new_n43873_ = ys__n47219 & ~new_n43803_;
  assign new_n43874_ = ~new_n43872_ & ~new_n43873_;
  assign ys__n31378 = ~new_n43806_ & ~new_n43874_;
  assign new_n43876_ = ys__n47287 & new_n43799_;
  assign new_n43877_ = ys__n47220 & ~new_n43803_;
  assign new_n43878_ = ~new_n43876_ & ~new_n43877_;
  assign ys__n31379 = ~new_n43806_ & ~new_n43878_;
  assign new_n43880_ = ys__n47288 & new_n43799_;
  assign new_n43881_ = ys__n47221 & ~new_n43803_;
  assign new_n43882_ = ~new_n43880_ & ~new_n43881_;
  assign ys__n31380 = ~new_n43806_ & ~new_n43882_;
  assign new_n43884_ = ys__n47289 & new_n43799_;
  assign new_n43885_ = ys__n47222 & ~new_n43803_;
  assign new_n43886_ = ~new_n43884_ & ~new_n43885_;
  assign ys__n31381 = ~new_n43806_ & ~new_n43886_;
  assign new_n43888_ = ys__n47290 & new_n43799_;
  assign new_n43889_ = ys__n47223 & ~new_n43803_;
  assign new_n43890_ = ~new_n43888_ & ~new_n43889_;
  assign ys__n31382 = ~new_n43806_ & ~new_n43890_;
  assign new_n43892_ = ys__n47291 & new_n43799_;
  assign new_n43893_ = ys__n47224 & ~new_n43803_;
  assign new_n43894_ = ~new_n43892_ & ~new_n43893_;
  assign ys__n31383 = ~new_n43806_ & ~new_n43894_;
  assign new_n43896_ = ys__n47292 & new_n43799_;
  assign new_n43897_ = ys__n47225 & ~new_n43803_;
  assign new_n43898_ = ~new_n43896_ & ~new_n43897_;
  assign ys__n31384 = ~new_n43806_ & ~new_n43898_;
  assign new_n43900_ = ys__n47293 & new_n43799_;
  assign new_n43901_ = ys__n47226 & ~new_n43803_;
  assign new_n43902_ = ~new_n43900_ & ~new_n43901_;
  assign ys__n31385 = ~new_n43806_ & ~new_n43902_;
  assign new_n43904_ = ys__n47294 & new_n43799_;
  assign new_n43905_ = ys__n47227 & ~new_n43803_;
  assign new_n43906_ = ~new_n43904_ & ~new_n43905_;
  assign ys__n31386 = ~new_n43806_ & ~new_n43906_;
  assign new_n43908_ = ys__n47295 & new_n43799_;
  assign new_n43909_ = ys__n47228 & ~new_n43803_;
  assign new_n43910_ = ~new_n43908_ & ~new_n43909_;
  assign ys__n31387 = ~new_n43806_ & ~new_n43910_;
  assign new_n43912_ = ys__n47296 & new_n43799_;
  assign new_n43913_ = ys__n47229 & ~new_n43803_;
  assign new_n43914_ = ~new_n43912_ & ~new_n43913_;
  assign ys__n31388 = ~new_n43806_ & ~new_n43914_;
  assign new_n43916_ = ys__n47297 & new_n43799_;
  assign new_n43917_ = ys__n47230 & ~new_n43803_;
  assign new_n43918_ = ~new_n43916_ & ~new_n43917_;
  assign ys__n31389 = ~new_n43806_ & ~new_n43918_;
  assign new_n43920_ = ys__n47298 & new_n43799_;
  assign new_n43921_ = ys__n47231 & ~new_n43803_;
  assign new_n43922_ = ~new_n43920_ & ~new_n43921_;
  assign ys__n31390 = ~new_n43806_ & ~new_n43922_;
  assign new_n43924_ = ys__n47299 & new_n43799_;
  assign new_n43925_ = ys__n47232 & ~new_n43803_;
  assign new_n43926_ = ~new_n43924_ & ~new_n43925_;
  assign ys__n31391 = ~new_n43806_ & ~new_n43926_;
  assign new_n43928_ = ys__n47300 & new_n43799_;
  assign new_n43929_ = ys__n47233 & ~new_n43803_;
  assign new_n43930_ = ~new_n43928_ & ~new_n43929_;
  assign ys__n31392 = ~new_n43806_ & ~new_n43930_;
  assign new_n43932_ = ys__n47301 & new_n43799_;
  assign new_n43933_ = ys__n18762 & ~new_n43803_;
  assign new_n43934_ = ~new_n43932_ & ~new_n43933_;
  assign ys__n31393 = ~new_n43806_ & ~new_n43934_;
  assign new_n43936_ = ys__n47302 & new_n43799_;
  assign new_n43937_ = ys__n18750 & ~new_n43803_;
  assign new_n43938_ = ~new_n43936_ & ~new_n43937_;
  assign ys__n31394 = ~new_n43806_ & ~new_n43938_;
  assign new_n43940_ = ys__n47303 & new_n43799_;
  assign new_n43941_ = ys__n18753 & ~new_n43803_;
  assign new_n43942_ = ~new_n43940_ & ~new_n43941_;
  assign ys__n31395 = ~new_n43806_ & ~new_n43942_;
  assign new_n43944_ = ys__n838 & new_n13240_;
  assign new_n43945_ = ys__n47305 & new_n43944_;
  assign new_n43946_ = ~ys__n840 & ~new_n13240_;
  assign new_n43947_ = ~ys__n838 & new_n13240_;
  assign new_n43948_ = ~new_n43946_ & ~new_n43947_;
  assign new_n43949_ = ys__n47202 & ~new_n43948_;
  assign new_n43950_ = ~new_n43945_ & ~new_n43949_;
  assign new_n43951_ = ~new_n43944_ & new_n43948_;
  assign ys__n31397 = ~new_n43950_ & ~new_n43951_;
  assign new_n43953_ = ys__n47306 & new_n43944_;
  assign new_n43954_ = ys__n47203 & ~new_n43948_;
  assign new_n43955_ = ~new_n43953_ & ~new_n43954_;
  assign ys__n31398 = ~new_n43951_ & ~new_n43955_;
  assign new_n43957_ = ys__n47307 & new_n43944_;
  assign new_n43958_ = ys__n47204 & ~new_n43948_;
  assign new_n43959_ = ~new_n43957_ & ~new_n43958_;
  assign ys__n31399 = ~new_n43951_ & ~new_n43959_;
  assign new_n43961_ = ys__n47308 & new_n43944_;
  assign new_n43962_ = ys__n47205 & ~new_n43948_;
  assign new_n43963_ = ~new_n43961_ & ~new_n43962_;
  assign ys__n31400 = ~new_n43951_ & ~new_n43963_;
  assign new_n43965_ = ys__n47309 & new_n43944_;
  assign new_n43966_ = ys__n47206 & ~new_n43948_;
  assign new_n43967_ = ~new_n43965_ & ~new_n43966_;
  assign ys__n31401 = ~new_n43951_ & ~new_n43967_;
  assign new_n43969_ = ys__n47310 & new_n43944_;
  assign new_n43970_ = ys__n47207 & ~new_n43948_;
  assign new_n43971_ = ~new_n43969_ & ~new_n43970_;
  assign ys__n31402 = ~new_n43951_ & ~new_n43971_;
  assign new_n43973_ = ys__n47311 & new_n43944_;
  assign new_n43974_ = ys__n47208 & ~new_n43948_;
  assign new_n43975_ = ~new_n43973_ & ~new_n43974_;
  assign ys__n31403 = ~new_n43951_ & ~new_n43975_;
  assign new_n43977_ = ys__n47312 & new_n43944_;
  assign new_n43978_ = ys__n47209 & ~new_n43948_;
  assign new_n43979_ = ~new_n43977_ & ~new_n43978_;
  assign ys__n31404 = ~new_n43951_ & ~new_n43979_;
  assign new_n43981_ = ys__n47313 & new_n43944_;
  assign new_n43982_ = ys__n47210 & ~new_n43948_;
  assign new_n43983_ = ~new_n43981_ & ~new_n43982_;
  assign ys__n31405 = ~new_n43951_ & ~new_n43983_;
  assign new_n43985_ = ys__n47314 & new_n43944_;
  assign new_n43986_ = ys__n47211 & ~new_n43948_;
  assign new_n43987_ = ~new_n43985_ & ~new_n43986_;
  assign ys__n31406 = ~new_n43951_ & ~new_n43987_;
  assign new_n43989_ = ys__n47315 & new_n43944_;
  assign new_n43990_ = ys__n47212 & ~new_n43948_;
  assign new_n43991_ = ~new_n43989_ & ~new_n43990_;
  assign ys__n31407 = ~new_n43951_ & ~new_n43991_;
  assign new_n43993_ = ys__n47316 & new_n43944_;
  assign new_n43994_ = ys__n47213 & ~new_n43948_;
  assign new_n43995_ = ~new_n43993_ & ~new_n43994_;
  assign ys__n31408 = ~new_n43951_ & ~new_n43995_;
  assign new_n43997_ = ys__n47317 & new_n43944_;
  assign new_n43998_ = ys__n47214 & ~new_n43948_;
  assign new_n43999_ = ~new_n43997_ & ~new_n43998_;
  assign ys__n31409 = ~new_n43951_ & ~new_n43999_;
  assign new_n44001_ = ys__n47318 & new_n43944_;
  assign new_n44002_ = ys__n47215 & ~new_n43948_;
  assign new_n44003_ = ~new_n44001_ & ~new_n44002_;
  assign ys__n31410 = ~new_n43951_ & ~new_n44003_;
  assign new_n44005_ = ys__n47319 & new_n43944_;
  assign new_n44006_ = ys__n47216 & ~new_n43948_;
  assign new_n44007_ = ~new_n44005_ & ~new_n44006_;
  assign ys__n31411 = ~new_n43951_ & ~new_n44007_;
  assign new_n44009_ = ys__n47320 & new_n43944_;
  assign new_n44010_ = ys__n47217 & ~new_n43948_;
  assign new_n44011_ = ~new_n44009_ & ~new_n44010_;
  assign ys__n31412 = ~new_n43951_ & ~new_n44011_;
  assign new_n44013_ = ys__n47321 & new_n43944_;
  assign new_n44014_ = ys__n47218 & ~new_n43948_;
  assign new_n44015_ = ~new_n44013_ & ~new_n44014_;
  assign ys__n31413 = ~new_n43951_ & ~new_n44015_;
  assign new_n44017_ = ys__n47322 & new_n43944_;
  assign new_n44018_ = ys__n47219 & ~new_n43948_;
  assign new_n44019_ = ~new_n44017_ & ~new_n44018_;
  assign ys__n31414 = ~new_n43951_ & ~new_n44019_;
  assign new_n44021_ = ys__n47323 & new_n43944_;
  assign new_n44022_ = ys__n47220 & ~new_n43948_;
  assign new_n44023_ = ~new_n44021_ & ~new_n44022_;
  assign ys__n31415 = ~new_n43951_ & ~new_n44023_;
  assign new_n44025_ = ys__n47324 & new_n43944_;
  assign new_n44026_ = ys__n47221 & ~new_n43948_;
  assign new_n44027_ = ~new_n44025_ & ~new_n44026_;
  assign ys__n31416 = ~new_n43951_ & ~new_n44027_;
  assign new_n44029_ = ys__n47325 & new_n43944_;
  assign new_n44030_ = ys__n47222 & ~new_n43948_;
  assign new_n44031_ = ~new_n44029_ & ~new_n44030_;
  assign ys__n31417 = ~new_n43951_ & ~new_n44031_;
  assign new_n44033_ = ys__n47326 & new_n43944_;
  assign new_n44034_ = ys__n47223 & ~new_n43948_;
  assign new_n44035_ = ~new_n44033_ & ~new_n44034_;
  assign ys__n31418 = ~new_n43951_ & ~new_n44035_;
  assign new_n44037_ = ys__n47327 & new_n43944_;
  assign new_n44038_ = ys__n47224 & ~new_n43948_;
  assign new_n44039_ = ~new_n44037_ & ~new_n44038_;
  assign ys__n31419 = ~new_n43951_ & ~new_n44039_;
  assign new_n44041_ = ys__n47328 & new_n43944_;
  assign new_n44042_ = ys__n47225 & ~new_n43948_;
  assign new_n44043_ = ~new_n44041_ & ~new_n44042_;
  assign ys__n31420 = ~new_n43951_ & ~new_n44043_;
  assign new_n44045_ = ys__n47329 & new_n43944_;
  assign new_n44046_ = ys__n47226 & ~new_n43948_;
  assign new_n44047_ = ~new_n44045_ & ~new_n44046_;
  assign ys__n31421 = ~new_n43951_ & ~new_n44047_;
  assign new_n44049_ = ys__n47330 & new_n43944_;
  assign new_n44050_ = ys__n47227 & ~new_n43948_;
  assign new_n44051_ = ~new_n44049_ & ~new_n44050_;
  assign ys__n31422 = ~new_n43951_ & ~new_n44051_;
  assign new_n44053_ = ys__n47331 & new_n43944_;
  assign new_n44054_ = ys__n47228 & ~new_n43948_;
  assign new_n44055_ = ~new_n44053_ & ~new_n44054_;
  assign ys__n31423 = ~new_n43951_ & ~new_n44055_;
  assign new_n44057_ = ys__n47332 & new_n43944_;
  assign new_n44058_ = ys__n47229 & ~new_n43948_;
  assign new_n44059_ = ~new_n44057_ & ~new_n44058_;
  assign ys__n31424 = ~new_n43951_ & ~new_n44059_;
  assign new_n44061_ = ys__n47333 & new_n43944_;
  assign new_n44062_ = ys__n47230 & ~new_n43948_;
  assign new_n44063_ = ~new_n44061_ & ~new_n44062_;
  assign ys__n31425 = ~new_n43951_ & ~new_n44063_;
  assign new_n44065_ = ys__n47334 & new_n43944_;
  assign new_n44066_ = ys__n47231 & ~new_n43948_;
  assign new_n44067_ = ~new_n44065_ & ~new_n44066_;
  assign ys__n31426 = ~new_n43951_ & ~new_n44067_;
  assign new_n44069_ = ys__n47335 & new_n43944_;
  assign new_n44070_ = ys__n47232 & ~new_n43948_;
  assign new_n44071_ = ~new_n44069_ & ~new_n44070_;
  assign ys__n31427 = ~new_n43951_ & ~new_n44071_;
  assign new_n44073_ = ys__n47336 & new_n43944_;
  assign new_n44074_ = ys__n47233 & ~new_n43948_;
  assign new_n44075_ = ~new_n44073_ & ~new_n44074_;
  assign ys__n31428 = ~new_n43951_ & ~new_n44075_;
  assign new_n44077_ = ys__n47337 & new_n43944_;
  assign new_n44078_ = ys__n18762 & ~new_n43948_;
  assign new_n44079_ = ~new_n44077_ & ~new_n44078_;
  assign ys__n31429 = ~new_n43951_ & ~new_n44079_;
  assign new_n44081_ = ys__n47338 & new_n43944_;
  assign new_n44082_ = ys__n18750 & ~new_n43948_;
  assign new_n44083_ = ~new_n44081_ & ~new_n44082_;
  assign ys__n31430 = ~new_n43951_ & ~new_n44083_;
  assign new_n44085_ = ys__n47339 & new_n43944_;
  assign new_n44086_ = ys__n18753 & ~new_n43948_;
  assign new_n44087_ = ~new_n44085_ & ~new_n44086_;
  assign ys__n31431 = ~new_n43951_ & ~new_n44087_;
  assign new_n44089_ = ys__n1386 & ys__n24188;
  assign new_n44090_ = ys__n47340 & ~ys__n2152;
  assign new_n44091_ = ys__n47342 & new_n36477_;
  assign new_n44092_ = ys__n47341 & new_n36479_;
  assign new_n44093_ = ~new_n44091_ & ~new_n44092_;
  assign new_n44094_ = ~ys__n182 & ~new_n36477_;
  assign new_n44095_ = ~new_n36479_ & new_n44094_;
  assign new_n44096_ = ~new_n44093_ & ~new_n44095_;
  assign new_n44097_ = new_n42891_ & new_n44096_;
  assign new_n44098_ = ~new_n44090_ & ~new_n44097_;
  assign new_n44099_ = ~new_n44089_ & new_n44098_;
  assign new_n44100_ = ys__n2152 & new_n42903_;
  assign ys__n33007 = ~new_n44099_ & ~new_n44100_;
  assign new_n44102_ = ~ys__n500 & new_n13763_;
  assign new_n44103_ = ~ys__n1386 & new_n44102_;
  assign new_n44104_ = ~ys__n1386 & ~new_n44103_;
  assign new_n44105_ = ys__n33007 & ~new_n44104_;
  assign new_n44106_ = ys__n502 & ~ys__n2152;
  assign new_n44107_ = ~ys__n504 & ~ys__n2152;
  assign new_n44108_ = ~ys__n502 & new_n44107_;
  assign new_n44109_ = ~new_n44106_ & ~new_n44108_;
  assign new_n44110_ = ys__n28787 & ~new_n44109_;
  assign new_n44111_ = ys__n504 & ~ys__n2152;
  assign new_n44112_ = ~ys__n502 & new_n44111_;
  assign new_n44113_ = ys__n47185 & new_n44112_;
  assign new_n44114_ = ys__n500 & new_n13763_;
  assign new_n44115_ = ~ys__n1386 & new_n44114_;
  assign new_n44116_ = ys__n47340 & new_n44115_;
  assign new_n44117_ = ~new_n44113_ & ~new_n44116_;
  assign new_n44118_ = ~new_n44110_ & new_n44117_;
  assign new_n44119_ = ~new_n44105_ & new_n44118_;
  assign new_n44120_ = new_n44104_ & ~new_n44115_;
  assign new_n44121_ = ~new_n44112_ & new_n44120_;
  assign new_n44122_ = new_n44109_ & new_n44121_;
  assign ys__n31432 = ~new_n44119_ & ~new_n44122_;
  assign new_n44124_ = ys__n1386 & ys__n24191;
  assign new_n44125_ = ys__n47341 & ~ys__n2152;
  assign new_n44126_ = ys__n47342 & new_n36479_;
  assign new_n44127_ = ~new_n44095_ & new_n44126_;
  assign new_n44128_ = new_n42891_ & new_n44127_;
  assign new_n44129_ = ~new_n44125_ & ~new_n44128_;
  assign new_n44130_ = ~new_n44124_ & new_n44129_;
  assign ys__n33008 = ~new_n44100_ & ~new_n44130_;
  assign new_n44132_ = ~new_n44104_ & ys__n33008;
  assign new_n44133_ = ys__n28788 & ~new_n44109_;
  assign new_n44134_ = ys__n47184 & new_n44112_;
  assign new_n44135_ = ys__n47341 & new_n44115_;
  assign new_n44136_ = ~new_n44134_ & ~new_n44135_;
  assign new_n44137_ = ~new_n44133_ & new_n44136_;
  assign new_n44138_ = ~new_n44132_ & new_n44137_;
  assign ys__n31433 = ~new_n44122_ & ~new_n44138_;
  assign new_n44140_ = ys__n47342 & ~ys__n2152;
  assign new_n44141_ = ys__n714 & ys__n1386;
  assign new_n44142_ = ~new_n44140_ & ~new_n44141_;
  assign ys__n33009 = ~new_n44100_ & ~new_n44142_;
  assign new_n44144_ = ~new_n44104_ & ys__n33009;
  assign new_n44145_ = ys__n28789 & ~new_n44109_;
  assign new_n44146_ = ys__n46956 & new_n44112_;
  assign new_n44147_ = ys__n47342 & new_n44115_;
  assign new_n44148_ = ~new_n44146_ & ~new_n44147_;
  assign new_n44149_ = ~new_n44145_ & new_n44148_;
  assign new_n44150_ = ~new_n44144_ & new_n44149_;
  assign ys__n31434 = ~new_n44122_ & ~new_n44150_;
  assign new_n44152_ = ys__n46957 & new_n44112_;
  assign new_n44153_ = ys__n28790 & ~new_n44109_;
  assign new_n44154_ = ~new_n44152_ & ~new_n44153_;
  assign ys__n31435 = ~new_n44122_ & ~new_n44154_;
  assign new_n44156_ = ys__n46958 & new_n44112_;
  assign new_n44157_ = ys__n28791 & ~new_n44109_;
  assign new_n44158_ = ~new_n44156_ & ~new_n44157_;
  assign ys__n31436 = ~new_n44122_ & ~new_n44158_;
  assign new_n44160_ = ys__n46959 & new_n44112_;
  assign new_n44161_ = ys__n28792 & ~new_n44109_;
  assign new_n44162_ = ~new_n44160_ & ~new_n44161_;
  assign ys__n31437 = ~new_n44122_ & ~new_n44162_;
  assign new_n44164_ = ys__n46960 & new_n44112_;
  assign new_n44165_ = ys__n28793 & ~new_n44109_;
  assign new_n44166_ = ~new_n44164_ & ~new_n44165_;
  assign ys__n31438 = ~new_n44122_ & ~new_n44166_;
  assign new_n44168_ = ys__n46961 & new_n44112_;
  assign new_n44169_ = ys__n28794 & ~new_n44109_;
  assign new_n44170_ = ~new_n44168_ & ~new_n44169_;
  assign ys__n31439 = ~new_n44122_ & ~new_n44170_;
  assign new_n44172_ = ys__n836 & new_n13240_;
  assign new_n44173_ = ys__n47343 & new_n44172_;
  assign new_n44174_ = ~ys__n838 & ~new_n13240_;
  assign new_n44175_ = ~ys__n836 & new_n13240_;
  assign new_n44176_ = ~new_n44174_ & ~new_n44175_;
  assign new_n44177_ = ys__n47202 & ~new_n44176_;
  assign new_n44178_ = ~new_n44173_ & ~new_n44177_;
  assign new_n44179_ = ~new_n44172_ & new_n44176_;
  assign ys__n31440 = ~new_n44178_ & ~new_n44179_;
  assign new_n44181_ = ys__n47344 & new_n44172_;
  assign new_n44182_ = ys__n47203 & ~new_n44176_;
  assign new_n44183_ = ~new_n44181_ & ~new_n44182_;
  assign ys__n31441 = ~new_n44179_ & ~new_n44183_;
  assign new_n44185_ = ys__n47345 & new_n44172_;
  assign new_n44186_ = ys__n47204 & ~new_n44176_;
  assign new_n44187_ = ~new_n44185_ & ~new_n44186_;
  assign ys__n31442 = ~new_n44179_ & ~new_n44187_;
  assign new_n44189_ = ys__n47346 & new_n44172_;
  assign new_n44190_ = ys__n47205 & ~new_n44176_;
  assign new_n44191_ = ~new_n44189_ & ~new_n44190_;
  assign ys__n31443 = ~new_n44179_ & ~new_n44191_;
  assign new_n44193_ = ys__n47347 & new_n44172_;
  assign new_n44194_ = ys__n47206 & ~new_n44176_;
  assign new_n44195_ = ~new_n44193_ & ~new_n44194_;
  assign ys__n31444 = ~new_n44179_ & ~new_n44195_;
  assign new_n44197_ = ys__n47348 & new_n44172_;
  assign new_n44198_ = ys__n47207 & ~new_n44176_;
  assign new_n44199_ = ~new_n44197_ & ~new_n44198_;
  assign ys__n31445 = ~new_n44179_ & ~new_n44199_;
  assign new_n44201_ = ys__n47349 & new_n44172_;
  assign new_n44202_ = ys__n47208 & ~new_n44176_;
  assign new_n44203_ = ~new_n44201_ & ~new_n44202_;
  assign ys__n31446 = ~new_n44179_ & ~new_n44203_;
  assign new_n44205_ = ys__n47350 & new_n44172_;
  assign new_n44206_ = ys__n47209 & ~new_n44176_;
  assign new_n44207_ = ~new_n44205_ & ~new_n44206_;
  assign ys__n31447 = ~new_n44179_ & ~new_n44207_;
  assign new_n44209_ = ys__n47351 & new_n44172_;
  assign new_n44210_ = ys__n47210 & ~new_n44176_;
  assign new_n44211_ = ~new_n44209_ & ~new_n44210_;
  assign ys__n31448 = ~new_n44179_ & ~new_n44211_;
  assign new_n44213_ = ys__n47352 & new_n44172_;
  assign new_n44214_ = ys__n47211 & ~new_n44176_;
  assign new_n44215_ = ~new_n44213_ & ~new_n44214_;
  assign ys__n31449 = ~new_n44179_ & ~new_n44215_;
  assign new_n44217_ = ys__n47353 & new_n44172_;
  assign new_n44218_ = ys__n47212 & ~new_n44176_;
  assign new_n44219_ = ~new_n44217_ & ~new_n44218_;
  assign ys__n31450 = ~new_n44179_ & ~new_n44219_;
  assign new_n44221_ = ys__n47354 & new_n44172_;
  assign new_n44222_ = ys__n47213 & ~new_n44176_;
  assign new_n44223_ = ~new_n44221_ & ~new_n44222_;
  assign ys__n31451 = ~new_n44179_ & ~new_n44223_;
  assign new_n44225_ = ys__n47355 & new_n44172_;
  assign new_n44226_ = ys__n47214 & ~new_n44176_;
  assign new_n44227_ = ~new_n44225_ & ~new_n44226_;
  assign ys__n31452 = ~new_n44179_ & ~new_n44227_;
  assign new_n44229_ = ys__n47356 & new_n44172_;
  assign new_n44230_ = ys__n47215 & ~new_n44176_;
  assign new_n44231_ = ~new_n44229_ & ~new_n44230_;
  assign ys__n31453 = ~new_n44179_ & ~new_n44231_;
  assign new_n44233_ = ys__n47357 & new_n44172_;
  assign new_n44234_ = ys__n47216 & ~new_n44176_;
  assign new_n44235_ = ~new_n44233_ & ~new_n44234_;
  assign ys__n31454 = ~new_n44179_ & ~new_n44235_;
  assign new_n44237_ = ys__n47358 & new_n44172_;
  assign new_n44238_ = ys__n47217 & ~new_n44176_;
  assign new_n44239_ = ~new_n44237_ & ~new_n44238_;
  assign ys__n31455 = ~new_n44179_ & ~new_n44239_;
  assign new_n44241_ = ys__n47359 & new_n44172_;
  assign new_n44242_ = ys__n47218 & ~new_n44176_;
  assign new_n44243_ = ~new_n44241_ & ~new_n44242_;
  assign ys__n31456 = ~new_n44179_ & ~new_n44243_;
  assign new_n44245_ = ys__n47360 & new_n44172_;
  assign new_n44246_ = ys__n47219 & ~new_n44176_;
  assign new_n44247_ = ~new_n44245_ & ~new_n44246_;
  assign ys__n31457 = ~new_n44179_ & ~new_n44247_;
  assign new_n44249_ = ys__n47361 & new_n44172_;
  assign new_n44250_ = ys__n47220 & ~new_n44176_;
  assign new_n44251_ = ~new_n44249_ & ~new_n44250_;
  assign ys__n31458 = ~new_n44179_ & ~new_n44251_;
  assign new_n44253_ = ys__n47362 & new_n44172_;
  assign new_n44254_ = ys__n47221 & ~new_n44176_;
  assign new_n44255_ = ~new_n44253_ & ~new_n44254_;
  assign ys__n31459 = ~new_n44179_ & ~new_n44255_;
  assign new_n44257_ = ys__n47363 & new_n44172_;
  assign new_n44258_ = ys__n47222 & ~new_n44176_;
  assign new_n44259_ = ~new_n44257_ & ~new_n44258_;
  assign ys__n31460 = ~new_n44179_ & ~new_n44259_;
  assign new_n44261_ = ys__n47364 & new_n44172_;
  assign new_n44262_ = ys__n47223 & ~new_n44176_;
  assign new_n44263_ = ~new_n44261_ & ~new_n44262_;
  assign ys__n31461 = ~new_n44179_ & ~new_n44263_;
  assign new_n44265_ = ys__n47365 & new_n44172_;
  assign new_n44266_ = ys__n47224 & ~new_n44176_;
  assign new_n44267_ = ~new_n44265_ & ~new_n44266_;
  assign ys__n31462 = ~new_n44179_ & ~new_n44267_;
  assign new_n44269_ = ys__n47366 & new_n44172_;
  assign new_n44270_ = ys__n47225 & ~new_n44176_;
  assign new_n44271_ = ~new_n44269_ & ~new_n44270_;
  assign ys__n31463 = ~new_n44179_ & ~new_n44271_;
  assign new_n44273_ = ys__n47367 & new_n44172_;
  assign new_n44274_ = ys__n47226 & ~new_n44176_;
  assign new_n44275_ = ~new_n44273_ & ~new_n44274_;
  assign ys__n31464 = ~new_n44179_ & ~new_n44275_;
  assign new_n44277_ = ys__n47368 & new_n44172_;
  assign new_n44278_ = ys__n47227 & ~new_n44176_;
  assign new_n44279_ = ~new_n44277_ & ~new_n44278_;
  assign ys__n31465 = ~new_n44179_ & ~new_n44279_;
  assign new_n44281_ = ys__n47369 & new_n44172_;
  assign new_n44282_ = ys__n47228 & ~new_n44176_;
  assign new_n44283_ = ~new_n44281_ & ~new_n44282_;
  assign ys__n31466 = ~new_n44179_ & ~new_n44283_;
  assign new_n44285_ = ys__n47370 & new_n44172_;
  assign new_n44286_ = ys__n47229 & ~new_n44176_;
  assign new_n44287_ = ~new_n44285_ & ~new_n44286_;
  assign ys__n31467 = ~new_n44179_ & ~new_n44287_;
  assign new_n44289_ = ys__n47371 & new_n44172_;
  assign new_n44290_ = ys__n47230 & ~new_n44176_;
  assign new_n44291_ = ~new_n44289_ & ~new_n44290_;
  assign ys__n31468 = ~new_n44179_ & ~new_n44291_;
  assign new_n44293_ = ys__n47372 & new_n44172_;
  assign new_n44294_ = ys__n47231 & ~new_n44176_;
  assign new_n44295_ = ~new_n44293_ & ~new_n44294_;
  assign ys__n31469 = ~new_n44179_ & ~new_n44295_;
  assign new_n44297_ = ys__n47373 & new_n44172_;
  assign new_n44298_ = ys__n47232 & ~new_n44176_;
  assign new_n44299_ = ~new_n44297_ & ~new_n44298_;
  assign ys__n31470 = ~new_n44179_ & ~new_n44299_;
  assign new_n44301_ = ys__n47374 & new_n44172_;
  assign new_n44302_ = ys__n47233 & ~new_n44176_;
  assign new_n44303_ = ~new_n44301_ & ~new_n44302_;
  assign ys__n31471 = ~new_n44179_ & ~new_n44303_;
  assign new_n44305_ = ys__n47375 & new_n44172_;
  assign new_n44306_ = ys__n18762 & ~new_n44176_;
  assign new_n44307_ = ~new_n44305_ & ~new_n44306_;
  assign ys__n31472 = ~new_n44179_ & ~new_n44307_;
  assign new_n44309_ = ys__n47376 & new_n44172_;
  assign new_n44310_ = ys__n18750 & ~new_n44176_;
  assign new_n44311_ = ~new_n44309_ & ~new_n44310_;
  assign ys__n31473 = ~new_n44179_ & ~new_n44311_;
  assign new_n44313_ = ys__n47377 & new_n44172_;
  assign new_n44314_ = ys__n18753 & ~new_n44176_;
  assign new_n44315_ = ~new_n44313_ & ~new_n44314_;
  assign ys__n31474 = ~new_n44179_ & ~new_n44315_;
  assign new_n44317_ = ys__n832 & new_n13240_;
  assign new_n44318_ = ys__n47378 & new_n44317_;
  assign new_n44319_ = ~ys__n834 & ~new_n13240_;
  assign new_n44320_ = ~ys__n832 & new_n13240_;
  assign new_n44321_ = ~new_n44319_ & ~new_n44320_;
  assign new_n44322_ = ys__n47202 & ~new_n44321_;
  assign new_n44323_ = ~new_n44318_ & ~new_n44322_;
  assign new_n44324_ = ~new_n44317_ & new_n44321_;
  assign ys__n31475 = ~new_n44323_ & ~new_n44324_;
  assign new_n44326_ = ys__n47379 & new_n44317_;
  assign new_n44327_ = ys__n47203 & ~new_n44321_;
  assign new_n44328_ = ~new_n44326_ & ~new_n44327_;
  assign ys__n31476 = ~new_n44324_ & ~new_n44328_;
  assign new_n44330_ = ys__n47380 & new_n44317_;
  assign new_n44331_ = ys__n47204 & ~new_n44321_;
  assign new_n44332_ = ~new_n44330_ & ~new_n44331_;
  assign ys__n31477 = ~new_n44324_ & ~new_n44332_;
  assign new_n44334_ = ys__n47381 & new_n44317_;
  assign new_n44335_ = ys__n47205 & ~new_n44321_;
  assign new_n44336_ = ~new_n44334_ & ~new_n44335_;
  assign ys__n31478 = ~new_n44324_ & ~new_n44336_;
  assign new_n44338_ = ys__n47382 & new_n44317_;
  assign new_n44339_ = ys__n47206 & ~new_n44321_;
  assign new_n44340_ = ~new_n44338_ & ~new_n44339_;
  assign ys__n31479 = ~new_n44324_ & ~new_n44340_;
  assign new_n44342_ = ys__n47383 & new_n44317_;
  assign new_n44343_ = ys__n47207 & ~new_n44321_;
  assign new_n44344_ = ~new_n44342_ & ~new_n44343_;
  assign ys__n31480 = ~new_n44324_ & ~new_n44344_;
  assign new_n44346_ = ys__n47384 & new_n44317_;
  assign new_n44347_ = ys__n47208 & ~new_n44321_;
  assign new_n44348_ = ~new_n44346_ & ~new_n44347_;
  assign ys__n31481 = ~new_n44324_ & ~new_n44348_;
  assign new_n44350_ = ys__n47385 & new_n44317_;
  assign new_n44351_ = ys__n47209 & ~new_n44321_;
  assign new_n44352_ = ~new_n44350_ & ~new_n44351_;
  assign ys__n31482 = ~new_n44324_ & ~new_n44352_;
  assign new_n44354_ = ys__n47386 & new_n44317_;
  assign new_n44355_ = ys__n47210 & ~new_n44321_;
  assign new_n44356_ = ~new_n44354_ & ~new_n44355_;
  assign ys__n31483 = ~new_n44324_ & ~new_n44356_;
  assign new_n44358_ = ys__n47387 & new_n44317_;
  assign new_n44359_ = ys__n47211 & ~new_n44321_;
  assign new_n44360_ = ~new_n44358_ & ~new_n44359_;
  assign ys__n31484 = ~new_n44324_ & ~new_n44360_;
  assign new_n44362_ = ys__n47388 & new_n44317_;
  assign new_n44363_ = ys__n47212 & ~new_n44321_;
  assign new_n44364_ = ~new_n44362_ & ~new_n44363_;
  assign ys__n31485 = ~new_n44324_ & ~new_n44364_;
  assign new_n44366_ = ys__n47389 & new_n44317_;
  assign new_n44367_ = ys__n47213 & ~new_n44321_;
  assign new_n44368_ = ~new_n44366_ & ~new_n44367_;
  assign ys__n31486 = ~new_n44324_ & ~new_n44368_;
  assign new_n44370_ = ys__n47390 & new_n44317_;
  assign new_n44371_ = ys__n47214 & ~new_n44321_;
  assign new_n44372_ = ~new_n44370_ & ~new_n44371_;
  assign ys__n31487 = ~new_n44324_ & ~new_n44372_;
  assign new_n44374_ = ys__n47391 & new_n44317_;
  assign new_n44375_ = ys__n47215 & ~new_n44321_;
  assign new_n44376_ = ~new_n44374_ & ~new_n44375_;
  assign ys__n31488 = ~new_n44324_ & ~new_n44376_;
  assign new_n44378_ = ys__n47392 & new_n44317_;
  assign new_n44379_ = ys__n47216 & ~new_n44321_;
  assign new_n44380_ = ~new_n44378_ & ~new_n44379_;
  assign ys__n31489 = ~new_n44324_ & ~new_n44380_;
  assign new_n44382_ = ys__n47393 & new_n44317_;
  assign new_n44383_ = ys__n47217 & ~new_n44321_;
  assign new_n44384_ = ~new_n44382_ & ~new_n44383_;
  assign ys__n31490 = ~new_n44324_ & ~new_n44384_;
  assign new_n44386_ = ys__n47394 & new_n44317_;
  assign new_n44387_ = ys__n47218 & ~new_n44321_;
  assign new_n44388_ = ~new_n44386_ & ~new_n44387_;
  assign ys__n31491 = ~new_n44324_ & ~new_n44388_;
  assign new_n44390_ = ys__n47395 & new_n44317_;
  assign new_n44391_ = ys__n47219 & ~new_n44321_;
  assign new_n44392_ = ~new_n44390_ & ~new_n44391_;
  assign ys__n31492 = ~new_n44324_ & ~new_n44392_;
  assign new_n44394_ = ys__n47396 & new_n44317_;
  assign new_n44395_ = ys__n47220 & ~new_n44321_;
  assign new_n44396_ = ~new_n44394_ & ~new_n44395_;
  assign ys__n31493 = ~new_n44324_ & ~new_n44396_;
  assign new_n44398_ = ys__n47397 & new_n44317_;
  assign new_n44399_ = ys__n47221 & ~new_n44321_;
  assign new_n44400_ = ~new_n44398_ & ~new_n44399_;
  assign ys__n31494 = ~new_n44324_ & ~new_n44400_;
  assign new_n44402_ = ys__n47398 & new_n44317_;
  assign new_n44403_ = ys__n47222 & ~new_n44321_;
  assign new_n44404_ = ~new_n44402_ & ~new_n44403_;
  assign ys__n31495 = ~new_n44324_ & ~new_n44404_;
  assign new_n44406_ = ys__n47399 & new_n44317_;
  assign new_n44407_ = ys__n47223 & ~new_n44321_;
  assign new_n44408_ = ~new_n44406_ & ~new_n44407_;
  assign ys__n31496 = ~new_n44324_ & ~new_n44408_;
  assign new_n44410_ = ys__n47400 & new_n44317_;
  assign new_n44411_ = ys__n47224 & ~new_n44321_;
  assign new_n44412_ = ~new_n44410_ & ~new_n44411_;
  assign ys__n31497 = ~new_n44324_ & ~new_n44412_;
  assign new_n44414_ = ys__n47401 & new_n44317_;
  assign new_n44415_ = ys__n47225 & ~new_n44321_;
  assign new_n44416_ = ~new_n44414_ & ~new_n44415_;
  assign ys__n31498 = ~new_n44324_ & ~new_n44416_;
  assign new_n44418_ = ys__n47402 & new_n44317_;
  assign new_n44419_ = ys__n47226 & ~new_n44321_;
  assign new_n44420_ = ~new_n44418_ & ~new_n44419_;
  assign ys__n31499 = ~new_n44324_ & ~new_n44420_;
  assign new_n44422_ = ys__n47403 & new_n44317_;
  assign new_n44423_ = ys__n47227 & ~new_n44321_;
  assign new_n44424_ = ~new_n44422_ & ~new_n44423_;
  assign ys__n31500 = ~new_n44324_ & ~new_n44424_;
  assign new_n44426_ = ys__n47404 & new_n44317_;
  assign new_n44427_ = ys__n47228 & ~new_n44321_;
  assign new_n44428_ = ~new_n44426_ & ~new_n44427_;
  assign ys__n31501 = ~new_n44324_ & ~new_n44428_;
  assign new_n44430_ = ys__n47405 & new_n44317_;
  assign new_n44431_ = ys__n47229 & ~new_n44321_;
  assign new_n44432_ = ~new_n44430_ & ~new_n44431_;
  assign ys__n31502 = ~new_n44324_ & ~new_n44432_;
  assign new_n44434_ = ys__n47406 & new_n44317_;
  assign new_n44435_ = ys__n47230 & ~new_n44321_;
  assign new_n44436_ = ~new_n44434_ & ~new_n44435_;
  assign ys__n31503 = ~new_n44324_ & ~new_n44436_;
  assign new_n44438_ = ys__n47407 & new_n44317_;
  assign new_n44439_ = ys__n47231 & ~new_n44321_;
  assign new_n44440_ = ~new_n44438_ & ~new_n44439_;
  assign ys__n31504 = ~new_n44324_ & ~new_n44440_;
  assign new_n44442_ = ys__n47408 & new_n44317_;
  assign new_n44443_ = ys__n47232 & ~new_n44321_;
  assign new_n44444_ = ~new_n44442_ & ~new_n44443_;
  assign ys__n31505 = ~new_n44324_ & ~new_n44444_;
  assign new_n44446_ = ys__n47409 & new_n44317_;
  assign new_n44447_ = ys__n47233 & ~new_n44321_;
  assign new_n44448_ = ~new_n44446_ & ~new_n44447_;
  assign ys__n31506 = ~new_n44324_ & ~new_n44448_;
  assign new_n44450_ = ys__n47410 & new_n44317_;
  assign new_n44451_ = ys__n18762 & ~new_n44321_;
  assign new_n44452_ = ~new_n44450_ & ~new_n44451_;
  assign ys__n31507 = ~new_n44324_ & ~new_n44452_;
  assign new_n44454_ = ys__n47411 & new_n44317_;
  assign new_n44455_ = ys__n18750 & ~new_n44321_;
  assign new_n44456_ = ~new_n44454_ & ~new_n44455_;
  assign ys__n31508 = ~new_n44324_ & ~new_n44456_;
  assign new_n44458_ = ys__n47412 & new_n44317_;
  assign new_n44459_ = ys__n18753 & ~new_n44321_;
  assign new_n44460_ = ~new_n44458_ & ~new_n44459_;
  assign ys__n31509 = ~new_n44324_ & ~new_n44460_;
  assign new_n44462_ = ys__n834 & new_n13240_;
  assign new_n44463_ = ys__n47413 & new_n44462_;
  assign new_n44464_ = ~ys__n836 & ~new_n13240_;
  assign new_n44465_ = ~ys__n834 & new_n13240_;
  assign new_n44466_ = ~new_n44464_ & ~new_n44465_;
  assign new_n44467_ = ys__n47202 & ~new_n44466_;
  assign new_n44468_ = ~new_n44463_ & ~new_n44467_;
  assign new_n44469_ = ~new_n44462_ & new_n44466_;
  assign ys__n31510 = ~new_n44468_ & ~new_n44469_;
  assign new_n44471_ = ys__n47414 & new_n44462_;
  assign new_n44472_ = ys__n47203 & ~new_n44466_;
  assign new_n44473_ = ~new_n44471_ & ~new_n44472_;
  assign ys__n31511 = ~new_n44469_ & ~new_n44473_;
  assign new_n44475_ = ys__n47415 & new_n44462_;
  assign new_n44476_ = ys__n47204 & ~new_n44466_;
  assign new_n44477_ = ~new_n44475_ & ~new_n44476_;
  assign ys__n31512 = ~new_n44469_ & ~new_n44477_;
  assign new_n44479_ = ys__n47416 & new_n44462_;
  assign new_n44480_ = ys__n47205 & ~new_n44466_;
  assign new_n44481_ = ~new_n44479_ & ~new_n44480_;
  assign ys__n31513 = ~new_n44469_ & ~new_n44481_;
  assign new_n44483_ = ys__n47417 & new_n44462_;
  assign new_n44484_ = ys__n47206 & ~new_n44466_;
  assign new_n44485_ = ~new_n44483_ & ~new_n44484_;
  assign ys__n31514 = ~new_n44469_ & ~new_n44485_;
  assign new_n44487_ = ys__n47418 & new_n44462_;
  assign new_n44488_ = ys__n47207 & ~new_n44466_;
  assign new_n44489_ = ~new_n44487_ & ~new_n44488_;
  assign ys__n31515 = ~new_n44469_ & ~new_n44489_;
  assign new_n44491_ = ys__n47419 & new_n44462_;
  assign new_n44492_ = ys__n47208 & ~new_n44466_;
  assign new_n44493_ = ~new_n44491_ & ~new_n44492_;
  assign ys__n31516 = ~new_n44469_ & ~new_n44493_;
  assign new_n44495_ = ys__n47420 & new_n44462_;
  assign new_n44496_ = ys__n47209 & ~new_n44466_;
  assign new_n44497_ = ~new_n44495_ & ~new_n44496_;
  assign ys__n31517 = ~new_n44469_ & ~new_n44497_;
  assign new_n44499_ = ys__n47421 & new_n44462_;
  assign new_n44500_ = ys__n47210 & ~new_n44466_;
  assign new_n44501_ = ~new_n44499_ & ~new_n44500_;
  assign ys__n31518 = ~new_n44469_ & ~new_n44501_;
  assign new_n44503_ = ys__n47422 & new_n44462_;
  assign new_n44504_ = ys__n47211 & ~new_n44466_;
  assign new_n44505_ = ~new_n44503_ & ~new_n44504_;
  assign ys__n31519 = ~new_n44469_ & ~new_n44505_;
  assign new_n44507_ = ys__n47423 & new_n44462_;
  assign new_n44508_ = ys__n47212 & ~new_n44466_;
  assign new_n44509_ = ~new_n44507_ & ~new_n44508_;
  assign ys__n31520 = ~new_n44469_ & ~new_n44509_;
  assign new_n44511_ = ys__n47424 & new_n44462_;
  assign new_n44512_ = ys__n47213 & ~new_n44466_;
  assign new_n44513_ = ~new_n44511_ & ~new_n44512_;
  assign ys__n31521 = ~new_n44469_ & ~new_n44513_;
  assign new_n44515_ = ys__n47425 & new_n44462_;
  assign new_n44516_ = ys__n47214 & ~new_n44466_;
  assign new_n44517_ = ~new_n44515_ & ~new_n44516_;
  assign ys__n31522 = ~new_n44469_ & ~new_n44517_;
  assign new_n44519_ = ys__n47426 & new_n44462_;
  assign new_n44520_ = ys__n47215 & ~new_n44466_;
  assign new_n44521_ = ~new_n44519_ & ~new_n44520_;
  assign ys__n31523 = ~new_n44469_ & ~new_n44521_;
  assign new_n44523_ = ys__n47427 & new_n44462_;
  assign new_n44524_ = ys__n47216 & ~new_n44466_;
  assign new_n44525_ = ~new_n44523_ & ~new_n44524_;
  assign ys__n31524 = ~new_n44469_ & ~new_n44525_;
  assign new_n44527_ = ys__n47428 & new_n44462_;
  assign new_n44528_ = ys__n47217 & ~new_n44466_;
  assign new_n44529_ = ~new_n44527_ & ~new_n44528_;
  assign ys__n31525 = ~new_n44469_ & ~new_n44529_;
  assign new_n44531_ = ys__n47429 & new_n44462_;
  assign new_n44532_ = ys__n47218 & ~new_n44466_;
  assign new_n44533_ = ~new_n44531_ & ~new_n44532_;
  assign ys__n31526 = ~new_n44469_ & ~new_n44533_;
  assign new_n44535_ = ys__n47430 & new_n44462_;
  assign new_n44536_ = ys__n47219 & ~new_n44466_;
  assign new_n44537_ = ~new_n44535_ & ~new_n44536_;
  assign ys__n31527 = ~new_n44469_ & ~new_n44537_;
  assign new_n44539_ = ys__n47431 & new_n44462_;
  assign new_n44540_ = ys__n47220 & ~new_n44466_;
  assign new_n44541_ = ~new_n44539_ & ~new_n44540_;
  assign ys__n31528 = ~new_n44469_ & ~new_n44541_;
  assign new_n44543_ = ys__n47432 & new_n44462_;
  assign new_n44544_ = ys__n47221 & ~new_n44466_;
  assign new_n44545_ = ~new_n44543_ & ~new_n44544_;
  assign ys__n31529 = ~new_n44469_ & ~new_n44545_;
  assign new_n44547_ = ys__n47433 & new_n44462_;
  assign new_n44548_ = ys__n47222 & ~new_n44466_;
  assign new_n44549_ = ~new_n44547_ & ~new_n44548_;
  assign ys__n31530 = ~new_n44469_ & ~new_n44549_;
  assign new_n44551_ = ys__n47434 & new_n44462_;
  assign new_n44552_ = ys__n47223 & ~new_n44466_;
  assign new_n44553_ = ~new_n44551_ & ~new_n44552_;
  assign ys__n31531 = ~new_n44469_ & ~new_n44553_;
  assign new_n44555_ = ys__n47435 & new_n44462_;
  assign new_n44556_ = ys__n47224 & ~new_n44466_;
  assign new_n44557_ = ~new_n44555_ & ~new_n44556_;
  assign ys__n31532 = ~new_n44469_ & ~new_n44557_;
  assign new_n44559_ = ys__n47436 & new_n44462_;
  assign new_n44560_ = ys__n47225 & ~new_n44466_;
  assign new_n44561_ = ~new_n44559_ & ~new_n44560_;
  assign ys__n31533 = ~new_n44469_ & ~new_n44561_;
  assign new_n44563_ = ys__n47437 & new_n44462_;
  assign new_n44564_ = ys__n47226 & ~new_n44466_;
  assign new_n44565_ = ~new_n44563_ & ~new_n44564_;
  assign ys__n31534 = ~new_n44469_ & ~new_n44565_;
  assign new_n44567_ = ys__n47438 & new_n44462_;
  assign new_n44568_ = ys__n47227 & ~new_n44466_;
  assign new_n44569_ = ~new_n44567_ & ~new_n44568_;
  assign ys__n31535 = ~new_n44469_ & ~new_n44569_;
  assign new_n44571_ = ys__n47439 & new_n44462_;
  assign new_n44572_ = ys__n47228 & ~new_n44466_;
  assign new_n44573_ = ~new_n44571_ & ~new_n44572_;
  assign ys__n31536 = ~new_n44469_ & ~new_n44573_;
  assign new_n44575_ = ys__n47440 & new_n44462_;
  assign new_n44576_ = ys__n47229 & ~new_n44466_;
  assign new_n44577_ = ~new_n44575_ & ~new_n44576_;
  assign ys__n31537 = ~new_n44469_ & ~new_n44577_;
  assign new_n44579_ = ys__n47441 & new_n44462_;
  assign new_n44580_ = ys__n47230 & ~new_n44466_;
  assign new_n44581_ = ~new_n44579_ & ~new_n44580_;
  assign ys__n31538 = ~new_n44469_ & ~new_n44581_;
  assign new_n44583_ = ys__n47442 & new_n44462_;
  assign new_n44584_ = ys__n47231 & ~new_n44466_;
  assign new_n44585_ = ~new_n44583_ & ~new_n44584_;
  assign ys__n31539 = ~new_n44469_ & ~new_n44585_;
  assign new_n44587_ = ys__n47443 & new_n44462_;
  assign new_n44588_ = ys__n47232 & ~new_n44466_;
  assign new_n44589_ = ~new_n44587_ & ~new_n44588_;
  assign ys__n31540 = ~new_n44469_ & ~new_n44589_;
  assign new_n44591_ = ys__n47444 & new_n44462_;
  assign new_n44592_ = ys__n47233 & ~new_n44466_;
  assign new_n44593_ = ~new_n44591_ & ~new_n44592_;
  assign ys__n31541 = ~new_n44469_ & ~new_n44593_;
  assign new_n44595_ = ys__n47445 & new_n44462_;
  assign new_n44596_ = ys__n18762 & ~new_n44466_;
  assign new_n44597_ = ~new_n44595_ & ~new_n44596_;
  assign ys__n31542 = ~new_n44469_ & ~new_n44597_;
  assign new_n44599_ = ys__n47446 & new_n44462_;
  assign new_n44600_ = ys__n18750 & ~new_n44466_;
  assign new_n44601_ = ~new_n44599_ & ~new_n44600_;
  assign ys__n31543 = ~new_n44469_ & ~new_n44601_;
  assign new_n44603_ = ys__n47447 & new_n44462_;
  assign new_n44604_ = ys__n18753 & ~new_n44466_;
  assign new_n44605_ = ~new_n44603_ & ~new_n44604_;
  assign ys__n31544 = ~new_n44469_ & ~new_n44605_;
  assign new_n44607_ = ys__n35057 & ~ys__n35059;
  assign new_n44608_ = ~ys__n488 & ys__n490;
  assign new_n44609_ = ~new_n44607_ & new_n44608_;
  assign new_n44610_ = ~ys__n35057 & ~ys__n35059;
  assign new_n44611_ = ~ys__n488 & ~ys__n490;
  assign new_n44612_ = ~new_n44610_ & new_n44611_;
  assign new_n44613_ = ~new_n44609_ & ~new_n44612_;
  assign new_n44614_ = ys__n488 & ys__n490;
  assign new_n44615_ = ~new_n44608_ & ~new_n44614_;
  assign new_n44616_ = ys__n488 & ~ys__n490;
  assign new_n44617_ = ~new_n44611_ & ~new_n44616_;
  assign new_n44618_ = new_n44615_ & new_n44617_;
  assign ys__n31559 = ~new_n44613_ & ~new_n44618_;
  assign new_n44620_ = ~ys__n35057 & ys__n35059;
  assign new_n44621_ = new_n44616_ & ~new_n44620_;
  assign new_n44622_ = ~new_n44609_ & ~new_n44621_;
  assign ys__n31560 = ~new_n44618_ & ~new_n44622_;
  assign new_n44624_ = ~new_n44610_ & ~new_n44620_;
  assign new_n44625_ = new_n44611_ & ~new_n44624_;
  assign new_n44626_ = ys__n35057 & ys__n35059;
  assign new_n44627_ = new_n44608_ & new_n44626_;
  assign new_n44628_ = new_n44607_ & new_n44616_;
  assign new_n44629_ = ~new_n44627_ & ~new_n44628_;
  assign new_n44630_ = ~new_n44625_ & new_n44629_;
  assign ys__n31562 = ~new_n44618_ & ~new_n44630_;
  assign new_n44632_ = new_n44616_ & new_n44620_;
  assign ys__n31564 = ~new_n44618_ & new_n44632_;
  assign new_n44634_ = new_n44607_ & new_n44608_;
  assign ys__n31567 = ~new_n44618_ & new_n44634_;
  assign new_n44636_ = ~new_n44611_ & ~new_n44614_;
  assign new_n44637_ = ~new_n44608_ & ~new_n44616_;
  assign new_n44638_ = new_n44636_ & new_n44637_;
  assign new_n44639_ = new_n44626_ & ~new_n44636_;
  assign ys__n31571 = ~new_n44638_ & new_n44639_;
  assign new_n44641_ = ys__n830 & new_n13240_;
  assign new_n44642_ = ys__n47449 & new_n44641_;
  assign new_n44643_ = ~ys__n832 & ~new_n13240_;
  assign new_n44644_ = ~ys__n830 & new_n13240_;
  assign new_n44645_ = ~new_n44643_ & ~new_n44644_;
  assign new_n44646_ = ys__n47202 & ~new_n44645_;
  assign new_n44647_ = ~new_n44642_ & ~new_n44646_;
  assign new_n44648_ = ~new_n44641_ & new_n44645_;
  assign ys__n31740 = ~new_n44647_ & ~new_n44648_;
  assign new_n44650_ = ys__n47450 & new_n44641_;
  assign new_n44651_ = ys__n47203 & ~new_n44645_;
  assign new_n44652_ = ~new_n44650_ & ~new_n44651_;
  assign ys__n31741 = ~new_n44648_ & ~new_n44652_;
  assign new_n44654_ = ys__n47451 & new_n44641_;
  assign new_n44655_ = ys__n47204 & ~new_n44645_;
  assign new_n44656_ = ~new_n44654_ & ~new_n44655_;
  assign ys__n31742 = ~new_n44648_ & ~new_n44656_;
  assign new_n44658_ = ys__n47452 & new_n44641_;
  assign new_n44659_ = ys__n47205 & ~new_n44645_;
  assign new_n44660_ = ~new_n44658_ & ~new_n44659_;
  assign ys__n31743 = ~new_n44648_ & ~new_n44660_;
  assign new_n44662_ = ys__n47453 & new_n44641_;
  assign new_n44663_ = ys__n47206 & ~new_n44645_;
  assign new_n44664_ = ~new_n44662_ & ~new_n44663_;
  assign ys__n31744 = ~new_n44648_ & ~new_n44664_;
  assign new_n44666_ = ys__n47454 & new_n44641_;
  assign new_n44667_ = ys__n47207 & ~new_n44645_;
  assign new_n44668_ = ~new_n44666_ & ~new_n44667_;
  assign ys__n31745 = ~new_n44648_ & ~new_n44668_;
  assign new_n44670_ = ys__n47455 & new_n44641_;
  assign new_n44671_ = ys__n47208 & ~new_n44645_;
  assign new_n44672_ = ~new_n44670_ & ~new_n44671_;
  assign ys__n31746 = ~new_n44648_ & ~new_n44672_;
  assign new_n44674_ = ys__n47456 & new_n44641_;
  assign new_n44675_ = ys__n47209 & ~new_n44645_;
  assign new_n44676_ = ~new_n44674_ & ~new_n44675_;
  assign ys__n31747 = ~new_n44648_ & ~new_n44676_;
  assign new_n44678_ = ys__n47457 & new_n44641_;
  assign new_n44679_ = ys__n47210 & ~new_n44645_;
  assign new_n44680_ = ~new_n44678_ & ~new_n44679_;
  assign ys__n31748 = ~new_n44648_ & ~new_n44680_;
  assign new_n44682_ = ys__n47458 & new_n44641_;
  assign new_n44683_ = ys__n47211 & ~new_n44645_;
  assign new_n44684_ = ~new_n44682_ & ~new_n44683_;
  assign ys__n31749 = ~new_n44648_ & ~new_n44684_;
  assign new_n44686_ = ys__n47459 & new_n44641_;
  assign new_n44687_ = ys__n47212 & ~new_n44645_;
  assign new_n44688_ = ~new_n44686_ & ~new_n44687_;
  assign ys__n31750 = ~new_n44648_ & ~new_n44688_;
  assign new_n44690_ = ys__n47460 & new_n44641_;
  assign new_n44691_ = ys__n47213 & ~new_n44645_;
  assign new_n44692_ = ~new_n44690_ & ~new_n44691_;
  assign ys__n31751 = ~new_n44648_ & ~new_n44692_;
  assign new_n44694_ = ys__n47461 & new_n44641_;
  assign new_n44695_ = ys__n47214 & ~new_n44645_;
  assign new_n44696_ = ~new_n44694_ & ~new_n44695_;
  assign ys__n31752 = ~new_n44648_ & ~new_n44696_;
  assign new_n44698_ = ys__n47462 & new_n44641_;
  assign new_n44699_ = ys__n47215 & ~new_n44645_;
  assign new_n44700_ = ~new_n44698_ & ~new_n44699_;
  assign ys__n31753 = ~new_n44648_ & ~new_n44700_;
  assign new_n44702_ = ys__n47463 & new_n44641_;
  assign new_n44703_ = ys__n47216 & ~new_n44645_;
  assign new_n44704_ = ~new_n44702_ & ~new_n44703_;
  assign ys__n31754 = ~new_n44648_ & ~new_n44704_;
  assign new_n44706_ = ys__n47464 & new_n44641_;
  assign new_n44707_ = ys__n47217 & ~new_n44645_;
  assign new_n44708_ = ~new_n44706_ & ~new_n44707_;
  assign ys__n31755 = ~new_n44648_ & ~new_n44708_;
  assign new_n44710_ = ys__n47465 & new_n44641_;
  assign new_n44711_ = ys__n47218 & ~new_n44645_;
  assign new_n44712_ = ~new_n44710_ & ~new_n44711_;
  assign ys__n31756 = ~new_n44648_ & ~new_n44712_;
  assign new_n44714_ = ys__n47466 & new_n44641_;
  assign new_n44715_ = ys__n47219 & ~new_n44645_;
  assign new_n44716_ = ~new_n44714_ & ~new_n44715_;
  assign ys__n31757 = ~new_n44648_ & ~new_n44716_;
  assign new_n44718_ = ys__n47467 & new_n44641_;
  assign new_n44719_ = ys__n47220 & ~new_n44645_;
  assign new_n44720_ = ~new_n44718_ & ~new_n44719_;
  assign ys__n31758 = ~new_n44648_ & ~new_n44720_;
  assign new_n44722_ = ys__n47468 & new_n44641_;
  assign new_n44723_ = ys__n47221 & ~new_n44645_;
  assign new_n44724_ = ~new_n44722_ & ~new_n44723_;
  assign ys__n31759 = ~new_n44648_ & ~new_n44724_;
  assign new_n44726_ = ys__n47469 & new_n44641_;
  assign new_n44727_ = ys__n47222 & ~new_n44645_;
  assign new_n44728_ = ~new_n44726_ & ~new_n44727_;
  assign ys__n31760 = ~new_n44648_ & ~new_n44728_;
  assign new_n44730_ = ys__n47470 & new_n44641_;
  assign new_n44731_ = ys__n47223 & ~new_n44645_;
  assign new_n44732_ = ~new_n44730_ & ~new_n44731_;
  assign ys__n31761 = ~new_n44648_ & ~new_n44732_;
  assign new_n44734_ = ys__n47471 & new_n44641_;
  assign new_n44735_ = ys__n47224 & ~new_n44645_;
  assign new_n44736_ = ~new_n44734_ & ~new_n44735_;
  assign ys__n31762 = ~new_n44648_ & ~new_n44736_;
  assign new_n44738_ = ys__n47472 & new_n44641_;
  assign new_n44739_ = ys__n47225 & ~new_n44645_;
  assign new_n44740_ = ~new_n44738_ & ~new_n44739_;
  assign ys__n31763 = ~new_n44648_ & ~new_n44740_;
  assign new_n44742_ = ys__n47473 & new_n44641_;
  assign new_n44743_ = ys__n47226 & ~new_n44645_;
  assign new_n44744_ = ~new_n44742_ & ~new_n44743_;
  assign ys__n31764 = ~new_n44648_ & ~new_n44744_;
  assign new_n44746_ = ys__n47474 & new_n44641_;
  assign new_n44747_ = ys__n47227 & ~new_n44645_;
  assign new_n44748_ = ~new_n44746_ & ~new_n44747_;
  assign ys__n31765 = ~new_n44648_ & ~new_n44748_;
  assign new_n44750_ = ys__n47475 & new_n44641_;
  assign new_n44751_ = ys__n47228 & ~new_n44645_;
  assign new_n44752_ = ~new_n44750_ & ~new_n44751_;
  assign ys__n31766 = ~new_n44648_ & ~new_n44752_;
  assign new_n44754_ = ys__n47476 & new_n44641_;
  assign new_n44755_ = ys__n47229 & ~new_n44645_;
  assign new_n44756_ = ~new_n44754_ & ~new_n44755_;
  assign ys__n31767 = ~new_n44648_ & ~new_n44756_;
  assign new_n44758_ = ys__n47477 & new_n44641_;
  assign new_n44759_ = ys__n47230 & ~new_n44645_;
  assign new_n44760_ = ~new_n44758_ & ~new_n44759_;
  assign ys__n31768 = ~new_n44648_ & ~new_n44760_;
  assign new_n44762_ = ys__n47478 & new_n44641_;
  assign new_n44763_ = ys__n47231 & ~new_n44645_;
  assign new_n44764_ = ~new_n44762_ & ~new_n44763_;
  assign ys__n31769 = ~new_n44648_ & ~new_n44764_;
  assign new_n44766_ = ys__n47479 & new_n44641_;
  assign new_n44767_ = ys__n47232 & ~new_n44645_;
  assign new_n44768_ = ~new_n44766_ & ~new_n44767_;
  assign ys__n31770 = ~new_n44648_ & ~new_n44768_;
  assign new_n44770_ = ys__n47480 & new_n44641_;
  assign new_n44771_ = ys__n47233 & ~new_n44645_;
  assign new_n44772_ = ~new_n44770_ & ~new_n44771_;
  assign ys__n31771 = ~new_n44648_ & ~new_n44772_;
  assign new_n44774_ = ys__n47481 & new_n44641_;
  assign new_n44775_ = ys__n18762 & ~new_n44645_;
  assign new_n44776_ = ~new_n44774_ & ~new_n44775_;
  assign ys__n31772 = ~new_n44648_ & ~new_n44776_;
  assign new_n44778_ = ys__n47482 & new_n44641_;
  assign new_n44779_ = ys__n18750 & ~new_n44645_;
  assign new_n44780_ = ~new_n44778_ & ~new_n44779_;
  assign ys__n31773 = ~new_n44648_ & ~new_n44780_;
  assign new_n44782_ = ys__n47483 & new_n44641_;
  assign new_n44783_ = ys__n18753 & ~new_n44645_;
  assign new_n44784_ = ~new_n44782_ & ~new_n44783_;
  assign ys__n31774 = ~new_n44648_ & ~new_n44784_;
  assign new_n44786_ = ys__n858 & new_n13240_;
  assign new_n44787_ = ys__n47484 & new_n44786_;
  assign new_n44788_ = ~ys__n830 & ~new_n13240_;
  assign new_n44789_ = ~ys__n858 & new_n13240_;
  assign new_n44790_ = ~new_n44788_ & ~new_n44789_;
  assign new_n44791_ = ys__n47202 & ~new_n44790_;
  assign new_n44792_ = ~new_n44787_ & ~new_n44791_;
  assign new_n44793_ = ~new_n44786_ & new_n44790_;
  assign ys__n31775 = ~new_n44792_ & ~new_n44793_;
  assign new_n44795_ = ys__n47485 & new_n44786_;
  assign new_n44796_ = ys__n47203 & ~new_n44790_;
  assign new_n44797_ = ~new_n44795_ & ~new_n44796_;
  assign ys__n31776 = ~new_n44793_ & ~new_n44797_;
  assign new_n44799_ = ys__n47486 & new_n44786_;
  assign new_n44800_ = ys__n47204 & ~new_n44790_;
  assign new_n44801_ = ~new_n44799_ & ~new_n44800_;
  assign ys__n31777 = ~new_n44793_ & ~new_n44801_;
  assign new_n44803_ = ys__n47487 & new_n44786_;
  assign new_n44804_ = ys__n47205 & ~new_n44790_;
  assign new_n44805_ = ~new_n44803_ & ~new_n44804_;
  assign ys__n31778 = ~new_n44793_ & ~new_n44805_;
  assign new_n44807_ = ys__n47488 & new_n44786_;
  assign new_n44808_ = ys__n47206 & ~new_n44790_;
  assign new_n44809_ = ~new_n44807_ & ~new_n44808_;
  assign ys__n31779 = ~new_n44793_ & ~new_n44809_;
  assign new_n44811_ = ys__n47489 & new_n44786_;
  assign new_n44812_ = ys__n47207 & ~new_n44790_;
  assign new_n44813_ = ~new_n44811_ & ~new_n44812_;
  assign ys__n31780 = ~new_n44793_ & ~new_n44813_;
  assign new_n44815_ = ys__n47490 & new_n44786_;
  assign new_n44816_ = ys__n47208 & ~new_n44790_;
  assign new_n44817_ = ~new_n44815_ & ~new_n44816_;
  assign ys__n31781 = ~new_n44793_ & ~new_n44817_;
  assign new_n44819_ = ys__n47491 & new_n44786_;
  assign new_n44820_ = ys__n47209 & ~new_n44790_;
  assign new_n44821_ = ~new_n44819_ & ~new_n44820_;
  assign ys__n31782 = ~new_n44793_ & ~new_n44821_;
  assign new_n44823_ = ys__n47492 & new_n44786_;
  assign new_n44824_ = ys__n47210 & ~new_n44790_;
  assign new_n44825_ = ~new_n44823_ & ~new_n44824_;
  assign ys__n31783 = ~new_n44793_ & ~new_n44825_;
  assign new_n44827_ = ys__n47493 & new_n44786_;
  assign new_n44828_ = ys__n47211 & ~new_n44790_;
  assign new_n44829_ = ~new_n44827_ & ~new_n44828_;
  assign ys__n31784 = ~new_n44793_ & ~new_n44829_;
  assign new_n44831_ = ys__n47494 & new_n44786_;
  assign new_n44832_ = ys__n47212 & ~new_n44790_;
  assign new_n44833_ = ~new_n44831_ & ~new_n44832_;
  assign ys__n31785 = ~new_n44793_ & ~new_n44833_;
  assign new_n44835_ = ys__n47495 & new_n44786_;
  assign new_n44836_ = ys__n47213 & ~new_n44790_;
  assign new_n44837_ = ~new_n44835_ & ~new_n44836_;
  assign ys__n31786 = ~new_n44793_ & ~new_n44837_;
  assign new_n44839_ = ys__n47496 & new_n44786_;
  assign new_n44840_ = ys__n47214 & ~new_n44790_;
  assign new_n44841_ = ~new_n44839_ & ~new_n44840_;
  assign ys__n31787 = ~new_n44793_ & ~new_n44841_;
  assign new_n44843_ = ys__n47497 & new_n44786_;
  assign new_n44844_ = ys__n47215 & ~new_n44790_;
  assign new_n44845_ = ~new_n44843_ & ~new_n44844_;
  assign ys__n31788 = ~new_n44793_ & ~new_n44845_;
  assign new_n44847_ = ys__n47498 & new_n44786_;
  assign new_n44848_ = ys__n47216 & ~new_n44790_;
  assign new_n44849_ = ~new_n44847_ & ~new_n44848_;
  assign ys__n31789 = ~new_n44793_ & ~new_n44849_;
  assign new_n44851_ = ys__n47499 & new_n44786_;
  assign new_n44852_ = ys__n47217 & ~new_n44790_;
  assign new_n44853_ = ~new_n44851_ & ~new_n44852_;
  assign ys__n31790 = ~new_n44793_ & ~new_n44853_;
  assign new_n44855_ = ys__n47500 & new_n44786_;
  assign new_n44856_ = ys__n47218 & ~new_n44790_;
  assign new_n44857_ = ~new_n44855_ & ~new_n44856_;
  assign ys__n31791 = ~new_n44793_ & ~new_n44857_;
  assign new_n44859_ = ys__n47501 & new_n44786_;
  assign new_n44860_ = ys__n47219 & ~new_n44790_;
  assign new_n44861_ = ~new_n44859_ & ~new_n44860_;
  assign ys__n31792 = ~new_n44793_ & ~new_n44861_;
  assign new_n44863_ = ys__n47502 & new_n44786_;
  assign new_n44864_ = ys__n47220 & ~new_n44790_;
  assign new_n44865_ = ~new_n44863_ & ~new_n44864_;
  assign ys__n31793 = ~new_n44793_ & ~new_n44865_;
  assign new_n44867_ = ys__n47503 & new_n44786_;
  assign new_n44868_ = ys__n47221 & ~new_n44790_;
  assign new_n44869_ = ~new_n44867_ & ~new_n44868_;
  assign ys__n31794 = ~new_n44793_ & ~new_n44869_;
  assign new_n44871_ = ys__n47504 & new_n44786_;
  assign new_n44872_ = ys__n47222 & ~new_n44790_;
  assign new_n44873_ = ~new_n44871_ & ~new_n44872_;
  assign ys__n31795 = ~new_n44793_ & ~new_n44873_;
  assign new_n44875_ = ys__n47505 & new_n44786_;
  assign new_n44876_ = ys__n47223 & ~new_n44790_;
  assign new_n44877_ = ~new_n44875_ & ~new_n44876_;
  assign ys__n31796 = ~new_n44793_ & ~new_n44877_;
  assign new_n44879_ = ys__n47506 & new_n44786_;
  assign new_n44880_ = ys__n47224 & ~new_n44790_;
  assign new_n44881_ = ~new_n44879_ & ~new_n44880_;
  assign ys__n31797 = ~new_n44793_ & ~new_n44881_;
  assign new_n44883_ = ys__n47507 & new_n44786_;
  assign new_n44884_ = ys__n47225 & ~new_n44790_;
  assign new_n44885_ = ~new_n44883_ & ~new_n44884_;
  assign ys__n31798 = ~new_n44793_ & ~new_n44885_;
  assign new_n44887_ = ys__n47508 & new_n44786_;
  assign new_n44888_ = ys__n47226 & ~new_n44790_;
  assign new_n44889_ = ~new_n44887_ & ~new_n44888_;
  assign ys__n31799 = ~new_n44793_ & ~new_n44889_;
  assign new_n44891_ = ys__n47509 & new_n44786_;
  assign new_n44892_ = ys__n47227 & ~new_n44790_;
  assign new_n44893_ = ~new_n44891_ & ~new_n44892_;
  assign ys__n31800 = ~new_n44793_ & ~new_n44893_;
  assign new_n44895_ = ys__n47510 & new_n44786_;
  assign new_n44896_ = ys__n47228 & ~new_n44790_;
  assign new_n44897_ = ~new_n44895_ & ~new_n44896_;
  assign ys__n31801 = ~new_n44793_ & ~new_n44897_;
  assign new_n44899_ = ys__n47511 & new_n44786_;
  assign new_n44900_ = ys__n47229 & ~new_n44790_;
  assign new_n44901_ = ~new_n44899_ & ~new_n44900_;
  assign ys__n31802 = ~new_n44793_ & ~new_n44901_;
  assign new_n44903_ = ys__n47512 & new_n44786_;
  assign new_n44904_ = ys__n47230 & ~new_n44790_;
  assign new_n44905_ = ~new_n44903_ & ~new_n44904_;
  assign ys__n31803 = ~new_n44793_ & ~new_n44905_;
  assign new_n44907_ = ys__n47513 & new_n44786_;
  assign new_n44908_ = ys__n47231 & ~new_n44790_;
  assign new_n44909_ = ~new_n44907_ & ~new_n44908_;
  assign ys__n31804 = ~new_n44793_ & ~new_n44909_;
  assign new_n44911_ = ys__n47514 & new_n44786_;
  assign new_n44912_ = ys__n47232 & ~new_n44790_;
  assign new_n44913_ = ~new_n44911_ & ~new_n44912_;
  assign ys__n31805 = ~new_n44793_ & ~new_n44913_;
  assign new_n44915_ = ys__n47515 & new_n44786_;
  assign new_n44916_ = ys__n47233 & ~new_n44790_;
  assign new_n44917_ = ~new_n44915_ & ~new_n44916_;
  assign ys__n31806 = ~new_n44793_ & ~new_n44917_;
  assign new_n44919_ = ys__n47516 & new_n44786_;
  assign new_n44920_ = ys__n18762 & ~new_n44790_;
  assign new_n44921_ = ~new_n44919_ & ~new_n44920_;
  assign ys__n31807 = ~new_n44793_ & ~new_n44921_;
  assign new_n44923_ = ys__n47517 & new_n44786_;
  assign new_n44924_ = ys__n18750 & ~new_n44790_;
  assign new_n44925_ = ~new_n44923_ & ~new_n44924_;
  assign ys__n31808 = ~new_n44793_ & ~new_n44925_;
  assign new_n44927_ = ys__n47518 & new_n44786_;
  assign new_n44928_ = ys__n18753 & ~new_n44790_;
  assign new_n44929_ = ~new_n44927_ & ~new_n44928_;
  assign ys__n31809 = ~new_n44793_ & ~new_n44929_;
  assign new_n44931_ = ys__n856 & new_n13240_;
  assign new_n44932_ = ys__n47519 & new_n44931_;
  assign new_n44933_ = ~ys__n858 & ~new_n13240_;
  assign new_n44934_ = ~ys__n856 & new_n13240_;
  assign new_n44935_ = ~new_n44933_ & ~new_n44934_;
  assign new_n44936_ = ys__n47202 & ~new_n44935_;
  assign new_n44937_ = ~new_n44932_ & ~new_n44936_;
  assign new_n44938_ = ~new_n44931_ & new_n44935_;
  assign ys__n31810 = ~new_n44937_ & ~new_n44938_;
  assign new_n44940_ = ys__n47520 & new_n44931_;
  assign new_n44941_ = ys__n47203 & ~new_n44935_;
  assign new_n44942_ = ~new_n44940_ & ~new_n44941_;
  assign ys__n31811 = ~new_n44938_ & ~new_n44942_;
  assign new_n44944_ = ys__n47521 & new_n44931_;
  assign new_n44945_ = ys__n47204 & ~new_n44935_;
  assign new_n44946_ = ~new_n44944_ & ~new_n44945_;
  assign ys__n31812 = ~new_n44938_ & ~new_n44946_;
  assign new_n44948_ = ys__n47522 & new_n44931_;
  assign new_n44949_ = ys__n47205 & ~new_n44935_;
  assign new_n44950_ = ~new_n44948_ & ~new_n44949_;
  assign ys__n31813 = ~new_n44938_ & ~new_n44950_;
  assign new_n44952_ = ys__n47523 & new_n44931_;
  assign new_n44953_ = ys__n47206 & ~new_n44935_;
  assign new_n44954_ = ~new_n44952_ & ~new_n44953_;
  assign ys__n31814 = ~new_n44938_ & ~new_n44954_;
  assign new_n44956_ = ys__n47524 & new_n44931_;
  assign new_n44957_ = ys__n47207 & ~new_n44935_;
  assign new_n44958_ = ~new_n44956_ & ~new_n44957_;
  assign ys__n31815 = ~new_n44938_ & ~new_n44958_;
  assign new_n44960_ = ys__n47525 & new_n44931_;
  assign new_n44961_ = ys__n47208 & ~new_n44935_;
  assign new_n44962_ = ~new_n44960_ & ~new_n44961_;
  assign ys__n31816 = ~new_n44938_ & ~new_n44962_;
  assign new_n44964_ = ys__n47526 & new_n44931_;
  assign new_n44965_ = ys__n47209 & ~new_n44935_;
  assign new_n44966_ = ~new_n44964_ & ~new_n44965_;
  assign ys__n31817 = ~new_n44938_ & ~new_n44966_;
  assign new_n44968_ = ys__n47527 & new_n44931_;
  assign new_n44969_ = ys__n47210 & ~new_n44935_;
  assign new_n44970_ = ~new_n44968_ & ~new_n44969_;
  assign ys__n31818 = ~new_n44938_ & ~new_n44970_;
  assign new_n44972_ = ys__n47528 & new_n44931_;
  assign new_n44973_ = ys__n47211 & ~new_n44935_;
  assign new_n44974_ = ~new_n44972_ & ~new_n44973_;
  assign ys__n31819 = ~new_n44938_ & ~new_n44974_;
  assign new_n44976_ = ys__n47529 & new_n44931_;
  assign new_n44977_ = ys__n47212 & ~new_n44935_;
  assign new_n44978_ = ~new_n44976_ & ~new_n44977_;
  assign ys__n31820 = ~new_n44938_ & ~new_n44978_;
  assign new_n44980_ = ys__n47530 & new_n44931_;
  assign new_n44981_ = ys__n47213 & ~new_n44935_;
  assign new_n44982_ = ~new_n44980_ & ~new_n44981_;
  assign ys__n31821 = ~new_n44938_ & ~new_n44982_;
  assign new_n44984_ = ys__n47531 & new_n44931_;
  assign new_n44985_ = ys__n47214 & ~new_n44935_;
  assign new_n44986_ = ~new_n44984_ & ~new_n44985_;
  assign ys__n31822 = ~new_n44938_ & ~new_n44986_;
  assign new_n44988_ = ys__n47532 & new_n44931_;
  assign new_n44989_ = ys__n47215 & ~new_n44935_;
  assign new_n44990_ = ~new_n44988_ & ~new_n44989_;
  assign ys__n31823 = ~new_n44938_ & ~new_n44990_;
  assign new_n44992_ = ys__n47533 & new_n44931_;
  assign new_n44993_ = ys__n47216 & ~new_n44935_;
  assign new_n44994_ = ~new_n44992_ & ~new_n44993_;
  assign ys__n31824 = ~new_n44938_ & ~new_n44994_;
  assign new_n44996_ = ys__n47534 & new_n44931_;
  assign new_n44997_ = ys__n47217 & ~new_n44935_;
  assign new_n44998_ = ~new_n44996_ & ~new_n44997_;
  assign ys__n31825 = ~new_n44938_ & ~new_n44998_;
  assign new_n45000_ = ys__n47535 & new_n44931_;
  assign new_n45001_ = ys__n47218 & ~new_n44935_;
  assign new_n45002_ = ~new_n45000_ & ~new_n45001_;
  assign ys__n31826 = ~new_n44938_ & ~new_n45002_;
  assign new_n45004_ = ys__n47536 & new_n44931_;
  assign new_n45005_ = ys__n47219 & ~new_n44935_;
  assign new_n45006_ = ~new_n45004_ & ~new_n45005_;
  assign ys__n31827 = ~new_n44938_ & ~new_n45006_;
  assign new_n45008_ = ys__n47537 & new_n44931_;
  assign new_n45009_ = ys__n47220 & ~new_n44935_;
  assign new_n45010_ = ~new_n45008_ & ~new_n45009_;
  assign ys__n31828 = ~new_n44938_ & ~new_n45010_;
  assign new_n45012_ = ys__n47538 & new_n44931_;
  assign new_n45013_ = ys__n47221 & ~new_n44935_;
  assign new_n45014_ = ~new_n45012_ & ~new_n45013_;
  assign ys__n31829 = ~new_n44938_ & ~new_n45014_;
  assign new_n45016_ = ys__n47539 & new_n44931_;
  assign new_n45017_ = ys__n47222 & ~new_n44935_;
  assign new_n45018_ = ~new_n45016_ & ~new_n45017_;
  assign ys__n31830 = ~new_n44938_ & ~new_n45018_;
  assign new_n45020_ = ys__n47540 & new_n44931_;
  assign new_n45021_ = ys__n47223 & ~new_n44935_;
  assign new_n45022_ = ~new_n45020_ & ~new_n45021_;
  assign ys__n31831 = ~new_n44938_ & ~new_n45022_;
  assign new_n45024_ = ys__n47541 & new_n44931_;
  assign new_n45025_ = ys__n47224 & ~new_n44935_;
  assign new_n45026_ = ~new_n45024_ & ~new_n45025_;
  assign ys__n31832 = ~new_n44938_ & ~new_n45026_;
  assign new_n45028_ = ys__n47542 & new_n44931_;
  assign new_n45029_ = ys__n47225 & ~new_n44935_;
  assign new_n45030_ = ~new_n45028_ & ~new_n45029_;
  assign ys__n31833 = ~new_n44938_ & ~new_n45030_;
  assign new_n45032_ = ys__n47543 & new_n44931_;
  assign new_n45033_ = ys__n47226 & ~new_n44935_;
  assign new_n45034_ = ~new_n45032_ & ~new_n45033_;
  assign ys__n31834 = ~new_n44938_ & ~new_n45034_;
  assign new_n45036_ = ys__n47544 & new_n44931_;
  assign new_n45037_ = ys__n47227 & ~new_n44935_;
  assign new_n45038_ = ~new_n45036_ & ~new_n45037_;
  assign ys__n31835 = ~new_n44938_ & ~new_n45038_;
  assign new_n45040_ = ys__n47545 & new_n44931_;
  assign new_n45041_ = ys__n47228 & ~new_n44935_;
  assign new_n45042_ = ~new_n45040_ & ~new_n45041_;
  assign ys__n31836 = ~new_n44938_ & ~new_n45042_;
  assign new_n45044_ = ys__n47546 & new_n44931_;
  assign new_n45045_ = ys__n47229 & ~new_n44935_;
  assign new_n45046_ = ~new_n45044_ & ~new_n45045_;
  assign ys__n31837 = ~new_n44938_ & ~new_n45046_;
  assign new_n45048_ = ys__n47547 & new_n44931_;
  assign new_n45049_ = ys__n47230 & ~new_n44935_;
  assign new_n45050_ = ~new_n45048_ & ~new_n45049_;
  assign ys__n31838 = ~new_n44938_ & ~new_n45050_;
  assign new_n45052_ = ys__n47548 & new_n44931_;
  assign new_n45053_ = ys__n47231 & ~new_n44935_;
  assign new_n45054_ = ~new_n45052_ & ~new_n45053_;
  assign ys__n31839 = ~new_n44938_ & ~new_n45054_;
  assign new_n45056_ = ys__n47549 & new_n44931_;
  assign new_n45057_ = ys__n47232 & ~new_n44935_;
  assign new_n45058_ = ~new_n45056_ & ~new_n45057_;
  assign ys__n31840 = ~new_n44938_ & ~new_n45058_;
  assign new_n45060_ = ys__n47550 & new_n44931_;
  assign new_n45061_ = ys__n47233 & ~new_n44935_;
  assign new_n45062_ = ~new_n45060_ & ~new_n45061_;
  assign ys__n31841 = ~new_n44938_ & ~new_n45062_;
  assign new_n45064_ = ys__n47551 & new_n44931_;
  assign new_n45065_ = ys__n18762 & ~new_n44935_;
  assign new_n45066_ = ~new_n45064_ & ~new_n45065_;
  assign ys__n31842 = ~new_n44938_ & ~new_n45066_;
  assign new_n45068_ = ys__n47552 & new_n44931_;
  assign new_n45069_ = ys__n18750 & ~new_n44935_;
  assign new_n45070_ = ~new_n45068_ & ~new_n45069_;
  assign ys__n31843 = ~new_n44938_ & ~new_n45070_;
  assign new_n45072_ = ys__n47553 & new_n44931_;
  assign new_n45073_ = ys__n18753 & ~new_n44935_;
  assign new_n45074_ = ~new_n45072_ & ~new_n45073_;
  assign ys__n31844 = ~new_n44938_ & ~new_n45074_;
  assign new_n45076_ = ys__n854 & new_n13240_;
  assign new_n45077_ = ys__n47554 & new_n45076_;
  assign new_n45078_ = ~ys__n856 & ~new_n13240_;
  assign new_n45079_ = ~ys__n854 & new_n13240_;
  assign new_n45080_ = ~new_n45078_ & ~new_n45079_;
  assign new_n45081_ = ys__n47202 & ~new_n45080_;
  assign new_n45082_ = ~new_n45077_ & ~new_n45081_;
  assign new_n45083_ = ~new_n45076_ & new_n45080_;
  assign ys__n31845 = ~new_n45082_ & ~new_n45083_;
  assign new_n45085_ = ys__n47555 & new_n45076_;
  assign new_n45086_ = ys__n47203 & ~new_n45080_;
  assign new_n45087_ = ~new_n45085_ & ~new_n45086_;
  assign ys__n31846 = ~new_n45083_ & ~new_n45087_;
  assign new_n45089_ = ys__n47556 & new_n45076_;
  assign new_n45090_ = ys__n47204 & ~new_n45080_;
  assign new_n45091_ = ~new_n45089_ & ~new_n45090_;
  assign ys__n31847 = ~new_n45083_ & ~new_n45091_;
  assign new_n45093_ = ys__n47557 & new_n45076_;
  assign new_n45094_ = ys__n47205 & ~new_n45080_;
  assign new_n45095_ = ~new_n45093_ & ~new_n45094_;
  assign ys__n31848 = ~new_n45083_ & ~new_n45095_;
  assign new_n45097_ = ys__n47558 & new_n45076_;
  assign new_n45098_ = ys__n47206 & ~new_n45080_;
  assign new_n45099_ = ~new_n45097_ & ~new_n45098_;
  assign ys__n31849 = ~new_n45083_ & ~new_n45099_;
  assign new_n45101_ = ys__n47559 & new_n45076_;
  assign new_n45102_ = ys__n47207 & ~new_n45080_;
  assign new_n45103_ = ~new_n45101_ & ~new_n45102_;
  assign ys__n31850 = ~new_n45083_ & ~new_n45103_;
  assign new_n45105_ = ys__n47560 & new_n45076_;
  assign new_n45106_ = ys__n47208 & ~new_n45080_;
  assign new_n45107_ = ~new_n45105_ & ~new_n45106_;
  assign ys__n31851 = ~new_n45083_ & ~new_n45107_;
  assign new_n45109_ = ys__n47561 & new_n45076_;
  assign new_n45110_ = ys__n47209 & ~new_n45080_;
  assign new_n45111_ = ~new_n45109_ & ~new_n45110_;
  assign ys__n31852 = ~new_n45083_ & ~new_n45111_;
  assign new_n45113_ = ys__n47562 & new_n45076_;
  assign new_n45114_ = ys__n47210 & ~new_n45080_;
  assign new_n45115_ = ~new_n45113_ & ~new_n45114_;
  assign ys__n31853 = ~new_n45083_ & ~new_n45115_;
  assign new_n45117_ = ys__n47563 & new_n45076_;
  assign new_n45118_ = ys__n47211 & ~new_n45080_;
  assign new_n45119_ = ~new_n45117_ & ~new_n45118_;
  assign ys__n31854 = ~new_n45083_ & ~new_n45119_;
  assign new_n45121_ = ys__n47564 & new_n45076_;
  assign new_n45122_ = ys__n47212 & ~new_n45080_;
  assign new_n45123_ = ~new_n45121_ & ~new_n45122_;
  assign ys__n31855 = ~new_n45083_ & ~new_n45123_;
  assign new_n45125_ = ys__n47565 & new_n45076_;
  assign new_n45126_ = ys__n47213 & ~new_n45080_;
  assign new_n45127_ = ~new_n45125_ & ~new_n45126_;
  assign ys__n31856 = ~new_n45083_ & ~new_n45127_;
  assign new_n45129_ = ys__n47566 & new_n45076_;
  assign new_n45130_ = ys__n47214 & ~new_n45080_;
  assign new_n45131_ = ~new_n45129_ & ~new_n45130_;
  assign ys__n31857 = ~new_n45083_ & ~new_n45131_;
  assign new_n45133_ = ys__n47567 & new_n45076_;
  assign new_n45134_ = ys__n47215 & ~new_n45080_;
  assign new_n45135_ = ~new_n45133_ & ~new_n45134_;
  assign ys__n31858 = ~new_n45083_ & ~new_n45135_;
  assign new_n45137_ = ys__n47568 & new_n45076_;
  assign new_n45138_ = ys__n47216 & ~new_n45080_;
  assign new_n45139_ = ~new_n45137_ & ~new_n45138_;
  assign ys__n31859 = ~new_n45083_ & ~new_n45139_;
  assign new_n45141_ = ys__n47569 & new_n45076_;
  assign new_n45142_ = ys__n47217 & ~new_n45080_;
  assign new_n45143_ = ~new_n45141_ & ~new_n45142_;
  assign ys__n31860 = ~new_n45083_ & ~new_n45143_;
  assign new_n45145_ = ys__n47570 & new_n45076_;
  assign new_n45146_ = ys__n47218 & ~new_n45080_;
  assign new_n45147_ = ~new_n45145_ & ~new_n45146_;
  assign ys__n31861 = ~new_n45083_ & ~new_n45147_;
  assign new_n45149_ = ys__n47571 & new_n45076_;
  assign new_n45150_ = ys__n47219 & ~new_n45080_;
  assign new_n45151_ = ~new_n45149_ & ~new_n45150_;
  assign ys__n31862 = ~new_n45083_ & ~new_n45151_;
  assign new_n45153_ = ys__n47572 & new_n45076_;
  assign new_n45154_ = ys__n47220 & ~new_n45080_;
  assign new_n45155_ = ~new_n45153_ & ~new_n45154_;
  assign ys__n31863 = ~new_n45083_ & ~new_n45155_;
  assign new_n45157_ = ys__n47573 & new_n45076_;
  assign new_n45158_ = ys__n47221 & ~new_n45080_;
  assign new_n45159_ = ~new_n45157_ & ~new_n45158_;
  assign ys__n31864 = ~new_n45083_ & ~new_n45159_;
  assign new_n45161_ = ys__n47574 & new_n45076_;
  assign new_n45162_ = ys__n47222 & ~new_n45080_;
  assign new_n45163_ = ~new_n45161_ & ~new_n45162_;
  assign ys__n31865 = ~new_n45083_ & ~new_n45163_;
  assign new_n45165_ = ys__n47575 & new_n45076_;
  assign new_n45166_ = ys__n47223 & ~new_n45080_;
  assign new_n45167_ = ~new_n45165_ & ~new_n45166_;
  assign ys__n31866 = ~new_n45083_ & ~new_n45167_;
  assign new_n45169_ = ys__n47576 & new_n45076_;
  assign new_n45170_ = ys__n47224 & ~new_n45080_;
  assign new_n45171_ = ~new_n45169_ & ~new_n45170_;
  assign ys__n31867 = ~new_n45083_ & ~new_n45171_;
  assign new_n45173_ = ys__n47577 & new_n45076_;
  assign new_n45174_ = ys__n47225 & ~new_n45080_;
  assign new_n45175_ = ~new_n45173_ & ~new_n45174_;
  assign ys__n31868 = ~new_n45083_ & ~new_n45175_;
  assign new_n45177_ = ys__n47578 & new_n45076_;
  assign new_n45178_ = ys__n47226 & ~new_n45080_;
  assign new_n45179_ = ~new_n45177_ & ~new_n45178_;
  assign ys__n31869 = ~new_n45083_ & ~new_n45179_;
  assign new_n45181_ = ys__n47579 & new_n45076_;
  assign new_n45182_ = ys__n47227 & ~new_n45080_;
  assign new_n45183_ = ~new_n45181_ & ~new_n45182_;
  assign ys__n31870 = ~new_n45083_ & ~new_n45183_;
  assign new_n45185_ = ys__n47580 & new_n45076_;
  assign new_n45186_ = ys__n47228 & ~new_n45080_;
  assign new_n45187_ = ~new_n45185_ & ~new_n45186_;
  assign ys__n31871 = ~new_n45083_ & ~new_n45187_;
  assign new_n45189_ = ys__n47581 & new_n45076_;
  assign new_n45190_ = ys__n47229 & ~new_n45080_;
  assign new_n45191_ = ~new_n45189_ & ~new_n45190_;
  assign ys__n31872 = ~new_n45083_ & ~new_n45191_;
  assign new_n45193_ = ys__n47582 & new_n45076_;
  assign new_n45194_ = ys__n47230 & ~new_n45080_;
  assign new_n45195_ = ~new_n45193_ & ~new_n45194_;
  assign ys__n31873 = ~new_n45083_ & ~new_n45195_;
  assign new_n45197_ = ys__n47583 & new_n45076_;
  assign new_n45198_ = ys__n47231 & ~new_n45080_;
  assign new_n45199_ = ~new_n45197_ & ~new_n45198_;
  assign ys__n31874 = ~new_n45083_ & ~new_n45199_;
  assign new_n45201_ = ys__n47584 & new_n45076_;
  assign new_n45202_ = ys__n47232 & ~new_n45080_;
  assign new_n45203_ = ~new_n45201_ & ~new_n45202_;
  assign ys__n31875 = ~new_n45083_ & ~new_n45203_;
  assign new_n45205_ = ys__n47585 & new_n45076_;
  assign new_n45206_ = ys__n47233 & ~new_n45080_;
  assign new_n45207_ = ~new_n45205_ & ~new_n45206_;
  assign ys__n31876 = ~new_n45083_ & ~new_n45207_;
  assign new_n45209_ = ys__n47586 & new_n45076_;
  assign new_n45210_ = ys__n18762 & ~new_n45080_;
  assign new_n45211_ = ~new_n45209_ & ~new_n45210_;
  assign ys__n31877 = ~new_n45083_ & ~new_n45211_;
  assign new_n45213_ = ys__n47587 & new_n45076_;
  assign new_n45214_ = ys__n18750 & ~new_n45080_;
  assign new_n45215_ = ~new_n45213_ & ~new_n45214_;
  assign ys__n31878 = ~new_n45083_ & ~new_n45215_;
  assign new_n45217_ = ys__n47588 & new_n45076_;
  assign new_n45218_ = ys__n18753 & ~new_n45080_;
  assign new_n45219_ = ~new_n45217_ & ~new_n45218_;
  assign ys__n31879 = ~new_n45083_ & ~new_n45219_;
  assign new_n45221_ = ys__n852 & new_n13240_;
  assign new_n45222_ = ys__n47589 & new_n45221_;
  assign new_n45223_ = ~ys__n854 & ~new_n13240_;
  assign new_n45224_ = ~ys__n852 & new_n13240_;
  assign new_n45225_ = ~new_n45223_ & ~new_n45224_;
  assign new_n45226_ = ys__n47202 & ~new_n45225_;
  assign new_n45227_ = ~new_n45222_ & ~new_n45226_;
  assign new_n45228_ = ~new_n45221_ & new_n45225_;
  assign ys__n31880 = ~new_n45227_ & ~new_n45228_;
  assign new_n45230_ = ys__n47590 & new_n45221_;
  assign new_n45231_ = ys__n47203 & ~new_n45225_;
  assign new_n45232_ = ~new_n45230_ & ~new_n45231_;
  assign ys__n31881 = ~new_n45228_ & ~new_n45232_;
  assign new_n45234_ = ys__n47591 & new_n45221_;
  assign new_n45235_ = ys__n47204 & ~new_n45225_;
  assign new_n45236_ = ~new_n45234_ & ~new_n45235_;
  assign ys__n31882 = ~new_n45228_ & ~new_n45236_;
  assign new_n45238_ = ys__n47592 & new_n45221_;
  assign new_n45239_ = ys__n47205 & ~new_n45225_;
  assign new_n45240_ = ~new_n45238_ & ~new_n45239_;
  assign ys__n31883 = ~new_n45228_ & ~new_n45240_;
  assign new_n45242_ = ys__n47593 & new_n45221_;
  assign new_n45243_ = ys__n47206 & ~new_n45225_;
  assign new_n45244_ = ~new_n45242_ & ~new_n45243_;
  assign ys__n31884 = ~new_n45228_ & ~new_n45244_;
  assign new_n45246_ = ys__n47594 & new_n45221_;
  assign new_n45247_ = ys__n47207 & ~new_n45225_;
  assign new_n45248_ = ~new_n45246_ & ~new_n45247_;
  assign ys__n31885 = ~new_n45228_ & ~new_n45248_;
  assign new_n45250_ = ys__n47595 & new_n45221_;
  assign new_n45251_ = ys__n47208 & ~new_n45225_;
  assign new_n45252_ = ~new_n45250_ & ~new_n45251_;
  assign ys__n31886 = ~new_n45228_ & ~new_n45252_;
  assign new_n45254_ = ys__n47596 & new_n45221_;
  assign new_n45255_ = ys__n47209 & ~new_n45225_;
  assign new_n45256_ = ~new_n45254_ & ~new_n45255_;
  assign ys__n31887 = ~new_n45228_ & ~new_n45256_;
  assign new_n45258_ = ys__n47597 & new_n45221_;
  assign new_n45259_ = ys__n47210 & ~new_n45225_;
  assign new_n45260_ = ~new_n45258_ & ~new_n45259_;
  assign ys__n31888 = ~new_n45228_ & ~new_n45260_;
  assign new_n45262_ = ys__n47598 & new_n45221_;
  assign new_n45263_ = ys__n47211 & ~new_n45225_;
  assign new_n45264_ = ~new_n45262_ & ~new_n45263_;
  assign ys__n31889 = ~new_n45228_ & ~new_n45264_;
  assign new_n45266_ = ys__n47599 & new_n45221_;
  assign new_n45267_ = ys__n47212 & ~new_n45225_;
  assign new_n45268_ = ~new_n45266_ & ~new_n45267_;
  assign ys__n31890 = ~new_n45228_ & ~new_n45268_;
  assign new_n45270_ = ys__n47600 & new_n45221_;
  assign new_n45271_ = ys__n47213 & ~new_n45225_;
  assign new_n45272_ = ~new_n45270_ & ~new_n45271_;
  assign ys__n31891 = ~new_n45228_ & ~new_n45272_;
  assign new_n45274_ = ys__n47601 & new_n45221_;
  assign new_n45275_ = ys__n47214 & ~new_n45225_;
  assign new_n45276_ = ~new_n45274_ & ~new_n45275_;
  assign ys__n31892 = ~new_n45228_ & ~new_n45276_;
  assign new_n45278_ = ys__n47602 & new_n45221_;
  assign new_n45279_ = ys__n47215 & ~new_n45225_;
  assign new_n45280_ = ~new_n45278_ & ~new_n45279_;
  assign ys__n31893 = ~new_n45228_ & ~new_n45280_;
  assign new_n45282_ = ys__n47603 & new_n45221_;
  assign new_n45283_ = ys__n47216 & ~new_n45225_;
  assign new_n45284_ = ~new_n45282_ & ~new_n45283_;
  assign ys__n31894 = ~new_n45228_ & ~new_n45284_;
  assign new_n45286_ = ys__n47604 & new_n45221_;
  assign new_n45287_ = ys__n47217 & ~new_n45225_;
  assign new_n45288_ = ~new_n45286_ & ~new_n45287_;
  assign ys__n31895 = ~new_n45228_ & ~new_n45288_;
  assign new_n45290_ = ys__n47605 & new_n45221_;
  assign new_n45291_ = ys__n47218 & ~new_n45225_;
  assign new_n45292_ = ~new_n45290_ & ~new_n45291_;
  assign ys__n31896 = ~new_n45228_ & ~new_n45292_;
  assign new_n45294_ = ys__n47606 & new_n45221_;
  assign new_n45295_ = ys__n47219 & ~new_n45225_;
  assign new_n45296_ = ~new_n45294_ & ~new_n45295_;
  assign ys__n31897 = ~new_n45228_ & ~new_n45296_;
  assign new_n45298_ = ys__n47607 & new_n45221_;
  assign new_n45299_ = ys__n47220 & ~new_n45225_;
  assign new_n45300_ = ~new_n45298_ & ~new_n45299_;
  assign ys__n31898 = ~new_n45228_ & ~new_n45300_;
  assign new_n45302_ = ys__n47608 & new_n45221_;
  assign new_n45303_ = ys__n47221 & ~new_n45225_;
  assign new_n45304_ = ~new_n45302_ & ~new_n45303_;
  assign ys__n31899 = ~new_n45228_ & ~new_n45304_;
  assign new_n45306_ = ys__n47609 & new_n45221_;
  assign new_n45307_ = ys__n47222 & ~new_n45225_;
  assign new_n45308_ = ~new_n45306_ & ~new_n45307_;
  assign ys__n31900 = ~new_n45228_ & ~new_n45308_;
  assign new_n45310_ = ys__n47610 & new_n45221_;
  assign new_n45311_ = ys__n47223 & ~new_n45225_;
  assign new_n45312_ = ~new_n45310_ & ~new_n45311_;
  assign ys__n31901 = ~new_n45228_ & ~new_n45312_;
  assign new_n45314_ = ys__n47611 & new_n45221_;
  assign new_n45315_ = ys__n47224 & ~new_n45225_;
  assign new_n45316_ = ~new_n45314_ & ~new_n45315_;
  assign ys__n31902 = ~new_n45228_ & ~new_n45316_;
  assign new_n45318_ = ys__n47612 & new_n45221_;
  assign new_n45319_ = ys__n47225 & ~new_n45225_;
  assign new_n45320_ = ~new_n45318_ & ~new_n45319_;
  assign ys__n31903 = ~new_n45228_ & ~new_n45320_;
  assign new_n45322_ = ys__n47613 & new_n45221_;
  assign new_n45323_ = ys__n47226 & ~new_n45225_;
  assign new_n45324_ = ~new_n45322_ & ~new_n45323_;
  assign ys__n31904 = ~new_n45228_ & ~new_n45324_;
  assign new_n45326_ = ys__n47614 & new_n45221_;
  assign new_n45327_ = ys__n47227 & ~new_n45225_;
  assign new_n45328_ = ~new_n45326_ & ~new_n45327_;
  assign ys__n31905 = ~new_n45228_ & ~new_n45328_;
  assign new_n45330_ = ys__n47615 & new_n45221_;
  assign new_n45331_ = ys__n47228 & ~new_n45225_;
  assign new_n45332_ = ~new_n45330_ & ~new_n45331_;
  assign ys__n31906 = ~new_n45228_ & ~new_n45332_;
  assign new_n45334_ = ys__n47616 & new_n45221_;
  assign new_n45335_ = ys__n47229 & ~new_n45225_;
  assign new_n45336_ = ~new_n45334_ & ~new_n45335_;
  assign ys__n31907 = ~new_n45228_ & ~new_n45336_;
  assign new_n45338_ = ys__n47617 & new_n45221_;
  assign new_n45339_ = ys__n47230 & ~new_n45225_;
  assign new_n45340_ = ~new_n45338_ & ~new_n45339_;
  assign ys__n31908 = ~new_n45228_ & ~new_n45340_;
  assign new_n45342_ = ys__n47618 & new_n45221_;
  assign new_n45343_ = ys__n47231 & ~new_n45225_;
  assign new_n45344_ = ~new_n45342_ & ~new_n45343_;
  assign ys__n31909 = ~new_n45228_ & ~new_n45344_;
  assign new_n45346_ = ys__n47619 & new_n45221_;
  assign new_n45347_ = ys__n47232 & ~new_n45225_;
  assign new_n45348_ = ~new_n45346_ & ~new_n45347_;
  assign ys__n31910 = ~new_n45228_ & ~new_n45348_;
  assign new_n45350_ = ys__n47620 & new_n45221_;
  assign new_n45351_ = ys__n47233 & ~new_n45225_;
  assign new_n45352_ = ~new_n45350_ & ~new_n45351_;
  assign ys__n31911 = ~new_n45228_ & ~new_n45352_;
  assign new_n45354_ = ys__n47621 & new_n45221_;
  assign new_n45355_ = ys__n18762 & ~new_n45225_;
  assign new_n45356_ = ~new_n45354_ & ~new_n45355_;
  assign ys__n31912 = ~new_n45228_ & ~new_n45356_;
  assign new_n45358_ = ys__n47622 & new_n45221_;
  assign new_n45359_ = ys__n18750 & ~new_n45225_;
  assign new_n45360_ = ~new_n45358_ & ~new_n45359_;
  assign ys__n31913 = ~new_n45228_ & ~new_n45360_;
  assign new_n45362_ = ys__n47623 & new_n45221_;
  assign new_n45363_ = ys__n18753 & ~new_n45225_;
  assign new_n45364_ = ~new_n45362_ & ~new_n45363_;
  assign ys__n31914 = ~new_n45228_ & ~new_n45364_;
  assign new_n45366_ = ys__n850 & new_n13240_;
  assign new_n45367_ = ys__n47624 & new_n45366_;
  assign new_n45368_ = ~ys__n852 & ~new_n13240_;
  assign new_n45369_ = ~ys__n850 & new_n13240_;
  assign new_n45370_ = ~new_n45368_ & ~new_n45369_;
  assign new_n45371_ = ys__n47202 & ~new_n45370_;
  assign new_n45372_ = ~new_n45367_ & ~new_n45371_;
  assign new_n45373_ = ~new_n45366_ & new_n45370_;
  assign ys__n31915 = ~new_n45372_ & ~new_n45373_;
  assign new_n45375_ = ys__n47625 & new_n45366_;
  assign new_n45376_ = ys__n47203 & ~new_n45370_;
  assign new_n45377_ = ~new_n45375_ & ~new_n45376_;
  assign ys__n31916 = ~new_n45373_ & ~new_n45377_;
  assign new_n45379_ = ys__n47626 & new_n45366_;
  assign new_n45380_ = ys__n47204 & ~new_n45370_;
  assign new_n45381_ = ~new_n45379_ & ~new_n45380_;
  assign ys__n31917 = ~new_n45373_ & ~new_n45381_;
  assign new_n45383_ = ys__n47627 & new_n45366_;
  assign new_n45384_ = ys__n47205 & ~new_n45370_;
  assign new_n45385_ = ~new_n45383_ & ~new_n45384_;
  assign ys__n31918 = ~new_n45373_ & ~new_n45385_;
  assign new_n45387_ = ys__n47628 & new_n45366_;
  assign new_n45388_ = ys__n47206 & ~new_n45370_;
  assign new_n45389_ = ~new_n45387_ & ~new_n45388_;
  assign ys__n31919 = ~new_n45373_ & ~new_n45389_;
  assign new_n45391_ = ys__n47629 & new_n45366_;
  assign new_n45392_ = ys__n47207 & ~new_n45370_;
  assign new_n45393_ = ~new_n45391_ & ~new_n45392_;
  assign ys__n31920 = ~new_n45373_ & ~new_n45393_;
  assign new_n45395_ = ys__n47630 & new_n45366_;
  assign new_n45396_ = ys__n47208 & ~new_n45370_;
  assign new_n45397_ = ~new_n45395_ & ~new_n45396_;
  assign ys__n31921 = ~new_n45373_ & ~new_n45397_;
  assign new_n45399_ = ys__n47631 & new_n45366_;
  assign new_n45400_ = ys__n47209 & ~new_n45370_;
  assign new_n45401_ = ~new_n45399_ & ~new_n45400_;
  assign ys__n31922 = ~new_n45373_ & ~new_n45401_;
  assign new_n45403_ = ys__n47632 & new_n45366_;
  assign new_n45404_ = ys__n47210 & ~new_n45370_;
  assign new_n45405_ = ~new_n45403_ & ~new_n45404_;
  assign ys__n31923 = ~new_n45373_ & ~new_n45405_;
  assign new_n45407_ = ys__n47633 & new_n45366_;
  assign new_n45408_ = ys__n47211 & ~new_n45370_;
  assign new_n45409_ = ~new_n45407_ & ~new_n45408_;
  assign ys__n31924 = ~new_n45373_ & ~new_n45409_;
  assign new_n45411_ = ys__n47634 & new_n45366_;
  assign new_n45412_ = ys__n47212 & ~new_n45370_;
  assign new_n45413_ = ~new_n45411_ & ~new_n45412_;
  assign ys__n31925 = ~new_n45373_ & ~new_n45413_;
  assign new_n45415_ = ys__n47635 & new_n45366_;
  assign new_n45416_ = ys__n47213 & ~new_n45370_;
  assign new_n45417_ = ~new_n45415_ & ~new_n45416_;
  assign ys__n31926 = ~new_n45373_ & ~new_n45417_;
  assign new_n45419_ = ys__n47636 & new_n45366_;
  assign new_n45420_ = ys__n47214 & ~new_n45370_;
  assign new_n45421_ = ~new_n45419_ & ~new_n45420_;
  assign ys__n31927 = ~new_n45373_ & ~new_n45421_;
  assign new_n45423_ = ys__n47637 & new_n45366_;
  assign new_n45424_ = ys__n47215 & ~new_n45370_;
  assign new_n45425_ = ~new_n45423_ & ~new_n45424_;
  assign ys__n31928 = ~new_n45373_ & ~new_n45425_;
  assign new_n45427_ = ys__n47638 & new_n45366_;
  assign new_n45428_ = ys__n47216 & ~new_n45370_;
  assign new_n45429_ = ~new_n45427_ & ~new_n45428_;
  assign ys__n31929 = ~new_n45373_ & ~new_n45429_;
  assign new_n45431_ = ys__n47639 & new_n45366_;
  assign new_n45432_ = ys__n47217 & ~new_n45370_;
  assign new_n45433_ = ~new_n45431_ & ~new_n45432_;
  assign ys__n31930 = ~new_n45373_ & ~new_n45433_;
  assign new_n45435_ = ys__n47640 & new_n45366_;
  assign new_n45436_ = ys__n47218 & ~new_n45370_;
  assign new_n45437_ = ~new_n45435_ & ~new_n45436_;
  assign ys__n31931 = ~new_n45373_ & ~new_n45437_;
  assign new_n45439_ = ys__n47641 & new_n45366_;
  assign new_n45440_ = ys__n47219 & ~new_n45370_;
  assign new_n45441_ = ~new_n45439_ & ~new_n45440_;
  assign ys__n31932 = ~new_n45373_ & ~new_n45441_;
  assign new_n45443_ = ys__n47642 & new_n45366_;
  assign new_n45444_ = ys__n47220 & ~new_n45370_;
  assign new_n45445_ = ~new_n45443_ & ~new_n45444_;
  assign ys__n31933 = ~new_n45373_ & ~new_n45445_;
  assign new_n45447_ = ys__n47643 & new_n45366_;
  assign new_n45448_ = ys__n47221 & ~new_n45370_;
  assign new_n45449_ = ~new_n45447_ & ~new_n45448_;
  assign ys__n31934 = ~new_n45373_ & ~new_n45449_;
  assign new_n45451_ = ys__n47644 & new_n45366_;
  assign new_n45452_ = ys__n47222 & ~new_n45370_;
  assign new_n45453_ = ~new_n45451_ & ~new_n45452_;
  assign ys__n31935 = ~new_n45373_ & ~new_n45453_;
  assign new_n45455_ = ys__n47645 & new_n45366_;
  assign new_n45456_ = ys__n47223 & ~new_n45370_;
  assign new_n45457_ = ~new_n45455_ & ~new_n45456_;
  assign ys__n31936 = ~new_n45373_ & ~new_n45457_;
  assign new_n45459_ = ys__n47646 & new_n45366_;
  assign new_n45460_ = ys__n47224 & ~new_n45370_;
  assign new_n45461_ = ~new_n45459_ & ~new_n45460_;
  assign ys__n31937 = ~new_n45373_ & ~new_n45461_;
  assign new_n45463_ = ys__n47647 & new_n45366_;
  assign new_n45464_ = ys__n47225 & ~new_n45370_;
  assign new_n45465_ = ~new_n45463_ & ~new_n45464_;
  assign ys__n31938 = ~new_n45373_ & ~new_n45465_;
  assign new_n45467_ = ys__n47648 & new_n45366_;
  assign new_n45468_ = ys__n47226 & ~new_n45370_;
  assign new_n45469_ = ~new_n45467_ & ~new_n45468_;
  assign ys__n31939 = ~new_n45373_ & ~new_n45469_;
  assign new_n45471_ = ys__n47649 & new_n45366_;
  assign new_n45472_ = ys__n47227 & ~new_n45370_;
  assign new_n45473_ = ~new_n45471_ & ~new_n45472_;
  assign ys__n31940 = ~new_n45373_ & ~new_n45473_;
  assign new_n45475_ = ys__n47650 & new_n45366_;
  assign new_n45476_ = ys__n47228 & ~new_n45370_;
  assign new_n45477_ = ~new_n45475_ & ~new_n45476_;
  assign ys__n31941 = ~new_n45373_ & ~new_n45477_;
  assign new_n45479_ = ys__n47651 & new_n45366_;
  assign new_n45480_ = ys__n47229 & ~new_n45370_;
  assign new_n45481_ = ~new_n45479_ & ~new_n45480_;
  assign ys__n31942 = ~new_n45373_ & ~new_n45481_;
  assign new_n45483_ = ys__n47652 & new_n45366_;
  assign new_n45484_ = ys__n47230 & ~new_n45370_;
  assign new_n45485_ = ~new_n45483_ & ~new_n45484_;
  assign ys__n31943 = ~new_n45373_ & ~new_n45485_;
  assign new_n45487_ = ys__n47653 & new_n45366_;
  assign new_n45488_ = ys__n47231 & ~new_n45370_;
  assign new_n45489_ = ~new_n45487_ & ~new_n45488_;
  assign ys__n31944 = ~new_n45373_ & ~new_n45489_;
  assign new_n45491_ = ys__n47654 & new_n45366_;
  assign new_n45492_ = ys__n47232 & ~new_n45370_;
  assign new_n45493_ = ~new_n45491_ & ~new_n45492_;
  assign ys__n31945 = ~new_n45373_ & ~new_n45493_;
  assign new_n45495_ = ys__n47655 & new_n45366_;
  assign new_n45496_ = ys__n47233 & ~new_n45370_;
  assign new_n45497_ = ~new_n45495_ & ~new_n45496_;
  assign ys__n31946 = ~new_n45373_ & ~new_n45497_;
  assign new_n45499_ = ys__n47656 & new_n45366_;
  assign new_n45500_ = ys__n18762 & ~new_n45370_;
  assign new_n45501_ = ~new_n45499_ & ~new_n45500_;
  assign ys__n31947 = ~new_n45373_ & ~new_n45501_;
  assign new_n45503_ = ys__n47657 & new_n45366_;
  assign new_n45504_ = ys__n18750 & ~new_n45370_;
  assign new_n45505_ = ~new_n45503_ & ~new_n45504_;
  assign ys__n31948 = ~new_n45373_ & ~new_n45505_;
  assign new_n45507_ = ys__n47658 & new_n45366_;
  assign new_n45508_ = ys__n18753 & ~new_n45370_;
  assign new_n45509_ = ~new_n45507_ & ~new_n45508_;
  assign ys__n31949 = ~new_n45373_ & ~new_n45509_;
  assign new_n45511_ = ~ys__n556 & ys__n558;
  assign new_n45512_ = ~ys__n935 & ~ys__n1802;
  assign new_n45513_ = new_n45511_ & new_n45512_;
  assign new_n45514_ = ys__n556 & ~ys__n935;
  assign new_n45515_ = ~ys__n1802 & new_n45514_;
  assign new_n45516_ = ~new_n45513_ & ~new_n45515_;
  assign new_n45517_ = ~ys__n556 & ~ys__n558;
  assign new_n45518_ = ys__n935 & ~ys__n1802;
  assign new_n45519_ = new_n45517_ & new_n45518_;
  assign new_n45520_ = ys__n556 & ys__n935;
  assign new_n45521_ = ~ys__n1802 & new_n45520_;
  assign new_n45522_ = ~ys__n1802 & ~new_n45521_;
  assign new_n45523_ = ~new_n45519_ & new_n45522_;
  assign new_n45524_ = new_n45511_ & new_n45518_;
  assign new_n45525_ = new_n45512_ & new_n45517_;
  assign new_n45526_ = ~new_n45524_ & ~new_n45525_;
  assign new_n45527_ = new_n45523_ & new_n45526_;
  assign new_n45528_ = new_n45516_ & new_n45527_;
  assign new_n45529_ = new_n13717_ & ~new_n45516_;
  assign new_n45530_ = ~new_n45528_ & new_n45529_;
  assign new_n45531_ = ys__n556 & ~ys__n1802;
  assign new_n45532_ = ys__n178 & new_n12124_;
  assign new_n45533_ = ~ys__n176 & ~ys__n558;
  assign new_n45534_ = new_n45532_ & new_n45533_;
  assign new_n45535_ = new_n45531_ & new_n45534_;
  assign new_n45536_ = ys__n178 & ~new_n12124_;
  assign new_n45537_ = new_n45533_ & new_n45536_;
  assign new_n45538_ = new_n45531_ & new_n45537_;
  assign new_n45539_ = ~new_n45535_ & ~new_n45538_;
  assign new_n45540_ = ~ys__n176 & ys__n558;
  assign new_n45541_ = new_n45532_ & new_n45540_;
  assign new_n45542_ = new_n45531_ & new_n45541_;
  assign new_n45543_ = new_n45536_ & new_n45540_;
  assign new_n45544_ = new_n45531_ & new_n45543_;
  assign new_n45545_ = ~new_n45542_ & ~new_n45544_;
  assign new_n45546_ = new_n45539_ & new_n45545_;
  assign new_n45547_ = new_n12127_ & new_n45511_;
  assign new_n45548_ = ~ys__n1802 & new_n45547_;
  assign new_n45549_ = ys__n556 & ~ys__n558;
  assign new_n45550_ = new_n12127_ & new_n45549_;
  assign new_n45551_ = ~ys__n1802 & new_n45550_;
  assign new_n45552_ = ~new_n45548_ & ~new_n45551_;
  assign new_n45553_ = ys__n556 & ys__n558;
  assign new_n45554_ = new_n12135_ & new_n45553_;
  assign new_n45555_ = ~ys__n1802 & new_n45554_;
  assign new_n45556_ = new_n12134_ & new_n45553_;
  assign new_n45557_ = ~ys__n1802 & new_n45556_;
  assign new_n45558_ = new_n12127_ & new_n45553_;
  assign new_n45559_ = ~ys__n1802 & new_n45558_;
  assign new_n45560_ = ~new_n45557_ & ~new_n45559_;
  assign new_n45561_ = ~new_n45555_ & new_n45560_;
  assign new_n45562_ = new_n45552_ & new_n45561_;
  assign new_n45563_ = ~ys__n556 & ~ys__n1802;
  assign new_n45564_ = new_n45541_ & new_n45563_;
  assign new_n45565_ = new_n45543_ & new_n45563_;
  assign new_n45566_ = ~new_n45564_ & ~new_n45565_;
  assign new_n45567_ = new_n45562_ & new_n45566_;
  assign new_n45568_ = new_n45546_ & new_n45567_;
  assign new_n45569_ = new_n12134_ & new_n45511_;
  assign new_n45570_ = ~ys__n1802 & new_n45569_;
  assign new_n45571_ = new_n12135_ & new_n45511_;
  assign new_n45572_ = ~ys__n1802 & new_n45571_;
  assign new_n45573_ = ~new_n45570_ & ~new_n45572_;
  assign new_n45574_ = new_n12134_ & new_n45549_;
  assign new_n45575_ = ~ys__n1802 & new_n45574_;
  assign new_n45576_ = new_n12135_ & new_n45549_;
  assign new_n45577_ = ~ys__n1802 & new_n45576_;
  assign new_n45578_ = ~new_n45575_ & ~new_n45577_;
  assign new_n45579_ = new_n45573_ & new_n45578_;
  assign new_n45580_ = new_n12134_ & new_n45517_;
  assign new_n45581_ = ~ys__n1802 & new_n45580_;
  assign new_n45582_ = ~ys__n1802 & ~new_n45581_;
  assign new_n45583_ = new_n12127_ & new_n45517_;
  assign new_n45584_ = ~ys__n1802 & new_n45583_;
  assign new_n45585_ = new_n12135_ & new_n45517_;
  assign new_n45586_ = ~ys__n1802 & new_n45585_;
  assign new_n45587_ = ~new_n45584_ & ~new_n45586_;
  assign new_n45588_ = new_n45582_ & new_n45587_;
  assign new_n45589_ = new_n45579_ & new_n45588_;
  assign new_n45590_ = new_n45534_ & new_n45563_;
  assign new_n45591_ = new_n45537_ & new_n45563_;
  assign new_n45592_ = ~new_n45590_ & ~new_n45591_;
  assign new_n45593_ = new_n45589_ & new_n45592_;
  assign new_n45594_ = new_n45568_ & new_n45593_;
  assign new_n45595_ = new_n12140_ & ~new_n45568_;
  assign new_n45596_ = ~new_n45594_ & new_n45595_;
  assign new_n45597_ = ~new_n45530_ & ~new_n45596_;
  assign new_n45598_ = ~ys__n738 & ~new_n12140_;
  assign new_n45599_ = ~new_n13717_ & new_n45598_;
  assign ys__n31950 = ~new_n45597_ & ~new_n45599_;
  assign new_n45601_ = ~new_n45559_ & ~new_n45584_;
  assign new_n45602_ = new_n45552_ & new_n45601_;
  assign new_n45603_ = ~new_n45564_ & new_n45602_;
  assign new_n45604_ = ~new_n45535_ & ~new_n45542_;
  assign new_n45605_ = ~new_n45590_ & new_n45604_;
  assign new_n45606_ = new_n45603_ & new_n45605_;
  assign new_n45607_ = ~new_n45555_ & ~new_n45572_;
  assign new_n45608_ = ~new_n45577_ & new_n45607_;
  assign new_n45609_ = new_n45606_ & new_n45608_;
  assign new_n45610_ = ~new_n45538_ & ~new_n45565_;
  assign new_n45611_ = ~new_n45544_ & ~new_n45591_;
  assign new_n45612_ = new_n45610_ & new_n45611_;
  assign new_n45613_ = ~new_n45557_ & ~new_n45570_;
  assign new_n45614_ = ~new_n45575_ & new_n45613_;
  assign new_n45615_ = new_n45612_ & new_n45614_;
  assign new_n45616_ = ~new_n45581_ & ~new_n45586_;
  assign new_n45617_ = ~ys__n1802 & new_n45616_;
  assign new_n45618_ = new_n45615_ & new_n45617_;
  assign new_n45619_ = new_n45609_ & new_n45618_;
  assign new_n45620_ = new_n45615_ & new_n45616_;
  assign new_n45621_ = new_n12140_ & ~new_n45620_;
  assign new_n45622_ = ~new_n45619_ & new_n45621_;
  assign new_n45623_ = ~new_n45531_ & ~new_n45563_;
  assign new_n45624_ = ~ys__n1802 & new_n45623_;
  assign new_n45625_ = ys__n738 & new_n45563_;
  assign new_n45626_ = ~new_n45624_ & new_n45625_;
  assign new_n45627_ = new_n45516_ & ~new_n45525_;
  assign new_n45628_ = ~new_n45521_ & ~new_n45524_;
  assign new_n45629_ = ~ys__n1802 & ~new_n45519_;
  assign new_n45630_ = new_n45628_ & new_n45629_;
  assign new_n45631_ = new_n45627_ & new_n45630_;
  assign new_n45632_ = new_n13717_ & new_n45519_;
  assign new_n45633_ = ~new_n45631_ & new_n45632_;
  assign new_n45634_ = ~new_n45626_ & ~new_n45633_;
  assign new_n45635_ = ~new_n45622_ & new_n45634_;
  assign ys__n31953 = ~new_n45599_ & ~new_n45635_;
  assign new_n45637_ = new_n45609_ & new_n45616_;
  assign new_n45638_ = new_n12140_ & ~new_n45619_;
  assign new_n45639_ = ~new_n45637_ & new_n45638_;
  assign new_n45640_ = ys__n738 & ~new_n45623_;
  assign new_n45641_ = ~new_n45624_ & new_n45640_;
  assign new_n45642_ = ~new_n45519_ & new_n45628_;
  assign new_n45643_ = new_n13717_ & ~new_n45642_;
  assign new_n45644_ = ~new_n45631_ & new_n45643_;
  assign new_n45645_ = ~new_n45641_ & ~new_n45644_;
  assign new_n45646_ = ~new_n45639_ & new_n45645_;
  assign ys__n31954 = ~new_n45599_ & ~new_n45646_;
  assign new_n45648_ = ~new_n45586_ & new_n45612_;
  assign new_n45649_ = new_n45606_ & new_n45648_;
  assign new_n45650_ = new_n12140_ & ~new_n45649_;
  assign new_n45651_ = ~new_n45619_ & new_n45650_;
  assign new_n45652_ = ~new_n45519_ & new_n45627_;
  assign new_n45653_ = new_n13717_ & ~new_n45631_;
  assign new_n45654_ = ~new_n45652_ & new_n45653_;
  assign new_n45655_ = ~new_n45626_ & ~new_n45654_;
  assign new_n45656_ = ~new_n45651_ & new_n45655_;
  assign ys__n31955 = ~new_n45599_ & ~new_n45656_;
  assign new_n45658_ = ys__n29846 & new_n11735_;
  assign new_n45659_ = ~new_n11735_ & ys__n29847;
  assign new_n45660_ = ~new_n45658_ & ~new_n45659_;
  assign new_n45661_ = ~ys__n23764 & ~new_n45660_;
  assign new_n45662_ = ys__n29898 & ~new_n11737_;
  assign new_n45663_ = ~new_n11735_ & new_n45662_;
  assign new_n45664_ = ~ys__n22466 & new_n45663_;
  assign new_n45665_ = ys__n22466 & ~new_n45660_;
  assign new_n45666_ = ~new_n45664_ & ~new_n45665_;
  assign new_n45667_ = ys__n23764 & ~new_n45666_;
  assign new_n45668_ = ~new_n45661_ & ~new_n45667_;
  assign ys__n31965 = new_n12000_ & ~new_n45668_;
  assign new_n45670_ = ys__n29887 & ~new_n11737_;
  assign new_n45671_ = ~new_n11735_ & new_n45670_;
  assign new_n45672_ = ~ys__n23764 & new_n45671_;
  assign new_n45673_ = ys__n29903 & ~new_n11737_;
  assign new_n45674_ = ~new_n11735_ & new_n45673_;
  assign new_n45675_ = ~ys__n22466 & new_n45674_;
  assign new_n45676_ = ys__n22466 & new_n45671_;
  assign new_n45677_ = ~new_n45675_ & ~new_n45676_;
  assign new_n45678_ = ys__n23764 & ~new_n45677_;
  assign new_n45679_ = ~new_n45672_ & ~new_n45678_;
  assign ys__n31971 = new_n12000_ & ~new_n45679_;
  assign new_n45681_ = ys__n29888 & ~new_n11737_;
  assign new_n45682_ = ~new_n11735_ & new_n45681_;
  assign new_n45683_ = ~ys__n23764 & new_n45682_;
  assign new_n45684_ = ys__n29904 & ~new_n11737_;
  assign new_n45685_ = ~new_n11735_ & new_n45684_;
  assign new_n45686_ = ~ys__n22466 & new_n45685_;
  assign new_n45687_ = ys__n22466 & new_n45682_;
  assign new_n45688_ = ~new_n45686_ & ~new_n45687_;
  assign new_n45689_ = ys__n23764 & ~new_n45688_;
  assign new_n45690_ = ~new_n45683_ & ~new_n45689_;
  assign ys__n31973 = new_n12000_ & ~new_n45690_;
  assign new_n45692_ = ys__n29889 & ~new_n11737_;
  assign new_n45693_ = ~new_n11735_ & new_n45692_;
  assign new_n45694_ = ~ys__n23764 & new_n45693_;
  assign new_n45695_ = ys__n29905 & ~new_n11737_;
  assign new_n45696_ = ~new_n11735_ & new_n45695_;
  assign new_n45697_ = ~ys__n22466 & new_n45696_;
  assign new_n45698_ = ys__n22466 & new_n45693_;
  assign new_n45699_ = ~new_n45697_ & ~new_n45698_;
  assign new_n45700_ = ys__n23764 & ~new_n45699_;
  assign new_n45701_ = ~new_n45694_ & ~new_n45700_;
  assign ys__n31975 = new_n12000_ & ~new_n45701_;
  assign new_n45703_ = ys__n29890 & ~new_n11737_;
  assign new_n45704_ = ~new_n11735_ & new_n45703_;
  assign new_n45705_ = ~ys__n23764 & new_n45704_;
  assign new_n45706_ = ys__n29906 & ~new_n11737_;
  assign new_n45707_ = ~new_n11735_ & new_n45706_;
  assign new_n45708_ = ~ys__n22466 & new_n45707_;
  assign new_n45709_ = ys__n22466 & new_n45704_;
  assign new_n45710_ = ~new_n45708_ & ~new_n45709_;
  assign new_n45711_ = ys__n23764 & ~new_n45710_;
  assign new_n45712_ = ~new_n45705_ & ~new_n45711_;
  assign new_n45713_ = ~new_n11993_ & ~new_n45712_;
  assign new_n45714_ = ~new_n13198_ & ~new_n45713_;
  assign ys__n31976 = ~new_n11999_ & ~new_n45714_;
  assign new_n45716_ = ys__n29891 & ~new_n11737_;
  assign new_n45717_ = ~new_n11735_ & new_n45716_;
  assign new_n45718_ = ~ys__n23764 & new_n45717_;
  assign new_n45719_ = ys__n29907 & ~new_n11737_;
  assign new_n45720_ = ~new_n11735_ & new_n45719_;
  assign new_n45721_ = ~ys__n22466 & new_n45720_;
  assign new_n45722_ = ys__n22466 & new_n45717_;
  assign new_n45723_ = ~new_n45721_ & ~new_n45722_;
  assign new_n45724_ = ys__n23764 & ~new_n45723_;
  assign new_n45725_ = ~new_n45718_ & ~new_n45724_;
  assign ys__n31978 = new_n12000_ & ~new_n45725_;
  assign new_n45727_ = ys__n29892 & ~new_n11737_;
  assign new_n45728_ = ~new_n11735_ & new_n45727_;
  assign new_n45729_ = ~ys__n23764 & new_n45728_;
  assign new_n45730_ = ys__n29908 & ~new_n11737_;
  assign new_n45731_ = ~new_n11735_ & new_n45730_;
  assign new_n45732_ = ~ys__n22466 & new_n45731_;
  assign new_n45733_ = ys__n22466 & new_n45728_;
  assign new_n45734_ = ~new_n45732_ & ~new_n45733_;
  assign new_n45735_ = ys__n23764 & ~new_n45734_;
  assign new_n45736_ = ~new_n45729_ & ~new_n45735_;
  assign new_n45737_ = ~new_n11993_ & ~new_n45736_;
  assign new_n45738_ = ~new_n13198_ & ~new_n45737_;
  assign ys__n31979 = ~new_n11999_ & ~new_n45738_;
  assign new_n45740_ = ~ys__n23764 & ~new_n11993_;
  assign new_n45741_ = ~new_n11999_ & new_n45740_;
  assign ys__n31984 = new_n45663_ & new_n45741_;
  assign ys__n31986 = new_n27304_ & new_n45741_;
  assign ys__n31988 = new_n27315_ & new_n45741_;
  assign ys__n31990 = new_n27326_ & new_n45741_;
  assign ys__n31992 = new_n18026_ & new_n45741_;
  assign ys__n31994 = new_n45674_ & new_n45741_;
  assign ys__n31996 = new_n45685_ & new_n45741_;
  assign ys__n31998 = new_n45696_ & new_n45741_;
  assign ys__n32000 = new_n45707_ & new_n45741_;
  assign ys__n32002 = new_n45720_ & new_n45741_;
  assign new_n45752_ = ~ys__n23764 & new_n45731_;
  assign new_n45753_ = ~new_n18045_ & ~new_n45752_;
  assign ys__n32004 = new_n12000_ & ~new_n45753_;
  assign new_n45755_ = ~ys__n23764 & new_n18041_;
  assign new_n45756_ = ~new_n13271_ & ~new_n45755_;
  assign ys__n32006 = new_n12000_ & ~new_n45756_;
  assign new_n45758_ = ~ys__n23764 & new_n13267_;
  assign new_n45759_ = ~new_n13253_ & ~new_n45758_;
  assign new_n45760_ = ~new_n11993_ & ~new_n45759_;
  assign new_n45761_ = ~new_n13198_ & ~new_n45760_;
  assign ys__n32007 = ~new_n11999_ & ~new_n45761_;
  assign new_n45763_ = ~ys__n23764 & new_n13249_;
  assign new_n45764_ = ~new_n13195_ & ~new_n45763_;
  assign new_n45765_ = ~new_n11993_ & ~new_n45764_;
  assign new_n45766_ = ~new_n13198_ & ~new_n45765_;
  assign ys__n32008 = ~new_n11999_ & ~new_n45766_;
  assign ys__n32010 = new_n13191_ & new_n45741_;
  assign new_n45769_ = ~ys__n23764 & new_n11754_;
  assign new_n45770_ = ~new_n11761_ & ~new_n45769_;
  assign ys__n32012 = new_n12000_ & ~new_n45770_;
  assign new_n45772_ = new_n12457_ & new_n22631_;
  assign ys__n32014 = ~new_n22633_ & new_n45772_;
  assign new_n45774_ = new_n12477_ & new_n22631_;
  assign ys__n32016 = ~new_n22633_ & new_n45774_;
  assign new_n45776_ = new_n12453_ & new_n22631_;
  assign ys__n32018 = ~new_n22633_ & new_n45776_;
  assign new_n45778_ = ~ys__n23661 & ys__n23663;
  assign new_n45779_ = ~ys__n28459 & new_n45778_;
  assign new_n45780_ = ys__n23661 & ~ys__n28457;
  assign new_n45781_ = ~new_n45779_ & ~new_n45780_;
  assign new_n45782_ = ~ys__n23658 & ~new_n45781_;
  assign new_n45783_ = ys__n23658 & ~ys__n28455;
  assign new_n45784_ = ~new_n45782_ & ~new_n45783_;
  assign new_n45785_ = ~ys__n23655 & ~new_n45784_;
  assign new_n45786_ = ys__n23655 & ~ys__n28453;
  assign new_n45787_ = ys__n38315 & new_n45786_;
  assign new_n45788_ = ~new_n45785_ & ~new_n45787_;
  assign new_n45789_ = ~ys__n352 & ~ys__n19973;
  assign new_n45790_ = ys__n38424 & new_n45789_;
  assign new_n45791_ = new_n45788_ & ~new_n45790_;
  assign new_n45792_ = ys__n544 & ~ys__n546;
  assign new_n45793_ = new_n45791_ & new_n45792_;
  assign new_n45794_ = ~ys__n544 & ~ys__n546;
  assign new_n45795_ = ~new_n45790_ & new_n45794_;
  assign new_n45796_ = ~new_n45788_ & new_n45795_;
  assign new_n45797_ = ~new_n45793_ & ~new_n45796_;
  assign new_n45798_ = new_n45790_ & new_n45794_;
  assign new_n45799_ = new_n45788_ & new_n45798_;
  assign new_n45800_ = ~new_n45796_ & ~new_n45799_;
  assign new_n45801_ = ~ys__n544 & ys__n546;
  assign new_n45802_ = new_n45791_ & new_n45801_;
  assign new_n45803_ = ~new_n45793_ & ~new_n45802_;
  assign ys__n32024 = ~new_n45800_ | ~new_n45803_;
  assign ys__n32022 = ~new_n45797_ & ys__n32024;
  assign ys__n32023 = ~new_n45800_ & ys__n32024;
  assign new_n45807_ = ys__n47692 & ~new_n13759_;
  assign new_n45808_ = ys__n47723 & new_n13760_;
  assign new_n45809_ = ~new_n45807_ & ~new_n45808_;
  assign ys__n32025 = ~new_n13761_ & ~new_n45809_;
  assign new_n45811_ = ys__n47693 & ~new_n13759_;
  assign new_n45812_ = ys__n47724 & new_n13760_;
  assign new_n45813_ = ~new_n45811_ & ~new_n45812_;
  assign ys__n32026 = ~new_n13761_ & ~new_n45813_;
  assign new_n45815_ = ys__n47694 & ~new_n13759_;
  assign new_n45816_ = ys__n47725 & new_n13760_;
  assign new_n45817_ = ~new_n45815_ & ~new_n45816_;
  assign ys__n32027 = ~new_n13761_ & ~new_n45817_;
  assign new_n45819_ = ys__n47695 & ~new_n13759_;
  assign new_n45820_ = ys__n47726 & new_n13760_;
  assign new_n45821_ = ~new_n45819_ & ~new_n45820_;
  assign ys__n32028 = ~new_n13761_ & ~new_n45821_;
  assign new_n45823_ = ys__n47696 & ~new_n13759_;
  assign new_n45824_ = ys__n47727 & new_n13760_;
  assign new_n45825_ = ~new_n45823_ & ~new_n45824_;
  assign ys__n32029 = ~new_n13761_ & ~new_n45825_;
  assign new_n45827_ = ys__n47697 & ~new_n13759_;
  assign new_n45828_ = ys__n47728 & new_n13760_;
  assign new_n45829_ = ~new_n45827_ & ~new_n45828_;
  assign ys__n32030 = ~new_n13761_ & ~new_n45829_;
  assign new_n45831_ = ys__n47698 & ~new_n13759_;
  assign new_n45832_ = ys__n47729 & new_n13760_;
  assign new_n45833_ = ~new_n45831_ & ~new_n45832_;
  assign ys__n32031 = ~new_n13761_ & ~new_n45833_;
  assign new_n45835_ = ys__n47699 & ~new_n13759_;
  assign new_n45836_ = ys__n47730 & new_n13760_;
  assign new_n45837_ = ~new_n45835_ & ~new_n45836_;
  assign ys__n32032 = ~new_n13761_ & ~new_n45837_;
  assign new_n45839_ = ys__n47700 & ~new_n13759_;
  assign new_n45840_ = ys__n47731 & new_n13760_;
  assign new_n45841_ = ~new_n45839_ & ~new_n45840_;
  assign ys__n32033 = ~new_n13761_ & ~new_n45841_;
  assign new_n45843_ = ys__n47701 & ~new_n13759_;
  assign new_n45844_ = ys__n47732 & new_n13760_;
  assign new_n45845_ = ~new_n45843_ & ~new_n45844_;
  assign ys__n32034 = ~new_n13761_ & ~new_n45845_;
  assign new_n45847_ = ys__n47702 & ~new_n13759_;
  assign new_n45848_ = ys__n47733 & new_n13760_;
  assign new_n45849_ = ~new_n45847_ & ~new_n45848_;
  assign ys__n32035 = ~new_n13761_ & ~new_n45849_;
  assign new_n45851_ = ys__n47703 & ~new_n13759_;
  assign new_n45852_ = ys__n47734 & new_n13760_;
  assign new_n45853_ = ~new_n45851_ & ~new_n45852_;
  assign ys__n32036 = ~new_n13761_ & ~new_n45853_;
  assign new_n45855_ = ys__n47704 & ~new_n13759_;
  assign new_n45856_ = ys__n47735 & new_n13760_;
  assign new_n45857_ = ~new_n45855_ & ~new_n45856_;
  assign ys__n32037 = ~new_n13761_ & ~new_n45857_;
  assign new_n45859_ = ys__n47705 & ~new_n13759_;
  assign new_n45860_ = ys__n47736 & new_n13760_;
  assign new_n45861_ = ~new_n45859_ & ~new_n45860_;
  assign ys__n32038 = ~new_n13761_ & ~new_n45861_;
  assign new_n45863_ = ys__n47706 & ~new_n13759_;
  assign new_n45864_ = ys__n47737 & new_n13760_;
  assign new_n45865_ = ~new_n45863_ & ~new_n45864_;
  assign ys__n32039 = ~new_n13761_ & ~new_n45865_;
  assign new_n45867_ = ys__n47707 & ~new_n13759_;
  assign new_n45868_ = ys__n47738 & new_n13760_;
  assign new_n45869_ = ~new_n45867_ & ~new_n45868_;
  assign ys__n32040 = ~new_n13761_ & ~new_n45869_;
  assign new_n45871_ = ys__n47708 & ~new_n13759_;
  assign new_n45872_ = ys__n47739 & new_n13760_;
  assign new_n45873_ = ~new_n45871_ & ~new_n45872_;
  assign ys__n32041 = ~new_n13761_ & ~new_n45873_;
  assign new_n45875_ = ys__n47709 & ~new_n13759_;
  assign new_n45876_ = ys__n47740 & new_n13760_;
  assign new_n45877_ = ~new_n45875_ & ~new_n45876_;
  assign ys__n32042 = ~new_n13761_ & ~new_n45877_;
  assign new_n45879_ = ys__n47710 & ~new_n13759_;
  assign new_n45880_ = ys__n47741 & new_n13760_;
  assign new_n45881_ = ~new_n45879_ & ~new_n45880_;
  assign ys__n32043 = ~new_n13761_ & ~new_n45881_;
  assign new_n45883_ = ys__n47711 & ~new_n13759_;
  assign new_n45884_ = ys__n47742 & new_n13760_;
  assign new_n45885_ = ~new_n45883_ & ~new_n45884_;
  assign ys__n32044 = ~new_n13761_ & ~new_n45885_;
  assign new_n45887_ = ys__n47712 & ~new_n13759_;
  assign new_n45888_ = ys__n47743 & new_n13760_;
  assign new_n45889_ = ~new_n45887_ & ~new_n45888_;
  assign ys__n32045 = ~new_n13761_ & ~new_n45889_;
  assign new_n45891_ = ys__n47713 & ~new_n13759_;
  assign new_n45892_ = ys__n47744 & new_n13760_;
  assign new_n45893_ = ~new_n45891_ & ~new_n45892_;
  assign ys__n32046 = ~new_n13761_ & ~new_n45893_;
  assign new_n45895_ = ys__n47714 & ~new_n13759_;
  assign new_n45896_ = ys__n47745 & new_n13760_;
  assign new_n45897_ = ~new_n45895_ & ~new_n45896_;
  assign ys__n32047 = ~new_n13761_ & ~new_n45897_;
  assign new_n45899_ = ys__n47715 & ~new_n13759_;
  assign new_n45900_ = ys__n47746 & new_n13760_;
  assign new_n45901_ = ~new_n45899_ & ~new_n45900_;
  assign ys__n32048 = ~new_n13761_ & ~new_n45901_;
  assign new_n45903_ = ys__n47716 & ~new_n13759_;
  assign new_n45904_ = ys__n47747 & new_n13760_;
  assign new_n45905_ = ~new_n45903_ & ~new_n45904_;
  assign ys__n32049 = ~new_n13761_ & ~new_n45905_;
  assign new_n45907_ = ys__n47717 & ~new_n13759_;
  assign new_n45908_ = ys__n47748 & new_n13760_;
  assign new_n45909_ = ~new_n45907_ & ~new_n45908_;
  assign ys__n32050 = ~new_n13761_ & ~new_n45909_;
  assign new_n45911_ = ys__n47718 & ~new_n13759_;
  assign new_n45912_ = ys__n47749 & new_n13760_;
  assign new_n45913_ = ~new_n45911_ & ~new_n45912_;
  assign ys__n32051 = ~new_n13761_ & ~new_n45913_;
  assign new_n45915_ = ys__n47719 & ~new_n13759_;
  assign new_n45916_ = ys__n47750 & new_n13760_;
  assign new_n45917_ = ~new_n45915_ & ~new_n45916_;
  assign ys__n32052 = ~new_n13761_ & ~new_n45917_;
  assign new_n45919_ = ys__n47720 & ~new_n13759_;
  assign new_n45920_ = ys__n47751 & new_n13760_;
  assign new_n45921_ = ~new_n45919_ & ~new_n45920_;
  assign ys__n32053 = ~new_n13761_ & ~new_n45921_;
  assign new_n45923_ = ys__n47721 & ~new_n13759_;
  assign new_n45924_ = ys__n47752 & new_n13760_;
  assign new_n45925_ = ~new_n45923_ & ~new_n45924_;
  assign ys__n32054 = ~new_n13761_ & ~new_n45925_;
  assign new_n45927_ = ys__n47722 & ~new_n13759_;
  assign new_n45928_ = ys__n47753 & new_n13760_;
  assign new_n45929_ = ~new_n45927_ & ~new_n45928_;
  assign ys__n32055 = ~new_n13761_ & ~new_n45929_;
  assign new_n45931_ = ys__n38323 & ~new_n13759_;
  assign new_n45932_ = ys__n47754 & new_n13760_;
  assign new_n45933_ = ~new_n45931_ & ~new_n45932_;
  assign ys__n32056 = ~new_n13761_ & ~new_n45933_;
  assign new_n45935_ = ~ys__n935 & new_n13431_;
  assign new_n45936_ = ys__n28462 & new_n45935_;
  assign new_n45937_ = ~ys__n226 & ys__n935;
  assign new_n45938_ = new_n13437_ & new_n45937_;
  assign new_n45939_ = ys__n23077 & new_n45938_;
  assign new_n45940_ = ys__n226 & ys__n935;
  assign new_n45941_ = ys__n22918 & new_n45940_;
  assign new_n45942_ = ~new_n13437_ & new_n45937_;
  assign new_n45943_ = ys__n23014 & new_n45942_;
  assign new_n45944_ = ~new_n45941_ & ~new_n45943_;
  assign new_n45945_ = ~new_n45939_ & new_n45944_;
  assign new_n45946_ = ~new_n45936_ & new_n45945_;
  assign new_n45947_ = ~new_n45940_ & ~new_n45942_;
  assign new_n45948_ = ~new_n45938_ & new_n45947_;
  assign new_n45949_ = ~new_n45935_ & new_n45948_;
  assign ys__n32057 = ~new_n45946_ & ~new_n45949_;
  assign new_n45951_ = ys__n28464 & new_n45935_;
  assign new_n45952_ = ys__n23078 & new_n45938_;
  assign new_n45953_ = ys__n22921 & new_n45940_;
  assign new_n45954_ = ys__n23016 & new_n45942_;
  assign new_n45955_ = ~new_n45953_ & ~new_n45954_;
  assign new_n45956_ = ~new_n45952_ & new_n45955_;
  assign new_n45957_ = ~new_n45951_ & new_n45956_;
  assign ys__n32058 = ~new_n45949_ & ~new_n45957_;
  assign new_n45959_ = ys__n28466 & new_n45935_;
  assign new_n45960_ = ys__n23079 & new_n45938_;
  assign new_n45961_ = ys__n22924 & new_n45940_;
  assign new_n45962_ = ys__n23018 & new_n45942_;
  assign new_n45963_ = ~new_n45961_ & ~new_n45962_;
  assign new_n45964_ = ~new_n45960_ & new_n45963_;
  assign new_n45965_ = ~new_n45959_ & new_n45964_;
  assign ys__n32059 = ~new_n45949_ & ~new_n45965_;
  assign new_n45967_ = ys__n28468 & new_n45935_;
  assign new_n45968_ = ys__n23080 & new_n45938_;
  assign new_n45969_ = ys__n22927 & new_n45940_;
  assign new_n45970_ = ys__n23020 & new_n45942_;
  assign new_n45971_ = ~new_n45969_ & ~new_n45970_;
  assign new_n45972_ = ~new_n45968_ & new_n45971_;
  assign new_n45973_ = ~new_n45967_ & new_n45972_;
  assign ys__n32060 = ~new_n45949_ & ~new_n45973_;
  assign new_n45975_ = ys__n28470 & new_n45935_;
  assign new_n45976_ = ys__n23081 & new_n45938_;
  assign new_n45977_ = ys__n22930 & new_n45940_;
  assign new_n45978_ = ys__n23022 & new_n45942_;
  assign new_n45979_ = ~new_n45977_ & ~new_n45978_;
  assign new_n45980_ = ~new_n45976_ & new_n45979_;
  assign new_n45981_ = ~new_n45975_ & new_n45980_;
  assign ys__n32061 = ~new_n45949_ & ~new_n45981_;
  assign new_n45983_ = ys__n28472 & new_n45935_;
  assign new_n45984_ = ys__n23082 & new_n45938_;
  assign new_n45985_ = ys__n22933 & new_n45940_;
  assign new_n45986_ = ys__n23024 & new_n45942_;
  assign new_n45987_ = ~new_n45985_ & ~new_n45986_;
  assign new_n45988_ = ~new_n45984_ & new_n45987_;
  assign new_n45989_ = ~new_n45983_ & new_n45988_;
  assign ys__n32062 = ~new_n45949_ & ~new_n45989_;
  assign new_n45991_ = ys__n29558 & new_n45935_;
  assign new_n45992_ = ys__n23083 & new_n45938_;
  assign new_n45993_ = ys__n22936 & new_n45940_;
  assign new_n45994_ = ys__n23026 & new_n45942_;
  assign new_n45995_ = ~new_n45993_ & ~new_n45994_;
  assign new_n45996_ = ~new_n45992_ & new_n45995_;
  assign new_n45997_ = ~new_n45991_ & new_n45996_;
  assign ys__n32063 = ~new_n45949_ & ~new_n45997_;
  assign new_n45999_ = ys__n29560 & new_n45935_;
  assign new_n46000_ = ys__n23084 & new_n45938_;
  assign new_n46001_ = ys__n22939 & new_n45940_;
  assign new_n46002_ = ys__n23028 & new_n45942_;
  assign new_n46003_ = ~new_n46001_ & ~new_n46002_;
  assign new_n46004_ = ~new_n46000_ & new_n46003_;
  assign new_n46005_ = ~new_n45999_ & new_n46004_;
  assign ys__n32064 = ~new_n45949_ & ~new_n46005_;
  assign new_n46007_ = ys__n29562 & new_n45935_;
  assign new_n46008_ = ys__n23085 & new_n45938_;
  assign new_n46009_ = ys__n22942 & new_n45940_;
  assign new_n46010_ = ys__n23030 & new_n45942_;
  assign new_n46011_ = ~new_n46009_ & ~new_n46010_;
  assign new_n46012_ = ~new_n46008_ & new_n46011_;
  assign new_n46013_ = ~new_n46007_ & new_n46012_;
  assign ys__n32065 = ~new_n45949_ & ~new_n46013_;
  assign new_n46015_ = ys__n29564 & new_n45935_;
  assign new_n46016_ = ys__n23086 & new_n45938_;
  assign new_n46017_ = ys__n22945 & new_n45940_;
  assign new_n46018_ = ys__n23032 & new_n45942_;
  assign new_n46019_ = ~new_n46017_ & ~new_n46018_;
  assign new_n46020_ = ~new_n46016_ & new_n46019_;
  assign new_n46021_ = ~new_n46015_ & new_n46020_;
  assign ys__n32066 = ~new_n45949_ & ~new_n46021_;
  assign new_n46023_ = ys__n29566 & new_n45935_;
  assign new_n46024_ = ys__n23087 & new_n45938_;
  assign new_n46025_ = ys__n22948 & new_n45940_;
  assign new_n46026_ = ys__n23034 & new_n45942_;
  assign new_n46027_ = ~new_n46025_ & ~new_n46026_;
  assign new_n46028_ = ~new_n46024_ & new_n46027_;
  assign new_n46029_ = ~new_n46023_ & new_n46028_;
  assign ys__n32067 = ~new_n45949_ & ~new_n46029_;
  assign new_n46031_ = ys__n29568 & new_n45935_;
  assign new_n46032_ = ys__n23088 & new_n45938_;
  assign new_n46033_ = ys__n22951 & new_n45940_;
  assign new_n46034_ = ys__n23036 & new_n45942_;
  assign new_n46035_ = ~new_n46033_ & ~new_n46034_;
  assign new_n46036_ = ~new_n46032_ & new_n46035_;
  assign new_n46037_ = ~new_n46031_ & new_n46036_;
  assign ys__n32068 = ~new_n45949_ & ~new_n46037_;
  assign new_n46039_ = ys__n29570 & new_n45935_;
  assign new_n46040_ = ys__n23089 & new_n45938_;
  assign new_n46041_ = ys__n22954 & new_n45940_;
  assign new_n46042_ = ys__n23038 & new_n45942_;
  assign new_n46043_ = ~new_n46041_ & ~new_n46042_;
  assign new_n46044_ = ~new_n46040_ & new_n46043_;
  assign new_n46045_ = ~new_n46039_ & new_n46044_;
  assign ys__n32069 = ~new_n45949_ & ~new_n46045_;
  assign new_n46047_ = ys__n29572 & new_n45935_;
  assign new_n46048_ = ys__n23090 & new_n45938_;
  assign new_n46049_ = ys__n22957 & new_n45940_;
  assign new_n46050_ = ys__n23040 & new_n45942_;
  assign new_n46051_ = ~new_n46049_ & ~new_n46050_;
  assign new_n46052_ = ~new_n46048_ & new_n46051_;
  assign new_n46053_ = ~new_n46047_ & new_n46052_;
  assign ys__n32070 = ~new_n45949_ & ~new_n46053_;
  assign new_n46055_ = ys__n29574 & new_n45935_;
  assign new_n46056_ = ys__n23091 & new_n45938_;
  assign new_n46057_ = ys__n22960 & new_n45940_;
  assign new_n46058_ = ys__n23042 & new_n45942_;
  assign new_n46059_ = ~new_n46057_ & ~new_n46058_;
  assign new_n46060_ = ~new_n46056_ & new_n46059_;
  assign new_n46061_ = ~new_n46055_ & new_n46060_;
  assign ys__n32071 = ~new_n45949_ & ~new_n46061_;
  assign new_n46063_ = ys__n29576 & new_n45935_;
  assign new_n46064_ = ys__n23092 & new_n45938_;
  assign new_n46065_ = ys__n22963 & new_n45940_;
  assign new_n46066_ = ys__n23044 & new_n45942_;
  assign new_n46067_ = ~new_n46065_ & ~new_n46066_;
  assign new_n46068_ = ~new_n46064_ & new_n46067_;
  assign new_n46069_ = ~new_n46063_ & new_n46068_;
  assign ys__n32072 = ~new_n45949_ & ~new_n46069_;
  assign new_n46071_ = ys__n29578 & new_n45935_;
  assign new_n46072_ = ys__n23093 & new_n45938_;
  assign new_n46073_ = ys__n22966 & new_n45940_;
  assign new_n46074_ = ys__n23046 & new_n45942_;
  assign new_n46075_ = ~new_n46073_ & ~new_n46074_;
  assign new_n46076_ = ~new_n46072_ & new_n46075_;
  assign new_n46077_ = ~new_n46071_ & new_n46076_;
  assign ys__n32073 = ~new_n45949_ & ~new_n46077_;
  assign new_n46079_ = ys__n29580 & new_n45935_;
  assign new_n46080_ = ys__n23094 & new_n45938_;
  assign new_n46081_ = ys__n22969 & new_n45940_;
  assign new_n46082_ = ys__n23048 & new_n45942_;
  assign new_n46083_ = ~new_n46081_ & ~new_n46082_;
  assign new_n46084_ = ~new_n46080_ & new_n46083_;
  assign new_n46085_ = ~new_n46079_ & new_n46084_;
  assign ys__n32074 = ~new_n45949_ & ~new_n46085_;
  assign new_n46087_ = ys__n29582 & new_n45935_;
  assign new_n46088_ = ys__n23095 & new_n45938_;
  assign new_n46089_ = ys__n22972 & new_n45940_;
  assign new_n46090_ = ys__n23050 & new_n45942_;
  assign new_n46091_ = ~new_n46089_ & ~new_n46090_;
  assign new_n46092_ = ~new_n46088_ & new_n46091_;
  assign new_n46093_ = ~new_n46087_ & new_n46092_;
  assign ys__n32075 = ~new_n45949_ & ~new_n46093_;
  assign new_n46095_ = ys__n29584 & new_n45935_;
  assign new_n46096_ = ys__n23096 & new_n45938_;
  assign new_n46097_ = ys__n22975 & new_n45940_;
  assign new_n46098_ = ys__n23052 & new_n45942_;
  assign new_n46099_ = ~new_n46097_ & ~new_n46098_;
  assign new_n46100_ = ~new_n46096_ & new_n46099_;
  assign new_n46101_ = ~new_n46095_ & new_n46100_;
  assign ys__n32076 = ~new_n45949_ & ~new_n46101_;
  assign new_n46103_ = ys__n29586 & new_n45935_;
  assign new_n46104_ = ys__n23097 & new_n45938_;
  assign new_n46105_ = ys__n22978 & new_n45940_;
  assign new_n46106_ = ys__n23054 & new_n45942_;
  assign new_n46107_ = ~new_n46105_ & ~new_n46106_;
  assign new_n46108_ = ~new_n46104_ & new_n46107_;
  assign new_n46109_ = ~new_n46103_ & new_n46108_;
  assign ys__n32077 = ~new_n45949_ & ~new_n46109_;
  assign new_n46111_ = ys__n29588 & new_n45935_;
  assign new_n46112_ = ys__n23098 & new_n45938_;
  assign new_n46113_ = ys__n22981 & new_n45940_;
  assign new_n46114_ = ys__n23056 & new_n45942_;
  assign new_n46115_ = ~new_n46113_ & ~new_n46114_;
  assign new_n46116_ = ~new_n46112_ & new_n46115_;
  assign new_n46117_ = ~new_n46111_ & new_n46116_;
  assign ys__n32078 = ~new_n45949_ & ~new_n46117_;
  assign new_n46119_ = ys__n29590 & new_n45935_;
  assign new_n46120_ = ys__n23099 & new_n45938_;
  assign new_n46121_ = ys__n22984 & new_n45940_;
  assign new_n46122_ = ys__n23058 & new_n45942_;
  assign new_n46123_ = ~new_n46121_ & ~new_n46122_;
  assign new_n46124_ = ~new_n46120_ & new_n46123_;
  assign new_n46125_ = ~new_n46119_ & new_n46124_;
  assign ys__n32079 = ~new_n45949_ & ~new_n46125_;
  assign new_n46127_ = ys__n29592 & new_n45935_;
  assign new_n46128_ = ys__n23100 & new_n45938_;
  assign new_n46129_ = ys__n22987 & new_n45940_;
  assign new_n46130_ = ys__n23060 & new_n45942_;
  assign new_n46131_ = ~new_n46129_ & ~new_n46130_;
  assign new_n46132_ = ~new_n46128_ & new_n46131_;
  assign new_n46133_ = ~new_n46127_ & new_n46132_;
  assign ys__n32080 = ~new_n45949_ & ~new_n46133_;
  assign new_n46135_ = ys__n29594 & new_n45935_;
  assign new_n46136_ = ys__n23101 & new_n45938_;
  assign new_n46137_ = ys__n22990 & new_n45940_;
  assign new_n46138_ = ys__n23062 & new_n45942_;
  assign new_n46139_ = ~new_n46137_ & ~new_n46138_;
  assign new_n46140_ = ~new_n46136_ & new_n46139_;
  assign new_n46141_ = ~new_n46135_ & new_n46140_;
  assign ys__n32081 = ~new_n45949_ & ~new_n46141_;
  assign new_n46143_ = ys__n29596 & new_n45935_;
  assign new_n46144_ = ys__n23102 & new_n45938_;
  assign new_n46145_ = ys__n22993 & new_n45940_;
  assign new_n46146_ = ys__n23064 & new_n45942_;
  assign new_n46147_ = ~new_n46145_ & ~new_n46146_;
  assign new_n46148_ = ~new_n46144_ & new_n46147_;
  assign new_n46149_ = ~new_n46143_ & new_n46148_;
  assign ys__n32082 = ~new_n45949_ & ~new_n46149_;
  assign new_n46151_ = ys__n29598 & new_n45935_;
  assign new_n46152_ = ys__n23103 & new_n45938_;
  assign new_n46153_ = ys__n22996 & new_n45940_;
  assign new_n46154_ = ys__n23066 & new_n45942_;
  assign new_n46155_ = ~new_n46153_ & ~new_n46154_;
  assign new_n46156_ = ~new_n46152_ & new_n46155_;
  assign new_n46157_ = ~new_n46151_ & new_n46156_;
  assign ys__n32083 = ~new_n45949_ & ~new_n46157_;
  assign new_n46159_ = ys__n29600 & new_n45935_;
  assign new_n46160_ = ys__n23104 & new_n45938_;
  assign new_n46161_ = ys__n22999 & new_n45940_;
  assign new_n46162_ = ys__n23068 & new_n45942_;
  assign new_n46163_ = ~new_n46161_ & ~new_n46162_;
  assign new_n46164_ = ~new_n46160_ & new_n46163_;
  assign new_n46165_ = ~new_n46159_ & new_n46164_;
  assign ys__n32084 = ~new_n45949_ & ~new_n46165_;
  assign new_n46167_ = ys__n29602 & new_n45935_;
  assign new_n46168_ = ys__n23105 & new_n45938_;
  assign new_n46169_ = ys__n23002 & new_n45940_;
  assign new_n46170_ = ys__n23070 & new_n45942_;
  assign new_n46171_ = ~new_n46169_ & ~new_n46170_;
  assign new_n46172_ = ~new_n46168_ & new_n46171_;
  assign new_n46173_ = ~new_n46167_ & new_n46172_;
  assign ys__n32085 = ~new_n45949_ & ~new_n46173_;
  assign new_n46175_ = ys__n29604 & new_n45935_;
  assign new_n46176_ = ys__n23106 & new_n45938_;
  assign new_n46177_ = ys__n23005 & new_n45940_;
  assign new_n46178_ = ys__n23072 & new_n45942_;
  assign new_n46179_ = ~new_n46177_ & ~new_n46178_;
  assign new_n46180_ = ~new_n46176_ & new_n46179_;
  assign new_n46181_ = ~new_n46175_ & new_n46180_;
  assign ys__n32086 = ~new_n45949_ & ~new_n46181_;
  assign new_n46183_ = ys__n29606 & new_n45935_;
  assign new_n46184_ = ys__n23107 & new_n45938_;
  assign new_n46185_ = ys__n23008 & new_n45940_;
  assign new_n46186_ = ys__n23074 & new_n45942_;
  assign new_n46187_ = ~new_n46185_ & ~new_n46186_;
  assign new_n46188_ = ~new_n46184_ & new_n46187_;
  assign new_n46189_ = ~new_n46183_ & new_n46188_;
  assign ys__n32087 = ~new_n45949_ & ~new_n46189_;
  assign new_n46191_ = ys__n29608 & new_n45935_;
  assign new_n46192_ = ys__n23108 & new_n45938_;
  assign new_n46193_ = ys__n23011 & new_n45940_;
  assign new_n46194_ = ys__n23076 & new_n45942_;
  assign new_n46195_ = ~new_n46193_ & ~new_n46194_;
  assign new_n46196_ = ~new_n46192_ & new_n46195_;
  assign new_n46197_ = ~new_n46191_ & new_n46196_;
  assign ys__n32088 = ~new_n45949_ & ~new_n46197_;
  assign new_n46199_ = ~new_n23757_ & ~new_n38778_;
  assign new_n46200_ = ~new_n24252_ & ~new_n46199_;
  assign new_n46201_ = ys__n38486 & new_n23752_;
  assign new_n46202_ = ~new_n46200_ & ~new_n46201_;
  assign new_n46203_ = ys__n27743 & new_n46201_;
  assign new_n46204_ = ~new_n46202_ & ~new_n46203_;
  assign new_n46205_ = ~ys__n278 & ~ys__n814;
  assign new_n46206_ = new_n13700_ & new_n46205_;
  assign new_n46207_ = ys__n20273 & ~ys__n250;
  assign new_n46208_ = ~ys__n252 & new_n46207_;
  assign new_n46209_ = new_n46206_ & new_n46208_;
  assign new_n46210_ = ys__n254 & new_n46209_;
  assign new_n46211_ = ~new_n46204_ & new_n46210_;
  assign new_n46212_ = ys__n20273 & ys__n250;
  assign new_n46213_ = new_n46206_ & new_n46212_;
  assign new_n46214_ = new_n13698_ & new_n46213_;
  assign new_n46215_ = ys__n19878 & new_n46214_;
  assign new_n46216_ = ys__n20956 & ~ys__n28243;
  assign new_n46217_ = ys__n21276 & ys__n28243;
  assign new_n46218_ = ~new_n46216_ & ~new_n46217_;
  assign new_n46219_ = ys__n28243 & ~new_n46218_;
  assign new_n46220_ = ~ys__n28243 & new_n46219_;
  assign new_n46221_ = ys__n21500 & ~ys__n28243;
  assign new_n46222_ = ys__n21820 & ys__n28243;
  assign new_n46223_ = ~new_n46221_ & ~new_n46222_;
  assign new_n46224_ = ~ys__n28243 & ~new_n46223_;
  assign new_n46225_ = ys__n21980 & ~ys__n28243;
  assign new_n46226_ = ys__n22300 & ys__n28243;
  assign new_n46227_ = ~new_n46225_ & ~new_n46226_;
  assign new_n46228_ = ys__n28243 & ~new_n46227_;
  assign new_n46229_ = ~new_n46224_ & ~new_n46228_;
  assign new_n46230_ = ys__n28243 & ~new_n46229_;
  assign new_n46231_ = ~new_n46220_ & ~new_n46230_;
  assign new_n46232_ = ys__n20273 & ~ys__n814;
  assign new_n46233_ = ys__n278 & new_n46232_;
  assign new_n46234_ = new_n13700_ & new_n46233_;
  assign new_n46235_ = new_n13699_ & new_n46234_;
  assign new_n46236_ = ~new_n46231_ & new_n46235_;
  assign new_n46237_ = ys__n252 & new_n46207_;
  assign new_n46238_ = new_n46206_ & new_n46237_;
  assign new_n46239_ = ~ys__n254 & new_n46238_;
  assign new_n46240_ = ys__n47791 & new_n46239_;
  assign new_n46241_ = ~new_n46236_ & ~new_n46240_;
  assign new_n46242_ = ys__n20273 & ~ys__n246;
  assign new_n46243_ = ys__n270 & new_n46242_;
  assign new_n46244_ = new_n46205_ & new_n46243_;
  assign new_n46245_ = new_n13699_ & new_n46244_;
  assign new_n46246_ = ys__n47759 & new_n46245_;
  assign new_n46247_ = ys__n464 & ~ys__n28243;
  assign new_n46248_ = ys__n28288 & ys__n28296;
  assign new_n46249_ = ys__n28243 & new_n46248_;
  assign new_n46250_ = ~new_n46247_ & ~new_n46249_;
  assign new_n46251_ = ys__n20273 & ys__n246;
  assign new_n46252_ = ~ys__n270 & new_n46251_;
  assign new_n46253_ = new_n46205_ & new_n46252_;
  assign new_n46254_ = new_n13699_ & new_n46253_;
  assign new_n46255_ = ~new_n46250_ & new_n46254_;
  assign new_n46256_ = ~new_n46246_ & ~new_n46255_;
  assign new_n46257_ = new_n46241_ & new_n46256_;
  assign new_n46258_ = ~new_n46215_ & new_n46257_;
  assign new_n46259_ = ~new_n46211_ & new_n46258_;
  assign new_n46260_ = ~new_n46210_ & ~new_n46239_;
  assign new_n46261_ = ~new_n46214_ & new_n46260_;
  assign new_n46262_ = ~new_n46235_ & new_n46261_;
  assign new_n46263_ = ~ys__n20273 & new_n46206_;
  assign new_n46264_ = new_n13699_ & new_n46263_;
  assign new_n46265_ = ~new_n46245_ & ~new_n46254_;
  assign new_n46266_ = ~new_n46264_ & new_n46265_;
  assign new_n46267_ = new_n46262_ & new_n46266_;
  assign ys__n32124 = ~new_n46259_ & ~new_n46267_;
  assign new_n46269_ = ~new_n23757_ & ~new_n38787_;
  assign new_n46270_ = ~new_n24271_ & ~new_n46269_;
  assign new_n46271_ = ~new_n46201_ & ~new_n46270_;
  assign new_n46272_ = ys__n27747 & new_n46201_;
  assign new_n46273_ = ~new_n46271_ & ~new_n46272_;
  assign new_n46274_ = new_n46210_ & ~new_n46273_;
  assign new_n46275_ = ys__n19881 & new_n46214_;
  assign new_n46276_ = ys__n20958 & ~ys__n28243;
  assign new_n46277_ = ys__n21278 & ys__n28243;
  assign new_n46278_ = ~new_n46276_ & ~new_n46277_;
  assign new_n46279_ = ys__n28243 & ~new_n46278_;
  assign new_n46280_ = ~ys__n28243 & new_n46279_;
  assign new_n46281_ = ys__n21502 & ~ys__n28243;
  assign new_n46282_ = ys__n21822 & ys__n28243;
  assign new_n46283_ = ~new_n46281_ & ~new_n46282_;
  assign new_n46284_ = ~ys__n28243 & ~new_n46283_;
  assign new_n46285_ = ys__n21982 & ~ys__n28243;
  assign new_n46286_ = ys__n22302 & ys__n28243;
  assign new_n46287_ = ~new_n46285_ & ~new_n46286_;
  assign new_n46288_ = ys__n28243 & ~new_n46287_;
  assign new_n46289_ = ~new_n46284_ & ~new_n46288_;
  assign new_n46290_ = ys__n28243 & ~new_n46289_;
  assign new_n46291_ = ~new_n46280_ & ~new_n46290_;
  assign new_n46292_ = new_n46235_ & ~new_n46291_;
  assign new_n46293_ = ys__n47792 & new_n46239_;
  assign new_n46294_ = ~new_n46292_ & ~new_n46293_;
  assign new_n46295_ = ys__n47760 & new_n46245_;
  assign new_n46296_ = ys__n4340 & ~ys__n28243;
  assign new_n46297_ = ys__n28287 & ys__n28288;
  assign new_n46298_ = ys__n28243 & new_n46297_;
  assign new_n46299_ = ~new_n46296_ & ~new_n46298_;
  assign new_n46300_ = new_n46254_ & ~new_n46299_;
  assign new_n46301_ = ~new_n46295_ & ~new_n46300_;
  assign new_n46302_ = new_n46294_ & new_n46301_;
  assign new_n46303_ = ~new_n46275_ & new_n46302_;
  assign new_n46304_ = ~new_n46274_ & new_n46303_;
  assign ys__n32125 = ~new_n46267_ & ~new_n46304_;
  assign new_n46306_ = ~new_n23757_ & ~new_n38795_;
  assign new_n46307_ = ~new_n24290_ & ~new_n46306_;
  assign new_n46308_ = ~new_n46201_ & ~new_n46307_;
  assign new_n46309_ = ys__n27750 & new_n46201_;
  assign new_n46310_ = ~new_n46308_ & ~new_n46309_;
  assign new_n46311_ = new_n46210_ & ~new_n46310_;
  assign new_n46312_ = ys__n19884 & new_n46214_;
  assign new_n46313_ = ys__n20960 & ~ys__n28243;
  assign new_n46314_ = ys__n21280 & ys__n28243;
  assign new_n46315_ = ~new_n46313_ & ~new_n46314_;
  assign new_n46316_ = ys__n28243 & ~new_n46315_;
  assign new_n46317_ = ~ys__n28243 & new_n46316_;
  assign new_n46318_ = ys__n21504 & ~ys__n28243;
  assign new_n46319_ = ys__n21824 & ys__n28243;
  assign new_n46320_ = ~new_n46318_ & ~new_n46319_;
  assign new_n46321_ = ~ys__n28243 & ~new_n46320_;
  assign new_n46322_ = ys__n21984 & ~ys__n28243;
  assign new_n46323_ = ys__n22304 & ys__n28243;
  assign new_n46324_ = ~new_n46322_ & ~new_n46323_;
  assign new_n46325_ = ys__n28243 & ~new_n46324_;
  assign new_n46326_ = ~new_n46321_ & ~new_n46325_;
  assign new_n46327_ = ys__n28243 & ~new_n46326_;
  assign new_n46328_ = ~new_n46317_ & ~new_n46327_;
  assign new_n46329_ = new_n46235_ & ~new_n46328_;
  assign new_n46330_ = ys__n47793 & new_n46239_;
  assign new_n46331_ = ~new_n46329_ & ~new_n46330_;
  assign new_n46332_ = ys__n47761 & new_n46245_;
  assign new_n46333_ = ys__n240 & ~ys__n28243;
  assign new_n46334_ = ys__n464 & ~ys__n28288;
  assign new_n46335_ = ys__n28288 & ys__n28290;
  assign new_n46336_ = ~new_n46334_ & ~new_n46335_;
  assign new_n46337_ = ys__n28243 & ~new_n46336_;
  assign new_n46338_ = ~new_n46333_ & ~new_n46337_;
  assign new_n46339_ = new_n46254_ & ~new_n46338_;
  assign new_n46340_ = ~new_n46332_ & ~new_n46339_;
  assign new_n46341_ = new_n46331_ & new_n46340_;
  assign new_n46342_ = ~new_n46312_ & new_n46341_;
  assign new_n46343_ = ~new_n46311_ & new_n46342_;
  assign ys__n32126 = ~new_n46267_ & ~new_n46343_;
  assign new_n46345_ = ~new_n23757_ & ~new_n38803_;
  assign new_n46346_ = ~new_n24309_ & ~new_n46345_;
  assign new_n46347_ = ~new_n46201_ & ~new_n46346_;
  assign new_n46348_ = ys__n27753 & new_n46201_;
  assign new_n46349_ = ~new_n46347_ & ~new_n46348_;
  assign new_n46350_ = new_n46210_ & ~new_n46349_;
  assign new_n46351_ = ys__n19887 & new_n46214_;
  assign new_n46352_ = ys__n20962 & ~ys__n28243;
  assign new_n46353_ = ys__n21282 & ys__n28243;
  assign new_n46354_ = ~new_n46352_ & ~new_n46353_;
  assign new_n46355_ = ys__n28243 & ~new_n46354_;
  assign new_n46356_ = ~ys__n28243 & new_n46355_;
  assign new_n46357_ = ys__n21506 & ~ys__n28243;
  assign new_n46358_ = ys__n21826 & ys__n28243;
  assign new_n46359_ = ~new_n46357_ & ~new_n46358_;
  assign new_n46360_ = ~ys__n28243 & ~new_n46359_;
  assign new_n46361_ = ys__n21986 & ~ys__n28243;
  assign new_n46362_ = ys__n22306 & ys__n28243;
  assign new_n46363_ = ~new_n46361_ & ~new_n46362_;
  assign new_n46364_ = ys__n28243 & ~new_n46363_;
  assign new_n46365_ = ~new_n46360_ & ~new_n46364_;
  assign new_n46366_ = ys__n28243 & ~new_n46365_;
  assign new_n46367_ = ~new_n46356_ & ~new_n46366_;
  assign new_n46368_ = new_n46235_ & ~new_n46367_;
  assign new_n46369_ = ys__n47794 & new_n46239_;
  assign new_n46370_ = ~new_n46368_ & ~new_n46369_;
  assign new_n46371_ = ys__n47762 & new_n46245_;
  assign new_n46372_ = ys__n238 & ~ys__n28243;
  assign new_n46373_ = ys__n4340 & ~ys__n28288;
  assign new_n46374_ = ys__n28288 & ys__n28292;
  assign new_n46375_ = ~new_n46373_ & ~new_n46374_;
  assign new_n46376_ = ys__n28243 & ~new_n46375_;
  assign new_n46377_ = ~new_n46372_ & ~new_n46376_;
  assign new_n46378_ = new_n46254_ & ~new_n46377_;
  assign new_n46379_ = ~new_n46371_ & ~new_n46378_;
  assign new_n46380_ = new_n46370_ & new_n46379_;
  assign new_n46381_ = ~new_n46351_ & new_n46380_;
  assign new_n46382_ = ~new_n46350_ & new_n46381_;
  assign ys__n32127 = ~new_n46267_ & ~new_n46382_;
  assign new_n46384_ = ~new_n23757_ & ~new_n38811_;
  assign new_n46385_ = ~new_n24328_ & ~new_n46384_;
  assign new_n46386_ = ~new_n46201_ & ~new_n46385_;
  assign new_n46387_ = ys__n27756 & new_n46201_;
  assign new_n46388_ = ~new_n46386_ & ~new_n46387_;
  assign new_n46389_ = new_n46210_ & ~new_n46388_;
  assign new_n46390_ = ys__n19890 & new_n46214_;
  assign new_n46391_ = ys__n20964 & ~ys__n28243;
  assign new_n46392_ = ys__n21284 & ys__n28243;
  assign new_n46393_ = ~new_n46391_ & ~new_n46392_;
  assign new_n46394_ = ys__n28243 & ~new_n46393_;
  assign new_n46395_ = ~ys__n28243 & new_n46394_;
  assign new_n46396_ = ys__n21508 & ~ys__n28243;
  assign new_n46397_ = ys__n21828 & ys__n28243;
  assign new_n46398_ = ~new_n46396_ & ~new_n46397_;
  assign new_n46399_ = ~ys__n28243 & ~new_n46398_;
  assign new_n46400_ = ys__n21988 & ~ys__n28243;
  assign new_n46401_ = ys__n22308 & ys__n28243;
  assign new_n46402_ = ~new_n46400_ & ~new_n46401_;
  assign new_n46403_ = ys__n28243 & ~new_n46402_;
  assign new_n46404_ = ~new_n46399_ & ~new_n46403_;
  assign new_n46405_ = ys__n28243 & ~new_n46404_;
  assign new_n46406_ = ~new_n46395_ & ~new_n46405_;
  assign new_n46407_ = new_n46235_ & ~new_n46406_;
  assign new_n46408_ = ys__n47795 & new_n46239_;
  assign new_n46409_ = ~new_n46407_ & ~new_n46408_;
  assign new_n46410_ = ys__n47763 & new_n46245_;
  assign new_n46411_ = ys__n242 & ~ys__n28243;
  assign new_n46412_ = ys__n28288 & ys__n28294;
  assign new_n46413_ = ys__n28243 & new_n46412_;
  assign new_n46414_ = ~new_n46411_ & ~new_n46413_;
  assign new_n46415_ = new_n46254_ & ~new_n46414_;
  assign new_n46416_ = ~new_n46410_ & ~new_n46415_;
  assign new_n46417_ = new_n46409_ & new_n46416_;
  assign new_n46418_ = ~new_n46390_ & new_n46417_;
  assign new_n46419_ = ~new_n46389_ & new_n46418_;
  assign ys__n32128 = ~new_n46267_ & ~new_n46419_;
  assign new_n46421_ = ~new_n23757_ & ~new_n38819_;
  assign new_n46422_ = ~new_n24347_ & ~new_n46421_;
  assign new_n46423_ = ~new_n46201_ & ~new_n46422_;
  assign new_n46424_ = ys__n27759 & new_n46201_;
  assign new_n46425_ = ~new_n46423_ & ~new_n46424_;
  assign new_n46426_ = new_n46210_ & ~new_n46425_;
  assign new_n46427_ = ys__n19893 & new_n46214_;
  assign new_n46428_ = ys__n47764 & new_n46245_;
  assign new_n46429_ = ys__n20966 & ~ys__n28243;
  assign new_n46430_ = ys__n21286 & ys__n28243;
  assign new_n46431_ = ~new_n46429_ & ~new_n46430_;
  assign new_n46432_ = ys__n28243 & ~new_n46431_;
  assign new_n46433_ = ~ys__n28243 & new_n46432_;
  assign new_n46434_ = ys__n21510 & ~ys__n28243;
  assign new_n46435_ = ys__n21830 & ys__n28243;
  assign new_n46436_ = ~new_n46434_ & ~new_n46435_;
  assign new_n46437_ = ~ys__n28243 & ~new_n46436_;
  assign new_n46438_ = ys__n21990 & ~ys__n28243;
  assign new_n46439_ = ys__n22310 & ys__n28243;
  assign new_n46440_ = ~new_n46438_ & ~new_n46439_;
  assign new_n46441_ = ys__n28243 & ~new_n46440_;
  assign new_n46442_ = ~new_n46437_ & ~new_n46441_;
  assign new_n46443_ = ys__n28243 & ~new_n46442_;
  assign new_n46444_ = ~new_n46433_ & ~new_n46443_;
  assign new_n46445_ = new_n46235_ & ~new_n46444_;
  assign new_n46446_ = ys__n47796 & new_n46239_;
  assign new_n46447_ = ~new_n46445_ & ~new_n46446_;
  assign new_n46448_ = ~new_n46428_ & new_n46447_;
  assign new_n46449_ = ~new_n46427_ & new_n46448_;
  assign new_n46450_ = ~new_n46426_ & new_n46449_;
  assign ys__n32129 = ~new_n46267_ & ~new_n46450_;
  assign new_n46452_ = ~new_n23757_ & ~new_n38827_;
  assign new_n46453_ = ~new_n24366_ & ~new_n46452_;
  assign new_n46454_ = ~new_n46201_ & ~new_n46453_;
  assign new_n46455_ = ys__n27762 & new_n46201_;
  assign new_n46456_ = ~new_n46454_ & ~new_n46455_;
  assign new_n46457_ = new_n46210_ & ~new_n46456_;
  assign new_n46458_ = ys__n19896 & new_n46214_;
  assign new_n46459_ = ys__n47765 & new_n46245_;
  assign new_n46460_ = ys__n20968 & ~ys__n28243;
  assign new_n46461_ = ys__n21288 & ys__n28243;
  assign new_n46462_ = ~new_n46460_ & ~new_n46461_;
  assign new_n46463_ = ys__n28243 & ~new_n46462_;
  assign new_n46464_ = ~ys__n28243 & new_n46463_;
  assign new_n46465_ = ys__n21512 & ~ys__n28243;
  assign new_n46466_ = ys__n21832 & ys__n28243;
  assign new_n46467_ = ~new_n46465_ & ~new_n46466_;
  assign new_n46468_ = ~ys__n28243 & ~new_n46467_;
  assign new_n46469_ = ys__n21992 & ~ys__n28243;
  assign new_n46470_ = ys__n22312 & ys__n28243;
  assign new_n46471_ = ~new_n46469_ & ~new_n46470_;
  assign new_n46472_ = ys__n28243 & ~new_n46471_;
  assign new_n46473_ = ~new_n46468_ & ~new_n46472_;
  assign new_n46474_ = ys__n28243 & ~new_n46473_;
  assign new_n46475_ = ~new_n46464_ & ~new_n46474_;
  assign new_n46476_ = new_n46235_ & ~new_n46475_;
  assign new_n46477_ = ys__n47797 & new_n46239_;
  assign new_n46478_ = ~new_n46476_ & ~new_n46477_;
  assign new_n46479_ = ~new_n46459_ & new_n46478_;
  assign new_n46480_ = ~new_n46458_ & new_n46479_;
  assign new_n46481_ = ~new_n46457_ & new_n46480_;
  assign ys__n32130 = ~new_n46267_ & ~new_n46481_;
  assign new_n46483_ = ~new_n23757_ & ~new_n38835_;
  assign new_n46484_ = ~new_n24385_ & ~new_n46483_;
  assign new_n46485_ = ~new_n46201_ & ~new_n46484_;
  assign new_n46486_ = ys__n27765 & new_n46201_;
  assign new_n46487_ = ~new_n46485_ & ~new_n46486_;
  assign new_n46488_ = new_n46210_ & ~new_n46487_;
  assign new_n46489_ = ys__n19899 & new_n46214_;
  assign new_n46490_ = ys__n47766 & new_n46245_;
  assign new_n46491_ = ys__n20970 & ~ys__n28243;
  assign new_n46492_ = ys__n21290 & ys__n28243;
  assign new_n46493_ = ~new_n46491_ & ~new_n46492_;
  assign new_n46494_ = ys__n28243 & ~new_n46493_;
  assign new_n46495_ = ~ys__n28243 & new_n46494_;
  assign new_n46496_ = ys__n21514 & ~ys__n28243;
  assign new_n46497_ = ys__n21834 & ys__n28243;
  assign new_n46498_ = ~new_n46496_ & ~new_n46497_;
  assign new_n46499_ = ~ys__n28243 & ~new_n46498_;
  assign new_n46500_ = ys__n21994 & ~ys__n28243;
  assign new_n46501_ = ys__n22314 & ys__n28243;
  assign new_n46502_ = ~new_n46500_ & ~new_n46501_;
  assign new_n46503_ = ys__n28243 & ~new_n46502_;
  assign new_n46504_ = ~new_n46499_ & ~new_n46503_;
  assign new_n46505_ = ys__n28243 & ~new_n46504_;
  assign new_n46506_ = ~new_n46495_ & ~new_n46505_;
  assign new_n46507_ = new_n46235_ & ~new_n46506_;
  assign new_n46508_ = ys__n47798 & new_n46239_;
  assign new_n46509_ = ~new_n46507_ & ~new_n46508_;
  assign new_n46510_ = ~new_n46490_ & new_n46509_;
  assign new_n46511_ = ~new_n46489_ & new_n46510_;
  assign new_n46512_ = ~new_n46488_ & new_n46511_;
  assign ys__n32131 = ~new_n46267_ & ~new_n46512_;
  assign new_n46514_ = ~new_n23757_ & ~new_n38843_;
  assign new_n46515_ = ~new_n24066_ & ~new_n46514_;
  assign new_n46516_ = ~new_n46201_ & ~new_n46515_;
  assign new_n46517_ = ys__n27768 & new_n46201_;
  assign new_n46518_ = ~new_n46516_ & ~new_n46517_;
  assign new_n46519_ = new_n46210_ & ~new_n46518_;
  assign new_n46520_ = ys__n19902 & new_n46214_;
  assign new_n46521_ = ys__n47767 & new_n46245_;
  assign new_n46522_ = ys__n20972 & ~ys__n28243;
  assign new_n46523_ = ys__n21292 & ys__n28243;
  assign new_n46524_ = ~new_n46522_ & ~new_n46523_;
  assign new_n46525_ = ys__n28243 & ~new_n46524_;
  assign new_n46526_ = ~ys__n28243 & new_n46525_;
  assign new_n46527_ = ys__n21516 & ~ys__n28243;
  assign new_n46528_ = ys__n21836 & ys__n28243;
  assign new_n46529_ = ~new_n46527_ & ~new_n46528_;
  assign new_n46530_ = ~ys__n28243 & ~new_n46529_;
  assign new_n46531_ = ys__n21996 & ~ys__n28243;
  assign new_n46532_ = ys__n22316 & ys__n28243;
  assign new_n46533_ = ~new_n46531_ & ~new_n46532_;
  assign new_n46534_ = ys__n28243 & ~new_n46533_;
  assign new_n46535_ = ~new_n46530_ & ~new_n46534_;
  assign new_n46536_ = ys__n28243 & ~new_n46535_;
  assign new_n46537_ = ~new_n46526_ & ~new_n46536_;
  assign new_n46538_ = new_n46235_ & ~new_n46537_;
  assign new_n46539_ = ys__n47799 & new_n46239_;
  assign new_n46540_ = ~new_n46538_ & ~new_n46539_;
  assign new_n46541_ = ~new_n46521_ & new_n46540_;
  assign new_n46542_ = ~new_n46520_ & new_n46541_;
  assign new_n46543_ = ~new_n46519_ & new_n46542_;
  assign ys__n32132 = ~new_n46267_ & ~new_n46543_;
  assign new_n46545_ = ~new_n23757_ & ~new_n38851_;
  assign new_n46546_ = ~new_n24084_ & ~new_n46545_;
  assign new_n46547_ = ~new_n46201_ & ~new_n46546_;
  assign new_n46548_ = ys__n27771 & new_n46201_;
  assign new_n46549_ = ~new_n46547_ & ~new_n46548_;
  assign new_n46550_ = new_n46210_ & ~new_n46549_;
  assign new_n46551_ = ys__n19905 & new_n46214_;
  assign new_n46552_ = ys__n47768 & new_n46245_;
  assign new_n46553_ = ys__n20974 & ~ys__n28243;
  assign new_n46554_ = ys__n21294 & ys__n28243;
  assign new_n46555_ = ~new_n46553_ & ~new_n46554_;
  assign new_n46556_ = ys__n28243 & ~new_n46555_;
  assign new_n46557_ = ~ys__n28243 & new_n46556_;
  assign new_n46558_ = ys__n21518 & ~ys__n28243;
  assign new_n46559_ = ys__n21838 & ys__n28243;
  assign new_n46560_ = ~new_n46558_ & ~new_n46559_;
  assign new_n46561_ = ~ys__n28243 & ~new_n46560_;
  assign new_n46562_ = ys__n21998 & ~ys__n28243;
  assign new_n46563_ = ys__n22318 & ys__n28243;
  assign new_n46564_ = ~new_n46562_ & ~new_n46563_;
  assign new_n46565_ = ys__n28243 & ~new_n46564_;
  assign new_n46566_ = ~new_n46561_ & ~new_n46565_;
  assign new_n46567_ = ys__n28243 & ~new_n46566_;
  assign new_n46568_ = ~new_n46557_ & ~new_n46567_;
  assign new_n46569_ = new_n46235_ & ~new_n46568_;
  assign new_n46570_ = ys__n47800 & new_n46239_;
  assign new_n46571_ = ~new_n46569_ & ~new_n46570_;
  assign new_n46572_ = ~new_n46552_ & new_n46571_;
  assign new_n46573_ = ~new_n46551_ & new_n46572_;
  assign new_n46574_ = ~new_n46550_ & new_n46573_;
  assign ys__n32133 = ~new_n46267_ & ~new_n46574_;
  assign new_n46576_ = ~new_n23757_ & ~new_n38859_;
  assign new_n46577_ = ~new_n24102_ & ~new_n46576_;
  assign new_n46578_ = ~new_n46201_ & ~new_n46577_;
  assign new_n46579_ = ys__n27774 & new_n46201_;
  assign new_n46580_ = ~new_n46578_ & ~new_n46579_;
  assign new_n46581_ = new_n46210_ & ~new_n46580_;
  assign new_n46582_ = ys__n19908 & new_n46214_;
  assign new_n46583_ = ys__n47769 & new_n46245_;
  assign new_n46584_ = ys__n20976 & ~ys__n28243;
  assign new_n46585_ = ys__n21296 & ys__n28243;
  assign new_n46586_ = ~new_n46584_ & ~new_n46585_;
  assign new_n46587_ = ys__n28243 & ~new_n46586_;
  assign new_n46588_ = ~ys__n28243 & new_n46587_;
  assign new_n46589_ = ys__n21520 & ~ys__n28243;
  assign new_n46590_ = ys__n21840 & ys__n28243;
  assign new_n46591_ = ~new_n46589_ & ~new_n46590_;
  assign new_n46592_ = ~ys__n28243 & ~new_n46591_;
  assign new_n46593_ = ys__n22000 & ~ys__n28243;
  assign new_n46594_ = ys__n22320 & ys__n28243;
  assign new_n46595_ = ~new_n46593_ & ~new_n46594_;
  assign new_n46596_ = ys__n28243 & ~new_n46595_;
  assign new_n46597_ = ~new_n46592_ & ~new_n46596_;
  assign new_n46598_ = ys__n28243 & ~new_n46597_;
  assign new_n46599_ = ~new_n46588_ & ~new_n46598_;
  assign new_n46600_ = new_n46235_ & ~new_n46599_;
  assign new_n46601_ = ys__n47801 & new_n46239_;
  assign new_n46602_ = ~new_n46600_ & ~new_n46601_;
  assign new_n46603_ = ~new_n46583_ & new_n46602_;
  assign new_n46604_ = ~new_n46582_ & new_n46603_;
  assign new_n46605_ = ~new_n46581_ & new_n46604_;
  assign ys__n32134 = ~new_n46267_ & ~new_n46605_;
  assign new_n46607_ = ~new_n23757_ & ~new_n38867_;
  assign new_n46608_ = ~new_n24120_ & ~new_n46607_;
  assign new_n46609_ = ~new_n46201_ & ~new_n46608_;
  assign new_n46610_ = ys__n27777 & new_n46201_;
  assign new_n46611_ = ~new_n46609_ & ~new_n46610_;
  assign new_n46612_ = new_n46210_ & ~new_n46611_;
  assign new_n46613_ = ys__n19911 & new_n46214_;
  assign new_n46614_ = ys__n47770 & new_n46245_;
  assign new_n46615_ = ys__n20978 & ~ys__n28243;
  assign new_n46616_ = ys__n21298 & ys__n28243;
  assign new_n46617_ = ~new_n46615_ & ~new_n46616_;
  assign new_n46618_ = ys__n28243 & ~new_n46617_;
  assign new_n46619_ = ~ys__n28243 & new_n46618_;
  assign new_n46620_ = ys__n21522 & ~ys__n28243;
  assign new_n46621_ = ys__n21842 & ys__n28243;
  assign new_n46622_ = ~new_n46620_ & ~new_n46621_;
  assign new_n46623_ = ~ys__n28243 & ~new_n46622_;
  assign new_n46624_ = ys__n22002 & ~ys__n28243;
  assign new_n46625_ = ys__n22322 & ys__n28243;
  assign new_n46626_ = ~new_n46624_ & ~new_n46625_;
  assign new_n46627_ = ys__n28243 & ~new_n46626_;
  assign new_n46628_ = ~new_n46623_ & ~new_n46627_;
  assign new_n46629_ = ys__n28243 & ~new_n46628_;
  assign new_n46630_ = ~new_n46619_ & ~new_n46629_;
  assign new_n46631_ = new_n46235_ & ~new_n46630_;
  assign new_n46632_ = ys__n47802 & new_n46239_;
  assign new_n46633_ = ~new_n46631_ & ~new_n46632_;
  assign new_n46634_ = ~new_n46614_ & new_n46633_;
  assign new_n46635_ = ~new_n46613_ & new_n46634_;
  assign new_n46636_ = ~new_n46612_ & new_n46635_;
  assign ys__n32135 = ~new_n46267_ & ~new_n46636_;
  assign new_n46638_ = ~new_n23757_ & ~new_n38875_;
  assign new_n46639_ = ~new_n24138_ & ~new_n46638_;
  assign new_n46640_ = ~new_n46201_ & ~new_n46639_;
  assign new_n46641_ = ys__n27780 & new_n46201_;
  assign new_n46642_ = ~new_n46640_ & ~new_n46641_;
  assign new_n46643_ = new_n46210_ & ~new_n46642_;
  assign new_n46644_ = ys__n19914 & new_n46214_;
  assign new_n46645_ = ys__n47771 & new_n46245_;
  assign new_n46646_ = ys__n20980 & ~ys__n28243;
  assign new_n46647_ = ys__n21300 & ys__n28243;
  assign new_n46648_ = ~new_n46646_ & ~new_n46647_;
  assign new_n46649_ = ys__n28243 & ~new_n46648_;
  assign new_n46650_ = ~ys__n28243 & new_n46649_;
  assign new_n46651_ = ys__n21524 & ~ys__n28243;
  assign new_n46652_ = ys__n21844 & ys__n28243;
  assign new_n46653_ = ~new_n46651_ & ~new_n46652_;
  assign new_n46654_ = ~ys__n28243 & ~new_n46653_;
  assign new_n46655_ = ys__n22004 & ~ys__n28243;
  assign new_n46656_ = ys__n22324 & ys__n28243;
  assign new_n46657_ = ~new_n46655_ & ~new_n46656_;
  assign new_n46658_ = ys__n28243 & ~new_n46657_;
  assign new_n46659_ = ~new_n46654_ & ~new_n46658_;
  assign new_n46660_ = ys__n28243 & ~new_n46659_;
  assign new_n46661_ = ~new_n46650_ & ~new_n46660_;
  assign new_n46662_ = new_n46235_ & ~new_n46661_;
  assign new_n46663_ = ys__n47803 & new_n46239_;
  assign new_n46664_ = ~new_n46662_ & ~new_n46663_;
  assign new_n46665_ = ~new_n46645_ & new_n46664_;
  assign new_n46666_ = ~new_n46644_ & new_n46665_;
  assign new_n46667_ = ~new_n46643_ & new_n46666_;
  assign ys__n32136 = ~new_n46267_ & ~new_n46667_;
  assign new_n46669_ = ~new_n23757_ & ~new_n38883_;
  assign new_n46670_ = ~new_n24156_ & ~new_n46669_;
  assign new_n46671_ = ~new_n46201_ & ~new_n46670_;
  assign new_n46672_ = ys__n27783 & new_n46201_;
  assign new_n46673_ = ~new_n46671_ & ~new_n46672_;
  assign new_n46674_ = new_n46210_ & ~new_n46673_;
  assign new_n46675_ = ys__n19917 & new_n46214_;
  assign new_n46676_ = ys__n47772 & new_n46245_;
  assign new_n46677_ = ys__n20982 & ~ys__n28243;
  assign new_n46678_ = ys__n21302 & ys__n28243;
  assign new_n46679_ = ~new_n46677_ & ~new_n46678_;
  assign new_n46680_ = ys__n28243 & ~new_n46679_;
  assign new_n46681_ = ~ys__n28243 & new_n46680_;
  assign new_n46682_ = ys__n21526 & ~ys__n28243;
  assign new_n46683_ = ys__n21846 & ys__n28243;
  assign new_n46684_ = ~new_n46682_ & ~new_n46683_;
  assign new_n46685_ = ~ys__n28243 & ~new_n46684_;
  assign new_n46686_ = ys__n22006 & ~ys__n28243;
  assign new_n46687_ = ys__n22326 & ys__n28243;
  assign new_n46688_ = ~new_n46686_ & ~new_n46687_;
  assign new_n46689_ = ys__n28243 & ~new_n46688_;
  assign new_n46690_ = ~new_n46685_ & ~new_n46689_;
  assign new_n46691_ = ys__n28243 & ~new_n46690_;
  assign new_n46692_ = ~new_n46681_ & ~new_n46691_;
  assign new_n46693_ = new_n46235_ & ~new_n46692_;
  assign new_n46694_ = ys__n47804 & new_n46239_;
  assign new_n46695_ = ~new_n46693_ & ~new_n46694_;
  assign new_n46696_ = ~new_n46676_ & new_n46695_;
  assign new_n46697_ = ~new_n46675_ & new_n46696_;
  assign new_n46698_ = ~new_n46674_ & new_n46697_;
  assign ys__n32137 = ~new_n46267_ & ~new_n46698_;
  assign new_n46700_ = ~new_n23757_ & ~new_n38891_;
  assign new_n46701_ = ~new_n24174_ & ~new_n46700_;
  assign new_n46702_ = ~new_n46201_ & ~new_n46701_;
  assign new_n46703_ = ys__n27786 & new_n46201_;
  assign new_n46704_ = ~new_n46702_ & ~new_n46703_;
  assign new_n46705_ = new_n46210_ & ~new_n46704_;
  assign new_n46706_ = ys__n19920 & new_n46214_;
  assign new_n46707_ = ys__n47773 & new_n46245_;
  assign new_n46708_ = ys__n20984 & ~ys__n28243;
  assign new_n46709_ = ys__n21304 & ys__n28243;
  assign new_n46710_ = ~new_n46708_ & ~new_n46709_;
  assign new_n46711_ = ys__n28243 & ~new_n46710_;
  assign new_n46712_ = ~ys__n28243 & new_n46711_;
  assign new_n46713_ = ys__n21528 & ~ys__n28243;
  assign new_n46714_ = ys__n21848 & ys__n28243;
  assign new_n46715_ = ~new_n46713_ & ~new_n46714_;
  assign new_n46716_ = ~ys__n28243 & ~new_n46715_;
  assign new_n46717_ = ys__n22008 & ~ys__n28243;
  assign new_n46718_ = ys__n22328 & ys__n28243;
  assign new_n46719_ = ~new_n46717_ & ~new_n46718_;
  assign new_n46720_ = ys__n28243 & ~new_n46719_;
  assign new_n46721_ = ~new_n46716_ & ~new_n46720_;
  assign new_n46722_ = ys__n28243 & ~new_n46721_;
  assign new_n46723_ = ~new_n46712_ & ~new_n46722_;
  assign new_n46724_ = new_n46235_ & ~new_n46723_;
  assign new_n46725_ = ys__n47805 & new_n46239_;
  assign new_n46726_ = ~new_n46724_ & ~new_n46725_;
  assign new_n46727_ = ~new_n46707_ & new_n46726_;
  assign new_n46728_ = ~new_n46706_ & new_n46727_;
  assign new_n46729_ = ~new_n46705_ & new_n46728_;
  assign ys__n32138 = ~new_n46267_ & ~new_n46729_;
  assign new_n46731_ = ~new_n23757_ & ~new_n38899_;
  assign new_n46732_ = ~new_n24192_ & ~new_n46731_;
  assign new_n46733_ = ~new_n46201_ & ~new_n46732_;
  assign new_n46734_ = ys__n27789 & new_n46201_;
  assign new_n46735_ = ~new_n46733_ & ~new_n46734_;
  assign new_n46736_ = new_n46210_ & ~new_n46735_;
  assign new_n46737_ = ys__n19923 & new_n46214_;
  assign new_n46738_ = ys__n47774 & new_n46245_;
  assign new_n46739_ = ys__n20986 & ~ys__n28243;
  assign new_n46740_ = ys__n21306 & ys__n28243;
  assign new_n46741_ = ~new_n46739_ & ~new_n46740_;
  assign new_n46742_ = ys__n28243 & ~new_n46741_;
  assign new_n46743_ = ~ys__n28243 & new_n46742_;
  assign new_n46744_ = ys__n21530 & ~ys__n28243;
  assign new_n46745_ = ys__n21850 & ys__n28243;
  assign new_n46746_ = ~new_n46744_ & ~new_n46745_;
  assign new_n46747_ = ~ys__n28243 & ~new_n46746_;
  assign new_n46748_ = ys__n22010 & ~ys__n28243;
  assign new_n46749_ = ys__n22330 & ys__n28243;
  assign new_n46750_ = ~new_n46748_ & ~new_n46749_;
  assign new_n46751_ = ys__n28243 & ~new_n46750_;
  assign new_n46752_ = ~new_n46747_ & ~new_n46751_;
  assign new_n46753_ = ys__n28243 & ~new_n46752_;
  assign new_n46754_ = ~new_n46743_ & ~new_n46753_;
  assign new_n46755_ = new_n46235_ & ~new_n46754_;
  assign new_n46756_ = ys__n47806 & new_n46239_;
  assign new_n46757_ = ~new_n46755_ & ~new_n46756_;
  assign new_n46758_ = ~new_n46738_ & new_n46757_;
  assign new_n46759_ = ~new_n46737_ & new_n46758_;
  assign new_n46760_ = ~new_n46736_ & new_n46759_;
  assign ys__n32139 = ~new_n46267_ & ~new_n46760_;
  assign new_n46762_ = ~new_n23757_ & ~new_n38907_;
  assign new_n46763_ = ~new_n23906_ & ~new_n46762_;
  assign new_n46764_ = ~new_n46201_ & ~new_n46763_;
  assign new_n46765_ = ys__n27792 & new_n46201_;
  assign new_n46766_ = ~new_n46764_ & ~new_n46765_;
  assign new_n46767_ = new_n46210_ & ~new_n46766_;
  assign new_n46768_ = ys__n19926 & new_n46214_;
  assign new_n46769_ = ys__n47775 & new_n46245_;
  assign new_n46770_ = ys__n20988 & ~ys__n28243;
  assign new_n46771_ = ys__n21308 & ys__n28243;
  assign new_n46772_ = ~new_n46770_ & ~new_n46771_;
  assign new_n46773_ = ys__n28243 & ~new_n46772_;
  assign new_n46774_ = ~ys__n28243 & new_n46773_;
  assign new_n46775_ = ys__n21532 & ~ys__n28243;
  assign new_n46776_ = ys__n21852 & ys__n28243;
  assign new_n46777_ = ~new_n46775_ & ~new_n46776_;
  assign new_n46778_ = ~ys__n28243 & ~new_n46777_;
  assign new_n46779_ = ys__n22012 & ~ys__n28243;
  assign new_n46780_ = ys__n22332 & ys__n28243;
  assign new_n46781_ = ~new_n46779_ & ~new_n46780_;
  assign new_n46782_ = ys__n28243 & ~new_n46781_;
  assign new_n46783_ = ~new_n46778_ & ~new_n46782_;
  assign new_n46784_ = ys__n28243 & ~new_n46783_;
  assign new_n46785_ = ~new_n46774_ & ~new_n46784_;
  assign new_n46786_ = new_n46235_ & ~new_n46785_;
  assign new_n46787_ = ys__n47807 & new_n46239_;
  assign new_n46788_ = ~new_n46786_ & ~new_n46787_;
  assign new_n46789_ = ~new_n46769_ & new_n46788_;
  assign new_n46790_ = ~new_n46768_ & new_n46789_;
  assign new_n46791_ = ~new_n46767_ & new_n46790_;
  assign ys__n32140 = ~new_n46267_ & ~new_n46791_;
  assign new_n46793_ = ~new_n23757_ & ~new_n38915_;
  assign new_n46794_ = ~new_n23921_ & ~new_n46793_;
  assign new_n46795_ = ~new_n46201_ & ~new_n46794_;
  assign new_n46796_ = ys__n27795 & new_n46201_;
  assign new_n46797_ = ~new_n46795_ & ~new_n46796_;
  assign new_n46798_ = new_n46210_ & ~new_n46797_;
  assign new_n46799_ = ys__n19929 & new_n46214_;
  assign new_n46800_ = ys__n47776 & new_n46245_;
  assign new_n46801_ = ys__n20990 & ~ys__n28243;
  assign new_n46802_ = ys__n21310 & ys__n28243;
  assign new_n46803_ = ~new_n46801_ & ~new_n46802_;
  assign new_n46804_ = ys__n28243 & ~new_n46803_;
  assign new_n46805_ = ~ys__n28243 & new_n46804_;
  assign new_n46806_ = ys__n21534 & ~ys__n28243;
  assign new_n46807_ = ys__n21854 & ys__n28243;
  assign new_n46808_ = ~new_n46806_ & ~new_n46807_;
  assign new_n46809_ = ~ys__n28243 & ~new_n46808_;
  assign new_n46810_ = ys__n22014 & ~ys__n28243;
  assign new_n46811_ = ys__n22334 & ys__n28243;
  assign new_n46812_ = ~new_n46810_ & ~new_n46811_;
  assign new_n46813_ = ys__n28243 & ~new_n46812_;
  assign new_n46814_ = ~new_n46809_ & ~new_n46813_;
  assign new_n46815_ = ys__n28243 & ~new_n46814_;
  assign new_n46816_ = ~new_n46805_ & ~new_n46815_;
  assign new_n46817_ = new_n46235_ & ~new_n46816_;
  assign new_n46818_ = ys__n47808 & new_n46239_;
  assign new_n46819_ = ~new_n46817_ & ~new_n46818_;
  assign new_n46820_ = ~new_n46800_ & new_n46819_;
  assign new_n46821_ = ~new_n46799_ & new_n46820_;
  assign new_n46822_ = ~new_n46798_ & new_n46821_;
  assign ys__n32141 = ~new_n46267_ & ~new_n46822_;
  assign new_n46824_ = ~new_n23757_ & ~new_n38923_;
  assign new_n46825_ = ~new_n23936_ & ~new_n46824_;
  assign new_n46826_ = ~new_n46201_ & ~new_n46825_;
  assign new_n46827_ = ys__n27798 & new_n46201_;
  assign new_n46828_ = ~new_n46826_ & ~new_n46827_;
  assign new_n46829_ = new_n46210_ & ~new_n46828_;
  assign new_n46830_ = ys__n19932 & new_n46214_;
  assign new_n46831_ = ys__n47777 & new_n46245_;
  assign new_n46832_ = ys__n20992 & ~ys__n28243;
  assign new_n46833_ = ys__n21312 & ys__n28243;
  assign new_n46834_ = ~new_n46832_ & ~new_n46833_;
  assign new_n46835_ = ys__n28243 & ~new_n46834_;
  assign new_n46836_ = ~ys__n28243 & new_n46835_;
  assign new_n46837_ = ys__n21536 & ~ys__n28243;
  assign new_n46838_ = ys__n21856 & ys__n28243;
  assign new_n46839_ = ~new_n46837_ & ~new_n46838_;
  assign new_n46840_ = ~ys__n28243 & ~new_n46839_;
  assign new_n46841_ = ys__n22016 & ~ys__n28243;
  assign new_n46842_ = ys__n22336 & ys__n28243;
  assign new_n46843_ = ~new_n46841_ & ~new_n46842_;
  assign new_n46844_ = ys__n28243 & ~new_n46843_;
  assign new_n46845_ = ~new_n46840_ & ~new_n46844_;
  assign new_n46846_ = ys__n28243 & ~new_n46845_;
  assign new_n46847_ = ~new_n46836_ & ~new_n46846_;
  assign new_n46848_ = new_n46235_ & ~new_n46847_;
  assign new_n46849_ = ys__n47809 & new_n46239_;
  assign new_n46850_ = ~new_n46848_ & ~new_n46849_;
  assign new_n46851_ = ~new_n46831_ & new_n46850_;
  assign new_n46852_ = ~new_n46830_ & new_n46851_;
  assign new_n46853_ = ~new_n46829_ & new_n46852_;
  assign ys__n32142 = ~new_n46267_ & ~new_n46853_;
  assign new_n46855_ = ~new_n23757_ & ~new_n38931_;
  assign new_n46856_ = ~new_n23951_ & ~new_n46855_;
  assign new_n46857_ = ~new_n46201_ & ~new_n46856_;
  assign new_n46858_ = ys__n27801 & new_n46201_;
  assign new_n46859_ = ~new_n46857_ & ~new_n46858_;
  assign new_n46860_ = new_n46210_ & ~new_n46859_;
  assign new_n46861_ = ys__n19935 & new_n46214_;
  assign new_n46862_ = ys__n47778 & new_n46245_;
  assign new_n46863_ = ys__n20994 & ~ys__n28243;
  assign new_n46864_ = ys__n21314 & ys__n28243;
  assign new_n46865_ = ~new_n46863_ & ~new_n46864_;
  assign new_n46866_ = ys__n28243 & ~new_n46865_;
  assign new_n46867_ = ~ys__n28243 & new_n46866_;
  assign new_n46868_ = ys__n21538 & ~ys__n28243;
  assign new_n46869_ = ys__n21858 & ys__n28243;
  assign new_n46870_ = ~new_n46868_ & ~new_n46869_;
  assign new_n46871_ = ~ys__n28243 & ~new_n46870_;
  assign new_n46872_ = ys__n22018 & ~ys__n28243;
  assign new_n46873_ = ys__n22338 & ys__n28243;
  assign new_n46874_ = ~new_n46872_ & ~new_n46873_;
  assign new_n46875_ = ys__n28243 & ~new_n46874_;
  assign new_n46876_ = ~new_n46871_ & ~new_n46875_;
  assign new_n46877_ = ys__n28243 & ~new_n46876_;
  assign new_n46878_ = ~new_n46867_ & ~new_n46877_;
  assign new_n46879_ = new_n46235_ & ~new_n46878_;
  assign new_n46880_ = ys__n47810 & new_n46239_;
  assign new_n46881_ = ~new_n46879_ & ~new_n46880_;
  assign new_n46882_ = ~new_n46862_ & new_n46881_;
  assign new_n46883_ = ~new_n46861_ & new_n46882_;
  assign new_n46884_ = ~new_n46860_ & new_n46883_;
  assign ys__n32143 = ~new_n46267_ & ~new_n46884_;
  assign new_n46886_ = ~new_n23757_ & ~new_n38939_;
  assign new_n46887_ = ~new_n23966_ & ~new_n46886_;
  assign new_n46888_ = ~new_n46201_ & ~new_n46887_;
  assign new_n46889_ = ys__n27804 & new_n46201_;
  assign new_n46890_ = ~new_n46888_ & ~new_n46889_;
  assign new_n46891_ = new_n46210_ & ~new_n46890_;
  assign new_n46892_ = ys__n19938 & new_n46214_;
  assign new_n46893_ = ys__n47779 & new_n46245_;
  assign new_n46894_ = ys__n20996 & ~ys__n28243;
  assign new_n46895_ = ys__n21316 & ys__n28243;
  assign new_n46896_ = ~new_n46894_ & ~new_n46895_;
  assign new_n46897_ = ys__n28243 & ~new_n46896_;
  assign new_n46898_ = ~ys__n28243 & new_n46897_;
  assign new_n46899_ = ys__n21540 & ~ys__n28243;
  assign new_n46900_ = ys__n21860 & ys__n28243;
  assign new_n46901_ = ~new_n46899_ & ~new_n46900_;
  assign new_n46902_ = ~ys__n28243 & ~new_n46901_;
  assign new_n46903_ = ys__n22020 & ~ys__n28243;
  assign new_n46904_ = ys__n22340 & ys__n28243;
  assign new_n46905_ = ~new_n46903_ & ~new_n46904_;
  assign new_n46906_ = ys__n28243 & ~new_n46905_;
  assign new_n46907_ = ~new_n46902_ & ~new_n46906_;
  assign new_n46908_ = ys__n28243 & ~new_n46907_;
  assign new_n46909_ = ~new_n46898_ & ~new_n46908_;
  assign new_n46910_ = new_n46235_ & ~new_n46909_;
  assign new_n46911_ = ys__n47811 & new_n46239_;
  assign new_n46912_ = ~new_n46910_ & ~new_n46911_;
  assign new_n46913_ = ~new_n46893_ & new_n46912_;
  assign new_n46914_ = ~new_n46892_ & new_n46913_;
  assign new_n46915_ = ~new_n46891_ & new_n46914_;
  assign ys__n32144 = ~new_n46267_ & ~new_n46915_;
  assign new_n46917_ = ~new_n23757_ & ~new_n38947_;
  assign new_n46918_ = ~new_n23981_ & ~new_n46917_;
  assign new_n46919_ = ~new_n46201_ & ~new_n46918_;
  assign new_n46920_ = ys__n27807 & new_n46201_;
  assign new_n46921_ = ~new_n46919_ & ~new_n46920_;
  assign new_n46922_ = new_n46210_ & ~new_n46921_;
  assign new_n46923_ = ys__n19941 & new_n46214_;
  assign new_n46924_ = ys__n47780 & new_n46245_;
  assign new_n46925_ = ys__n20998 & ~ys__n28243;
  assign new_n46926_ = ys__n21318 & ys__n28243;
  assign new_n46927_ = ~new_n46925_ & ~new_n46926_;
  assign new_n46928_ = ys__n28243 & ~new_n46927_;
  assign new_n46929_ = ~ys__n28243 & new_n46928_;
  assign new_n46930_ = ys__n21542 & ~ys__n28243;
  assign new_n46931_ = ys__n21862 & ys__n28243;
  assign new_n46932_ = ~new_n46930_ & ~new_n46931_;
  assign new_n46933_ = ~ys__n28243 & ~new_n46932_;
  assign new_n46934_ = ys__n22022 & ~ys__n28243;
  assign new_n46935_ = ys__n22342 & ys__n28243;
  assign new_n46936_ = ~new_n46934_ & ~new_n46935_;
  assign new_n46937_ = ys__n28243 & ~new_n46936_;
  assign new_n46938_ = ~new_n46933_ & ~new_n46937_;
  assign new_n46939_ = ys__n28243 & ~new_n46938_;
  assign new_n46940_ = ~new_n46929_ & ~new_n46939_;
  assign new_n46941_ = new_n46235_ & ~new_n46940_;
  assign new_n46942_ = ys__n47812 & new_n46239_;
  assign new_n46943_ = ~new_n46941_ & ~new_n46942_;
  assign new_n46944_ = ~new_n46924_ & new_n46943_;
  assign new_n46945_ = ~new_n46923_ & new_n46944_;
  assign new_n46946_ = ~new_n46922_ & new_n46945_;
  assign ys__n32145 = ~new_n46267_ & ~new_n46946_;
  assign new_n46948_ = ~new_n23757_ & ~new_n38955_;
  assign new_n46949_ = ~new_n23996_ & ~new_n46948_;
  assign new_n46950_ = ~new_n46201_ & ~new_n46949_;
  assign new_n46951_ = ys__n27810 & new_n46201_;
  assign new_n46952_ = ~new_n46950_ & ~new_n46951_;
  assign new_n46953_ = new_n46210_ & ~new_n46952_;
  assign new_n46954_ = ys__n19944 & new_n46214_;
  assign new_n46955_ = ys__n47781 & new_n46245_;
  assign new_n46956_ = ys__n21000 & ~ys__n28243;
  assign new_n46957_ = ys__n21320 & ys__n28243;
  assign new_n46958_ = ~new_n46956_ & ~new_n46957_;
  assign new_n46959_ = ys__n28243 & ~new_n46958_;
  assign new_n46960_ = ~ys__n28243 & new_n46959_;
  assign new_n46961_ = ys__n21544 & ~ys__n28243;
  assign new_n46962_ = ys__n21864 & ys__n28243;
  assign new_n46963_ = ~new_n46961_ & ~new_n46962_;
  assign new_n46964_ = ~ys__n28243 & ~new_n46963_;
  assign new_n46965_ = ys__n22024 & ~ys__n28243;
  assign new_n46966_ = ys__n22344 & ys__n28243;
  assign new_n46967_ = ~new_n46965_ & ~new_n46966_;
  assign new_n46968_ = ys__n28243 & ~new_n46967_;
  assign new_n46969_ = ~new_n46964_ & ~new_n46968_;
  assign new_n46970_ = ys__n28243 & ~new_n46969_;
  assign new_n46971_ = ~new_n46960_ & ~new_n46970_;
  assign new_n46972_ = new_n46235_ & ~new_n46971_;
  assign new_n46973_ = ys__n47813 & new_n46239_;
  assign new_n46974_ = ~new_n46972_ & ~new_n46973_;
  assign new_n46975_ = ~new_n46955_ & new_n46974_;
  assign new_n46976_ = ~new_n46954_ & new_n46975_;
  assign new_n46977_ = ~new_n46953_ & new_n46976_;
  assign ys__n32146 = ~new_n46267_ & ~new_n46977_;
  assign new_n46979_ = ys__n19947 & new_n46214_;
  assign new_n46980_ = ~new_n23757_ & ~new_n38963_;
  assign new_n46981_ = ~new_n24011_ & ~new_n46980_;
  assign new_n46982_ = ~new_n46201_ & ~new_n46981_;
  assign new_n46983_ = ys__n27813 & new_n46201_;
  assign new_n46984_ = ~new_n46982_ & ~new_n46983_;
  assign new_n46985_ = new_n46210_ & ~new_n46984_;
  assign new_n46986_ = ys__n47782 & new_n46245_;
  assign new_n46987_ = ys__n21002 & ~ys__n28243;
  assign new_n46988_ = ys__n21322 & ys__n28243;
  assign new_n46989_ = ~new_n46987_ & ~new_n46988_;
  assign new_n46990_ = ys__n28243 & ~new_n46989_;
  assign new_n46991_ = ~ys__n28243 & new_n46990_;
  assign new_n46992_ = ys__n21546 & ~ys__n28243;
  assign new_n46993_ = ys__n21866 & ys__n28243;
  assign new_n46994_ = ~new_n46992_ & ~new_n46993_;
  assign new_n46995_ = ~ys__n28243 & ~new_n46994_;
  assign new_n46996_ = ys__n22026 & ~ys__n28243;
  assign new_n46997_ = ys__n22346 & ys__n28243;
  assign new_n46998_ = ~new_n46996_ & ~new_n46997_;
  assign new_n46999_ = ys__n28243 & ~new_n46998_;
  assign new_n47000_ = ~new_n46995_ & ~new_n46999_;
  assign new_n47001_ = ys__n28243 & ~new_n47000_;
  assign new_n47002_ = ~new_n46991_ & ~new_n47001_;
  assign new_n47003_ = new_n46235_ & ~new_n47002_;
  assign new_n47004_ = ys__n47814 & new_n46239_;
  assign new_n47005_ = ~new_n47003_ & ~new_n47004_;
  assign new_n47006_ = ~new_n46986_ & new_n47005_;
  assign new_n47007_ = ~new_n46985_ & new_n47006_;
  assign new_n47008_ = ~new_n46979_ & new_n47007_;
  assign ys__n32147 = ~new_n46267_ & ~new_n47008_;
  assign new_n47010_ = ~new_n23757_ & ~new_n38971_;
  assign new_n47011_ = ~new_n23758_ & ~new_n47010_;
  assign new_n47012_ = ~new_n46201_ & ~new_n47011_;
  assign new_n47013_ = ys__n27816 & new_n46201_;
  assign new_n47014_ = ~new_n47012_ & ~new_n47013_;
  assign new_n47015_ = new_n46210_ & ~new_n47014_;
  assign new_n47016_ = ys__n19950 & new_n46214_;
  assign new_n47017_ = ys__n47783 & new_n46245_;
  assign new_n47018_ = ys__n21004 & ~ys__n28243;
  assign new_n47019_ = ys__n21324 & ys__n28243;
  assign new_n47020_ = ~new_n47018_ & ~new_n47019_;
  assign new_n47021_ = ys__n28243 & ~new_n47020_;
  assign new_n47022_ = ~ys__n28243 & new_n47021_;
  assign new_n47023_ = ys__n21548 & ~ys__n28243;
  assign new_n47024_ = ys__n21868 & ys__n28243;
  assign new_n47025_ = ~new_n47023_ & ~new_n47024_;
  assign new_n47026_ = ~ys__n28243 & ~new_n47025_;
  assign new_n47027_ = ys__n22028 & ~ys__n28243;
  assign new_n47028_ = ys__n22348 & ys__n28243;
  assign new_n47029_ = ~new_n47027_ & ~new_n47028_;
  assign new_n47030_ = ys__n28243 & ~new_n47029_;
  assign new_n47031_ = ~new_n47026_ & ~new_n47030_;
  assign new_n47032_ = ys__n28243 & ~new_n47031_;
  assign new_n47033_ = ~new_n47022_ & ~new_n47032_;
  assign new_n47034_ = new_n46235_ & ~new_n47033_;
  assign new_n47035_ = ys__n47815 & new_n46239_;
  assign new_n47036_ = ~new_n47034_ & ~new_n47035_;
  assign new_n47037_ = ~new_n47017_ & new_n47036_;
  assign new_n47038_ = ~new_n47016_ & new_n47037_;
  assign new_n47039_ = ~new_n47015_ & new_n47038_;
  assign ys__n32148 = ~new_n46267_ & ~new_n47039_;
  assign new_n47041_ = ~new_n23757_ & ~new_n38979_;
  assign new_n47042_ = ~new_n23773_ & ~new_n47041_;
  assign new_n47043_ = ~new_n46201_ & ~new_n47042_;
  assign new_n47044_ = ys__n27819 & new_n46201_;
  assign new_n47045_ = ~new_n47043_ & ~new_n47044_;
  assign new_n47046_ = new_n46210_ & ~new_n47045_;
  assign new_n47047_ = ys__n19953 & new_n46214_;
  assign new_n47048_ = ys__n47784 & new_n46245_;
  assign new_n47049_ = ys__n21006 & ~ys__n28243;
  assign new_n47050_ = ys__n21326 & ys__n28243;
  assign new_n47051_ = ~new_n47049_ & ~new_n47050_;
  assign new_n47052_ = ys__n28243 & ~new_n47051_;
  assign new_n47053_ = ~ys__n28243 & new_n47052_;
  assign new_n47054_ = ys__n21550 & ~ys__n28243;
  assign new_n47055_ = ys__n21870 & ys__n28243;
  assign new_n47056_ = ~new_n47054_ & ~new_n47055_;
  assign new_n47057_ = ~ys__n28243 & ~new_n47056_;
  assign new_n47058_ = ys__n22030 & ~ys__n28243;
  assign new_n47059_ = ys__n22350 & ys__n28243;
  assign new_n47060_ = ~new_n47058_ & ~new_n47059_;
  assign new_n47061_ = ys__n28243 & ~new_n47060_;
  assign new_n47062_ = ~new_n47057_ & ~new_n47061_;
  assign new_n47063_ = ys__n28243 & ~new_n47062_;
  assign new_n47064_ = ~new_n47053_ & ~new_n47063_;
  assign new_n47065_ = new_n46235_ & ~new_n47064_;
  assign new_n47066_ = ys__n47816 & new_n46239_;
  assign new_n47067_ = ~new_n47065_ & ~new_n47066_;
  assign new_n47068_ = ~new_n47048_ & new_n47067_;
  assign new_n47069_ = ~new_n47047_ & new_n47068_;
  assign new_n47070_ = ~new_n47046_ & new_n47069_;
  assign ys__n32149 = ~new_n46267_ & ~new_n47070_;
  assign new_n47072_ = ~new_n23757_ & ~new_n38987_;
  assign new_n47073_ = ~new_n23788_ & ~new_n47072_;
  assign new_n47074_ = ~new_n46201_ & ~new_n47073_;
  assign new_n47075_ = ys__n27822 & new_n46201_;
  assign new_n47076_ = ~new_n47074_ & ~new_n47075_;
  assign new_n47077_ = new_n46210_ & ~new_n47076_;
  assign new_n47078_ = ys__n19956 & new_n46214_;
  assign new_n47079_ = ys__n47785 & new_n46245_;
  assign new_n47080_ = ys__n21008 & ~ys__n28243;
  assign new_n47081_ = ys__n21328 & ys__n28243;
  assign new_n47082_ = ~new_n47080_ & ~new_n47081_;
  assign new_n47083_ = ys__n28243 & ~new_n47082_;
  assign new_n47084_ = ~ys__n28243 & new_n47083_;
  assign new_n47085_ = ys__n21552 & ~ys__n28243;
  assign new_n47086_ = ys__n21872 & ys__n28243;
  assign new_n47087_ = ~new_n47085_ & ~new_n47086_;
  assign new_n47088_ = ~ys__n28243 & ~new_n47087_;
  assign new_n47089_ = ys__n22032 & ~ys__n28243;
  assign new_n47090_ = ys__n22352 & ys__n28243;
  assign new_n47091_ = ~new_n47089_ & ~new_n47090_;
  assign new_n47092_ = ys__n28243 & ~new_n47091_;
  assign new_n47093_ = ~new_n47088_ & ~new_n47092_;
  assign new_n47094_ = ys__n28243 & ~new_n47093_;
  assign new_n47095_ = ~new_n47084_ & ~new_n47094_;
  assign new_n47096_ = new_n46235_ & ~new_n47095_;
  assign new_n47097_ = ys__n47817 & new_n46239_;
  assign new_n47098_ = ~new_n47096_ & ~new_n47097_;
  assign new_n47099_ = ~new_n47079_ & new_n47098_;
  assign new_n47100_ = ~new_n47078_ & new_n47099_;
  assign new_n47101_ = ~new_n47077_ & new_n47100_;
  assign ys__n32150 = ~new_n46267_ & ~new_n47101_;
  assign new_n47103_ = ys__n19959 & new_n46214_;
  assign new_n47104_ = ~new_n23757_ & ~new_n38995_;
  assign new_n47105_ = ~new_n23803_ & ~new_n47104_;
  assign new_n47106_ = ~new_n46201_ & ~new_n47105_;
  assign new_n47107_ = ys__n27825 & new_n46201_;
  assign new_n47108_ = ~new_n47106_ & ~new_n47107_;
  assign new_n47109_ = new_n46210_ & ~new_n47108_;
  assign new_n47110_ = ys__n47786 & new_n46245_;
  assign new_n47111_ = ys__n21010 & ~ys__n28243;
  assign new_n47112_ = ys__n21330 & ys__n28243;
  assign new_n47113_ = ~new_n47111_ & ~new_n47112_;
  assign new_n47114_ = ys__n28243 & ~new_n47113_;
  assign new_n47115_ = ~ys__n28243 & new_n47114_;
  assign new_n47116_ = ys__n21554 & ~ys__n28243;
  assign new_n47117_ = ys__n21874 & ys__n28243;
  assign new_n47118_ = ~new_n47116_ & ~new_n47117_;
  assign new_n47119_ = ~ys__n28243 & ~new_n47118_;
  assign new_n47120_ = ys__n22034 & ~ys__n28243;
  assign new_n47121_ = ys__n22354 & ys__n28243;
  assign new_n47122_ = ~new_n47120_ & ~new_n47121_;
  assign new_n47123_ = ys__n28243 & ~new_n47122_;
  assign new_n47124_ = ~new_n47119_ & ~new_n47123_;
  assign new_n47125_ = ys__n28243 & ~new_n47124_;
  assign new_n47126_ = ~new_n47115_ & ~new_n47125_;
  assign new_n47127_ = new_n46235_ & ~new_n47126_;
  assign new_n47128_ = ys__n47818 & new_n46239_;
  assign new_n47129_ = ~new_n47127_ & ~new_n47128_;
  assign new_n47130_ = ~new_n47110_ & new_n47129_;
  assign new_n47131_ = ~new_n47109_ & new_n47130_;
  assign new_n47132_ = ~new_n47103_ & new_n47131_;
  assign ys__n32151 = ~new_n46267_ & ~new_n47132_;
  assign new_n47134_ = ~new_n23757_ & ~new_n39003_;
  assign new_n47135_ = ~new_n23818_ & ~new_n47134_;
  assign new_n47136_ = ~new_n46201_ & ~new_n47135_;
  assign new_n47137_ = ys__n27828 & new_n46201_;
  assign new_n47138_ = ~new_n47136_ & ~new_n47137_;
  assign new_n47139_ = new_n46210_ & ~new_n47138_;
  assign new_n47140_ = ys__n19962 & new_n46214_;
  assign new_n47141_ = ys__n47787 & new_n46245_;
  assign new_n47142_ = ys__n21012 & ~ys__n28243;
  assign new_n47143_ = ys__n21332 & ys__n28243;
  assign new_n47144_ = ~new_n47142_ & ~new_n47143_;
  assign new_n47145_ = ys__n28243 & ~new_n47144_;
  assign new_n47146_ = ~ys__n28243 & new_n47145_;
  assign new_n47147_ = ys__n21556 & ~ys__n28243;
  assign new_n47148_ = ys__n21876 & ys__n28243;
  assign new_n47149_ = ~new_n47147_ & ~new_n47148_;
  assign new_n47150_ = ~ys__n28243 & ~new_n47149_;
  assign new_n47151_ = ys__n22036 & ~ys__n28243;
  assign new_n47152_ = ys__n22356 & ys__n28243;
  assign new_n47153_ = ~new_n47151_ & ~new_n47152_;
  assign new_n47154_ = ys__n28243 & ~new_n47153_;
  assign new_n47155_ = ~new_n47150_ & ~new_n47154_;
  assign new_n47156_ = ys__n28243 & ~new_n47155_;
  assign new_n47157_ = ~new_n47146_ & ~new_n47156_;
  assign new_n47158_ = new_n46235_ & ~new_n47157_;
  assign new_n47159_ = ys__n47819 & new_n46239_;
  assign new_n47160_ = ~new_n47158_ & ~new_n47159_;
  assign new_n47161_ = ~new_n47141_ & new_n47160_;
  assign new_n47162_ = ~new_n47140_ & new_n47161_;
  assign new_n47163_ = ~new_n47139_ & new_n47162_;
  assign ys__n32152 = ~new_n46267_ & ~new_n47163_;
  assign new_n47165_ = ys__n19965 & new_n46214_;
  assign new_n47166_ = ~new_n23757_ & ~new_n39011_;
  assign new_n47167_ = ~new_n23833_ & ~new_n47166_;
  assign new_n47168_ = ~new_n46201_ & ~new_n47167_;
  assign new_n47169_ = ys__n27831 & new_n46201_;
  assign new_n47170_ = ~new_n47168_ & ~new_n47169_;
  assign new_n47171_ = new_n46210_ & ~new_n47170_;
  assign new_n47172_ = ys__n47788 & new_n46245_;
  assign new_n47173_ = ys__n21014 & ~ys__n28243;
  assign new_n47174_ = ys__n21334 & ys__n28243;
  assign new_n47175_ = ~new_n47173_ & ~new_n47174_;
  assign new_n47176_ = ys__n28243 & ~new_n47175_;
  assign new_n47177_ = ~ys__n28243 & new_n47176_;
  assign new_n47178_ = ys__n21558 & ~ys__n28243;
  assign new_n47179_ = ys__n21878 & ys__n28243;
  assign new_n47180_ = ~new_n47178_ & ~new_n47179_;
  assign new_n47181_ = ~ys__n28243 & ~new_n47180_;
  assign new_n47182_ = ys__n22038 & ~ys__n28243;
  assign new_n47183_ = ys__n22358 & ys__n28243;
  assign new_n47184_ = ~new_n47182_ & ~new_n47183_;
  assign new_n47185_ = ys__n28243 & ~new_n47184_;
  assign new_n47186_ = ~new_n47181_ & ~new_n47185_;
  assign new_n47187_ = ys__n28243 & ~new_n47186_;
  assign new_n47188_ = ~new_n47177_ & ~new_n47187_;
  assign new_n47189_ = new_n46235_ & ~new_n47188_;
  assign new_n47190_ = ys__n47820 & new_n46239_;
  assign new_n47191_ = ~new_n47189_ & ~new_n47190_;
  assign new_n47192_ = ~new_n47172_ & new_n47191_;
  assign new_n47193_ = ~new_n47171_ & new_n47192_;
  assign new_n47194_ = ~new_n47165_ & new_n47193_;
  assign ys__n32153 = ~new_n46267_ & ~new_n47194_;
  assign new_n47196_ = ys__n19968 & new_n46214_;
  assign new_n47197_ = ~new_n23757_ & ~new_n39019_;
  assign new_n47198_ = ~new_n23848_ & ~new_n47197_;
  assign new_n47199_ = ~new_n46201_ & ~new_n47198_;
  assign new_n47200_ = ys__n27834 & new_n46201_;
  assign new_n47201_ = ~new_n47199_ & ~new_n47200_;
  assign new_n47202_ = new_n46210_ & ~new_n47201_;
  assign new_n47203_ = ys__n47789 & new_n46245_;
  assign new_n47204_ = ys__n21016 & ~ys__n28243;
  assign new_n47205_ = ys__n21336 & ys__n28243;
  assign new_n47206_ = ~new_n47204_ & ~new_n47205_;
  assign new_n47207_ = ys__n28243 & ~new_n47206_;
  assign new_n47208_ = ~ys__n28243 & new_n47207_;
  assign new_n47209_ = ys__n21560 & ~ys__n28243;
  assign new_n47210_ = ys__n21880 & ys__n28243;
  assign new_n47211_ = ~new_n47209_ & ~new_n47210_;
  assign new_n47212_ = ~ys__n28243 & ~new_n47211_;
  assign new_n47213_ = ys__n22040 & ~ys__n28243;
  assign new_n47214_ = ys__n22360 & ys__n28243;
  assign new_n47215_ = ~new_n47213_ & ~new_n47214_;
  assign new_n47216_ = ys__n28243 & ~new_n47215_;
  assign new_n47217_ = ~new_n47212_ & ~new_n47216_;
  assign new_n47218_ = ys__n28243 & ~new_n47217_;
  assign new_n47219_ = ~new_n47208_ & ~new_n47218_;
  assign new_n47220_ = new_n46235_ & ~new_n47219_;
  assign new_n47221_ = ys__n47821 & new_n46239_;
  assign new_n47222_ = ~new_n47220_ & ~new_n47221_;
  assign new_n47223_ = ~new_n47203_ & new_n47222_;
  assign new_n47224_ = ~new_n47202_ & new_n47223_;
  assign new_n47225_ = ~new_n47196_ & new_n47224_;
  assign ys__n32154 = ~new_n46267_ & ~new_n47225_;
  assign new_n47227_ = ys__n19971 & new_n46214_;
  assign new_n47228_ = ~new_n23757_ & ~new_n39027_;
  assign new_n47229_ = ~new_n23863_ & ~new_n47228_;
  assign new_n47230_ = ~new_n46201_ & ~new_n47229_;
  assign new_n47231_ = ys__n27837 & new_n46201_;
  assign new_n47232_ = ~new_n47230_ & ~new_n47231_;
  assign new_n47233_ = new_n46210_ & ~new_n47232_;
  assign new_n47234_ = ys__n47790 & new_n46245_;
  assign new_n47235_ = ys__n21018 & ~ys__n28243;
  assign new_n47236_ = ys__n21338 & ys__n28243;
  assign new_n47237_ = ~new_n47235_ & ~new_n47236_;
  assign new_n47238_ = ys__n28243 & ~new_n47237_;
  assign new_n47239_ = ~ys__n28243 & new_n47238_;
  assign new_n47240_ = ys__n21562 & ~ys__n28243;
  assign new_n47241_ = ys__n21882 & ys__n28243;
  assign new_n47242_ = ~new_n47240_ & ~new_n47241_;
  assign new_n47243_ = ~ys__n28243 & ~new_n47242_;
  assign new_n47244_ = ys__n22042 & ~ys__n28243;
  assign new_n47245_ = ys__n22362 & ys__n28243;
  assign new_n47246_ = ~new_n47244_ & ~new_n47245_;
  assign new_n47247_ = ys__n28243 & ~new_n47246_;
  assign new_n47248_ = ~new_n47243_ & ~new_n47247_;
  assign new_n47249_ = ys__n28243 & ~new_n47248_;
  assign new_n47250_ = ~new_n47239_ & ~new_n47249_;
  assign new_n47251_ = new_n46235_ & ~new_n47250_;
  assign new_n47252_ = ys__n47822 & new_n46239_;
  assign new_n47253_ = ~new_n47251_ & ~new_n47252_;
  assign new_n47254_ = ~new_n47234_ & new_n47253_;
  assign new_n47255_ = ~new_n47233_ & new_n47254_;
  assign new_n47256_ = ~new_n47227_ & new_n47255_;
  assign ys__n32155 = ~new_n46267_ & ~new_n47256_;
  assign new_n47258_ = ~ys__n310 & new_n12842_;
  assign new_n47259_ = new_n12212_ & new_n47258_;
  assign ys__n32158 = ~new_n15100_ & new_n47259_;
  assign new_n47261_ = ys__n308 & ys__n310;
  assign new_n47262_ = ~new_n12908_ & ~new_n47261_;
  assign new_n47263_ = new_n12212_ & new_n12842_;
  assign new_n47264_ = ~new_n47262_ & new_n47263_;
  assign new_n47265_ = ~new_n12205_ & ~new_n47264_;
  assign ys__n32159 = ~new_n15100_ & ~new_n47265_;
  assign new_n47267_ = ys__n1301 & ~new_n12860_;
  assign new_n47268_ = ys__n47823 & new_n47267_;
  assign new_n47269_ = ~ys__n816 & new_n12860_;
  assign new_n47270_ = ~ys__n1301 & ~new_n12860_;
  assign new_n47271_ = ~new_n47269_ & ~new_n47270_;
  assign new_n47272_ = ys__n47857 & ~new_n47271_;
  assign new_n47273_ = ~new_n47268_ & ~new_n47272_;
  assign new_n47274_ = ~new_n47267_ & new_n47271_;
  assign ys__n32160 = ~new_n47273_ & ~new_n47274_;
  assign new_n47276_ = ys__n47824 & new_n47267_;
  assign new_n47277_ = ys__n47858 & ~new_n47271_;
  assign new_n47278_ = ~new_n47276_ & ~new_n47277_;
  assign ys__n32161 = ~new_n47274_ & ~new_n47278_;
  assign new_n47280_ = ys__n47825 & new_n47267_;
  assign new_n47281_ = ys__n47859 & ~new_n47271_;
  assign new_n47282_ = ~new_n47280_ & ~new_n47281_;
  assign ys__n32162 = ~new_n47274_ & ~new_n47282_;
  assign new_n47284_ = ys__n47826 & new_n47267_;
  assign new_n47285_ = ys__n47860 & ~new_n47271_;
  assign new_n47286_ = ~new_n47284_ & ~new_n47285_;
  assign ys__n32163 = ~new_n47274_ & ~new_n47286_;
  assign new_n47288_ = ys__n47827 & new_n47267_;
  assign new_n47289_ = ys__n47861 & ~new_n47271_;
  assign new_n47290_ = ~new_n47288_ & ~new_n47289_;
  assign ys__n32164 = ~new_n47274_ & ~new_n47290_;
  assign new_n47292_ = ys__n47828 & new_n47267_;
  assign new_n47293_ = ys__n47862 & ~new_n47271_;
  assign new_n47294_ = ~new_n47292_ & ~new_n47293_;
  assign ys__n32165 = ~new_n47274_ & ~new_n47294_;
  assign new_n47296_ = ys__n47829 & new_n47267_;
  assign new_n47297_ = ys__n47863 & ~new_n47271_;
  assign new_n47298_ = ~new_n47296_ & ~new_n47297_;
  assign ys__n32166 = ~new_n47274_ & ~new_n47298_;
  assign new_n47300_ = ys__n47830 & new_n47267_;
  assign new_n47301_ = ys__n47864 & ~new_n47271_;
  assign new_n47302_ = ~new_n47300_ & ~new_n47301_;
  assign ys__n32167 = ~new_n47274_ & ~new_n47302_;
  assign new_n47304_ = ys__n47831 & new_n47267_;
  assign new_n47305_ = ys__n47865 & ~new_n47271_;
  assign new_n47306_ = ~new_n47304_ & ~new_n47305_;
  assign ys__n32168 = ~new_n47274_ & ~new_n47306_;
  assign new_n47308_ = ys__n47832 & new_n47267_;
  assign new_n47309_ = ys__n47866 & ~new_n47271_;
  assign new_n47310_ = ~new_n47308_ & ~new_n47309_;
  assign ys__n32169 = ~new_n47274_ & ~new_n47310_;
  assign new_n47312_ = ys__n47833 & new_n47267_;
  assign new_n47313_ = ys__n47867 & ~new_n47271_;
  assign new_n47314_ = ~new_n47312_ & ~new_n47313_;
  assign ys__n32170 = ~new_n47274_ & ~new_n47314_;
  assign new_n47316_ = ys__n47834 & new_n47267_;
  assign new_n47317_ = ys__n47868 & ~new_n47271_;
  assign new_n47318_ = ~new_n47316_ & ~new_n47317_;
  assign ys__n32171 = ~new_n47274_ & ~new_n47318_;
  assign new_n47320_ = ys__n47835 & new_n47267_;
  assign new_n47321_ = ys__n47869 & ~new_n47271_;
  assign new_n47322_ = ~new_n47320_ & ~new_n47321_;
  assign ys__n32172 = ~new_n47274_ & ~new_n47322_;
  assign new_n47324_ = ys__n47836 & new_n47267_;
  assign new_n47325_ = ys__n47870 & ~new_n47271_;
  assign new_n47326_ = ~new_n47324_ & ~new_n47325_;
  assign ys__n32173 = ~new_n47274_ & ~new_n47326_;
  assign new_n47328_ = ys__n47837 & new_n47267_;
  assign new_n47329_ = ys__n47871 & ~new_n47271_;
  assign new_n47330_ = ~new_n47328_ & ~new_n47329_;
  assign ys__n32174 = ~new_n47274_ & ~new_n47330_;
  assign new_n47332_ = ys__n47838 & new_n47267_;
  assign new_n47333_ = ys__n47872 & ~new_n47271_;
  assign new_n47334_ = ~new_n47332_ & ~new_n47333_;
  assign ys__n32175 = ~new_n47274_ & ~new_n47334_;
  assign new_n47336_ = ys__n47839 & new_n47267_;
  assign new_n47337_ = ys__n47873 & ~new_n47271_;
  assign new_n47338_ = ~new_n47336_ & ~new_n47337_;
  assign ys__n32176 = ~new_n47274_ & ~new_n47338_;
  assign new_n47340_ = ys__n47840 & new_n47267_;
  assign new_n47341_ = ys__n47874 & ~new_n47271_;
  assign new_n47342_ = ~new_n47340_ & ~new_n47341_;
  assign ys__n32177 = ~new_n47274_ & ~new_n47342_;
  assign new_n47344_ = ys__n47841 & new_n47267_;
  assign new_n47345_ = ys__n47875 & ~new_n47271_;
  assign new_n47346_ = ~new_n47344_ & ~new_n47345_;
  assign ys__n32178 = ~new_n47274_ & ~new_n47346_;
  assign new_n47348_ = ys__n47842 & new_n47267_;
  assign new_n47349_ = ys__n47876 & ~new_n47271_;
  assign new_n47350_ = ~new_n47348_ & ~new_n47349_;
  assign ys__n32179 = ~new_n47274_ & ~new_n47350_;
  assign new_n47352_ = ys__n47843 & new_n47267_;
  assign new_n47353_ = ys__n47877 & ~new_n47271_;
  assign new_n47354_ = ~new_n47352_ & ~new_n47353_;
  assign ys__n32180 = ~new_n47274_ & ~new_n47354_;
  assign new_n47356_ = ys__n47844 & new_n47267_;
  assign new_n47357_ = ys__n47878 & ~new_n47271_;
  assign new_n47358_ = ~new_n47356_ & ~new_n47357_;
  assign ys__n32181 = ~new_n47274_ & ~new_n47358_;
  assign new_n47360_ = ys__n47845 & new_n47267_;
  assign new_n47361_ = ys__n47879 & ~new_n47271_;
  assign new_n47362_ = ~new_n47360_ & ~new_n47361_;
  assign ys__n32182 = ~new_n47274_ & ~new_n47362_;
  assign new_n47364_ = ys__n47846 & new_n47267_;
  assign new_n47365_ = ys__n47880 & ~new_n47271_;
  assign new_n47366_ = ~new_n47364_ & ~new_n47365_;
  assign ys__n32183 = ~new_n47274_ & ~new_n47366_;
  assign new_n47368_ = ys__n47847 & new_n47267_;
  assign new_n47369_ = ys__n47881 & ~new_n47271_;
  assign new_n47370_ = ~new_n47368_ & ~new_n47369_;
  assign ys__n32184 = ~new_n47274_ & ~new_n47370_;
  assign new_n47372_ = ys__n47848 & new_n47267_;
  assign new_n47373_ = ys__n47882 & ~new_n47271_;
  assign new_n47374_ = ~new_n47372_ & ~new_n47373_;
  assign ys__n32185 = ~new_n47274_ & ~new_n47374_;
  assign new_n47376_ = ys__n47849 & new_n47267_;
  assign new_n47377_ = ys__n47883 & ~new_n47271_;
  assign new_n47378_ = ~new_n47376_ & ~new_n47377_;
  assign ys__n32186 = ~new_n47274_ & ~new_n47378_;
  assign new_n47380_ = ys__n47850 & new_n47267_;
  assign new_n47381_ = ys__n47884 & ~new_n47271_;
  assign new_n47382_ = ~new_n47380_ & ~new_n47381_;
  assign ys__n32187 = ~new_n47274_ & ~new_n47382_;
  assign new_n47384_ = ys__n47851 & new_n47267_;
  assign new_n47385_ = ys__n47885 & ~new_n47271_;
  assign new_n47386_ = ~new_n47384_ & ~new_n47385_;
  assign ys__n32188 = ~new_n47274_ & ~new_n47386_;
  assign new_n47388_ = ys__n47852 & new_n47267_;
  assign new_n47389_ = ys__n47886 & ~new_n47271_;
  assign new_n47390_ = ~new_n47388_ & ~new_n47389_;
  assign ys__n32189 = ~new_n47274_ & ~new_n47390_;
  assign new_n47392_ = ys__n47853 & new_n47267_;
  assign new_n47393_ = ys__n47887 & ~new_n47271_;
  assign new_n47394_ = ~new_n47392_ & ~new_n47393_;
  assign ys__n32190 = ~new_n47274_ & ~new_n47394_;
  assign new_n47396_ = ys__n47854 & new_n47267_;
  assign new_n47397_ = ys__n47888 & ~new_n47271_;
  assign new_n47398_ = ~new_n47396_ & ~new_n47397_;
  assign ys__n32191 = ~new_n47274_ & ~new_n47398_;
  assign new_n47400_ = ys__n47855 & new_n47267_;
  assign new_n47401_ = ys__n19215 & ~new_n47271_;
  assign new_n47402_ = ~new_n47400_ & ~new_n47401_;
  assign ys__n32192 = ~new_n47274_ & ~new_n47402_;
  assign new_n47404_ = ys__n47856 & new_n47267_;
  assign new_n47405_ = ys__n47889 & ~new_n47271_;
  assign new_n47406_ = ~new_n47404_ & ~new_n47405_;
  assign ys__n32193 = ~new_n47274_ & ~new_n47406_;
  assign new_n47408_ = ys__n816 & ~new_n12860_;
  assign new_n47409_ = ys__n47890 & new_n47408_;
  assign new_n47410_ = ~ys__n818 & new_n12860_;
  assign new_n47411_ = ~ys__n816 & ~new_n12860_;
  assign new_n47412_ = ~new_n47410_ & ~new_n47411_;
  assign new_n47413_ = ys__n47857 & ~new_n47412_;
  assign new_n47414_ = ~new_n47409_ & ~new_n47413_;
  assign new_n47415_ = ~new_n47408_ & new_n47412_;
  assign ys__n32194 = ~new_n47414_ & ~new_n47415_;
  assign new_n47417_ = ys__n47891 & new_n47408_;
  assign new_n47418_ = ys__n47858 & ~new_n47412_;
  assign new_n47419_ = ~new_n47417_ & ~new_n47418_;
  assign ys__n32195 = ~new_n47415_ & ~new_n47419_;
  assign new_n47421_ = ys__n47892 & new_n47408_;
  assign new_n47422_ = ys__n47859 & ~new_n47412_;
  assign new_n47423_ = ~new_n47421_ & ~new_n47422_;
  assign ys__n32196 = ~new_n47415_ & ~new_n47423_;
  assign new_n47425_ = ys__n47893 & new_n47408_;
  assign new_n47426_ = ys__n47860 & ~new_n47412_;
  assign new_n47427_ = ~new_n47425_ & ~new_n47426_;
  assign ys__n32197 = ~new_n47415_ & ~new_n47427_;
  assign new_n47429_ = ys__n47894 & new_n47408_;
  assign new_n47430_ = ys__n47861 & ~new_n47412_;
  assign new_n47431_ = ~new_n47429_ & ~new_n47430_;
  assign ys__n32198 = ~new_n47415_ & ~new_n47431_;
  assign new_n47433_ = ys__n47895 & new_n47408_;
  assign new_n47434_ = ys__n47862 & ~new_n47412_;
  assign new_n47435_ = ~new_n47433_ & ~new_n47434_;
  assign ys__n32199 = ~new_n47415_ & ~new_n47435_;
  assign new_n47437_ = ys__n47896 & new_n47408_;
  assign new_n47438_ = ys__n47863 & ~new_n47412_;
  assign new_n47439_ = ~new_n47437_ & ~new_n47438_;
  assign ys__n32200 = ~new_n47415_ & ~new_n47439_;
  assign new_n47441_ = ys__n47897 & new_n47408_;
  assign new_n47442_ = ys__n47864 & ~new_n47412_;
  assign new_n47443_ = ~new_n47441_ & ~new_n47442_;
  assign ys__n32201 = ~new_n47415_ & ~new_n47443_;
  assign new_n47445_ = ys__n47898 & new_n47408_;
  assign new_n47446_ = ys__n47865 & ~new_n47412_;
  assign new_n47447_ = ~new_n47445_ & ~new_n47446_;
  assign ys__n32202 = ~new_n47415_ & ~new_n47447_;
  assign new_n47449_ = ys__n47899 & new_n47408_;
  assign new_n47450_ = ys__n47866 & ~new_n47412_;
  assign new_n47451_ = ~new_n47449_ & ~new_n47450_;
  assign ys__n32203 = ~new_n47415_ & ~new_n47451_;
  assign new_n47453_ = ys__n47900 & new_n47408_;
  assign new_n47454_ = ys__n47867 & ~new_n47412_;
  assign new_n47455_ = ~new_n47453_ & ~new_n47454_;
  assign ys__n32204 = ~new_n47415_ & ~new_n47455_;
  assign new_n47457_ = ys__n47901 & new_n47408_;
  assign new_n47458_ = ys__n47868 & ~new_n47412_;
  assign new_n47459_ = ~new_n47457_ & ~new_n47458_;
  assign ys__n32205 = ~new_n47415_ & ~new_n47459_;
  assign new_n47461_ = ys__n47902 & new_n47408_;
  assign new_n47462_ = ys__n47869 & ~new_n47412_;
  assign new_n47463_ = ~new_n47461_ & ~new_n47462_;
  assign ys__n32206 = ~new_n47415_ & ~new_n47463_;
  assign new_n47465_ = ys__n47903 & new_n47408_;
  assign new_n47466_ = ys__n47870 & ~new_n47412_;
  assign new_n47467_ = ~new_n47465_ & ~new_n47466_;
  assign ys__n32207 = ~new_n47415_ & ~new_n47467_;
  assign new_n47469_ = ys__n47904 & new_n47408_;
  assign new_n47470_ = ys__n47871 & ~new_n47412_;
  assign new_n47471_ = ~new_n47469_ & ~new_n47470_;
  assign ys__n32208 = ~new_n47415_ & ~new_n47471_;
  assign new_n47473_ = ys__n47905 & new_n47408_;
  assign new_n47474_ = ys__n47872 & ~new_n47412_;
  assign new_n47475_ = ~new_n47473_ & ~new_n47474_;
  assign ys__n32209 = ~new_n47415_ & ~new_n47475_;
  assign new_n47477_ = ys__n47906 & new_n47408_;
  assign new_n47478_ = ys__n47873 & ~new_n47412_;
  assign new_n47479_ = ~new_n47477_ & ~new_n47478_;
  assign ys__n32210 = ~new_n47415_ & ~new_n47479_;
  assign new_n47481_ = ys__n47907 & new_n47408_;
  assign new_n47482_ = ys__n47874 & ~new_n47412_;
  assign new_n47483_ = ~new_n47481_ & ~new_n47482_;
  assign ys__n32211 = ~new_n47415_ & ~new_n47483_;
  assign new_n47485_ = ys__n47908 & new_n47408_;
  assign new_n47486_ = ys__n47875 & ~new_n47412_;
  assign new_n47487_ = ~new_n47485_ & ~new_n47486_;
  assign ys__n32212 = ~new_n47415_ & ~new_n47487_;
  assign new_n47489_ = ys__n47909 & new_n47408_;
  assign new_n47490_ = ys__n47876 & ~new_n47412_;
  assign new_n47491_ = ~new_n47489_ & ~new_n47490_;
  assign ys__n32213 = ~new_n47415_ & ~new_n47491_;
  assign new_n47493_ = ys__n47910 & new_n47408_;
  assign new_n47494_ = ys__n47877 & ~new_n47412_;
  assign new_n47495_ = ~new_n47493_ & ~new_n47494_;
  assign ys__n32214 = ~new_n47415_ & ~new_n47495_;
  assign new_n47497_ = ys__n47911 & new_n47408_;
  assign new_n47498_ = ys__n47878 & ~new_n47412_;
  assign new_n47499_ = ~new_n47497_ & ~new_n47498_;
  assign ys__n32215 = ~new_n47415_ & ~new_n47499_;
  assign new_n47501_ = ys__n47912 & new_n47408_;
  assign new_n47502_ = ys__n47879 & ~new_n47412_;
  assign new_n47503_ = ~new_n47501_ & ~new_n47502_;
  assign ys__n32216 = ~new_n47415_ & ~new_n47503_;
  assign new_n47505_ = ys__n47913 & new_n47408_;
  assign new_n47506_ = ys__n47880 & ~new_n47412_;
  assign new_n47507_ = ~new_n47505_ & ~new_n47506_;
  assign ys__n32217 = ~new_n47415_ & ~new_n47507_;
  assign new_n47509_ = ys__n47914 & new_n47408_;
  assign new_n47510_ = ys__n47881 & ~new_n47412_;
  assign new_n47511_ = ~new_n47509_ & ~new_n47510_;
  assign ys__n32218 = ~new_n47415_ & ~new_n47511_;
  assign new_n47513_ = ys__n47915 & new_n47408_;
  assign new_n47514_ = ys__n47882 & ~new_n47412_;
  assign new_n47515_ = ~new_n47513_ & ~new_n47514_;
  assign ys__n32219 = ~new_n47415_ & ~new_n47515_;
  assign new_n47517_ = ys__n47916 & new_n47408_;
  assign new_n47518_ = ys__n47883 & ~new_n47412_;
  assign new_n47519_ = ~new_n47517_ & ~new_n47518_;
  assign ys__n32220 = ~new_n47415_ & ~new_n47519_;
  assign new_n47521_ = ys__n47917 & new_n47408_;
  assign new_n47522_ = ys__n47884 & ~new_n47412_;
  assign new_n47523_ = ~new_n47521_ & ~new_n47522_;
  assign ys__n32221 = ~new_n47415_ & ~new_n47523_;
  assign new_n47525_ = ys__n47918 & new_n47408_;
  assign new_n47526_ = ys__n47885 & ~new_n47412_;
  assign new_n47527_ = ~new_n47525_ & ~new_n47526_;
  assign ys__n32222 = ~new_n47415_ & ~new_n47527_;
  assign new_n47529_ = ys__n47919 & new_n47408_;
  assign new_n47530_ = ys__n47886 & ~new_n47412_;
  assign new_n47531_ = ~new_n47529_ & ~new_n47530_;
  assign ys__n32223 = ~new_n47415_ & ~new_n47531_;
  assign new_n47533_ = ys__n47920 & new_n47408_;
  assign new_n47534_ = ys__n47887 & ~new_n47412_;
  assign new_n47535_ = ~new_n47533_ & ~new_n47534_;
  assign ys__n32224 = ~new_n47415_ & ~new_n47535_;
  assign new_n47537_ = ys__n47921 & new_n47408_;
  assign new_n47538_ = ys__n47888 & ~new_n47412_;
  assign new_n47539_ = ~new_n47537_ & ~new_n47538_;
  assign ys__n32225 = ~new_n47415_ & ~new_n47539_;
  assign new_n47541_ = ys__n47922 & new_n47408_;
  assign new_n47542_ = ys__n19215 & ~new_n47412_;
  assign new_n47543_ = ~new_n47541_ & ~new_n47542_;
  assign ys__n32226 = ~new_n47415_ & ~new_n47543_;
  assign new_n47545_ = ys__n47923 & new_n47408_;
  assign new_n47546_ = ys__n47889 & ~new_n47412_;
  assign new_n47547_ = ~new_n47545_ & ~new_n47546_;
  assign ys__n32227 = ~new_n47415_ & ~new_n47547_;
  assign new_n47549_ = ys__n818 & ~new_n12860_;
  assign new_n47550_ = ys__n47924 & new_n47549_;
  assign new_n47551_ = ~ys__n820 & new_n12860_;
  assign new_n47552_ = ~ys__n818 & ~new_n12860_;
  assign new_n47553_ = ~new_n47551_ & ~new_n47552_;
  assign new_n47554_ = ys__n47857 & ~new_n47553_;
  assign new_n47555_ = ~new_n47550_ & ~new_n47554_;
  assign new_n47556_ = ~new_n47549_ & new_n47553_;
  assign ys__n32228 = ~new_n47555_ & ~new_n47556_;
  assign new_n47558_ = ys__n47925 & new_n47549_;
  assign new_n47559_ = ys__n47858 & ~new_n47553_;
  assign new_n47560_ = ~new_n47558_ & ~new_n47559_;
  assign ys__n32229 = ~new_n47556_ & ~new_n47560_;
  assign new_n47562_ = ys__n47926 & new_n47549_;
  assign new_n47563_ = ys__n47859 & ~new_n47553_;
  assign new_n47564_ = ~new_n47562_ & ~new_n47563_;
  assign ys__n32230 = ~new_n47556_ & ~new_n47564_;
  assign new_n47566_ = ys__n47927 & new_n47549_;
  assign new_n47567_ = ys__n47860 & ~new_n47553_;
  assign new_n47568_ = ~new_n47566_ & ~new_n47567_;
  assign ys__n32231 = ~new_n47556_ & ~new_n47568_;
  assign new_n47570_ = ys__n47928 & new_n47549_;
  assign new_n47571_ = ys__n47861 & ~new_n47553_;
  assign new_n47572_ = ~new_n47570_ & ~new_n47571_;
  assign ys__n32232 = ~new_n47556_ & ~new_n47572_;
  assign new_n47574_ = ys__n47929 & new_n47549_;
  assign new_n47575_ = ys__n47862 & ~new_n47553_;
  assign new_n47576_ = ~new_n47574_ & ~new_n47575_;
  assign ys__n32233 = ~new_n47556_ & ~new_n47576_;
  assign new_n47578_ = ys__n47930 & new_n47549_;
  assign new_n47579_ = ys__n47863 & ~new_n47553_;
  assign new_n47580_ = ~new_n47578_ & ~new_n47579_;
  assign ys__n32234 = ~new_n47556_ & ~new_n47580_;
  assign new_n47582_ = ys__n47931 & new_n47549_;
  assign new_n47583_ = ys__n47864 & ~new_n47553_;
  assign new_n47584_ = ~new_n47582_ & ~new_n47583_;
  assign ys__n32235 = ~new_n47556_ & ~new_n47584_;
  assign new_n47586_ = ys__n47932 & new_n47549_;
  assign new_n47587_ = ys__n47865 & ~new_n47553_;
  assign new_n47588_ = ~new_n47586_ & ~new_n47587_;
  assign ys__n32236 = ~new_n47556_ & ~new_n47588_;
  assign new_n47590_ = ys__n47933 & new_n47549_;
  assign new_n47591_ = ys__n47866 & ~new_n47553_;
  assign new_n47592_ = ~new_n47590_ & ~new_n47591_;
  assign ys__n32237 = ~new_n47556_ & ~new_n47592_;
  assign new_n47594_ = ys__n47934 & new_n47549_;
  assign new_n47595_ = ys__n47867 & ~new_n47553_;
  assign new_n47596_ = ~new_n47594_ & ~new_n47595_;
  assign ys__n32238 = ~new_n47556_ & ~new_n47596_;
  assign new_n47598_ = ys__n47935 & new_n47549_;
  assign new_n47599_ = ys__n47868 & ~new_n47553_;
  assign new_n47600_ = ~new_n47598_ & ~new_n47599_;
  assign ys__n32239 = ~new_n47556_ & ~new_n47600_;
  assign new_n47602_ = ys__n47936 & new_n47549_;
  assign new_n47603_ = ys__n47869 & ~new_n47553_;
  assign new_n47604_ = ~new_n47602_ & ~new_n47603_;
  assign ys__n32240 = ~new_n47556_ & ~new_n47604_;
  assign new_n47606_ = ys__n47937 & new_n47549_;
  assign new_n47607_ = ys__n47870 & ~new_n47553_;
  assign new_n47608_ = ~new_n47606_ & ~new_n47607_;
  assign ys__n32241 = ~new_n47556_ & ~new_n47608_;
  assign new_n47610_ = ys__n47938 & new_n47549_;
  assign new_n47611_ = ys__n47871 & ~new_n47553_;
  assign new_n47612_ = ~new_n47610_ & ~new_n47611_;
  assign ys__n32242 = ~new_n47556_ & ~new_n47612_;
  assign new_n47614_ = ys__n47939 & new_n47549_;
  assign new_n47615_ = ys__n47872 & ~new_n47553_;
  assign new_n47616_ = ~new_n47614_ & ~new_n47615_;
  assign ys__n32243 = ~new_n47556_ & ~new_n47616_;
  assign new_n47618_ = ys__n47940 & new_n47549_;
  assign new_n47619_ = ys__n47873 & ~new_n47553_;
  assign new_n47620_ = ~new_n47618_ & ~new_n47619_;
  assign ys__n32244 = ~new_n47556_ & ~new_n47620_;
  assign new_n47622_ = ys__n47941 & new_n47549_;
  assign new_n47623_ = ys__n47874 & ~new_n47553_;
  assign new_n47624_ = ~new_n47622_ & ~new_n47623_;
  assign ys__n32245 = ~new_n47556_ & ~new_n47624_;
  assign new_n47626_ = ys__n47942 & new_n47549_;
  assign new_n47627_ = ys__n47875 & ~new_n47553_;
  assign new_n47628_ = ~new_n47626_ & ~new_n47627_;
  assign ys__n32246 = ~new_n47556_ & ~new_n47628_;
  assign new_n47630_ = ys__n47943 & new_n47549_;
  assign new_n47631_ = ys__n47876 & ~new_n47553_;
  assign new_n47632_ = ~new_n47630_ & ~new_n47631_;
  assign ys__n32247 = ~new_n47556_ & ~new_n47632_;
  assign new_n47634_ = ys__n47944 & new_n47549_;
  assign new_n47635_ = ys__n47877 & ~new_n47553_;
  assign new_n47636_ = ~new_n47634_ & ~new_n47635_;
  assign ys__n32248 = ~new_n47556_ & ~new_n47636_;
  assign new_n47638_ = ys__n47945 & new_n47549_;
  assign new_n47639_ = ys__n47878 & ~new_n47553_;
  assign new_n47640_ = ~new_n47638_ & ~new_n47639_;
  assign ys__n32249 = ~new_n47556_ & ~new_n47640_;
  assign new_n47642_ = ys__n47946 & new_n47549_;
  assign new_n47643_ = ys__n47879 & ~new_n47553_;
  assign new_n47644_ = ~new_n47642_ & ~new_n47643_;
  assign ys__n32250 = ~new_n47556_ & ~new_n47644_;
  assign new_n47646_ = ys__n47947 & new_n47549_;
  assign new_n47647_ = ys__n47880 & ~new_n47553_;
  assign new_n47648_ = ~new_n47646_ & ~new_n47647_;
  assign ys__n32251 = ~new_n47556_ & ~new_n47648_;
  assign new_n47650_ = ys__n47948 & new_n47549_;
  assign new_n47651_ = ys__n47881 & ~new_n47553_;
  assign new_n47652_ = ~new_n47650_ & ~new_n47651_;
  assign ys__n32252 = ~new_n47556_ & ~new_n47652_;
  assign new_n47654_ = ys__n47949 & new_n47549_;
  assign new_n47655_ = ys__n47882 & ~new_n47553_;
  assign new_n47656_ = ~new_n47654_ & ~new_n47655_;
  assign ys__n32253 = ~new_n47556_ & ~new_n47656_;
  assign new_n47658_ = ys__n47950 & new_n47549_;
  assign new_n47659_ = ys__n47883 & ~new_n47553_;
  assign new_n47660_ = ~new_n47658_ & ~new_n47659_;
  assign ys__n32254 = ~new_n47556_ & ~new_n47660_;
  assign new_n47662_ = ys__n47951 & new_n47549_;
  assign new_n47663_ = ys__n47884 & ~new_n47553_;
  assign new_n47664_ = ~new_n47662_ & ~new_n47663_;
  assign ys__n32255 = ~new_n47556_ & ~new_n47664_;
  assign new_n47666_ = ys__n47952 & new_n47549_;
  assign new_n47667_ = ys__n47885 & ~new_n47553_;
  assign new_n47668_ = ~new_n47666_ & ~new_n47667_;
  assign ys__n32256 = ~new_n47556_ & ~new_n47668_;
  assign new_n47670_ = ys__n47953 & new_n47549_;
  assign new_n47671_ = ys__n47886 & ~new_n47553_;
  assign new_n47672_ = ~new_n47670_ & ~new_n47671_;
  assign ys__n32257 = ~new_n47556_ & ~new_n47672_;
  assign new_n47674_ = ys__n47954 & new_n47549_;
  assign new_n47675_ = ys__n47887 & ~new_n47553_;
  assign new_n47676_ = ~new_n47674_ & ~new_n47675_;
  assign ys__n32258 = ~new_n47556_ & ~new_n47676_;
  assign new_n47678_ = ys__n47955 & new_n47549_;
  assign new_n47679_ = ys__n47888 & ~new_n47553_;
  assign new_n47680_ = ~new_n47678_ & ~new_n47679_;
  assign ys__n32259 = ~new_n47556_ & ~new_n47680_;
  assign new_n47682_ = ys__n47956 & new_n47549_;
  assign new_n47683_ = ys__n19215 & ~new_n47553_;
  assign new_n47684_ = ~new_n47682_ & ~new_n47683_;
  assign ys__n32260 = ~new_n47556_ & ~new_n47684_;
  assign new_n47686_ = ys__n47957 & new_n47549_;
  assign new_n47687_ = ys__n47889 & ~new_n47553_;
  assign new_n47688_ = ~new_n47686_ & ~new_n47687_;
  assign ys__n32261 = ~new_n47556_ & ~new_n47688_;
  assign new_n47690_ = ys__n820 & ~new_n12860_;
  assign new_n47691_ = ys__n47958 & new_n47690_;
  assign new_n47692_ = ~ys__n822 & new_n12860_;
  assign new_n47693_ = ~ys__n820 & ~new_n12860_;
  assign new_n47694_ = ~new_n47692_ & ~new_n47693_;
  assign new_n47695_ = ys__n47857 & ~new_n47694_;
  assign new_n47696_ = ~new_n47691_ & ~new_n47695_;
  assign new_n47697_ = ~new_n47690_ & new_n47694_;
  assign ys__n32262 = ~new_n47696_ & ~new_n47697_;
  assign new_n47699_ = ys__n47959 & new_n47690_;
  assign new_n47700_ = ys__n47858 & ~new_n47694_;
  assign new_n47701_ = ~new_n47699_ & ~new_n47700_;
  assign ys__n32263 = ~new_n47697_ & ~new_n47701_;
  assign new_n47703_ = ys__n47960 & new_n47690_;
  assign new_n47704_ = ys__n47859 & ~new_n47694_;
  assign new_n47705_ = ~new_n47703_ & ~new_n47704_;
  assign ys__n32264 = ~new_n47697_ & ~new_n47705_;
  assign new_n47707_ = ys__n47961 & new_n47690_;
  assign new_n47708_ = ys__n47860 & ~new_n47694_;
  assign new_n47709_ = ~new_n47707_ & ~new_n47708_;
  assign ys__n32265 = ~new_n47697_ & ~new_n47709_;
  assign new_n47711_ = ys__n47962 & new_n47690_;
  assign new_n47712_ = ys__n47861 & ~new_n47694_;
  assign new_n47713_ = ~new_n47711_ & ~new_n47712_;
  assign ys__n32266 = ~new_n47697_ & ~new_n47713_;
  assign new_n47715_ = ys__n47963 & new_n47690_;
  assign new_n47716_ = ys__n47862 & ~new_n47694_;
  assign new_n47717_ = ~new_n47715_ & ~new_n47716_;
  assign ys__n32267 = ~new_n47697_ & ~new_n47717_;
  assign new_n47719_ = ys__n47964 & new_n47690_;
  assign new_n47720_ = ys__n47863 & ~new_n47694_;
  assign new_n47721_ = ~new_n47719_ & ~new_n47720_;
  assign ys__n32268 = ~new_n47697_ & ~new_n47721_;
  assign new_n47723_ = ys__n47965 & new_n47690_;
  assign new_n47724_ = ys__n47864 & ~new_n47694_;
  assign new_n47725_ = ~new_n47723_ & ~new_n47724_;
  assign ys__n32269 = ~new_n47697_ & ~new_n47725_;
  assign new_n47727_ = ys__n47966 & new_n47690_;
  assign new_n47728_ = ys__n47865 & ~new_n47694_;
  assign new_n47729_ = ~new_n47727_ & ~new_n47728_;
  assign ys__n32270 = ~new_n47697_ & ~new_n47729_;
  assign new_n47731_ = ys__n47967 & new_n47690_;
  assign new_n47732_ = ys__n47866 & ~new_n47694_;
  assign new_n47733_ = ~new_n47731_ & ~new_n47732_;
  assign ys__n32271 = ~new_n47697_ & ~new_n47733_;
  assign new_n47735_ = ys__n47968 & new_n47690_;
  assign new_n47736_ = ys__n47867 & ~new_n47694_;
  assign new_n47737_ = ~new_n47735_ & ~new_n47736_;
  assign ys__n32272 = ~new_n47697_ & ~new_n47737_;
  assign new_n47739_ = ys__n47969 & new_n47690_;
  assign new_n47740_ = ys__n47868 & ~new_n47694_;
  assign new_n47741_ = ~new_n47739_ & ~new_n47740_;
  assign ys__n32273 = ~new_n47697_ & ~new_n47741_;
  assign new_n47743_ = ys__n47970 & new_n47690_;
  assign new_n47744_ = ys__n47869 & ~new_n47694_;
  assign new_n47745_ = ~new_n47743_ & ~new_n47744_;
  assign ys__n32274 = ~new_n47697_ & ~new_n47745_;
  assign new_n47747_ = ys__n47971 & new_n47690_;
  assign new_n47748_ = ys__n47870 & ~new_n47694_;
  assign new_n47749_ = ~new_n47747_ & ~new_n47748_;
  assign ys__n32275 = ~new_n47697_ & ~new_n47749_;
  assign new_n47751_ = ys__n47972 & new_n47690_;
  assign new_n47752_ = ys__n47871 & ~new_n47694_;
  assign new_n47753_ = ~new_n47751_ & ~new_n47752_;
  assign ys__n32276 = ~new_n47697_ & ~new_n47753_;
  assign new_n47755_ = ys__n47973 & new_n47690_;
  assign new_n47756_ = ys__n47872 & ~new_n47694_;
  assign new_n47757_ = ~new_n47755_ & ~new_n47756_;
  assign ys__n32277 = ~new_n47697_ & ~new_n47757_;
  assign new_n47759_ = ys__n47974 & new_n47690_;
  assign new_n47760_ = ys__n47873 & ~new_n47694_;
  assign new_n47761_ = ~new_n47759_ & ~new_n47760_;
  assign ys__n32278 = ~new_n47697_ & ~new_n47761_;
  assign new_n47763_ = ys__n47975 & new_n47690_;
  assign new_n47764_ = ys__n47874 & ~new_n47694_;
  assign new_n47765_ = ~new_n47763_ & ~new_n47764_;
  assign ys__n32279 = ~new_n47697_ & ~new_n47765_;
  assign new_n47767_ = ys__n47976 & new_n47690_;
  assign new_n47768_ = ys__n47875 & ~new_n47694_;
  assign new_n47769_ = ~new_n47767_ & ~new_n47768_;
  assign ys__n32280 = ~new_n47697_ & ~new_n47769_;
  assign new_n47771_ = ys__n47977 & new_n47690_;
  assign new_n47772_ = ys__n47876 & ~new_n47694_;
  assign new_n47773_ = ~new_n47771_ & ~new_n47772_;
  assign ys__n32281 = ~new_n47697_ & ~new_n47773_;
  assign new_n47775_ = ys__n47978 & new_n47690_;
  assign new_n47776_ = ys__n47877 & ~new_n47694_;
  assign new_n47777_ = ~new_n47775_ & ~new_n47776_;
  assign ys__n32282 = ~new_n47697_ & ~new_n47777_;
  assign new_n47779_ = ys__n47979 & new_n47690_;
  assign new_n47780_ = ys__n47878 & ~new_n47694_;
  assign new_n47781_ = ~new_n47779_ & ~new_n47780_;
  assign ys__n32283 = ~new_n47697_ & ~new_n47781_;
  assign new_n47783_ = ys__n47980 & new_n47690_;
  assign new_n47784_ = ys__n47879 & ~new_n47694_;
  assign new_n47785_ = ~new_n47783_ & ~new_n47784_;
  assign ys__n32284 = ~new_n47697_ & ~new_n47785_;
  assign new_n47787_ = ys__n47981 & new_n47690_;
  assign new_n47788_ = ys__n47880 & ~new_n47694_;
  assign new_n47789_ = ~new_n47787_ & ~new_n47788_;
  assign ys__n32285 = ~new_n47697_ & ~new_n47789_;
  assign new_n47791_ = ys__n47982 & new_n47690_;
  assign new_n47792_ = ys__n47881 & ~new_n47694_;
  assign new_n47793_ = ~new_n47791_ & ~new_n47792_;
  assign ys__n32286 = ~new_n47697_ & ~new_n47793_;
  assign new_n47795_ = ys__n47983 & new_n47690_;
  assign new_n47796_ = ys__n47882 & ~new_n47694_;
  assign new_n47797_ = ~new_n47795_ & ~new_n47796_;
  assign ys__n32287 = ~new_n47697_ & ~new_n47797_;
  assign new_n47799_ = ys__n47984 & new_n47690_;
  assign new_n47800_ = ys__n47883 & ~new_n47694_;
  assign new_n47801_ = ~new_n47799_ & ~new_n47800_;
  assign ys__n32288 = ~new_n47697_ & ~new_n47801_;
  assign new_n47803_ = ys__n47985 & new_n47690_;
  assign new_n47804_ = ys__n47884 & ~new_n47694_;
  assign new_n47805_ = ~new_n47803_ & ~new_n47804_;
  assign ys__n32289 = ~new_n47697_ & ~new_n47805_;
  assign new_n47807_ = ys__n47986 & new_n47690_;
  assign new_n47808_ = ys__n47885 & ~new_n47694_;
  assign new_n47809_ = ~new_n47807_ & ~new_n47808_;
  assign ys__n32290 = ~new_n47697_ & ~new_n47809_;
  assign new_n47811_ = ys__n47987 & new_n47690_;
  assign new_n47812_ = ys__n47886 & ~new_n47694_;
  assign new_n47813_ = ~new_n47811_ & ~new_n47812_;
  assign ys__n32291 = ~new_n47697_ & ~new_n47813_;
  assign new_n47815_ = ys__n47988 & new_n47690_;
  assign new_n47816_ = ys__n47887 & ~new_n47694_;
  assign new_n47817_ = ~new_n47815_ & ~new_n47816_;
  assign ys__n32292 = ~new_n47697_ & ~new_n47817_;
  assign new_n47819_ = ys__n47989 & new_n47690_;
  assign new_n47820_ = ys__n47888 & ~new_n47694_;
  assign new_n47821_ = ~new_n47819_ & ~new_n47820_;
  assign ys__n32293 = ~new_n47697_ & ~new_n47821_;
  assign new_n47823_ = ys__n47990 & new_n47690_;
  assign new_n47824_ = ys__n19215 & ~new_n47694_;
  assign new_n47825_ = ~new_n47823_ & ~new_n47824_;
  assign ys__n32294 = ~new_n47697_ & ~new_n47825_;
  assign new_n47827_ = ys__n47991 & new_n47690_;
  assign new_n47828_ = ys__n47889 & ~new_n47694_;
  assign new_n47829_ = ~new_n47827_ & ~new_n47828_;
  assign ys__n32295 = ~new_n47697_ & ~new_n47829_;
  assign new_n47831_ = ys__n822 & ~new_n12860_;
  assign new_n47832_ = ys__n47992 & new_n47831_;
  assign new_n47833_ = ~ys__n824 & new_n12860_;
  assign new_n47834_ = ~ys__n822 & ~new_n12860_;
  assign new_n47835_ = ~new_n47833_ & ~new_n47834_;
  assign new_n47836_ = ys__n47857 & ~new_n47835_;
  assign new_n47837_ = ~new_n47832_ & ~new_n47836_;
  assign new_n47838_ = ~new_n47831_ & new_n47835_;
  assign ys__n32296 = ~new_n47837_ & ~new_n47838_;
  assign new_n47840_ = ys__n47993 & new_n47831_;
  assign new_n47841_ = ys__n47858 & ~new_n47835_;
  assign new_n47842_ = ~new_n47840_ & ~new_n47841_;
  assign ys__n32297 = ~new_n47838_ & ~new_n47842_;
  assign new_n47844_ = ys__n47994 & new_n47831_;
  assign new_n47845_ = ys__n47859 & ~new_n47835_;
  assign new_n47846_ = ~new_n47844_ & ~new_n47845_;
  assign ys__n32298 = ~new_n47838_ & ~new_n47846_;
  assign new_n47848_ = ys__n47995 & new_n47831_;
  assign new_n47849_ = ys__n47860 & ~new_n47835_;
  assign new_n47850_ = ~new_n47848_ & ~new_n47849_;
  assign ys__n32299 = ~new_n47838_ & ~new_n47850_;
  assign new_n47852_ = ys__n47996 & new_n47831_;
  assign new_n47853_ = ys__n47861 & ~new_n47835_;
  assign new_n47854_ = ~new_n47852_ & ~new_n47853_;
  assign ys__n32300 = ~new_n47838_ & ~new_n47854_;
  assign new_n47856_ = ys__n47997 & new_n47831_;
  assign new_n47857_ = ys__n47862 & ~new_n47835_;
  assign new_n47858_ = ~new_n47856_ & ~new_n47857_;
  assign ys__n32301 = ~new_n47838_ & ~new_n47858_;
  assign new_n47860_ = ys__n47998 & new_n47831_;
  assign new_n47861_ = ys__n47863 & ~new_n47835_;
  assign new_n47862_ = ~new_n47860_ & ~new_n47861_;
  assign ys__n32302 = ~new_n47838_ & ~new_n47862_;
  assign new_n47864_ = ys__n47999 & new_n47831_;
  assign new_n47865_ = ys__n47864 & ~new_n47835_;
  assign new_n47866_ = ~new_n47864_ & ~new_n47865_;
  assign ys__n32303 = ~new_n47838_ & ~new_n47866_;
  assign new_n47868_ = ys__n48000 & new_n47831_;
  assign new_n47869_ = ys__n47865 & ~new_n47835_;
  assign new_n47870_ = ~new_n47868_ & ~new_n47869_;
  assign ys__n32304 = ~new_n47838_ & ~new_n47870_;
  assign new_n47872_ = ys__n48001 & new_n47831_;
  assign new_n47873_ = ys__n47866 & ~new_n47835_;
  assign new_n47874_ = ~new_n47872_ & ~new_n47873_;
  assign ys__n32305 = ~new_n47838_ & ~new_n47874_;
  assign new_n47876_ = ys__n48002 & new_n47831_;
  assign new_n47877_ = ys__n47867 & ~new_n47835_;
  assign new_n47878_ = ~new_n47876_ & ~new_n47877_;
  assign ys__n32306 = ~new_n47838_ & ~new_n47878_;
  assign new_n47880_ = ys__n48003 & new_n47831_;
  assign new_n47881_ = ys__n47868 & ~new_n47835_;
  assign new_n47882_ = ~new_n47880_ & ~new_n47881_;
  assign ys__n32307 = ~new_n47838_ & ~new_n47882_;
  assign new_n47884_ = ys__n48004 & new_n47831_;
  assign new_n47885_ = ys__n47869 & ~new_n47835_;
  assign new_n47886_ = ~new_n47884_ & ~new_n47885_;
  assign ys__n32308 = ~new_n47838_ & ~new_n47886_;
  assign new_n47888_ = ys__n48005 & new_n47831_;
  assign new_n47889_ = ys__n47870 & ~new_n47835_;
  assign new_n47890_ = ~new_n47888_ & ~new_n47889_;
  assign ys__n32309 = ~new_n47838_ & ~new_n47890_;
  assign new_n47892_ = ys__n48006 & new_n47831_;
  assign new_n47893_ = ys__n47871 & ~new_n47835_;
  assign new_n47894_ = ~new_n47892_ & ~new_n47893_;
  assign ys__n32310 = ~new_n47838_ & ~new_n47894_;
  assign new_n47896_ = ys__n48007 & new_n47831_;
  assign new_n47897_ = ys__n47872 & ~new_n47835_;
  assign new_n47898_ = ~new_n47896_ & ~new_n47897_;
  assign ys__n32311 = ~new_n47838_ & ~new_n47898_;
  assign new_n47900_ = ys__n48008 & new_n47831_;
  assign new_n47901_ = ys__n47873 & ~new_n47835_;
  assign new_n47902_ = ~new_n47900_ & ~new_n47901_;
  assign ys__n32312 = ~new_n47838_ & ~new_n47902_;
  assign new_n47904_ = ys__n48009 & new_n47831_;
  assign new_n47905_ = ys__n47874 & ~new_n47835_;
  assign new_n47906_ = ~new_n47904_ & ~new_n47905_;
  assign ys__n32313 = ~new_n47838_ & ~new_n47906_;
  assign new_n47908_ = ys__n48010 & new_n47831_;
  assign new_n47909_ = ys__n47875 & ~new_n47835_;
  assign new_n47910_ = ~new_n47908_ & ~new_n47909_;
  assign ys__n32314 = ~new_n47838_ & ~new_n47910_;
  assign new_n47912_ = ys__n48011 & new_n47831_;
  assign new_n47913_ = ys__n47876 & ~new_n47835_;
  assign new_n47914_ = ~new_n47912_ & ~new_n47913_;
  assign ys__n32315 = ~new_n47838_ & ~new_n47914_;
  assign new_n47916_ = ys__n48012 & new_n47831_;
  assign new_n47917_ = ys__n47877 & ~new_n47835_;
  assign new_n47918_ = ~new_n47916_ & ~new_n47917_;
  assign ys__n32316 = ~new_n47838_ & ~new_n47918_;
  assign new_n47920_ = ys__n48013 & new_n47831_;
  assign new_n47921_ = ys__n47878 & ~new_n47835_;
  assign new_n47922_ = ~new_n47920_ & ~new_n47921_;
  assign ys__n32317 = ~new_n47838_ & ~new_n47922_;
  assign new_n47924_ = ys__n48014 & new_n47831_;
  assign new_n47925_ = ys__n47879 & ~new_n47835_;
  assign new_n47926_ = ~new_n47924_ & ~new_n47925_;
  assign ys__n32318 = ~new_n47838_ & ~new_n47926_;
  assign new_n47928_ = ys__n48015 & new_n47831_;
  assign new_n47929_ = ys__n47880 & ~new_n47835_;
  assign new_n47930_ = ~new_n47928_ & ~new_n47929_;
  assign ys__n32319 = ~new_n47838_ & ~new_n47930_;
  assign new_n47932_ = ys__n48016 & new_n47831_;
  assign new_n47933_ = ys__n47881 & ~new_n47835_;
  assign new_n47934_ = ~new_n47932_ & ~new_n47933_;
  assign ys__n32320 = ~new_n47838_ & ~new_n47934_;
  assign new_n47936_ = ys__n48017 & new_n47831_;
  assign new_n47937_ = ys__n47882 & ~new_n47835_;
  assign new_n47938_ = ~new_n47936_ & ~new_n47937_;
  assign ys__n32321 = ~new_n47838_ & ~new_n47938_;
  assign new_n47940_ = ys__n48018 & new_n47831_;
  assign new_n47941_ = ys__n47883 & ~new_n47835_;
  assign new_n47942_ = ~new_n47940_ & ~new_n47941_;
  assign ys__n32322 = ~new_n47838_ & ~new_n47942_;
  assign new_n47944_ = ys__n48019 & new_n47831_;
  assign new_n47945_ = ys__n47884 & ~new_n47835_;
  assign new_n47946_ = ~new_n47944_ & ~new_n47945_;
  assign ys__n32323 = ~new_n47838_ & ~new_n47946_;
  assign new_n47948_ = ys__n48020 & new_n47831_;
  assign new_n47949_ = ys__n47885 & ~new_n47835_;
  assign new_n47950_ = ~new_n47948_ & ~new_n47949_;
  assign ys__n32324 = ~new_n47838_ & ~new_n47950_;
  assign new_n47952_ = ys__n48021 & new_n47831_;
  assign new_n47953_ = ys__n47886 & ~new_n47835_;
  assign new_n47954_ = ~new_n47952_ & ~new_n47953_;
  assign ys__n32325 = ~new_n47838_ & ~new_n47954_;
  assign new_n47956_ = ys__n48022 & new_n47831_;
  assign new_n47957_ = ys__n47887 & ~new_n47835_;
  assign new_n47958_ = ~new_n47956_ & ~new_n47957_;
  assign ys__n32326 = ~new_n47838_ & ~new_n47958_;
  assign new_n47960_ = ys__n48023 & new_n47831_;
  assign new_n47961_ = ys__n47888 & ~new_n47835_;
  assign new_n47962_ = ~new_n47960_ & ~new_n47961_;
  assign ys__n32327 = ~new_n47838_ & ~new_n47962_;
  assign new_n47964_ = ys__n48024 & new_n47831_;
  assign new_n47965_ = ys__n19215 & ~new_n47835_;
  assign new_n47966_ = ~new_n47964_ & ~new_n47965_;
  assign ys__n32328 = ~new_n47838_ & ~new_n47966_;
  assign new_n47968_ = ys__n48025 & new_n47831_;
  assign new_n47969_ = ys__n47889 & ~new_n47835_;
  assign new_n47970_ = ~new_n47968_ & ~new_n47969_;
  assign ys__n32329 = ~new_n47838_ & ~new_n47970_;
  assign new_n47972_ = ys__n824 & ~new_n12860_;
  assign new_n47973_ = ys__n48026 & new_n47972_;
  assign new_n47974_ = ~ys__n826 & new_n12860_;
  assign new_n47975_ = ~ys__n824 & ~new_n12860_;
  assign new_n47976_ = ~new_n47974_ & ~new_n47975_;
  assign new_n47977_ = ys__n47857 & ~new_n47976_;
  assign new_n47978_ = ~new_n47973_ & ~new_n47977_;
  assign new_n47979_ = ~new_n47972_ & new_n47976_;
  assign ys__n32330 = ~new_n47978_ & ~new_n47979_;
  assign new_n47981_ = ys__n48027 & new_n47972_;
  assign new_n47982_ = ys__n47858 & ~new_n47976_;
  assign new_n47983_ = ~new_n47981_ & ~new_n47982_;
  assign ys__n32331 = ~new_n47979_ & ~new_n47983_;
  assign new_n47985_ = ys__n48028 & new_n47972_;
  assign new_n47986_ = ys__n47859 & ~new_n47976_;
  assign new_n47987_ = ~new_n47985_ & ~new_n47986_;
  assign ys__n32332 = ~new_n47979_ & ~new_n47987_;
  assign new_n47989_ = ys__n48029 & new_n47972_;
  assign new_n47990_ = ys__n47860 & ~new_n47976_;
  assign new_n47991_ = ~new_n47989_ & ~new_n47990_;
  assign ys__n32333 = ~new_n47979_ & ~new_n47991_;
  assign new_n47993_ = ys__n48030 & new_n47972_;
  assign new_n47994_ = ys__n47861 & ~new_n47976_;
  assign new_n47995_ = ~new_n47993_ & ~new_n47994_;
  assign ys__n32334 = ~new_n47979_ & ~new_n47995_;
  assign new_n47997_ = ys__n48031 & new_n47972_;
  assign new_n47998_ = ys__n47862 & ~new_n47976_;
  assign new_n47999_ = ~new_n47997_ & ~new_n47998_;
  assign ys__n32335 = ~new_n47979_ & ~new_n47999_;
  assign new_n48001_ = ys__n48032 & new_n47972_;
  assign new_n48002_ = ys__n47863 & ~new_n47976_;
  assign new_n48003_ = ~new_n48001_ & ~new_n48002_;
  assign ys__n32336 = ~new_n47979_ & ~new_n48003_;
  assign new_n48005_ = ys__n48033 & new_n47972_;
  assign new_n48006_ = ys__n47864 & ~new_n47976_;
  assign new_n48007_ = ~new_n48005_ & ~new_n48006_;
  assign ys__n32337 = ~new_n47979_ & ~new_n48007_;
  assign new_n48009_ = ys__n48034 & new_n47972_;
  assign new_n48010_ = ys__n47865 & ~new_n47976_;
  assign new_n48011_ = ~new_n48009_ & ~new_n48010_;
  assign ys__n32338 = ~new_n47979_ & ~new_n48011_;
  assign new_n48013_ = ys__n48035 & new_n47972_;
  assign new_n48014_ = ys__n47866 & ~new_n47976_;
  assign new_n48015_ = ~new_n48013_ & ~new_n48014_;
  assign ys__n32339 = ~new_n47979_ & ~new_n48015_;
  assign new_n48017_ = ys__n48036 & new_n47972_;
  assign new_n48018_ = ys__n47867 & ~new_n47976_;
  assign new_n48019_ = ~new_n48017_ & ~new_n48018_;
  assign ys__n32340 = ~new_n47979_ & ~new_n48019_;
  assign new_n48021_ = ys__n48037 & new_n47972_;
  assign new_n48022_ = ys__n47868 & ~new_n47976_;
  assign new_n48023_ = ~new_n48021_ & ~new_n48022_;
  assign ys__n32341 = ~new_n47979_ & ~new_n48023_;
  assign new_n48025_ = ys__n48038 & new_n47972_;
  assign new_n48026_ = ys__n47869 & ~new_n47976_;
  assign new_n48027_ = ~new_n48025_ & ~new_n48026_;
  assign ys__n32342 = ~new_n47979_ & ~new_n48027_;
  assign new_n48029_ = ys__n48039 & new_n47972_;
  assign new_n48030_ = ys__n47870 & ~new_n47976_;
  assign new_n48031_ = ~new_n48029_ & ~new_n48030_;
  assign ys__n32343 = ~new_n47979_ & ~new_n48031_;
  assign new_n48033_ = ys__n48040 & new_n47972_;
  assign new_n48034_ = ys__n47871 & ~new_n47976_;
  assign new_n48035_ = ~new_n48033_ & ~new_n48034_;
  assign ys__n32344 = ~new_n47979_ & ~new_n48035_;
  assign new_n48037_ = ys__n48041 & new_n47972_;
  assign new_n48038_ = ys__n47872 & ~new_n47976_;
  assign new_n48039_ = ~new_n48037_ & ~new_n48038_;
  assign ys__n32345 = ~new_n47979_ & ~new_n48039_;
  assign new_n48041_ = ys__n48042 & new_n47972_;
  assign new_n48042_ = ys__n47873 & ~new_n47976_;
  assign new_n48043_ = ~new_n48041_ & ~new_n48042_;
  assign ys__n32346 = ~new_n47979_ & ~new_n48043_;
  assign new_n48045_ = ys__n48043 & new_n47972_;
  assign new_n48046_ = ys__n47874 & ~new_n47976_;
  assign new_n48047_ = ~new_n48045_ & ~new_n48046_;
  assign ys__n32347 = ~new_n47979_ & ~new_n48047_;
  assign new_n48049_ = ys__n48044 & new_n47972_;
  assign new_n48050_ = ys__n47875 & ~new_n47976_;
  assign new_n48051_ = ~new_n48049_ & ~new_n48050_;
  assign ys__n32348 = ~new_n47979_ & ~new_n48051_;
  assign new_n48053_ = ys__n48045 & new_n47972_;
  assign new_n48054_ = ys__n47876 & ~new_n47976_;
  assign new_n48055_ = ~new_n48053_ & ~new_n48054_;
  assign ys__n32349 = ~new_n47979_ & ~new_n48055_;
  assign new_n48057_ = ys__n48046 & new_n47972_;
  assign new_n48058_ = ys__n47877 & ~new_n47976_;
  assign new_n48059_ = ~new_n48057_ & ~new_n48058_;
  assign ys__n32350 = ~new_n47979_ & ~new_n48059_;
  assign new_n48061_ = ys__n48047 & new_n47972_;
  assign new_n48062_ = ys__n47878 & ~new_n47976_;
  assign new_n48063_ = ~new_n48061_ & ~new_n48062_;
  assign ys__n32351 = ~new_n47979_ & ~new_n48063_;
  assign new_n48065_ = ys__n48048 & new_n47972_;
  assign new_n48066_ = ys__n47879 & ~new_n47976_;
  assign new_n48067_ = ~new_n48065_ & ~new_n48066_;
  assign ys__n32352 = ~new_n47979_ & ~new_n48067_;
  assign new_n48069_ = ys__n48049 & new_n47972_;
  assign new_n48070_ = ys__n47880 & ~new_n47976_;
  assign new_n48071_ = ~new_n48069_ & ~new_n48070_;
  assign ys__n32353 = ~new_n47979_ & ~new_n48071_;
  assign new_n48073_ = ys__n48050 & new_n47972_;
  assign new_n48074_ = ys__n47881 & ~new_n47976_;
  assign new_n48075_ = ~new_n48073_ & ~new_n48074_;
  assign ys__n32354 = ~new_n47979_ & ~new_n48075_;
  assign new_n48077_ = ys__n48051 & new_n47972_;
  assign new_n48078_ = ys__n47882 & ~new_n47976_;
  assign new_n48079_ = ~new_n48077_ & ~new_n48078_;
  assign ys__n32355 = ~new_n47979_ & ~new_n48079_;
  assign new_n48081_ = ys__n48052 & new_n47972_;
  assign new_n48082_ = ys__n47883 & ~new_n47976_;
  assign new_n48083_ = ~new_n48081_ & ~new_n48082_;
  assign ys__n32356 = ~new_n47979_ & ~new_n48083_;
  assign new_n48085_ = ys__n48053 & new_n47972_;
  assign new_n48086_ = ys__n47884 & ~new_n47976_;
  assign new_n48087_ = ~new_n48085_ & ~new_n48086_;
  assign ys__n32357 = ~new_n47979_ & ~new_n48087_;
  assign new_n48089_ = ys__n48054 & new_n47972_;
  assign new_n48090_ = ys__n47885 & ~new_n47976_;
  assign new_n48091_ = ~new_n48089_ & ~new_n48090_;
  assign ys__n32358 = ~new_n47979_ & ~new_n48091_;
  assign new_n48093_ = ys__n48055 & new_n47972_;
  assign new_n48094_ = ys__n47886 & ~new_n47976_;
  assign new_n48095_ = ~new_n48093_ & ~new_n48094_;
  assign ys__n32359 = ~new_n47979_ & ~new_n48095_;
  assign new_n48097_ = ys__n48056 & new_n47972_;
  assign new_n48098_ = ys__n47887 & ~new_n47976_;
  assign new_n48099_ = ~new_n48097_ & ~new_n48098_;
  assign ys__n32360 = ~new_n47979_ & ~new_n48099_;
  assign new_n48101_ = ys__n48057 & new_n47972_;
  assign new_n48102_ = ys__n47888 & ~new_n47976_;
  assign new_n48103_ = ~new_n48101_ & ~new_n48102_;
  assign ys__n32361 = ~new_n47979_ & ~new_n48103_;
  assign new_n48105_ = ys__n48058 & new_n47972_;
  assign new_n48106_ = ys__n19215 & ~new_n47976_;
  assign new_n48107_ = ~new_n48105_ & ~new_n48106_;
  assign ys__n32362 = ~new_n47979_ & ~new_n48107_;
  assign new_n48109_ = ys__n48059 & new_n47972_;
  assign new_n48110_ = ys__n47889 & ~new_n47976_;
  assign new_n48111_ = ~new_n48109_ & ~new_n48110_;
  assign ys__n32363 = ~new_n47979_ & ~new_n48111_;
  assign new_n48113_ = ys__n826 & ~new_n12860_;
  assign new_n48114_ = ys__n48060 & new_n48113_;
  assign new_n48115_ = ~ys__n828 & new_n12860_;
  assign new_n48116_ = ~ys__n826 & ~new_n12860_;
  assign new_n48117_ = ~new_n48115_ & ~new_n48116_;
  assign new_n48118_ = ys__n47857 & ~new_n48117_;
  assign new_n48119_ = ~new_n48114_ & ~new_n48118_;
  assign new_n48120_ = ~new_n48113_ & new_n48117_;
  assign ys__n32364 = ~new_n48119_ & ~new_n48120_;
  assign new_n48122_ = ys__n48061 & new_n48113_;
  assign new_n48123_ = ys__n47858 & ~new_n48117_;
  assign new_n48124_ = ~new_n48122_ & ~new_n48123_;
  assign ys__n32365 = ~new_n48120_ & ~new_n48124_;
  assign new_n48126_ = ys__n48062 & new_n48113_;
  assign new_n48127_ = ys__n47859 & ~new_n48117_;
  assign new_n48128_ = ~new_n48126_ & ~new_n48127_;
  assign ys__n32366 = ~new_n48120_ & ~new_n48128_;
  assign new_n48130_ = ys__n48063 & new_n48113_;
  assign new_n48131_ = ys__n47860 & ~new_n48117_;
  assign new_n48132_ = ~new_n48130_ & ~new_n48131_;
  assign ys__n32367 = ~new_n48120_ & ~new_n48132_;
  assign new_n48134_ = ys__n48064 & new_n48113_;
  assign new_n48135_ = ys__n47861 & ~new_n48117_;
  assign new_n48136_ = ~new_n48134_ & ~new_n48135_;
  assign ys__n32368 = ~new_n48120_ & ~new_n48136_;
  assign new_n48138_ = ys__n48065 & new_n48113_;
  assign new_n48139_ = ys__n47862 & ~new_n48117_;
  assign new_n48140_ = ~new_n48138_ & ~new_n48139_;
  assign ys__n32369 = ~new_n48120_ & ~new_n48140_;
  assign new_n48142_ = ys__n48066 & new_n48113_;
  assign new_n48143_ = ys__n47863 & ~new_n48117_;
  assign new_n48144_ = ~new_n48142_ & ~new_n48143_;
  assign ys__n32370 = ~new_n48120_ & ~new_n48144_;
  assign new_n48146_ = ys__n48067 & new_n48113_;
  assign new_n48147_ = ys__n47864 & ~new_n48117_;
  assign new_n48148_ = ~new_n48146_ & ~new_n48147_;
  assign ys__n32371 = ~new_n48120_ & ~new_n48148_;
  assign new_n48150_ = ys__n48068 & new_n48113_;
  assign new_n48151_ = ys__n47865 & ~new_n48117_;
  assign new_n48152_ = ~new_n48150_ & ~new_n48151_;
  assign ys__n32372 = ~new_n48120_ & ~new_n48152_;
  assign new_n48154_ = ys__n48069 & new_n48113_;
  assign new_n48155_ = ys__n47866 & ~new_n48117_;
  assign new_n48156_ = ~new_n48154_ & ~new_n48155_;
  assign ys__n32373 = ~new_n48120_ & ~new_n48156_;
  assign new_n48158_ = ys__n48070 & new_n48113_;
  assign new_n48159_ = ys__n47867 & ~new_n48117_;
  assign new_n48160_ = ~new_n48158_ & ~new_n48159_;
  assign ys__n32374 = ~new_n48120_ & ~new_n48160_;
  assign new_n48162_ = ys__n48071 & new_n48113_;
  assign new_n48163_ = ys__n47868 & ~new_n48117_;
  assign new_n48164_ = ~new_n48162_ & ~new_n48163_;
  assign ys__n32375 = ~new_n48120_ & ~new_n48164_;
  assign new_n48166_ = ys__n48072 & new_n48113_;
  assign new_n48167_ = ys__n47869 & ~new_n48117_;
  assign new_n48168_ = ~new_n48166_ & ~new_n48167_;
  assign ys__n32376 = ~new_n48120_ & ~new_n48168_;
  assign new_n48170_ = ys__n48073 & new_n48113_;
  assign new_n48171_ = ys__n47870 & ~new_n48117_;
  assign new_n48172_ = ~new_n48170_ & ~new_n48171_;
  assign ys__n32377 = ~new_n48120_ & ~new_n48172_;
  assign new_n48174_ = ys__n48074 & new_n48113_;
  assign new_n48175_ = ys__n47871 & ~new_n48117_;
  assign new_n48176_ = ~new_n48174_ & ~new_n48175_;
  assign ys__n32378 = ~new_n48120_ & ~new_n48176_;
  assign new_n48178_ = ys__n48075 & new_n48113_;
  assign new_n48179_ = ys__n47872 & ~new_n48117_;
  assign new_n48180_ = ~new_n48178_ & ~new_n48179_;
  assign ys__n32379 = ~new_n48120_ & ~new_n48180_;
  assign new_n48182_ = ys__n48076 & new_n48113_;
  assign new_n48183_ = ys__n47873 & ~new_n48117_;
  assign new_n48184_ = ~new_n48182_ & ~new_n48183_;
  assign ys__n32380 = ~new_n48120_ & ~new_n48184_;
  assign new_n48186_ = ys__n48077 & new_n48113_;
  assign new_n48187_ = ys__n47874 & ~new_n48117_;
  assign new_n48188_ = ~new_n48186_ & ~new_n48187_;
  assign ys__n32381 = ~new_n48120_ & ~new_n48188_;
  assign new_n48190_ = ys__n48078 & new_n48113_;
  assign new_n48191_ = ys__n47875 & ~new_n48117_;
  assign new_n48192_ = ~new_n48190_ & ~new_n48191_;
  assign ys__n32382 = ~new_n48120_ & ~new_n48192_;
  assign new_n48194_ = ys__n48079 & new_n48113_;
  assign new_n48195_ = ys__n47876 & ~new_n48117_;
  assign new_n48196_ = ~new_n48194_ & ~new_n48195_;
  assign ys__n32383 = ~new_n48120_ & ~new_n48196_;
  assign new_n48198_ = ys__n48080 & new_n48113_;
  assign new_n48199_ = ys__n47877 & ~new_n48117_;
  assign new_n48200_ = ~new_n48198_ & ~new_n48199_;
  assign ys__n32384 = ~new_n48120_ & ~new_n48200_;
  assign new_n48202_ = ys__n48081 & new_n48113_;
  assign new_n48203_ = ys__n47878 & ~new_n48117_;
  assign new_n48204_ = ~new_n48202_ & ~new_n48203_;
  assign ys__n32385 = ~new_n48120_ & ~new_n48204_;
  assign new_n48206_ = ys__n48082 & new_n48113_;
  assign new_n48207_ = ys__n47879 & ~new_n48117_;
  assign new_n48208_ = ~new_n48206_ & ~new_n48207_;
  assign ys__n32386 = ~new_n48120_ & ~new_n48208_;
  assign new_n48210_ = ys__n48083 & new_n48113_;
  assign new_n48211_ = ys__n47880 & ~new_n48117_;
  assign new_n48212_ = ~new_n48210_ & ~new_n48211_;
  assign ys__n32387 = ~new_n48120_ & ~new_n48212_;
  assign new_n48214_ = ys__n48084 & new_n48113_;
  assign new_n48215_ = ys__n47881 & ~new_n48117_;
  assign new_n48216_ = ~new_n48214_ & ~new_n48215_;
  assign ys__n32388 = ~new_n48120_ & ~new_n48216_;
  assign new_n48218_ = ys__n48085 & new_n48113_;
  assign new_n48219_ = ys__n47882 & ~new_n48117_;
  assign new_n48220_ = ~new_n48218_ & ~new_n48219_;
  assign ys__n32389 = ~new_n48120_ & ~new_n48220_;
  assign new_n48222_ = ys__n48086 & new_n48113_;
  assign new_n48223_ = ys__n47883 & ~new_n48117_;
  assign new_n48224_ = ~new_n48222_ & ~new_n48223_;
  assign ys__n32390 = ~new_n48120_ & ~new_n48224_;
  assign new_n48226_ = ys__n48087 & new_n48113_;
  assign new_n48227_ = ys__n47884 & ~new_n48117_;
  assign new_n48228_ = ~new_n48226_ & ~new_n48227_;
  assign ys__n32391 = ~new_n48120_ & ~new_n48228_;
  assign new_n48230_ = ys__n48088 & new_n48113_;
  assign new_n48231_ = ys__n47885 & ~new_n48117_;
  assign new_n48232_ = ~new_n48230_ & ~new_n48231_;
  assign ys__n32392 = ~new_n48120_ & ~new_n48232_;
  assign new_n48234_ = ys__n48089 & new_n48113_;
  assign new_n48235_ = ys__n47886 & ~new_n48117_;
  assign new_n48236_ = ~new_n48234_ & ~new_n48235_;
  assign ys__n32393 = ~new_n48120_ & ~new_n48236_;
  assign new_n48238_ = ys__n48090 & new_n48113_;
  assign new_n48239_ = ys__n47887 & ~new_n48117_;
  assign new_n48240_ = ~new_n48238_ & ~new_n48239_;
  assign ys__n32394 = ~new_n48120_ & ~new_n48240_;
  assign new_n48242_ = ys__n48091 & new_n48113_;
  assign new_n48243_ = ys__n47888 & ~new_n48117_;
  assign new_n48244_ = ~new_n48242_ & ~new_n48243_;
  assign ys__n32395 = ~new_n48120_ & ~new_n48244_;
  assign new_n48246_ = ys__n48092 & new_n48113_;
  assign new_n48247_ = ys__n19215 & ~new_n48117_;
  assign new_n48248_ = ~new_n48246_ & ~new_n48247_;
  assign ys__n32396 = ~new_n48120_ & ~new_n48248_;
  assign new_n48250_ = ys__n48093 & new_n48113_;
  assign new_n48251_ = ys__n47889 & ~new_n48117_;
  assign new_n48252_ = ~new_n48250_ & ~new_n48251_;
  assign ys__n32397 = ~new_n48120_ & ~new_n48252_;
  assign new_n48254_ = ys__n116 & new_n13240_;
  assign new_n48255_ = ys__n48094 & new_n48254_;
  assign new_n48256_ = ~ys__n846 & ~new_n13240_;
  assign new_n48257_ = ~ys__n116 & new_n13240_;
  assign new_n48258_ = ~new_n48256_ & ~new_n48257_;
  assign new_n48259_ = ys__n18654 & ~new_n48258_;
  assign new_n48260_ = ~new_n48255_ & ~new_n48259_;
  assign new_n48261_ = ~new_n48254_ & new_n48258_;
  assign ys__n32398 = ~new_n48260_ & ~new_n48261_;
  assign new_n48263_ = ys__n48095 & new_n48254_;
  assign new_n48264_ = ys__n18657 & ~new_n48258_;
  assign new_n48265_ = ~new_n48263_ & ~new_n48264_;
  assign ys__n32399 = ~new_n48261_ & ~new_n48265_;
  assign new_n48267_ = ys__n48096 & new_n48254_;
  assign new_n48268_ = ys__n18660 & ~new_n48258_;
  assign new_n48269_ = ~new_n48267_ & ~new_n48268_;
  assign ys__n32400 = ~new_n48261_ & ~new_n48269_;
  assign new_n48271_ = ys__n48097 & new_n48254_;
  assign new_n48272_ = ys__n18663 & ~new_n48258_;
  assign new_n48273_ = ~new_n48271_ & ~new_n48272_;
  assign ys__n32401 = ~new_n48261_ & ~new_n48273_;
  assign new_n48275_ = ys__n37758 & new_n48254_;
  assign new_n48276_ = ys__n18666 & ~new_n48258_;
  assign new_n48277_ = ~new_n48275_ & ~new_n48276_;
  assign ys__n32402 = ~new_n48261_ & ~new_n48277_;
  assign new_n48279_ = ys__n37759 & new_n48254_;
  assign new_n48280_ = ys__n18669 & ~new_n48258_;
  assign new_n48281_ = ~new_n48279_ & ~new_n48280_;
  assign ys__n32403 = ~new_n48261_ & ~new_n48281_;
  assign new_n48283_ = ys__n37760 & new_n48254_;
  assign new_n48284_ = ys__n18672 & ~new_n48258_;
  assign new_n48285_ = ~new_n48283_ & ~new_n48284_;
  assign ys__n32404 = ~new_n48261_ & ~new_n48285_;
  assign new_n48287_ = ys__n37761 & new_n48254_;
  assign new_n48288_ = ys__n18675 & ~new_n48258_;
  assign new_n48289_ = ~new_n48287_ & ~new_n48288_;
  assign ys__n32405 = ~new_n48261_ & ~new_n48289_;
  assign new_n48291_ = ys__n37762 & new_n48254_;
  assign new_n48292_ = ys__n18678 & ~new_n48258_;
  assign new_n48293_ = ~new_n48291_ & ~new_n48292_;
  assign ys__n32406 = ~new_n48261_ & ~new_n48293_;
  assign new_n48295_ = ys__n37763 & new_n48254_;
  assign new_n48296_ = ys__n18681 & ~new_n48258_;
  assign new_n48297_ = ~new_n48295_ & ~new_n48296_;
  assign ys__n32407 = ~new_n48261_ & ~new_n48297_;
  assign new_n48299_ = ys__n37764 & new_n48254_;
  assign new_n48300_ = ys__n18684 & ~new_n48258_;
  assign new_n48301_ = ~new_n48299_ & ~new_n48300_;
  assign ys__n32408 = ~new_n48261_ & ~new_n48301_;
  assign new_n48303_ = ys__n37765 & new_n48254_;
  assign new_n48304_ = ys__n18687 & ~new_n48258_;
  assign new_n48305_ = ~new_n48303_ & ~new_n48304_;
  assign ys__n32409 = ~new_n48261_ & ~new_n48305_;
  assign new_n48307_ = ys__n37766 & new_n48254_;
  assign new_n48308_ = ys__n18690 & ~new_n48258_;
  assign new_n48309_ = ~new_n48307_ & ~new_n48308_;
  assign ys__n32410 = ~new_n48261_ & ~new_n48309_;
  assign new_n48311_ = ys__n37767 & new_n48254_;
  assign new_n48312_ = ys__n18693 & ~new_n48258_;
  assign new_n48313_ = ~new_n48311_ & ~new_n48312_;
  assign ys__n32411 = ~new_n48261_ & ~new_n48313_;
  assign new_n48315_ = ys__n37768 & new_n48254_;
  assign new_n48316_ = ys__n18696 & ~new_n48258_;
  assign new_n48317_ = ~new_n48315_ & ~new_n48316_;
  assign ys__n32412 = ~new_n48261_ & ~new_n48317_;
  assign new_n48319_ = ys__n37769 & new_n48254_;
  assign new_n48320_ = ys__n18699 & ~new_n48258_;
  assign new_n48321_ = ~new_n48319_ & ~new_n48320_;
  assign ys__n32413 = ~new_n48261_ & ~new_n48321_;
  assign new_n48323_ = ys__n37770 & new_n48254_;
  assign new_n48324_ = ys__n18702 & ~new_n48258_;
  assign new_n48325_ = ~new_n48323_ & ~new_n48324_;
  assign ys__n32414 = ~new_n48261_ & ~new_n48325_;
  assign new_n48327_ = ys__n37771 & new_n48254_;
  assign new_n48328_ = ys__n18705 & ~new_n48258_;
  assign new_n48329_ = ~new_n48327_ & ~new_n48328_;
  assign ys__n32415 = ~new_n48261_ & ~new_n48329_;
  assign new_n48331_ = ys__n37772 & new_n48254_;
  assign new_n48332_ = ys__n18708 & ~new_n48258_;
  assign new_n48333_ = ~new_n48331_ & ~new_n48332_;
  assign ys__n32416 = ~new_n48261_ & ~new_n48333_;
  assign new_n48335_ = ys__n37773 & new_n48254_;
  assign new_n48336_ = ys__n18711 & ~new_n48258_;
  assign new_n48337_ = ~new_n48335_ & ~new_n48336_;
  assign ys__n32417 = ~new_n48261_ & ~new_n48337_;
  assign new_n48339_ = ys__n37774 & new_n48254_;
  assign new_n48340_ = ys__n18714 & ~new_n48258_;
  assign new_n48341_ = ~new_n48339_ & ~new_n48340_;
  assign ys__n32418 = ~new_n48261_ & ~new_n48341_;
  assign new_n48343_ = ys__n37775 & new_n48254_;
  assign new_n48344_ = ys__n18717 & ~new_n48258_;
  assign new_n48345_ = ~new_n48343_ & ~new_n48344_;
  assign ys__n32419 = ~new_n48261_ & ~new_n48345_;
  assign new_n48347_ = ys__n37776 & new_n48254_;
  assign new_n48348_ = ys__n18720 & ~new_n48258_;
  assign new_n48349_ = ~new_n48347_ & ~new_n48348_;
  assign ys__n32420 = ~new_n48261_ & ~new_n48349_;
  assign new_n48351_ = ys__n37777 & new_n48254_;
  assign new_n48352_ = ys__n18723 & ~new_n48258_;
  assign new_n48353_ = ~new_n48351_ & ~new_n48352_;
  assign ys__n32421 = ~new_n48261_ & ~new_n48353_;
  assign new_n48355_ = ys__n37778 & new_n48254_;
  assign new_n48356_ = ys__n18726 & ~new_n48258_;
  assign new_n48357_ = ~new_n48355_ & ~new_n48356_;
  assign ys__n32422 = ~new_n48261_ & ~new_n48357_;
  assign new_n48359_ = ys__n37779 & new_n48254_;
  assign new_n48360_ = ys__n18729 & ~new_n48258_;
  assign new_n48361_ = ~new_n48359_ & ~new_n48360_;
  assign ys__n32423 = ~new_n48261_ & ~new_n48361_;
  assign new_n48363_ = ys__n37780 & new_n48254_;
  assign new_n48364_ = ys__n18732 & ~new_n48258_;
  assign new_n48365_ = ~new_n48363_ & ~new_n48364_;
  assign ys__n32424 = ~new_n48261_ & ~new_n48365_;
  assign new_n48367_ = ys__n37781 & new_n48254_;
  assign new_n48368_ = ys__n18735 & ~new_n48258_;
  assign new_n48369_ = ~new_n48367_ & ~new_n48368_;
  assign ys__n32425 = ~new_n48261_ & ~new_n48369_;
  assign new_n48371_ = ys__n37782 & new_n48254_;
  assign new_n48372_ = ys__n18738 & ~new_n48258_;
  assign new_n48373_ = ~new_n48371_ & ~new_n48372_;
  assign ys__n32426 = ~new_n48261_ & ~new_n48373_;
  assign new_n48375_ = ys__n37783 & new_n48254_;
  assign new_n48376_ = ys__n18741 & ~new_n48258_;
  assign new_n48377_ = ~new_n48375_ & ~new_n48376_;
  assign ys__n32427 = ~new_n48261_ & ~new_n48377_;
  assign new_n48379_ = ys__n37784 & new_n48254_;
  assign new_n48380_ = ys__n18744 & ~new_n48258_;
  assign new_n48381_ = ~new_n48379_ & ~new_n48380_;
  assign ys__n32428 = ~new_n48261_ & ~new_n48381_;
  assign new_n48383_ = ys__n37785 & new_n48254_;
  assign new_n48384_ = ys__n18747 & ~new_n48258_;
  assign new_n48385_ = ~new_n48383_ & ~new_n48384_;
  assign ys__n32429 = ~new_n48261_ & ~new_n48385_;
  assign new_n48387_ = ys__n846 & new_n13240_;
  assign new_n48388_ = ys__n48098 & new_n48387_;
  assign new_n48389_ = ~ys__n848 & ~new_n13240_;
  assign new_n48390_ = ~ys__n846 & new_n13240_;
  assign new_n48391_ = ~new_n48389_ & ~new_n48390_;
  assign new_n48392_ = ys__n18654 & ~new_n48391_;
  assign new_n48393_ = ~new_n48388_ & ~new_n48392_;
  assign new_n48394_ = ~new_n48387_ & new_n48391_;
  assign ys__n32430 = ~new_n48393_ & ~new_n48394_;
  assign new_n48396_ = ys__n48099 & new_n48387_;
  assign new_n48397_ = ys__n18657 & ~new_n48391_;
  assign new_n48398_ = ~new_n48396_ & ~new_n48397_;
  assign ys__n32431 = ~new_n48394_ & ~new_n48398_;
  assign new_n48400_ = ys__n48100 & new_n48387_;
  assign new_n48401_ = ys__n18660 & ~new_n48391_;
  assign new_n48402_ = ~new_n48400_ & ~new_n48401_;
  assign ys__n32432 = ~new_n48394_ & ~new_n48402_;
  assign new_n48404_ = ys__n48101 & new_n48387_;
  assign new_n48405_ = ys__n18663 & ~new_n48391_;
  assign new_n48406_ = ~new_n48404_ & ~new_n48405_;
  assign ys__n32433 = ~new_n48394_ & ~new_n48406_;
  assign new_n48408_ = ys__n37786 & new_n48387_;
  assign new_n48409_ = ys__n18666 & ~new_n48391_;
  assign new_n48410_ = ~new_n48408_ & ~new_n48409_;
  assign ys__n32434 = ~new_n48394_ & ~new_n48410_;
  assign new_n48412_ = ys__n37787 & new_n48387_;
  assign new_n48413_ = ys__n18669 & ~new_n48391_;
  assign new_n48414_ = ~new_n48412_ & ~new_n48413_;
  assign ys__n32435 = ~new_n48394_ & ~new_n48414_;
  assign new_n48416_ = ys__n37788 & new_n48387_;
  assign new_n48417_ = ys__n18672 & ~new_n48391_;
  assign new_n48418_ = ~new_n48416_ & ~new_n48417_;
  assign ys__n32436 = ~new_n48394_ & ~new_n48418_;
  assign new_n48420_ = ys__n37789 & new_n48387_;
  assign new_n48421_ = ys__n18675 & ~new_n48391_;
  assign new_n48422_ = ~new_n48420_ & ~new_n48421_;
  assign ys__n32437 = ~new_n48394_ & ~new_n48422_;
  assign new_n48424_ = ys__n37790 & new_n48387_;
  assign new_n48425_ = ys__n18678 & ~new_n48391_;
  assign new_n48426_ = ~new_n48424_ & ~new_n48425_;
  assign ys__n32438 = ~new_n48394_ & ~new_n48426_;
  assign new_n48428_ = ys__n37791 & new_n48387_;
  assign new_n48429_ = ys__n18681 & ~new_n48391_;
  assign new_n48430_ = ~new_n48428_ & ~new_n48429_;
  assign ys__n32439 = ~new_n48394_ & ~new_n48430_;
  assign new_n48432_ = ys__n37792 & new_n48387_;
  assign new_n48433_ = ys__n18684 & ~new_n48391_;
  assign new_n48434_ = ~new_n48432_ & ~new_n48433_;
  assign ys__n32440 = ~new_n48394_ & ~new_n48434_;
  assign new_n48436_ = ys__n37793 & new_n48387_;
  assign new_n48437_ = ys__n18687 & ~new_n48391_;
  assign new_n48438_ = ~new_n48436_ & ~new_n48437_;
  assign ys__n32441 = ~new_n48394_ & ~new_n48438_;
  assign new_n48440_ = ys__n37794 & new_n48387_;
  assign new_n48441_ = ys__n18690 & ~new_n48391_;
  assign new_n48442_ = ~new_n48440_ & ~new_n48441_;
  assign ys__n32442 = ~new_n48394_ & ~new_n48442_;
  assign new_n48444_ = ys__n37795 & new_n48387_;
  assign new_n48445_ = ys__n18693 & ~new_n48391_;
  assign new_n48446_ = ~new_n48444_ & ~new_n48445_;
  assign ys__n32443 = ~new_n48394_ & ~new_n48446_;
  assign new_n48448_ = ys__n37796 & new_n48387_;
  assign new_n48449_ = ys__n18696 & ~new_n48391_;
  assign new_n48450_ = ~new_n48448_ & ~new_n48449_;
  assign ys__n32444 = ~new_n48394_ & ~new_n48450_;
  assign new_n48452_ = ys__n37797 & new_n48387_;
  assign new_n48453_ = ys__n18699 & ~new_n48391_;
  assign new_n48454_ = ~new_n48452_ & ~new_n48453_;
  assign ys__n32445 = ~new_n48394_ & ~new_n48454_;
  assign new_n48456_ = ys__n37798 & new_n48387_;
  assign new_n48457_ = ys__n18702 & ~new_n48391_;
  assign new_n48458_ = ~new_n48456_ & ~new_n48457_;
  assign ys__n32446 = ~new_n48394_ & ~new_n48458_;
  assign new_n48460_ = ys__n37799 & new_n48387_;
  assign new_n48461_ = ys__n18705 & ~new_n48391_;
  assign new_n48462_ = ~new_n48460_ & ~new_n48461_;
  assign ys__n32447 = ~new_n48394_ & ~new_n48462_;
  assign new_n48464_ = ys__n37800 & new_n48387_;
  assign new_n48465_ = ys__n18708 & ~new_n48391_;
  assign new_n48466_ = ~new_n48464_ & ~new_n48465_;
  assign ys__n32448 = ~new_n48394_ & ~new_n48466_;
  assign new_n48468_ = ys__n37801 & new_n48387_;
  assign new_n48469_ = ys__n18711 & ~new_n48391_;
  assign new_n48470_ = ~new_n48468_ & ~new_n48469_;
  assign ys__n32449 = ~new_n48394_ & ~new_n48470_;
  assign new_n48472_ = ys__n37802 & new_n48387_;
  assign new_n48473_ = ys__n18714 & ~new_n48391_;
  assign new_n48474_ = ~new_n48472_ & ~new_n48473_;
  assign ys__n32450 = ~new_n48394_ & ~new_n48474_;
  assign new_n48476_ = ys__n37803 & new_n48387_;
  assign new_n48477_ = ys__n18717 & ~new_n48391_;
  assign new_n48478_ = ~new_n48476_ & ~new_n48477_;
  assign ys__n32451 = ~new_n48394_ & ~new_n48478_;
  assign new_n48480_ = ys__n37804 & new_n48387_;
  assign new_n48481_ = ys__n18720 & ~new_n48391_;
  assign new_n48482_ = ~new_n48480_ & ~new_n48481_;
  assign ys__n32452 = ~new_n48394_ & ~new_n48482_;
  assign new_n48484_ = ys__n37805 & new_n48387_;
  assign new_n48485_ = ys__n18723 & ~new_n48391_;
  assign new_n48486_ = ~new_n48484_ & ~new_n48485_;
  assign ys__n32453 = ~new_n48394_ & ~new_n48486_;
  assign new_n48488_ = ys__n37806 & new_n48387_;
  assign new_n48489_ = ys__n18726 & ~new_n48391_;
  assign new_n48490_ = ~new_n48488_ & ~new_n48489_;
  assign ys__n32454 = ~new_n48394_ & ~new_n48490_;
  assign new_n48492_ = ys__n37807 & new_n48387_;
  assign new_n48493_ = ys__n18729 & ~new_n48391_;
  assign new_n48494_ = ~new_n48492_ & ~new_n48493_;
  assign ys__n32455 = ~new_n48394_ & ~new_n48494_;
  assign new_n48496_ = ys__n37808 & new_n48387_;
  assign new_n48497_ = ys__n18732 & ~new_n48391_;
  assign new_n48498_ = ~new_n48496_ & ~new_n48497_;
  assign ys__n32456 = ~new_n48394_ & ~new_n48498_;
  assign new_n48500_ = ys__n37809 & new_n48387_;
  assign new_n48501_ = ys__n18735 & ~new_n48391_;
  assign new_n48502_ = ~new_n48500_ & ~new_n48501_;
  assign ys__n32457 = ~new_n48394_ & ~new_n48502_;
  assign new_n48504_ = ys__n37810 & new_n48387_;
  assign new_n48505_ = ys__n18738 & ~new_n48391_;
  assign new_n48506_ = ~new_n48504_ & ~new_n48505_;
  assign ys__n32458 = ~new_n48394_ & ~new_n48506_;
  assign new_n48508_ = ys__n37811 & new_n48387_;
  assign new_n48509_ = ys__n18741 & ~new_n48391_;
  assign new_n48510_ = ~new_n48508_ & ~new_n48509_;
  assign ys__n32459 = ~new_n48394_ & ~new_n48510_;
  assign new_n48512_ = ys__n37812 & new_n48387_;
  assign new_n48513_ = ys__n18744 & ~new_n48391_;
  assign new_n48514_ = ~new_n48512_ & ~new_n48513_;
  assign ys__n32460 = ~new_n48394_ & ~new_n48514_;
  assign new_n48516_ = ys__n37813 & new_n48387_;
  assign new_n48517_ = ys__n18747 & ~new_n48391_;
  assign new_n48518_ = ~new_n48516_ & ~new_n48517_;
  assign ys__n32461 = ~new_n48394_ & ~new_n48518_;
  assign new_n48520_ = ys__n848 & new_n13240_;
  assign new_n48521_ = ys__n48102 & new_n48520_;
  assign new_n48522_ = ~ys__n850 & ~new_n13240_;
  assign new_n48523_ = ~ys__n848 & new_n13240_;
  assign new_n48524_ = ~new_n48522_ & ~new_n48523_;
  assign new_n48525_ = ys__n18654 & ~new_n48524_;
  assign new_n48526_ = ~new_n48521_ & ~new_n48525_;
  assign new_n48527_ = ~new_n48520_ & new_n48524_;
  assign ys__n32462 = ~new_n48526_ & ~new_n48527_;
  assign new_n48529_ = ys__n48103 & new_n48520_;
  assign new_n48530_ = ys__n18657 & ~new_n48524_;
  assign new_n48531_ = ~new_n48529_ & ~new_n48530_;
  assign ys__n32463 = ~new_n48527_ & ~new_n48531_;
  assign new_n48533_ = ys__n48104 & new_n48520_;
  assign new_n48534_ = ys__n18660 & ~new_n48524_;
  assign new_n48535_ = ~new_n48533_ & ~new_n48534_;
  assign ys__n32464 = ~new_n48527_ & ~new_n48535_;
  assign new_n48537_ = ys__n48105 & new_n48520_;
  assign new_n48538_ = ys__n18663 & ~new_n48524_;
  assign new_n48539_ = ~new_n48537_ & ~new_n48538_;
  assign ys__n32465 = ~new_n48527_ & ~new_n48539_;
  assign new_n48541_ = ys__n37814 & new_n48520_;
  assign new_n48542_ = ys__n18666 & ~new_n48524_;
  assign new_n48543_ = ~new_n48541_ & ~new_n48542_;
  assign ys__n32466 = ~new_n48527_ & ~new_n48543_;
  assign new_n48545_ = ys__n37815 & new_n48520_;
  assign new_n48546_ = ys__n18669 & ~new_n48524_;
  assign new_n48547_ = ~new_n48545_ & ~new_n48546_;
  assign ys__n32467 = ~new_n48527_ & ~new_n48547_;
  assign new_n48549_ = ys__n37816 & new_n48520_;
  assign new_n48550_ = ys__n18672 & ~new_n48524_;
  assign new_n48551_ = ~new_n48549_ & ~new_n48550_;
  assign ys__n32468 = ~new_n48527_ & ~new_n48551_;
  assign new_n48553_ = ys__n37817 & new_n48520_;
  assign new_n48554_ = ys__n18675 & ~new_n48524_;
  assign new_n48555_ = ~new_n48553_ & ~new_n48554_;
  assign ys__n32469 = ~new_n48527_ & ~new_n48555_;
  assign new_n48557_ = ys__n37818 & new_n48520_;
  assign new_n48558_ = ys__n18678 & ~new_n48524_;
  assign new_n48559_ = ~new_n48557_ & ~new_n48558_;
  assign ys__n32470 = ~new_n48527_ & ~new_n48559_;
  assign new_n48561_ = ys__n37819 & new_n48520_;
  assign new_n48562_ = ys__n18681 & ~new_n48524_;
  assign new_n48563_ = ~new_n48561_ & ~new_n48562_;
  assign ys__n32471 = ~new_n48527_ & ~new_n48563_;
  assign new_n48565_ = ys__n37820 & new_n48520_;
  assign new_n48566_ = ys__n18684 & ~new_n48524_;
  assign new_n48567_ = ~new_n48565_ & ~new_n48566_;
  assign ys__n32472 = ~new_n48527_ & ~new_n48567_;
  assign new_n48569_ = ys__n37821 & new_n48520_;
  assign new_n48570_ = ys__n18687 & ~new_n48524_;
  assign new_n48571_ = ~new_n48569_ & ~new_n48570_;
  assign ys__n32473 = ~new_n48527_ & ~new_n48571_;
  assign new_n48573_ = ys__n37822 & new_n48520_;
  assign new_n48574_ = ys__n18690 & ~new_n48524_;
  assign new_n48575_ = ~new_n48573_ & ~new_n48574_;
  assign ys__n32474 = ~new_n48527_ & ~new_n48575_;
  assign new_n48577_ = ys__n37823 & new_n48520_;
  assign new_n48578_ = ys__n18693 & ~new_n48524_;
  assign new_n48579_ = ~new_n48577_ & ~new_n48578_;
  assign ys__n32475 = ~new_n48527_ & ~new_n48579_;
  assign new_n48581_ = ys__n37824 & new_n48520_;
  assign new_n48582_ = ys__n18696 & ~new_n48524_;
  assign new_n48583_ = ~new_n48581_ & ~new_n48582_;
  assign ys__n32476 = ~new_n48527_ & ~new_n48583_;
  assign new_n48585_ = ys__n37825 & new_n48520_;
  assign new_n48586_ = ys__n18699 & ~new_n48524_;
  assign new_n48587_ = ~new_n48585_ & ~new_n48586_;
  assign ys__n32477 = ~new_n48527_ & ~new_n48587_;
  assign new_n48589_ = ys__n37826 & new_n48520_;
  assign new_n48590_ = ys__n18702 & ~new_n48524_;
  assign new_n48591_ = ~new_n48589_ & ~new_n48590_;
  assign ys__n32478 = ~new_n48527_ & ~new_n48591_;
  assign new_n48593_ = ys__n37827 & new_n48520_;
  assign new_n48594_ = ys__n18705 & ~new_n48524_;
  assign new_n48595_ = ~new_n48593_ & ~new_n48594_;
  assign ys__n32479 = ~new_n48527_ & ~new_n48595_;
  assign new_n48597_ = ys__n37828 & new_n48520_;
  assign new_n48598_ = ys__n18708 & ~new_n48524_;
  assign new_n48599_ = ~new_n48597_ & ~new_n48598_;
  assign ys__n32480 = ~new_n48527_ & ~new_n48599_;
  assign new_n48601_ = ys__n37829 & new_n48520_;
  assign new_n48602_ = ys__n18711 & ~new_n48524_;
  assign new_n48603_ = ~new_n48601_ & ~new_n48602_;
  assign ys__n32481 = ~new_n48527_ & ~new_n48603_;
  assign new_n48605_ = ys__n37830 & new_n48520_;
  assign new_n48606_ = ys__n18714 & ~new_n48524_;
  assign new_n48607_ = ~new_n48605_ & ~new_n48606_;
  assign ys__n32482 = ~new_n48527_ & ~new_n48607_;
  assign new_n48609_ = ys__n37831 & new_n48520_;
  assign new_n48610_ = ys__n18717 & ~new_n48524_;
  assign new_n48611_ = ~new_n48609_ & ~new_n48610_;
  assign ys__n32483 = ~new_n48527_ & ~new_n48611_;
  assign new_n48613_ = ys__n37832 & new_n48520_;
  assign new_n48614_ = ys__n18720 & ~new_n48524_;
  assign new_n48615_ = ~new_n48613_ & ~new_n48614_;
  assign ys__n32484 = ~new_n48527_ & ~new_n48615_;
  assign new_n48617_ = ys__n37833 & new_n48520_;
  assign new_n48618_ = ys__n18723 & ~new_n48524_;
  assign new_n48619_ = ~new_n48617_ & ~new_n48618_;
  assign ys__n32485 = ~new_n48527_ & ~new_n48619_;
  assign new_n48621_ = ys__n37834 & new_n48520_;
  assign new_n48622_ = ys__n18726 & ~new_n48524_;
  assign new_n48623_ = ~new_n48621_ & ~new_n48622_;
  assign ys__n32486 = ~new_n48527_ & ~new_n48623_;
  assign new_n48625_ = ys__n37835 & new_n48520_;
  assign new_n48626_ = ys__n18729 & ~new_n48524_;
  assign new_n48627_ = ~new_n48625_ & ~new_n48626_;
  assign ys__n32487 = ~new_n48527_ & ~new_n48627_;
  assign new_n48629_ = ys__n37836 & new_n48520_;
  assign new_n48630_ = ys__n18732 & ~new_n48524_;
  assign new_n48631_ = ~new_n48629_ & ~new_n48630_;
  assign ys__n32488 = ~new_n48527_ & ~new_n48631_;
  assign new_n48633_ = ys__n37837 & new_n48520_;
  assign new_n48634_ = ys__n18735 & ~new_n48524_;
  assign new_n48635_ = ~new_n48633_ & ~new_n48634_;
  assign ys__n32489 = ~new_n48527_ & ~new_n48635_;
  assign new_n48637_ = ys__n37838 & new_n48520_;
  assign new_n48638_ = ys__n18738 & ~new_n48524_;
  assign new_n48639_ = ~new_n48637_ & ~new_n48638_;
  assign ys__n32490 = ~new_n48527_ & ~new_n48639_;
  assign new_n48641_ = ys__n37839 & new_n48520_;
  assign new_n48642_ = ys__n18741 & ~new_n48524_;
  assign new_n48643_ = ~new_n48641_ & ~new_n48642_;
  assign ys__n32491 = ~new_n48527_ & ~new_n48643_;
  assign new_n48645_ = ys__n37840 & new_n48520_;
  assign new_n48646_ = ys__n18744 & ~new_n48524_;
  assign new_n48647_ = ~new_n48645_ & ~new_n48646_;
  assign ys__n32492 = ~new_n48527_ & ~new_n48647_;
  assign new_n48649_ = ys__n37841 & new_n48520_;
  assign new_n48650_ = ys__n18747 & ~new_n48524_;
  assign new_n48651_ = ~new_n48649_ & ~new_n48650_;
  assign ys__n32493 = ~new_n48527_ & ~new_n48651_;
  assign new_n48653_ = ys__n48106 & new_n45366_;
  assign new_n48654_ = ys__n18654 & ~new_n45370_;
  assign new_n48655_ = ~new_n48653_ & ~new_n48654_;
  assign ys__n32494 = ~new_n45373_ & ~new_n48655_;
  assign new_n48657_ = ys__n48107 & new_n45366_;
  assign new_n48658_ = ys__n18657 & ~new_n45370_;
  assign new_n48659_ = ~new_n48657_ & ~new_n48658_;
  assign ys__n32495 = ~new_n45373_ & ~new_n48659_;
  assign new_n48661_ = ys__n48108 & new_n45366_;
  assign new_n48662_ = ys__n18660 & ~new_n45370_;
  assign new_n48663_ = ~new_n48661_ & ~new_n48662_;
  assign ys__n32496 = ~new_n45373_ & ~new_n48663_;
  assign new_n48665_ = ys__n48109 & new_n45366_;
  assign new_n48666_ = ys__n18663 & ~new_n45370_;
  assign new_n48667_ = ~new_n48665_ & ~new_n48666_;
  assign ys__n32497 = ~new_n45373_ & ~new_n48667_;
  assign new_n48669_ = ys__n37842 & new_n45366_;
  assign new_n48670_ = ys__n18666 & ~new_n45370_;
  assign new_n48671_ = ~new_n48669_ & ~new_n48670_;
  assign ys__n32498 = ~new_n45373_ & ~new_n48671_;
  assign new_n48673_ = ys__n37843 & new_n45366_;
  assign new_n48674_ = ys__n18669 & ~new_n45370_;
  assign new_n48675_ = ~new_n48673_ & ~new_n48674_;
  assign ys__n32499 = ~new_n45373_ & ~new_n48675_;
  assign new_n48677_ = ys__n37844 & new_n45366_;
  assign new_n48678_ = ys__n18672 & ~new_n45370_;
  assign new_n48679_ = ~new_n48677_ & ~new_n48678_;
  assign ys__n32500 = ~new_n45373_ & ~new_n48679_;
  assign new_n48681_ = ys__n37845 & new_n45366_;
  assign new_n48682_ = ys__n18675 & ~new_n45370_;
  assign new_n48683_ = ~new_n48681_ & ~new_n48682_;
  assign ys__n32501 = ~new_n45373_ & ~new_n48683_;
  assign new_n48685_ = ys__n37846 & new_n45366_;
  assign new_n48686_ = ys__n18678 & ~new_n45370_;
  assign new_n48687_ = ~new_n48685_ & ~new_n48686_;
  assign ys__n32502 = ~new_n45373_ & ~new_n48687_;
  assign new_n48689_ = ys__n37847 & new_n45366_;
  assign new_n48690_ = ys__n18681 & ~new_n45370_;
  assign new_n48691_ = ~new_n48689_ & ~new_n48690_;
  assign ys__n32503 = ~new_n45373_ & ~new_n48691_;
  assign new_n48693_ = ys__n37848 & new_n45366_;
  assign new_n48694_ = ys__n18684 & ~new_n45370_;
  assign new_n48695_ = ~new_n48693_ & ~new_n48694_;
  assign ys__n32504 = ~new_n45373_ & ~new_n48695_;
  assign new_n48697_ = ys__n37849 & new_n45366_;
  assign new_n48698_ = ys__n18687 & ~new_n45370_;
  assign new_n48699_ = ~new_n48697_ & ~new_n48698_;
  assign ys__n32505 = ~new_n45373_ & ~new_n48699_;
  assign new_n48701_ = ys__n37850 & new_n45366_;
  assign new_n48702_ = ys__n18690 & ~new_n45370_;
  assign new_n48703_ = ~new_n48701_ & ~new_n48702_;
  assign ys__n32506 = ~new_n45373_ & ~new_n48703_;
  assign new_n48705_ = ys__n37851 & new_n45366_;
  assign new_n48706_ = ys__n18693 & ~new_n45370_;
  assign new_n48707_ = ~new_n48705_ & ~new_n48706_;
  assign ys__n32507 = ~new_n45373_ & ~new_n48707_;
  assign new_n48709_ = ys__n37852 & new_n45366_;
  assign new_n48710_ = ys__n18696 & ~new_n45370_;
  assign new_n48711_ = ~new_n48709_ & ~new_n48710_;
  assign ys__n32508 = ~new_n45373_ & ~new_n48711_;
  assign new_n48713_ = ys__n37853 & new_n45366_;
  assign new_n48714_ = ys__n18699 & ~new_n45370_;
  assign new_n48715_ = ~new_n48713_ & ~new_n48714_;
  assign ys__n32509 = ~new_n45373_ & ~new_n48715_;
  assign new_n48717_ = ys__n37854 & new_n45366_;
  assign new_n48718_ = ys__n18702 & ~new_n45370_;
  assign new_n48719_ = ~new_n48717_ & ~new_n48718_;
  assign ys__n32510 = ~new_n45373_ & ~new_n48719_;
  assign new_n48721_ = ys__n37855 & new_n45366_;
  assign new_n48722_ = ys__n18705 & ~new_n45370_;
  assign new_n48723_ = ~new_n48721_ & ~new_n48722_;
  assign ys__n32511 = ~new_n45373_ & ~new_n48723_;
  assign new_n48725_ = ys__n37856 & new_n45366_;
  assign new_n48726_ = ys__n18708 & ~new_n45370_;
  assign new_n48727_ = ~new_n48725_ & ~new_n48726_;
  assign ys__n32512 = ~new_n45373_ & ~new_n48727_;
  assign new_n48729_ = ys__n37857 & new_n45366_;
  assign new_n48730_ = ys__n18711 & ~new_n45370_;
  assign new_n48731_ = ~new_n48729_ & ~new_n48730_;
  assign ys__n32513 = ~new_n45373_ & ~new_n48731_;
  assign new_n48733_ = ys__n37858 & new_n45366_;
  assign new_n48734_ = ys__n18714 & ~new_n45370_;
  assign new_n48735_ = ~new_n48733_ & ~new_n48734_;
  assign ys__n32514 = ~new_n45373_ & ~new_n48735_;
  assign new_n48737_ = ys__n37859 & new_n45366_;
  assign new_n48738_ = ys__n18717 & ~new_n45370_;
  assign new_n48739_ = ~new_n48737_ & ~new_n48738_;
  assign ys__n32515 = ~new_n45373_ & ~new_n48739_;
  assign new_n48741_ = ys__n37860 & new_n45366_;
  assign new_n48742_ = ys__n18720 & ~new_n45370_;
  assign new_n48743_ = ~new_n48741_ & ~new_n48742_;
  assign ys__n32516 = ~new_n45373_ & ~new_n48743_;
  assign new_n48745_ = ys__n37861 & new_n45366_;
  assign new_n48746_ = ys__n18723 & ~new_n45370_;
  assign new_n48747_ = ~new_n48745_ & ~new_n48746_;
  assign ys__n32517 = ~new_n45373_ & ~new_n48747_;
  assign new_n48749_ = ys__n37862 & new_n45366_;
  assign new_n48750_ = ys__n18726 & ~new_n45370_;
  assign new_n48751_ = ~new_n48749_ & ~new_n48750_;
  assign ys__n32518 = ~new_n45373_ & ~new_n48751_;
  assign new_n48753_ = ys__n37863 & new_n45366_;
  assign new_n48754_ = ys__n18729 & ~new_n45370_;
  assign new_n48755_ = ~new_n48753_ & ~new_n48754_;
  assign ys__n32519 = ~new_n45373_ & ~new_n48755_;
  assign new_n48757_ = ys__n37864 & new_n45366_;
  assign new_n48758_ = ys__n18732 & ~new_n45370_;
  assign new_n48759_ = ~new_n48757_ & ~new_n48758_;
  assign ys__n32520 = ~new_n45373_ & ~new_n48759_;
  assign new_n48761_ = ys__n37865 & new_n45366_;
  assign new_n48762_ = ys__n18735 & ~new_n45370_;
  assign new_n48763_ = ~new_n48761_ & ~new_n48762_;
  assign ys__n32521 = ~new_n45373_ & ~new_n48763_;
  assign new_n48765_ = ys__n37866 & new_n45366_;
  assign new_n48766_ = ys__n18738 & ~new_n45370_;
  assign new_n48767_ = ~new_n48765_ & ~new_n48766_;
  assign ys__n32522 = ~new_n45373_ & ~new_n48767_;
  assign new_n48769_ = ys__n37867 & new_n45366_;
  assign new_n48770_ = ys__n18741 & ~new_n45370_;
  assign new_n48771_ = ~new_n48769_ & ~new_n48770_;
  assign ys__n32523 = ~new_n45373_ & ~new_n48771_;
  assign new_n48773_ = ys__n37868 & new_n45366_;
  assign new_n48774_ = ys__n18744 & ~new_n45370_;
  assign new_n48775_ = ~new_n48773_ & ~new_n48774_;
  assign ys__n32524 = ~new_n45373_ & ~new_n48775_;
  assign new_n48777_ = ys__n37869 & new_n45366_;
  assign new_n48778_ = ys__n18747 & ~new_n45370_;
  assign new_n48779_ = ~new_n48777_ & ~new_n48778_;
  assign ys__n32525 = ~new_n45373_ & ~new_n48779_;
  assign new_n48781_ = ys__n48110 & new_n45221_;
  assign new_n48782_ = ys__n18654 & ~new_n45225_;
  assign new_n48783_ = ~new_n48781_ & ~new_n48782_;
  assign ys__n32526 = ~new_n45228_ & ~new_n48783_;
  assign new_n48785_ = ys__n48111 & new_n45221_;
  assign new_n48786_ = ys__n18657 & ~new_n45225_;
  assign new_n48787_ = ~new_n48785_ & ~new_n48786_;
  assign ys__n32527 = ~new_n45228_ & ~new_n48787_;
  assign new_n48789_ = ys__n48112 & new_n45221_;
  assign new_n48790_ = ys__n18660 & ~new_n45225_;
  assign new_n48791_ = ~new_n48789_ & ~new_n48790_;
  assign ys__n32528 = ~new_n45228_ & ~new_n48791_;
  assign new_n48793_ = ys__n48113 & new_n45221_;
  assign new_n48794_ = ys__n18663 & ~new_n45225_;
  assign new_n48795_ = ~new_n48793_ & ~new_n48794_;
  assign ys__n32529 = ~new_n45228_ & ~new_n48795_;
  assign new_n48797_ = ys__n37870 & new_n45221_;
  assign new_n48798_ = ys__n18666 & ~new_n45225_;
  assign new_n48799_ = ~new_n48797_ & ~new_n48798_;
  assign ys__n32530 = ~new_n45228_ & ~new_n48799_;
  assign new_n48801_ = ys__n37871 & new_n45221_;
  assign new_n48802_ = ys__n18669 & ~new_n45225_;
  assign new_n48803_ = ~new_n48801_ & ~new_n48802_;
  assign ys__n32531 = ~new_n45228_ & ~new_n48803_;
  assign new_n48805_ = ys__n37872 & new_n45221_;
  assign new_n48806_ = ys__n18672 & ~new_n45225_;
  assign new_n48807_ = ~new_n48805_ & ~new_n48806_;
  assign ys__n32532 = ~new_n45228_ & ~new_n48807_;
  assign new_n48809_ = ys__n37873 & new_n45221_;
  assign new_n48810_ = ys__n18675 & ~new_n45225_;
  assign new_n48811_ = ~new_n48809_ & ~new_n48810_;
  assign ys__n32533 = ~new_n45228_ & ~new_n48811_;
  assign new_n48813_ = ys__n37874 & new_n45221_;
  assign new_n48814_ = ys__n18678 & ~new_n45225_;
  assign new_n48815_ = ~new_n48813_ & ~new_n48814_;
  assign ys__n32534 = ~new_n45228_ & ~new_n48815_;
  assign new_n48817_ = ys__n37875 & new_n45221_;
  assign new_n48818_ = ys__n18681 & ~new_n45225_;
  assign new_n48819_ = ~new_n48817_ & ~new_n48818_;
  assign ys__n32535 = ~new_n45228_ & ~new_n48819_;
  assign new_n48821_ = ys__n37876 & new_n45221_;
  assign new_n48822_ = ys__n18684 & ~new_n45225_;
  assign new_n48823_ = ~new_n48821_ & ~new_n48822_;
  assign ys__n32536 = ~new_n45228_ & ~new_n48823_;
  assign new_n48825_ = ys__n37877 & new_n45221_;
  assign new_n48826_ = ys__n18687 & ~new_n45225_;
  assign new_n48827_ = ~new_n48825_ & ~new_n48826_;
  assign ys__n32537 = ~new_n45228_ & ~new_n48827_;
  assign new_n48829_ = ys__n37878 & new_n45221_;
  assign new_n48830_ = ys__n18690 & ~new_n45225_;
  assign new_n48831_ = ~new_n48829_ & ~new_n48830_;
  assign ys__n32538 = ~new_n45228_ & ~new_n48831_;
  assign new_n48833_ = ys__n37879 & new_n45221_;
  assign new_n48834_ = ys__n18693 & ~new_n45225_;
  assign new_n48835_ = ~new_n48833_ & ~new_n48834_;
  assign ys__n32539 = ~new_n45228_ & ~new_n48835_;
  assign new_n48837_ = ys__n37880 & new_n45221_;
  assign new_n48838_ = ys__n18696 & ~new_n45225_;
  assign new_n48839_ = ~new_n48837_ & ~new_n48838_;
  assign ys__n32540 = ~new_n45228_ & ~new_n48839_;
  assign new_n48841_ = ys__n37881 & new_n45221_;
  assign new_n48842_ = ys__n18699 & ~new_n45225_;
  assign new_n48843_ = ~new_n48841_ & ~new_n48842_;
  assign ys__n32541 = ~new_n45228_ & ~new_n48843_;
  assign new_n48845_ = ys__n37882 & new_n45221_;
  assign new_n48846_ = ys__n18702 & ~new_n45225_;
  assign new_n48847_ = ~new_n48845_ & ~new_n48846_;
  assign ys__n32542 = ~new_n45228_ & ~new_n48847_;
  assign new_n48849_ = ys__n37883 & new_n45221_;
  assign new_n48850_ = ys__n18705 & ~new_n45225_;
  assign new_n48851_ = ~new_n48849_ & ~new_n48850_;
  assign ys__n32543 = ~new_n45228_ & ~new_n48851_;
  assign new_n48853_ = ys__n37884 & new_n45221_;
  assign new_n48854_ = ys__n18708 & ~new_n45225_;
  assign new_n48855_ = ~new_n48853_ & ~new_n48854_;
  assign ys__n32544 = ~new_n45228_ & ~new_n48855_;
  assign new_n48857_ = ys__n37885 & new_n45221_;
  assign new_n48858_ = ys__n18711 & ~new_n45225_;
  assign new_n48859_ = ~new_n48857_ & ~new_n48858_;
  assign ys__n32545 = ~new_n45228_ & ~new_n48859_;
  assign new_n48861_ = ys__n37886 & new_n45221_;
  assign new_n48862_ = ys__n18714 & ~new_n45225_;
  assign new_n48863_ = ~new_n48861_ & ~new_n48862_;
  assign ys__n32546 = ~new_n45228_ & ~new_n48863_;
  assign new_n48865_ = ys__n37887 & new_n45221_;
  assign new_n48866_ = ys__n18717 & ~new_n45225_;
  assign new_n48867_ = ~new_n48865_ & ~new_n48866_;
  assign ys__n32547 = ~new_n45228_ & ~new_n48867_;
  assign new_n48869_ = ys__n37888 & new_n45221_;
  assign new_n48870_ = ys__n18720 & ~new_n45225_;
  assign new_n48871_ = ~new_n48869_ & ~new_n48870_;
  assign ys__n32548 = ~new_n45228_ & ~new_n48871_;
  assign new_n48873_ = ys__n37889 & new_n45221_;
  assign new_n48874_ = ys__n18723 & ~new_n45225_;
  assign new_n48875_ = ~new_n48873_ & ~new_n48874_;
  assign ys__n32549 = ~new_n45228_ & ~new_n48875_;
  assign new_n48877_ = ys__n37890 & new_n45221_;
  assign new_n48878_ = ys__n18726 & ~new_n45225_;
  assign new_n48879_ = ~new_n48877_ & ~new_n48878_;
  assign ys__n32550 = ~new_n45228_ & ~new_n48879_;
  assign new_n48881_ = ys__n37891 & new_n45221_;
  assign new_n48882_ = ys__n18729 & ~new_n45225_;
  assign new_n48883_ = ~new_n48881_ & ~new_n48882_;
  assign ys__n32551 = ~new_n45228_ & ~new_n48883_;
  assign new_n48885_ = ys__n37892 & new_n45221_;
  assign new_n48886_ = ys__n18732 & ~new_n45225_;
  assign new_n48887_ = ~new_n48885_ & ~new_n48886_;
  assign ys__n32552 = ~new_n45228_ & ~new_n48887_;
  assign new_n48889_ = ys__n37893 & new_n45221_;
  assign new_n48890_ = ys__n18735 & ~new_n45225_;
  assign new_n48891_ = ~new_n48889_ & ~new_n48890_;
  assign ys__n32553 = ~new_n45228_ & ~new_n48891_;
  assign new_n48893_ = ys__n37894 & new_n45221_;
  assign new_n48894_ = ys__n18738 & ~new_n45225_;
  assign new_n48895_ = ~new_n48893_ & ~new_n48894_;
  assign ys__n32554 = ~new_n45228_ & ~new_n48895_;
  assign new_n48897_ = ys__n37895 & new_n45221_;
  assign new_n48898_ = ys__n18741 & ~new_n45225_;
  assign new_n48899_ = ~new_n48897_ & ~new_n48898_;
  assign ys__n32555 = ~new_n45228_ & ~new_n48899_;
  assign new_n48901_ = ys__n37896 & new_n45221_;
  assign new_n48902_ = ys__n18744 & ~new_n45225_;
  assign new_n48903_ = ~new_n48901_ & ~new_n48902_;
  assign ys__n32556 = ~new_n45228_ & ~new_n48903_;
  assign new_n48905_ = ys__n37897 & new_n45221_;
  assign new_n48906_ = ys__n18747 & ~new_n45225_;
  assign new_n48907_ = ~new_n48905_ & ~new_n48906_;
  assign ys__n32557 = ~new_n45228_ & ~new_n48907_;
  assign new_n48909_ = ys__n48114 & new_n45076_;
  assign new_n48910_ = ys__n18654 & ~new_n45080_;
  assign new_n48911_ = ~new_n48909_ & ~new_n48910_;
  assign ys__n32558 = ~new_n45083_ & ~new_n48911_;
  assign new_n48913_ = ys__n48115 & new_n45076_;
  assign new_n48914_ = ys__n18657 & ~new_n45080_;
  assign new_n48915_ = ~new_n48913_ & ~new_n48914_;
  assign ys__n32559 = ~new_n45083_ & ~new_n48915_;
  assign new_n48917_ = ys__n48116 & new_n45076_;
  assign new_n48918_ = ys__n18660 & ~new_n45080_;
  assign new_n48919_ = ~new_n48917_ & ~new_n48918_;
  assign ys__n32560 = ~new_n45083_ & ~new_n48919_;
  assign new_n48921_ = ys__n48117 & new_n45076_;
  assign new_n48922_ = ys__n18663 & ~new_n45080_;
  assign new_n48923_ = ~new_n48921_ & ~new_n48922_;
  assign ys__n32561 = ~new_n45083_ & ~new_n48923_;
  assign new_n48925_ = ys__n37898 & new_n45076_;
  assign new_n48926_ = ys__n18666 & ~new_n45080_;
  assign new_n48927_ = ~new_n48925_ & ~new_n48926_;
  assign ys__n32562 = ~new_n45083_ & ~new_n48927_;
  assign new_n48929_ = ys__n37899 & new_n45076_;
  assign new_n48930_ = ys__n18669 & ~new_n45080_;
  assign new_n48931_ = ~new_n48929_ & ~new_n48930_;
  assign ys__n32563 = ~new_n45083_ & ~new_n48931_;
  assign new_n48933_ = ys__n37900 & new_n45076_;
  assign new_n48934_ = ys__n18672 & ~new_n45080_;
  assign new_n48935_ = ~new_n48933_ & ~new_n48934_;
  assign ys__n32564 = ~new_n45083_ & ~new_n48935_;
  assign new_n48937_ = ys__n37901 & new_n45076_;
  assign new_n48938_ = ys__n18675 & ~new_n45080_;
  assign new_n48939_ = ~new_n48937_ & ~new_n48938_;
  assign ys__n32565 = ~new_n45083_ & ~new_n48939_;
  assign new_n48941_ = ys__n37902 & new_n45076_;
  assign new_n48942_ = ys__n18678 & ~new_n45080_;
  assign new_n48943_ = ~new_n48941_ & ~new_n48942_;
  assign ys__n32566 = ~new_n45083_ & ~new_n48943_;
  assign new_n48945_ = ys__n37903 & new_n45076_;
  assign new_n48946_ = ys__n18681 & ~new_n45080_;
  assign new_n48947_ = ~new_n48945_ & ~new_n48946_;
  assign ys__n32567 = ~new_n45083_ & ~new_n48947_;
  assign new_n48949_ = ys__n37904 & new_n45076_;
  assign new_n48950_ = ys__n18684 & ~new_n45080_;
  assign new_n48951_ = ~new_n48949_ & ~new_n48950_;
  assign ys__n32568 = ~new_n45083_ & ~new_n48951_;
  assign new_n48953_ = ys__n37905 & new_n45076_;
  assign new_n48954_ = ys__n18687 & ~new_n45080_;
  assign new_n48955_ = ~new_n48953_ & ~new_n48954_;
  assign ys__n32569 = ~new_n45083_ & ~new_n48955_;
  assign new_n48957_ = ys__n37906 & new_n45076_;
  assign new_n48958_ = ys__n18690 & ~new_n45080_;
  assign new_n48959_ = ~new_n48957_ & ~new_n48958_;
  assign ys__n32570 = ~new_n45083_ & ~new_n48959_;
  assign new_n48961_ = ys__n37907 & new_n45076_;
  assign new_n48962_ = ys__n18693 & ~new_n45080_;
  assign new_n48963_ = ~new_n48961_ & ~new_n48962_;
  assign ys__n32571 = ~new_n45083_ & ~new_n48963_;
  assign new_n48965_ = ys__n37908 & new_n45076_;
  assign new_n48966_ = ys__n18696 & ~new_n45080_;
  assign new_n48967_ = ~new_n48965_ & ~new_n48966_;
  assign ys__n32572 = ~new_n45083_ & ~new_n48967_;
  assign new_n48969_ = ys__n37909 & new_n45076_;
  assign new_n48970_ = ys__n18699 & ~new_n45080_;
  assign new_n48971_ = ~new_n48969_ & ~new_n48970_;
  assign ys__n32573 = ~new_n45083_ & ~new_n48971_;
  assign new_n48973_ = ys__n37910 & new_n45076_;
  assign new_n48974_ = ys__n18702 & ~new_n45080_;
  assign new_n48975_ = ~new_n48973_ & ~new_n48974_;
  assign ys__n32574 = ~new_n45083_ & ~new_n48975_;
  assign new_n48977_ = ys__n37911 & new_n45076_;
  assign new_n48978_ = ys__n18705 & ~new_n45080_;
  assign new_n48979_ = ~new_n48977_ & ~new_n48978_;
  assign ys__n32575 = ~new_n45083_ & ~new_n48979_;
  assign new_n48981_ = ys__n37912 & new_n45076_;
  assign new_n48982_ = ys__n18708 & ~new_n45080_;
  assign new_n48983_ = ~new_n48981_ & ~new_n48982_;
  assign ys__n32576 = ~new_n45083_ & ~new_n48983_;
  assign new_n48985_ = ys__n37913 & new_n45076_;
  assign new_n48986_ = ys__n18711 & ~new_n45080_;
  assign new_n48987_ = ~new_n48985_ & ~new_n48986_;
  assign ys__n32577 = ~new_n45083_ & ~new_n48987_;
  assign new_n48989_ = ys__n37914 & new_n45076_;
  assign new_n48990_ = ys__n18714 & ~new_n45080_;
  assign new_n48991_ = ~new_n48989_ & ~new_n48990_;
  assign ys__n32578 = ~new_n45083_ & ~new_n48991_;
  assign new_n48993_ = ys__n37915 & new_n45076_;
  assign new_n48994_ = ys__n18717 & ~new_n45080_;
  assign new_n48995_ = ~new_n48993_ & ~new_n48994_;
  assign ys__n32579 = ~new_n45083_ & ~new_n48995_;
  assign new_n48997_ = ys__n37916 & new_n45076_;
  assign new_n48998_ = ys__n18720 & ~new_n45080_;
  assign new_n48999_ = ~new_n48997_ & ~new_n48998_;
  assign ys__n32580 = ~new_n45083_ & ~new_n48999_;
  assign new_n49001_ = ys__n37917 & new_n45076_;
  assign new_n49002_ = ys__n18723 & ~new_n45080_;
  assign new_n49003_ = ~new_n49001_ & ~new_n49002_;
  assign ys__n32581 = ~new_n45083_ & ~new_n49003_;
  assign new_n49005_ = ys__n37918 & new_n45076_;
  assign new_n49006_ = ys__n18726 & ~new_n45080_;
  assign new_n49007_ = ~new_n49005_ & ~new_n49006_;
  assign ys__n32582 = ~new_n45083_ & ~new_n49007_;
  assign new_n49009_ = ys__n37919 & new_n45076_;
  assign new_n49010_ = ys__n18729 & ~new_n45080_;
  assign new_n49011_ = ~new_n49009_ & ~new_n49010_;
  assign ys__n32583 = ~new_n45083_ & ~new_n49011_;
  assign new_n49013_ = ys__n37920 & new_n45076_;
  assign new_n49014_ = ys__n18732 & ~new_n45080_;
  assign new_n49015_ = ~new_n49013_ & ~new_n49014_;
  assign ys__n32584 = ~new_n45083_ & ~new_n49015_;
  assign new_n49017_ = ys__n37921 & new_n45076_;
  assign new_n49018_ = ys__n18735 & ~new_n45080_;
  assign new_n49019_ = ~new_n49017_ & ~new_n49018_;
  assign ys__n32585 = ~new_n45083_ & ~new_n49019_;
  assign new_n49021_ = ys__n37922 & new_n45076_;
  assign new_n49022_ = ys__n18738 & ~new_n45080_;
  assign new_n49023_ = ~new_n49021_ & ~new_n49022_;
  assign ys__n32586 = ~new_n45083_ & ~new_n49023_;
  assign new_n49025_ = ys__n37923 & new_n45076_;
  assign new_n49026_ = ys__n18741 & ~new_n45080_;
  assign new_n49027_ = ~new_n49025_ & ~new_n49026_;
  assign ys__n32587 = ~new_n45083_ & ~new_n49027_;
  assign new_n49029_ = ys__n37924 & new_n45076_;
  assign new_n49030_ = ys__n18744 & ~new_n45080_;
  assign new_n49031_ = ~new_n49029_ & ~new_n49030_;
  assign ys__n32588 = ~new_n45083_ & ~new_n49031_;
  assign new_n49033_ = ys__n37925 & new_n45076_;
  assign new_n49034_ = ys__n18747 & ~new_n45080_;
  assign new_n49035_ = ~new_n49033_ & ~new_n49034_;
  assign ys__n32589 = ~new_n45083_ & ~new_n49035_;
  assign new_n49037_ = ys__n48118 & new_n44931_;
  assign new_n49038_ = ys__n18654 & ~new_n44935_;
  assign new_n49039_ = ~new_n49037_ & ~new_n49038_;
  assign ys__n32590 = ~new_n44938_ & ~new_n49039_;
  assign new_n49041_ = ys__n48119 & new_n44931_;
  assign new_n49042_ = ys__n18657 & ~new_n44935_;
  assign new_n49043_ = ~new_n49041_ & ~new_n49042_;
  assign ys__n32591 = ~new_n44938_ & ~new_n49043_;
  assign new_n49045_ = ys__n48120 & new_n44931_;
  assign new_n49046_ = ys__n18660 & ~new_n44935_;
  assign new_n49047_ = ~new_n49045_ & ~new_n49046_;
  assign ys__n32592 = ~new_n44938_ & ~new_n49047_;
  assign new_n49049_ = ys__n48121 & new_n44931_;
  assign new_n49050_ = ys__n18663 & ~new_n44935_;
  assign new_n49051_ = ~new_n49049_ & ~new_n49050_;
  assign ys__n32593 = ~new_n44938_ & ~new_n49051_;
  assign new_n49053_ = ys__n37926 & new_n44931_;
  assign new_n49054_ = ys__n18666 & ~new_n44935_;
  assign new_n49055_ = ~new_n49053_ & ~new_n49054_;
  assign ys__n32594 = ~new_n44938_ & ~new_n49055_;
  assign new_n49057_ = ys__n37927 & new_n44931_;
  assign new_n49058_ = ys__n18669 & ~new_n44935_;
  assign new_n49059_ = ~new_n49057_ & ~new_n49058_;
  assign ys__n32595 = ~new_n44938_ & ~new_n49059_;
  assign new_n49061_ = ys__n37928 & new_n44931_;
  assign new_n49062_ = ys__n18672 & ~new_n44935_;
  assign new_n49063_ = ~new_n49061_ & ~new_n49062_;
  assign ys__n32596 = ~new_n44938_ & ~new_n49063_;
  assign new_n49065_ = ys__n37929 & new_n44931_;
  assign new_n49066_ = ys__n18675 & ~new_n44935_;
  assign new_n49067_ = ~new_n49065_ & ~new_n49066_;
  assign ys__n32597 = ~new_n44938_ & ~new_n49067_;
  assign new_n49069_ = ys__n37930 & new_n44931_;
  assign new_n49070_ = ys__n18678 & ~new_n44935_;
  assign new_n49071_ = ~new_n49069_ & ~new_n49070_;
  assign ys__n32598 = ~new_n44938_ & ~new_n49071_;
  assign new_n49073_ = ys__n37931 & new_n44931_;
  assign new_n49074_ = ys__n18681 & ~new_n44935_;
  assign new_n49075_ = ~new_n49073_ & ~new_n49074_;
  assign ys__n32599 = ~new_n44938_ & ~new_n49075_;
  assign new_n49077_ = ys__n37932 & new_n44931_;
  assign new_n49078_ = ys__n18684 & ~new_n44935_;
  assign new_n49079_ = ~new_n49077_ & ~new_n49078_;
  assign ys__n32600 = ~new_n44938_ & ~new_n49079_;
  assign new_n49081_ = ys__n37933 & new_n44931_;
  assign new_n49082_ = ys__n18687 & ~new_n44935_;
  assign new_n49083_ = ~new_n49081_ & ~new_n49082_;
  assign ys__n32601 = ~new_n44938_ & ~new_n49083_;
  assign new_n49085_ = ys__n37934 & new_n44931_;
  assign new_n49086_ = ys__n18690 & ~new_n44935_;
  assign new_n49087_ = ~new_n49085_ & ~new_n49086_;
  assign ys__n32602 = ~new_n44938_ & ~new_n49087_;
  assign new_n49089_ = ys__n37935 & new_n44931_;
  assign new_n49090_ = ys__n18693 & ~new_n44935_;
  assign new_n49091_ = ~new_n49089_ & ~new_n49090_;
  assign ys__n32603 = ~new_n44938_ & ~new_n49091_;
  assign new_n49093_ = ys__n37936 & new_n44931_;
  assign new_n49094_ = ys__n18696 & ~new_n44935_;
  assign new_n49095_ = ~new_n49093_ & ~new_n49094_;
  assign ys__n32604 = ~new_n44938_ & ~new_n49095_;
  assign new_n49097_ = ys__n37937 & new_n44931_;
  assign new_n49098_ = ys__n18699 & ~new_n44935_;
  assign new_n49099_ = ~new_n49097_ & ~new_n49098_;
  assign ys__n32605 = ~new_n44938_ & ~new_n49099_;
  assign new_n49101_ = ys__n37938 & new_n44931_;
  assign new_n49102_ = ys__n18702 & ~new_n44935_;
  assign new_n49103_ = ~new_n49101_ & ~new_n49102_;
  assign ys__n32606 = ~new_n44938_ & ~new_n49103_;
  assign new_n49105_ = ys__n37939 & new_n44931_;
  assign new_n49106_ = ys__n18705 & ~new_n44935_;
  assign new_n49107_ = ~new_n49105_ & ~new_n49106_;
  assign ys__n32607 = ~new_n44938_ & ~new_n49107_;
  assign new_n49109_ = ys__n37940 & new_n44931_;
  assign new_n49110_ = ys__n18708 & ~new_n44935_;
  assign new_n49111_ = ~new_n49109_ & ~new_n49110_;
  assign ys__n32608 = ~new_n44938_ & ~new_n49111_;
  assign new_n49113_ = ys__n37941 & new_n44931_;
  assign new_n49114_ = ys__n18711 & ~new_n44935_;
  assign new_n49115_ = ~new_n49113_ & ~new_n49114_;
  assign ys__n32609 = ~new_n44938_ & ~new_n49115_;
  assign new_n49117_ = ys__n37942 & new_n44931_;
  assign new_n49118_ = ys__n18714 & ~new_n44935_;
  assign new_n49119_ = ~new_n49117_ & ~new_n49118_;
  assign ys__n32610 = ~new_n44938_ & ~new_n49119_;
  assign new_n49121_ = ys__n37943 & new_n44931_;
  assign new_n49122_ = ys__n18717 & ~new_n44935_;
  assign new_n49123_ = ~new_n49121_ & ~new_n49122_;
  assign ys__n32611 = ~new_n44938_ & ~new_n49123_;
  assign new_n49125_ = ys__n37944 & new_n44931_;
  assign new_n49126_ = ys__n18720 & ~new_n44935_;
  assign new_n49127_ = ~new_n49125_ & ~new_n49126_;
  assign ys__n32612 = ~new_n44938_ & ~new_n49127_;
  assign new_n49129_ = ys__n37945 & new_n44931_;
  assign new_n49130_ = ys__n18723 & ~new_n44935_;
  assign new_n49131_ = ~new_n49129_ & ~new_n49130_;
  assign ys__n32613 = ~new_n44938_ & ~new_n49131_;
  assign new_n49133_ = ys__n37946 & new_n44931_;
  assign new_n49134_ = ys__n18726 & ~new_n44935_;
  assign new_n49135_ = ~new_n49133_ & ~new_n49134_;
  assign ys__n32614 = ~new_n44938_ & ~new_n49135_;
  assign new_n49137_ = ys__n37947 & new_n44931_;
  assign new_n49138_ = ys__n18729 & ~new_n44935_;
  assign new_n49139_ = ~new_n49137_ & ~new_n49138_;
  assign ys__n32615 = ~new_n44938_ & ~new_n49139_;
  assign new_n49141_ = ys__n37948 & new_n44931_;
  assign new_n49142_ = ys__n18732 & ~new_n44935_;
  assign new_n49143_ = ~new_n49141_ & ~new_n49142_;
  assign ys__n32616 = ~new_n44938_ & ~new_n49143_;
  assign new_n49145_ = ys__n37949 & new_n44931_;
  assign new_n49146_ = ys__n18735 & ~new_n44935_;
  assign new_n49147_ = ~new_n49145_ & ~new_n49146_;
  assign ys__n32617 = ~new_n44938_ & ~new_n49147_;
  assign new_n49149_ = ys__n37950 & new_n44931_;
  assign new_n49150_ = ys__n18738 & ~new_n44935_;
  assign new_n49151_ = ~new_n49149_ & ~new_n49150_;
  assign ys__n32618 = ~new_n44938_ & ~new_n49151_;
  assign new_n49153_ = ys__n37951 & new_n44931_;
  assign new_n49154_ = ys__n18741 & ~new_n44935_;
  assign new_n49155_ = ~new_n49153_ & ~new_n49154_;
  assign ys__n32619 = ~new_n44938_ & ~new_n49155_;
  assign new_n49157_ = ys__n37952 & new_n44931_;
  assign new_n49158_ = ys__n18744 & ~new_n44935_;
  assign new_n49159_ = ~new_n49157_ & ~new_n49158_;
  assign ys__n32620 = ~new_n44938_ & ~new_n49159_;
  assign new_n49161_ = ys__n37953 & new_n44931_;
  assign new_n49162_ = ys__n18747 & ~new_n44935_;
  assign new_n49163_ = ~new_n49161_ & ~new_n49162_;
  assign ys__n32621 = ~new_n44938_ & ~new_n49163_;
  assign new_n49165_ = ys__n48122 & new_n44786_;
  assign new_n49166_ = ys__n18654 & ~new_n44790_;
  assign new_n49167_ = ~new_n49165_ & ~new_n49166_;
  assign ys__n32622 = ~new_n44793_ & ~new_n49167_;
  assign new_n49169_ = ys__n48123 & new_n44786_;
  assign new_n49170_ = ys__n18657 & ~new_n44790_;
  assign new_n49171_ = ~new_n49169_ & ~new_n49170_;
  assign ys__n32623 = ~new_n44793_ & ~new_n49171_;
  assign new_n49173_ = ys__n48124 & new_n44786_;
  assign new_n49174_ = ys__n18660 & ~new_n44790_;
  assign new_n49175_ = ~new_n49173_ & ~new_n49174_;
  assign ys__n32624 = ~new_n44793_ & ~new_n49175_;
  assign new_n49177_ = ys__n48125 & new_n44786_;
  assign new_n49178_ = ys__n18663 & ~new_n44790_;
  assign new_n49179_ = ~new_n49177_ & ~new_n49178_;
  assign ys__n32625 = ~new_n44793_ & ~new_n49179_;
  assign new_n49181_ = ys__n37954 & new_n44786_;
  assign new_n49182_ = ys__n18666 & ~new_n44790_;
  assign new_n49183_ = ~new_n49181_ & ~new_n49182_;
  assign ys__n32626 = ~new_n44793_ & ~new_n49183_;
  assign new_n49185_ = ys__n37955 & new_n44786_;
  assign new_n49186_ = ys__n18669 & ~new_n44790_;
  assign new_n49187_ = ~new_n49185_ & ~new_n49186_;
  assign ys__n32627 = ~new_n44793_ & ~new_n49187_;
  assign new_n49189_ = ys__n37956 & new_n44786_;
  assign new_n49190_ = ys__n18672 & ~new_n44790_;
  assign new_n49191_ = ~new_n49189_ & ~new_n49190_;
  assign ys__n32628 = ~new_n44793_ & ~new_n49191_;
  assign new_n49193_ = ys__n37957 & new_n44786_;
  assign new_n49194_ = ys__n18675 & ~new_n44790_;
  assign new_n49195_ = ~new_n49193_ & ~new_n49194_;
  assign ys__n32629 = ~new_n44793_ & ~new_n49195_;
  assign new_n49197_ = ys__n37958 & new_n44786_;
  assign new_n49198_ = ys__n18678 & ~new_n44790_;
  assign new_n49199_ = ~new_n49197_ & ~new_n49198_;
  assign ys__n32630 = ~new_n44793_ & ~new_n49199_;
  assign new_n49201_ = ys__n37959 & new_n44786_;
  assign new_n49202_ = ys__n18681 & ~new_n44790_;
  assign new_n49203_ = ~new_n49201_ & ~new_n49202_;
  assign ys__n32631 = ~new_n44793_ & ~new_n49203_;
  assign new_n49205_ = ys__n37960 & new_n44786_;
  assign new_n49206_ = ys__n18684 & ~new_n44790_;
  assign new_n49207_ = ~new_n49205_ & ~new_n49206_;
  assign ys__n32632 = ~new_n44793_ & ~new_n49207_;
  assign new_n49209_ = ys__n37961 & new_n44786_;
  assign new_n49210_ = ys__n18687 & ~new_n44790_;
  assign new_n49211_ = ~new_n49209_ & ~new_n49210_;
  assign ys__n32633 = ~new_n44793_ & ~new_n49211_;
  assign new_n49213_ = ys__n37962 & new_n44786_;
  assign new_n49214_ = ys__n18690 & ~new_n44790_;
  assign new_n49215_ = ~new_n49213_ & ~new_n49214_;
  assign ys__n32634 = ~new_n44793_ & ~new_n49215_;
  assign new_n49217_ = ys__n37963 & new_n44786_;
  assign new_n49218_ = ys__n18693 & ~new_n44790_;
  assign new_n49219_ = ~new_n49217_ & ~new_n49218_;
  assign ys__n32635 = ~new_n44793_ & ~new_n49219_;
  assign new_n49221_ = ys__n37964 & new_n44786_;
  assign new_n49222_ = ys__n18696 & ~new_n44790_;
  assign new_n49223_ = ~new_n49221_ & ~new_n49222_;
  assign ys__n32636 = ~new_n44793_ & ~new_n49223_;
  assign new_n49225_ = ys__n37965 & new_n44786_;
  assign new_n49226_ = ys__n18699 & ~new_n44790_;
  assign new_n49227_ = ~new_n49225_ & ~new_n49226_;
  assign ys__n32637 = ~new_n44793_ & ~new_n49227_;
  assign new_n49229_ = ys__n37966 & new_n44786_;
  assign new_n49230_ = ys__n18702 & ~new_n44790_;
  assign new_n49231_ = ~new_n49229_ & ~new_n49230_;
  assign ys__n32638 = ~new_n44793_ & ~new_n49231_;
  assign new_n49233_ = ys__n37967 & new_n44786_;
  assign new_n49234_ = ys__n18705 & ~new_n44790_;
  assign new_n49235_ = ~new_n49233_ & ~new_n49234_;
  assign ys__n32639 = ~new_n44793_ & ~new_n49235_;
  assign new_n49237_ = ys__n37968 & new_n44786_;
  assign new_n49238_ = ys__n18708 & ~new_n44790_;
  assign new_n49239_ = ~new_n49237_ & ~new_n49238_;
  assign ys__n32640 = ~new_n44793_ & ~new_n49239_;
  assign new_n49241_ = ys__n37969 & new_n44786_;
  assign new_n49242_ = ys__n18711 & ~new_n44790_;
  assign new_n49243_ = ~new_n49241_ & ~new_n49242_;
  assign ys__n32641 = ~new_n44793_ & ~new_n49243_;
  assign new_n49245_ = ys__n37970 & new_n44786_;
  assign new_n49246_ = ys__n18714 & ~new_n44790_;
  assign new_n49247_ = ~new_n49245_ & ~new_n49246_;
  assign ys__n32642 = ~new_n44793_ & ~new_n49247_;
  assign new_n49249_ = ys__n37971 & new_n44786_;
  assign new_n49250_ = ys__n18717 & ~new_n44790_;
  assign new_n49251_ = ~new_n49249_ & ~new_n49250_;
  assign ys__n32643 = ~new_n44793_ & ~new_n49251_;
  assign new_n49253_ = ys__n37972 & new_n44786_;
  assign new_n49254_ = ys__n18720 & ~new_n44790_;
  assign new_n49255_ = ~new_n49253_ & ~new_n49254_;
  assign ys__n32644 = ~new_n44793_ & ~new_n49255_;
  assign new_n49257_ = ys__n37973 & new_n44786_;
  assign new_n49258_ = ys__n18723 & ~new_n44790_;
  assign new_n49259_ = ~new_n49257_ & ~new_n49258_;
  assign ys__n32645 = ~new_n44793_ & ~new_n49259_;
  assign new_n49261_ = ys__n37974 & new_n44786_;
  assign new_n49262_ = ys__n18726 & ~new_n44790_;
  assign new_n49263_ = ~new_n49261_ & ~new_n49262_;
  assign ys__n32646 = ~new_n44793_ & ~new_n49263_;
  assign new_n49265_ = ys__n37975 & new_n44786_;
  assign new_n49266_ = ys__n18729 & ~new_n44790_;
  assign new_n49267_ = ~new_n49265_ & ~new_n49266_;
  assign ys__n32647 = ~new_n44793_ & ~new_n49267_;
  assign new_n49269_ = ys__n37976 & new_n44786_;
  assign new_n49270_ = ys__n18732 & ~new_n44790_;
  assign new_n49271_ = ~new_n49269_ & ~new_n49270_;
  assign ys__n32648 = ~new_n44793_ & ~new_n49271_;
  assign new_n49273_ = ys__n37977 & new_n44786_;
  assign new_n49274_ = ys__n18735 & ~new_n44790_;
  assign new_n49275_ = ~new_n49273_ & ~new_n49274_;
  assign ys__n32649 = ~new_n44793_ & ~new_n49275_;
  assign new_n49277_ = ys__n37978 & new_n44786_;
  assign new_n49278_ = ys__n18738 & ~new_n44790_;
  assign new_n49279_ = ~new_n49277_ & ~new_n49278_;
  assign ys__n32650 = ~new_n44793_ & ~new_n49279_;
  assign new_n49281_ = ys__n37979 & new_n44786_;
  assign new_n49282_ = ys__n18741 & ~new_n44790_;
  assign new_n49283_ = ~new_n49281_ & ~new_n49282_;
  assign ys__n32651 = ~new_n44793_ & ~new_n49283_;
  assign new_n49285_ = ys__n37980 & new_n44786_;
  assign new_n49286_ = ys__n18744 & ~new_n44790_;
  assign new_n49287_ = ~new_n49285_ & ~new_n49286_;
  assign ys__n32652 = ~new_n44793_ & ~new_n49287_;
  assign new_n49289_ = ys__n37981 & new_n44786_;
  assign new_n49290_ = ys__n18747 & ~new_n44790_;
  assign new_n49291_ = ~new_n49289_ & ~new_n49290_;
  assign ys__n32653 = ~new_n44793_ & ~new_n49291_;
  assign new_n49293_ = ys__n48126 & new_n44641_;
  assign new_n49294_ = ys__n18654 & ~new_n44645_;
  assign new_n49295_ = ~new_n49293_ & ~new_n49294_;
  assign ys__n32654 = ~new_n44648_ & ~new_n49295_;
  assign new_n49297_ = ys__n48127 & new_n44641_;
  assign new_n49298_ = ys__n18657 & ~new_n44645_;
  assign new_n49299_ = ~new_n49297_ & ~new_n49298_;
  assign ys__n32655 = ~new_n44648_ & ~new_n49299_;
  assign new_n49301_ = ys__n48128 & new_n44641_;
  assign new_n49302_ = ys__n18660 & ~new_n44645_;
  assign new_n49303_ = ~new_n49301_ & ~new_n49302_;
  assign ys__n32656 = ~new_n44648_ & ~new_n49303_;
  assign new_n49305_ = ys__n48129 & new_n44641_;
  assign new_n49306_ = ys__n18663 & ~new_n44645_;
  assign new_n49307_ = ~new_n49305_ & ~new_n49306_;
  assign ys__n32657 = ~new_n44648_ & ~new_n49307_;
  assign new_n49309_ = ys__n37982 & new_n44641_;
  assign new_n49310_ = ys__n18666 & ~new_n44645_;
  assign new_n49311_ = ~new_n49309_ & ~new_n49310_;
  assign ys__n32658 = ~new_n44648_ & ~new_n49311_;
  assign new_n49313_ = ys__n37983 & new_n44641_;
  assign new_n49314_ = ys__n18669 & ~new_n44645_;
  assign new_n49315_ = ~new_n49313_ & ~new_n49314_;
  assign ys__n32659 = ~new_n44648_ & ~new_n49315_;
  assign new_n49317_ = ys__n37984 & new_n44641_;
  assign new_n49318_ = ys__n18672 & ~new_n44645_;
  assign new_n49319_ = ~new_n49317_ & ~new_n49318_;
  assign ys__n32660 = ~new_n44648_ & ~new_n49319_;
  assign new_n49321_ = ys__n37985 & new_n44641_;
  assign new_n49322_ = ys__n18675 & ~new_n44645_;
  assign new_n49323_ = ~new_n49321_ & ~new_n49322_;
  assign ys__n32661 = ~new_n44648_ & ~new_n49323_;
  assign new_n49325_ = ys__n37986 & new_n44641_;
  assign new_n49326_ = ys__n18678 & ~new_n44645_;
  assign new_n49327_ = ~new_n49325_ & ~new_n49326_;
  assign ys__n32662 = ~new_n44648_ & ~new_n49327_;
  assign new_n49329_ = ys__n37987 & new_n44641_;
  assign new_n49330_ = ys__n18681 & ~new_n44645_;
  assign new_n49331_ = ~new_n49329_ & ~new_n49330_;
  assign ys__n32663 = ~new_n44648_ & ~new_n49331_;
  assign new_n49333_ = ys__n37988 & new_n44641_;
  assign new_n49334_ = ys__n18684 & ~new_n44645_;
  assign new_n49335_ = ~new_n49333_ & ~new_n49334_;
  assign ys__n32664 = ~new_n44648_ & ~new_n49335_;
  assign new_n49337_ = ys__n37989 & new_n44641_;
  assign new_n49338_ = ys__n18687 & ~new_n44645_;
  assign new_n49339_ = ~new_n49337_ & ~new_n49338_;
  assign ys__n32665 = ~new_n44648_ & ~new_n49339_;
  assign new_n49341_ = ys__n37990 & new_n44641_;
  assign new_n49342_ = ys__n18690 & ~new_n44645_;
  assign new_n49343_ = ~new_n49341_ & ~new_n49342_;
  assign ys__n32666 = ~new_n44648_ & ~new_n49343_;
  assign new_n49345_ = ys__n37991 & new_n44641_;
  assign new_n49346_ = ys__n18693 & ~new_n44645_;
  assign new_n49347_ = ~new_n49345_ & ~new_n49346_;
  assign ys__n32667 = ~new_n44648_ & ~new_n49347_;
  assign new_n49349_ = ys__n37992 & new_n44641_;
  assign new_n49350_ = ys__n18696 & ~new_n44645_;
  assign new_n49351_ = ~new_n49349_ & ~new_n49350_;
  assign ys__n32668 = ~new_n44648_ & ~new_n49351_;
  assign new_n49353_ = ys__n37993 & new_n44641_;
  assign new_n49354_ = ys__n18699 & ~new_n44645_;
  assign new_n49355_ = ~new_n49353_ & ~new_n49354_;
  assign ys__n32669 = ~new_n44648_ & ~new_n49355_;
  assign new_n49357_ = ys__n37994 & new_n44641_;
  assign new_n49358_ = ys__n18702 & ~new_n44645_;
  assign new_n49359_ = ~new_n49357_ & ~new_n49358_;
  assign ys__n32670 = ~new_n44648_ & ~new_n49359_;
  assign new_n49361_ = ys__n37995 & new_n44641_;
  assign new_n49362_ = ys__n18705 & ~new_n44645_;
  assign new_n49363_ = ~new_n49361_ & ~new_n49362_;
  assign ys__n32671 = ~new_n44648_ & ~new_n49363_;
  assign new_n49365_ = ys__n37996 & new_n44641_;
  assign new_n49366_ = ys__n18708 & ~new_n44645_;
  assign new_n49367_ = ~new_n49365_ & ~new_n49366_;
  assign ys__n32672 = ~new_n44648_ & ~new_n49367_;
  assign new_n49369_ = ys__n37997 & new_n44641_;
  assign new_n49370_ = ys__n18711 & ~new_n44645_;
  assign new_n49371_ = ~new_n49369_ & ~new_n49370_;
  assign ys__n32673 = ~new_n44648_ & ~new_n49371_;
  assign new_n49373_ = ys__n37998 & new_n44641_;
  assign new_n49374_ = ys__n18714 & ~new_n44645_;
  assign new_n49375_ = ~new_n49373_ & ~new_n49374_;
  assign ys__n32674 = ~new_n44648_ & ~new_n49375_;
  assign new_n49377_ = ys__n37999 & new_n44641_;
  assign new_n49378_ = ys__n18717 & ~new_n44645_;
  assign new_n49379_ = ~new_n49377_ & ~new_n49378_;
  assign ys__n32675 = ~new_n44648_ & ~new_n49379_;
  assign new_n49381_ = ys__n38000 & new_n44641_;
  assign new_n49382_ = ys__n18720 & ~new_n44645_;
  assign new_n49383_ = ~new_n49381_ & ~new_n49382_;
  assign ys__n32676 = ~new_n44648_ & ~new_n49383_;
  assign new_n49385_ = ys__n38001 & new_n44641_;
  assign new_n49386_ = ys__n18723 & ~new_n44645_;
  assign new_n49387_ = ~new_n49385_ & ~new_n49386_;
  assign ys__n32677 = ~new_n44648_ & ~new_n49387_;
  assign new_n49389_ = ys__n38002 & new_n44641_;
  assign new_n49390_ = ys__n18726 & ~new_n44645_;
  assign new_n49391_ = ~new_n49389_ & ~new_n49390_;
  assign ys__n32678 = ~new_n44648_ & ~new_n49391_;
  assign new_n49393_ = ys__n38003 & new_n44641_;
  assign new_n49394_ = ys__n18729 & ~new_n44645_;
  assign new_n49395_ = ~new_n49393_ & ~new_n49394_;
  assign ys__n32679 = ~new_n44648_ & ~new_n49395_;
  assign new_n49397_ = ys__n38004 & new_n44641_;
  assign new_n49398_ = ys__n18732 & ~new_n44645_;
  assign new_n49399_ = ~new_n49397_ & ~new_n49398_;
  assign ys__n32680 = ~new_n44648_ & ~new_n49399_;
  assign new_n49401_ = ys__n38005 & new_n44641_;
  assign new_n49402_ = ys__n18735 & ~new_n44645_;
  assign new_n49403_ = ~new_n49401_ & ~new_n49402_;
  assign ys__n32681 = ~new_n44648_ & ~new_n49403_;
  assign new_n49405_ = ys__n38006 & new_n44641_;
  assign new_n49406_ = ys__n18738 & ~new_n44645_;
  assign new_n49407_ = ~new_n49405_ & ~new_n49406_;
  assign ys__n32682 = ~new_n44648_ & ~new_n49407_;
  assign new_n49409_ = ys__n38007 & new_n44641_;
  assign new_n49410_ = ys__n18741 & ~new_n44645_;
  assign new_n49411_ = ~new_n49409_ & ~new_n49410_;
  assign ys__n32683 = ~new_n44648_ & ~new_n49411_;
  assign new_n49413_ = ys__n38008 & new_n44641_;
  assign new_n49414_ = ys__n18744 & ~new_n44645_;
  assign new_n49415_ = ~new_n49413_ & ~new_n49414_;
  assign ys__n32684 = ~new_n44648_ & ~new_n49415_;
  assign new_n49417_ = ys__n38009 & new_n44641_;
  assign new_n49418_ = ys__n18747 & ~new_n44645_;
  assign new_n49419_ = ~new_n49417_ & ~new_n49418_;
  assign ys__n32685 = ~new_n44648_ & ~new_n49419_;
  assign new_n49421_ = ys__n48130 & new_n44317_;
  assign new_n49422_ = ys__n18654 & ~new_n44321_;
  assign new_n49423_ = ~new_n49421_ & ~new_n49422_;
  assign ys__n32686 = ~new_n44324_ & ~new_n49423_;
  assign new_n49425_ = ys__n48131 & new_n44317_;
  assign new_n49426_ = ys__n18657 & ~new_n44321_;
  assign new_n49427_ = ~new_n49425_ & ~new_n49426_;
  assign ys__n32687 = ~new_n44324_ & ~new_n49427_;
  assign new_n49429_ = ys__n48132 & new_n44317_;
  assign new_n49430_ = ys__n18660 & ~new_n44321_;
  assign new_n49431_ = ~new_n49429_ & ~new_n49430_;
  assign ys__n32688 = ~new_n44324_ & ~new_n49431_;
  assign new_n49433_ = ys__n48133 & new_n44317_;
  assign new_n49434_ = ys__n18663 & ~new_n44321_;
  assign new_n49435_ = ~new_n49433_ & ~new_n49434_;
  assign ys__n32689 = ~new_n44324_ & ~new_n49435_;
  assign new_n49437_ = ys__n38010 & new_n44317_;
  assign new_n49438_ = ys__n18666 & ~new_n44321_;
  assign new_n49439_ = ~new_n49437_ & ~new_n49438_;
  assign ys__n32690 = ~new_n44324_ & ~new_n49439_;
  assign new_n49441_ = ys__n38011 & new_n44317_;
  assign new_n49442_ = ys__n18669 & ~new_n44321_;
  assign new_n49443_ = ~new_n49441_ & ~new_n49442_;
  assign ys__n32691 = ~new_n44324_ & ~new_n49443_;
  assign new_n49445_ = ys__n38012 & new_n44317_;
  assign new_n49446_ = ys__n18672 & ~new_n44321_;
  assign new_n49447_ = ~new_n49445_ & ~new_n49446_;
  assign ys__n32692 = ~new_n44324_ & ~new_n49447_;
  assign new_n49449_ = ys__n38013 & new_n44317_;
  assign new_n49450_ = ys__n18675 & ~new_n44321_;
  assign new_n49451_ = ~new_n49449_ & ~new_n49450_;
  assign ys__n32693 = ~new_n44324_ & ~new_n49451_;
  assign new_n49453_ = ys__n38014 & new_n44317_;
  assign new_n49454_ = ys__n18678 & ~new_n44321_;
  assign new_n49455_ = ~new_n49453_ & ~new_n49454_;
  assign ys__n32694 = ~new_n44324_ & ~new_n49455_;
  assign new_n49457_ = ys__n38015 & new_n44317_;
  assign new_n49458_ = ys__n18681 & ~new_n44321_;
  assign new_n49459_ = ~new_n49457_ & ~new_n49458_;
  assign ys__n32695 = ~new_n44324_ & ~new_n49459_;
  assign new_n49461_ = ys__n38016 & new_n44317_;
  assign new_n49462_ = ys__n18684 & ~new_n44321_;
  assign new_n49463_ = ~new_n49461_ & ~new_n49462_;
  assign ys__n32696 = ~new_n44324_ & ~new_n49463_;
  assign new_n49465_ = ys__n38017 & new_n44317_;
  assign new_n49466_ = ys__n18687 & ~new_n44321_;
  assign new_n49467_ = ~new_n49465_ & ~new_n49466_;
  assign ys__n32697 = ~new_n44324_ & ~new_n49467_;
  assign new_n49469_ = ys__n38018 & new_n44317_;
  assign new_n49470_ = ys__n18690 & ~new_n44321_;
  assign new_n49471_ = ~new_n49469_ & ~new_n49470_;
  assign ys__n32698 = ~new_n44324_ & ~new_n49471_;
  assign new_n49473_ = ys__n38019 & new_n44317_;
  assign new_n49474_ = ys__n18693 & ~new_n44321_;
  assign new_n49475_ = ~new_n49473_ & ~new_n49474_;
  assign ys__n32699 = ~new_n44324_ & ~new_n49475_;
  assign new_n49477_ = ys__n38020 & new_n44317_;
  assign new_n49478_ = ys__n18696 & ~new_n44321_;
  assign new_n49479_ = ~new_n49477_ & ~new_n49478_;
  assign ys__n32700 = ~new_n44324_ & ~new_n49479_;
  assign new_n49481_ = ys__n38021 & new_n44317_;
  assign new_n49482_ = ys__n18699 & ~new_n44321_;
  assign new_n49483_ = ~new_n49481_ & ~new_n49482_;
  assign ys__n32701 = ~new_n44324_ & ~new_n49483_;
  assign new_n49485_ = ys__n38022 & new_n44317_;
  assign new_n49486_ = ys__n18702 & ~new_n44321_;
  assign new_n49487_ = ~new_n49485_ & ~new_n49486_;
  assign ys__n32702 = ~new_n44324_ & ~new_n49487_;
  assign new_n49489_ = ys__n38023 & new_n44317_;
  assign new_n49490_ = ys__n18705 & ~new_n44321_;
  assign new_n49491_ = ~new_n49489_ & ~new_n49490_;
  assign ys__n32703 = ~new_n44324_ & ~new_n49491_;
  assign new_n49493_ = ys__n38024 & new_n44317_;
  assign new_n49494_ = ys__n18708 & ~new_n44321_;
  assign new_n49495_ = ~new_n49493_ & ~new_n49494_;
  assign ys__n32704 = ~new_n44324_ & ~new_n49495_;
  assign new_n49497_ = ys__n38025 & new_n44317_;
  assign new_n49498_ = ys__n18711 & ~new_n44321_;
  assign new_n49499_ = ~new_n49497_ & ~new_n49498_;
  assign ys__n32705 = ~new_n44324_ & ~new_n49499_;
  assign new_n49501_ = ys__n38026 & new_n44317_;
  assign new_n49502_ = ys__n18714 & ~new_n44321_;
  assign new_n49503_ = ~new_n49501_ & ~new_n49502_;
  assign ys__n32706 = ~new_n44324_ & ~new_n49503_;
  assign new_n49505_ = ys__n38027 & new_n44317_;
  assign new_n49506_ = ys__n18717 & ~new_n44321_;
  assign new_n49507_ = ~new_n49505_ & ~new_n49506_;
  assign ys__n32707 = ~new_n44324_ & ~new_n49507_;
  assign new_n49509_ = ys__n38028 & new_n44317_;
  assign new_n49510_ = ys__n18720 & ~new_n44321_;
  assign new_n49511_ = ~new_n49509_ & ~new_n49510_;
  assign ys__n32708 = ~new_n44324_ & ~new_n49511_;
  assign new_n49513_ = ys__n38029 & new_n44317_;
  assign new_n49514_ = ys__n18723 & ~new_n44321_;
  assign new_n49515_ = ~new_n49513_ & ~new_n49514_;
  assign ys__n32709 = ~new_n44324_ & ~new_n49515_;
  assign new_n49517_ = ys__n38030 & new_n44317_;
  assign new_n49518_ = ys__n18726 & ~new_n44321_;
  assign new_n49519_ = ~new_n49517_ & ~new_n49518_;
  assign ys__n32710 = ~new_n44324_ & ~new_n49519_;
  assign new_n49521_ = ys__n38031 & new_n44317_;
  assign new_n49522_ = ys__n18729 & ~new_n44321_;
  assign new_n49523_ = ~new_n49521_ & ~new_n49522_;
  assign ys__n32711 = ~new_n44324_ & ~new_n49523_;
  assign new_n49525_ = ys__n38032 & new_n44317_;
  assign new_n49526_ = ys__n18732 & ~new_n44321_;
  assign new_n49527_ = ~new_n49525_ & ~new_n49526_;
  assign ys__n32712 = ~new_n44324_ & ~new_n49527_;
  assign new_n49529_ = ys__n38033 & new_n44317_;
  assign new_n49530_ = ys__n18735 & ~new_n44321_;
  assign new_n49531_ = ~new_n49529_ & ~new_n49530_;
  assign ys__n32713 = ~new_n44324_ & ~new_n49531_;
  assign new_n49533_ = ys__n38034 & new_n44317_;
  assign new_n49534_ = ys__n18738 & ~new_n44321_;
  assign new_n49535_ = ~new_n49533_ & ~new_n49534_;
  assign ys__n32714 = ~new_n44324_ & ~new_n49535_;
  assign new_n49537_ = ys__n38035 & new_n44317_;
  assign new_n49538_ = ys__n18741 & ~new_n44321_;
  assign new_n49539_ = ~new_n49537_ & ~new_n49538_;
  assign ys__n32715 = ~new_n44324_ & ~new_n49539_;
  assign new_n49541_ = ys__n38036 & new_n44317_;
  assign new_n49542_ = ys__n18744 & ~new_n44321_;
  assign new_n49543_ = ~new_n49541_ & ~new_n49542_;
  assign ys__n32716 = ~new_n44324_ & ~new_n49543_;
  assign new_n49545_ = ys__n38037 & new_n44317_;
  assign new_n49546_ = ys__n18747 & ~new_n44321_;
  assign new_n49547_ = ~new_n49545_ & ~new_n49546_;
  assign ys__n32717 = ~new_n44324_ & ~new_n49547_;
  assign new_n49549_ = ys__n48134 & new_n44462_;
  assign new_n49550_ = ys__n18654 & ~new_n44466_;
  assign new_n49551_ = ~new_n49549_ & ~new_n49550_;
  assign ys__n32718 = ~new_n44469_ & ~new_n49551_;
  assign new_n49553_ = ys__n48135 & new_n44462_;
  assign new_n49554_ = ys__n18657 & ~new_n44466_;
  assign new_n49555_ = ~new_n49553_ & ~new_n49554_;
  assign ys__n32719 = ~new_n44469_ & ~new_n49555_;
  assign new_n49557_ = ys__n48136 & new_n44462_;
  assign new_n49558_ = ys__n18660 & ~new_n44466_;
  assign new_n49559_ = ~new_n49557_ & ~new_n49558_;
  assign ys__n32720 = ~new_n44469_ & ~new_n49559_;
  assign new_n49561_ = ys__n48137 & new_n44462_;
  assign new_n49562_ = ys__n18663 & ~new_n44466_;
  assign new_n49563_ = ~new_n49561_ & ~new_n49562_;
  assign ys__n32721 = ~new_n44469_ & ~new_n49563_;
  assign new_n49565_ = ys__n38038 & new_n44462_;
  assign new_n49566_ = ys__n18666 & ~new_n44466_;
  assign new_n49567_ = ~new_n49565_ & ~new_n49566_;
  assign ys__n32722 = ~new_n44469_ & ~new_n49567_;
  assign new_n49569_ = ys__n38039 & new_n44462_;
  assign new_n49570_ = ys__n18669 & ~new_n44466_;
  assign new_n49571_ = ~new_n49569_ & ~new_n49570_;
  assign ys__n32723 = ~new_n44469_ & ~new_n49571_;
  assign new_n49573_ = ys__n38040 & new_n44462_;
  assign new_n49574_ = ys__n18672 & ~new_n44466_;
  assign new_n49575_ = ~new_n49573_ & ~new_n49574_;
  assign ys__n32724 = ~new_n44469_ & ~new_n49575_;
  assign new_n49577_ = ys__n38041 & new_n44462_;
  assign new_n49578_ = ys__n18675 & ~new_n44466_;
  assign new_n49579_ = ~new_n49577_ & ~new_n49578_;
  assign ys__n32725 = ~new_n44469_ & ~new_n49579_;
  assign new_n49581_ = ys__n38042 & new_n44462_;
  assign new_n49582_ = ys__n18678 & ~new_n44466_;
  assign new_n49583_ = ~new_n49581_ & ~new_n49582_;
  assign ys__n32726 = ~new_n44469_ & ~new_n49583_;
  assign new_n49585_ = ys__n38043 & new_n44462_;
  assign new_n49586_ = ys__n18681 & ~new_n44466_;
  assign new_n49587_ = ~new_n49585_ & ~new_n49586_;
  assign ys__n32727 = ~new_n44469_ & ~new_n49587_;
  assign new_n49589_ = ys__n38044 & new_n44462_;
  assign new_n49590_ = ys__n18684 & ~new_n44466_;
  assign new_n49591_ = ~new_n49589_ & ~new_n49590_;
  assign ys__n32728 = ~new_n44469_ & ~new_n49591_;
  assign new_n49593_ = ys__n38045 & new_n44462_;
  assign new_n49594_ = ys__n18687 & ~new_n44466_;
  assign new_n49595_ = ~new_n49593_ & ~new_n49594_;
  assign ys__n32729 = ~new_n44469_ & ~new_n49595_;
  assign new_n49597_ = ys__n38046 & new_n44462_;
  assign new_n49598_ = ys__n18690 & ~new_n44466_;
  assign new_n49599_ = ~new_n49597_ & ~new_n49598_;
  assign ys__n32730 = ~new_n44469_ & ~new_n49599_;
  assign new_n49601_ = ys__n38047 & new_n44462_;
  assign new_n49602_ = ys__n18693 & ~new_n44466_;
  assign new_n49603_ = ~new_n49601_ & ~new_n49602_;
  assign ys__n32731 = ~new_n44469_ & ~new_n49603_;
  assign new_n49605_ = ys__n38048 & new_n44462_;
  assign new_n49606_ = ys__n18696 & ~new_n44466_;
  assign new_n49607_ = ~new_n49605_ & ~new_n49606_;
  assign ys__n32732 = ~new_n44469_ & ~new_n49607_;
  assign new_n49609_ = ys__n38049 & new_n44462_;
  assign new_n49610_ = ys__n18699 & ~new_n44466_;
  assign new_n49611_ = ~new_n49609_ & ~new_n49610_;
  assign ys__n32733 = ~new_n44469_ & ~new_n49611_;
  assign new_n49613_ = ys__n38050 & new_n44462_;
  assign new_n49614_ = ys__n18702 & ~new_n44466_;
  assign new_n49615_ = ~new_n49613_ & ~new_n49614_;
  assign ys__n32734 = ~new_n44469_ & ~new_n49615_;
  assign new_n49617_ = ys__n38051 & new_n44462_;
  assign new_n49618_ = ys__n18705 & ~new_n44466_;
  assign new_n49619_ = ~new_n49617_ & ~new_n49618_;
  assign ys__n32735 = ~new_n44469_ & ~new_n49619_;
  assign new_n49621_ = ys__n38052 & new_n44462_;
  assign new_n49622_ = ys__n18708 & ~new_n44466_;
  assign new_n49623_ = ~new_n49621_ & ~new_n49622_;
  assign ys__n32736 = ~new_n44469_ & ~new_n49623_;
  assign new_n49625_ = ys__n38053 & new_n44462_;
  assign new_n49626_ = ys__n18711 & ~new_n44466_;
  assign new_n49627_ = ~new_n49625_ & ~new_n49626_;
  assign ys__n32737 = ~new_n44469_ & ~new_n49627_;
  assign new_n49629_ = ys__n38054 & new_n44462_;
  assign new_n49630_ = ys__n18714 & ~new_n44466_;
  assign new_n49631_ = ~new_n49629_ & ~new_n49630_;
  assign ys__n32738 = ~new_n44469_ & ~new_n49631_;
  assign new_n49633_ = ys__n38055 & new_n44462_;
  assign new_n49634_ = ys__n18717 & ~new_n44466_;
  assign new_n49635_ = ~new_n49633_ & ~new_n49634_;
  assign ys__n32739 = ~new_n44469_ & ~new_n49635_;
  assign new_n49637_ = ys__n38056 & new_n44462_;
  assign new_n49638_ = ys__n18720 & ~new_n44466_;
  assign new_n49639_ = ~new_n49637_ & ~new_n49638_;
  assign ys__n32740 = ~new_n44469_ & ~new_n49639_;
  assign new_n49641_ = ys__n38057 & new_n44462_;
  assign new_n49642_ = ys__n18723 & ~new_n44466_;
  assign new_n49643_ = ~new_n49641_ & ~new_n49642_;
  assign ys__n32741 = ~new_n44469_ & ~new_n49643_;
  assign new_n49645_ = ys__n38058 & new_n44462_;
  assign new_n49646_ = ys__n18726 & ~new_n44466_;
  assign new_n49647_ = ~new_n49645_ & ~new_n49646_;
  assign ys__n32742 = ~new_n44469_ & ~new_n49647_;
  assign new_n49649_ = ys__n38059 & new_n44462_;
  assign new_n49650_ = ys__n18729 & ~new_n44466_;
  assign new_n49651_ = ~new_n49649_ & ~new_n49650_;
  assign ys__n32743 = ~new_n44469_ & ~new_n49651_;
  assign new_n49653_ = ys__n38060 & new_n44462_;
  assign new_n49654_ = ys__n18732 & ~new_n44466_;
  assign new_n49655_ = ~new_n49653_ & ~new_n49654_;
  assign ys__n32744 = ~new_n44469_ & ~new_n49655_;
  assign new_n49657_ = ys__n38061 & new_n44462_;
  assign new_n49658_ = ys__n18735 & ~new_n44466_;
  assign new_n49659_ = ~new_n49657_ & ~new_n49658_;
  assign ys__n32745 = ~new_n44469_ & ~new_n49659_;
  assign new_n49661_ = ys__n38062 & new_n44462_;
  assign new_n49662_ = ys__n18738 & ~new_n44466_;
  assign new_n49663_ = ~new_n49661_ & ~new_n49662_;
  assign ys__n32746 = ~new_n44469_ & ~new_n49663_;
  assign new_n49665_ = ys__n38063 & new_n44462_;
  assign new_n49666_ = ys__n18741 & ~new_n44466_;
  assign new_n49667_ = ~new_n49665_ & ~new_n49666_;
  assign ys__n32747 = ~new_n44469_ & ~new_n49667_;
  assign new_n49669_ = ys__n38064 & new_n44462_;
  assign new_n49670_ = ys__n18744 & ~new_n44466_;
  assign new_n49671_ = ~new_n49669_ & ~new_n49670_;
  assign ys__n32748 = ~new_n44469_ & ~new_n49671_;
  assign new_n49673_ = ys__n38065 & new_n44462_;
  assign new_n49674_ = ys__n18747 & ~new_n44466_;
  assign new_n49675_ = ~new_n49673_ & ~new_n49674_;
  assign ys__n32749 = ~new_n44469_ & ~new_n49675_;
  assign new_n49677_ = ys__n48138 & new_n44172_;
  assign new_n49678_ = ys__n18654 & ~new_n44176_;
  assign new_n49679_ = ~new_n49677_ & ~new_n49678_;
  assign ys__n32750 = ~new_n44179_ & ~new_n49679_;
  assign new_n49681_ = ys__n48139 & new_n44172_;
  assign new_n49682_ = ys__n18657 & ~new_n44176_;
  assign new_n49683_ = ~new_n49681_ & ~new_n49682_;
  assign ys__n32751 = ~new_n44179_ & ~new_n49683_;
  assign new_n49685_ = ys__n48140 & new_n44172_;
  assign new_n49686_ = ys__n18660 & ~new_n44176_;
  assign new_n49687_ = ~new_n49685_ & ~new_n49686_;
  assign ys__n32752 = ~new_n44179_ & ~new_n49687_;
  assign new_n49689_ = ys__n48141 & new_n44172_;
  assign new_n49690_ = ys__n18663 & ~new_n44176_;
  assign new_n49691_ = ~new_n49689_ & ~new_n49690_;
  assign ys__n32753 = ~new_n44179_ & ~new_n49691_;
  assign new_n49693_ = ys__n38066 & new_n44172_;
  assign new_n49694_ = ys__n18666 & ~new_n44176_;
  assign new_n49695_ = ~new_n49693_ & ~new_n49694_;
  assign ys__n32754 = ~new_n44179_ & ~new_n49695_;
  assign new_n49697_ = ys__n38067 & new_n44172_;
  assign new_n49698_ = ys__n18669 & ~new_n44176_;
  assign new_n49699_ = ~new_n49697_ & ~new_n49698_;
  assign ys__n32755 = ~new_n44179_ & ~new_n49699_;
  assign new_n49701_ = ys__n38068 & new_n44172_;
  assign new_n49702_ = ys__n18672 & ~new_n44176_;
  assign new_n49703_ = ~new_n49701_ & ~new_n49702_;
  assign ys__n32756 = ~new_n44179_ & ~new_n49703_;
  assign new_n49705_ = ys__n38069 & new_n44172_;
  assign new_n49706_ = ys__n18675 & ~new_n44176_;
  assign new_n49707_ = ~new_n49705_ & ~new_n49706_;
  assign ys__n32757 = ~new_n44179_ & ~new_n49707_;
  assign new_n49709_ = ys__n38070 & new_n44172_;
  assign new_n49710_ = ys__n18678 & ~new_n44176_;
  assign new_n49711_ = ~new_n49709_ & ~new_n49710_;
  assign ys__n32758 = ~new_n44179_ & ~new_n49711_;
  assign new_n49713_ = ys__n38071 & new_n44172_;
  assign new_n49714_ = ys__n18681 & ~new_n44176_;
  assign new_n49715_ = ~new_n49713_ & ~new_n49714_;
  assign ys__n32759 = ~new_n44179_ & ~new_n49715_;
  assign new_n49717_ = ys__n38072 & new_n44172_;
  assign new_n49718_ = ys__n18684 & ~new_n44176_;
  assign new_n49719_ = ~new_n49717_ & ~new_n49718_;
  assign ys__n32760 = ~new_n44179_ & ~new_n49719_;
  assign new_n49721_ = ys__n38073 & new_n44172_;
  assign new_n49722_ = ys__n18687 & ~new_n44176_;
  assign new_n49723_ = ~new_n49721_ & ~new_n49722_;
  assign ys__n32761 = ~new_n44179_ & ~new_n49723_;
  assign new_n49725_ = ys__n38074 & new_n44172_;
  assign new_n49726_ = ys__n18690 & ~new_n44176_;
  assign new_n49727_ = ~new_n49725_ & ~new_n49726_;
  assign ys__n32762 = ~new_n44179_ & ~new_n49727_;
  assign new_n49729_ = ys__n38075 & new_n44172_;
  assign new_n49730_ = ys__n18693 & ~new_n44176_;
  assign new_n49731_ = ~new_n49729_ & ~new_n49730_;
  assign ys__n32763 = ~new_n44179_ & ~new_n49731_;
  assign new_n49733_ = ys__n38076 & new_n44172_;
  assign new_n49734_ = ys__n18696 & ~new_n44176_;
  assign new_n49735_ = ~new_n49733_ & ~new_n49734_;
  assign ys__n32764 = ~new_n44179_ & ~new_n49735_;
  assign new_n49737_ = ys__n38077 & new_n44172_;
  assign new_n49738_ = ys__n18699 & ~new_n44176_;
  assign new_n49739_ = ~new_n49737_ & ~new_n49738_;
  assign ys__n32765 = ~new_n44179_ & ~new_n49739_;
  assign new_n49741_ = ys__n38078 & new_n44172_;
  assign new_n49742_ = ys__n18702 & ~new_n44176_;
  assign new_n49743_ = ~new_n49741_ & ~new_n49742_;
  assign ys__n32766 = ~new_n44179_ & ~new_n49743_;
  assign new_n49745_ = ys__n38079 & new_n44172_;
  assign new_n49746_ = ys__n18705 & ~new_n44176_;
  assign new_n49747_ = ~new_n49745_ & ~new_n49746_;
  assign ys__n32767 = ~new_n44179_ & ~new_n49747_;
  assign new_n49749_ = ys__n38080 & new_n44172_;
  assign new_n49750_ = ys__n18708 & ~new_n44176_;
  assign new_n49751_ = ~new_n49749_ & ~new_n49750_;
  assign ys__n32768 = ~new_n44179_ & ~new_n49751_;
  assign new_n49753_ = ys__n38081 & new_n44172_;
  assign new_n49754_ = ys__n18711 & ~new_n44176_;
  assign new_n49755_ = ~new_n49753_ & ~new_n49754_;
  assign ys__n32769 = ~new_n44179_ & ~new_n49755_;
  assign new_n49757_ = ys__n38082 & new_n44172_;
  assign new_n49758_ = ys__n18714 & ~new_n44176_;
  assign new_n49759_ = ~new_n49757_ & ~new_n49758_;
  assign ys__n32770 = ~new_n44179_ & ~new_n49759_;
  assign new_n49761_ = ys__n38083 & new_n44172_;
  assign new_n49762_ = ys__n18717 & ~new_n44176_;
  assign new_n49763_ = ~new_n49761_ & ~new_n49762_;
  assign ys__n32771 = ~new_n44179_ & ~new_n49763_;
  assign new_n49765_ = ys__n38084 & new_n44172_;
  assign new_n49766_ = ys__n18720 & ~new_n44176_;
  assign new_n49767_ = ~new_n49765_ & ~new_n49766_;
  assign ys__n32772 = ~new_n44179_ & ~new_n49767_;
  assign new_n49769_ = ys__n38085 & new_n44172_;
  assign new_n49770_ = ys__n18723 & ~new_n44176_;
  assign new_n49771_ = ~new_n49769_ & ~new_n49770_;
  assign ys__n32773 = ~new_n44179_ & ~new_n49771_;
  assign new_n49773_ = ys__n38086 & new_n44172_;
  assign new_n49774_ = ys__n18726 & ~new_n44176_;
  assign new_n49775_ = ~new_n49773_ & ~new_n49774_;
  assign ys__n32774 = ~new_n44179_ & ~new_n49775_;
  assign new_n49777_ = ys__n38087 & new_n44172_;
  assign new_n49778_ = ys__n18729 & ~new_n44176_;
  assign new_n49779_ = ~new_n49777_ & ~new_n49778_;
  assign ys__n32775 = ~new_n44179_ & ~new_n49779_;
  assign new_n49781_ = ys__n38088 & new_n44172_;
  assign new_n49782_ = ys__n18732 & ~new_n44176_;
  assign new_n49783_ = ~new_n49781_ & ~new_n49782_;
  assign ys__n32776 = ~new_n44179_ & ~new_n49783_;
  assign new_n49785_ = ys__n38089 & new_n44172_;
  assign new_n49786_ = ys__n18735 & ~new_n44176_;
  assign new_n49787_ = ~new_n49785_ & ~new_n49786_;
  assign ys__n32777 = ~new_n44179_ & ~new_n49787_;
  assign new_n49789_ = ys__n38090 & new_n44172_;
  assign new_n49790_ = ys__n18738 & ~new_n44176_;
  assign new_n49791_ = ~new_n49789_ & ~new_n49790_;
  assign ys__n32778 = ~new_n44179_ & ~new_n49791_;
  assign new_n49793_ = ys__n38091 & new_n44172_;
  assign new_n49794_ = ys__n18741 & ~new_n44176_;
  assign new_n49795_ = ~new_n49793_ & ~new_n49794_;
  assign ys__n32779 = ~new_n44179_ & ~new_n49795_;
  assign new_n49797_ = ys__n38092 & new_n44172_;
  assign new_n49798_ = ys__n18744 & ~new_n44176_;
  assign new_n49799_ = ~new_n49797_ & ~new_n49798_;
  assign ys__n32780 = ~new_n44179_ & ~new_n49799_;
  assign new_n49801_ = ys__n38093 & new_n44172_;
  assign new_n49802_ = ys__n18747 & ~new_n44176_;
  assign new_n49803_ = ~new_n49801_ & ~new_n49802_;
  assign ys__n32781 = ~new_n44179_ & ~new_n49803_;
  assign new_n49805_ = ys__n48142 & new_n43944_;
  assign new_n49806_ = ys__n18654 & ~new_n43948_;
  assign new_n49807_ = ~new_n49805_ & ~new_n49806_;
  assign ys__n32782 = ~new_n43951_ & ~new_n49807_;
  assign new_n49809_ = ys__n48143 & new_n43944_;
  assign new_n49810_ = ys__n18657 & ~new_n43948_;
  assign new_n49811_ = ~new_n49809_ & ~new_n49810_;
  assign ys__n32783 = ~new_n43951_ & ~new_n49811_;
  assign new_n49813_ = ys__n48144 & new_n43944_;
  assign new_n49814_ = ys__n18660 & ~new_n43948_;
  assign new_n49815_ = ~new_n49813_ & ~new_n49814_;
  assign ys__n32784 = ~new_n43951_ & ~new_n49815_;
  assign new_n49817_ = ys__n48145 & new_n43944_;
  assign new_n49818_ = ys__n18663 & ~new_n43948_;
  assign new_n49819_ = ~new_n49817_ & ~new_n49818_;
  assign ys__n32785 = ~new_n43951_ & ~new_n49819_;
  assign new_n49821_ = ys__n38094 & new_n43944_;
  assign new_n49822_ = ys__n18666 & ~new_n43948_;
  assign new_n49823_ = ~new_n49821_ & ~new_n49822_;
  assign ys__n32786 = ~new_n43951_ & ~new_n49823_;
  assign new_n49825_ = ys__n38095 & new_n43944_;
  assign new_n49826_ = ys__n18669 & ~new_n43948_;
  assign new_n49827_ = ~new_n49825_ & ~new_n49826_;
  assign ys__n32787 = ~new_n43951_ & ~new_n49827_;
  assign new_n49829_ = ys__n38096 & new_n43944_;
  assign new_n49830_ = ys__n18672 & ~new_n43948_;
  assign new_n49831_ = ~new_n49829_ & ~new_n49830_;
  assign ys__n32788 = ~new_n43951_ & ~new_n49831_;
  assign new_n49833_ = ys__n38097 & new_n43944_;
  assign new_n49834_ = ys__n18675 & ~new_n43948_;
  assign new_n49835_ = ~new_n49833_ & ~new_n49834_;
  assign ys__n32789 = ~new_n43951_ & ~new_n49835_;
  assign new_n49837_ = ys__n38098 & new_n43944_;
  assign new_n49838_ = ys__n18678 & ~new_n43948_;
  assign new_n49839_ = ~new_n49837_ & ~new_n49838_;
  assign ys__n32790 = ~new_n43951_ & ~new_n49839_;
  assign new_n49841_ = ys__n38099 & new_n43944_;
  assign new_n49842_ = ys__n18681 & ~new_n43948_;
  assign new_n49843_ = ~new_n49841_ & ~new_n49842_;
  assign ys__n32791 = ~new_n43951_ & ~new_n49843_;
  assign new_n49845_ = ys__n38100 & new_n43944_;
  assign new_n49846_ = ys__n18684 & ~new_n43948_;
  assign new_n49847_ = ~new_n49845_ & ~new_n49846_;
  assign ys__n32792 = ~new_n43951_ & ~new_n49847_;
  assign new_n49849_ = ys__n38101 & new_n43944_;
  assign new_n49850_ = ys__n18687 & ~new_n43948_;
  assign new_n49851_ = ~new_n49849_ & ~new_n49850_;
  assign ys__n32793 = ~new_n43951_ & ~new_n49851_;
  assign new_n49853_ = ys__n38102 & new_n43944_;
  assign new_n49854_ = ys__n18690 & ~new_n43948_;
  assign new_n49855_ = ~new_n49853_ & ~new_n49854_;
  assign ys__n32794 = ~new_n43951_ & ~new_n49855_;
  assign new_n49857_ = ys__n38103 & new_n43944_;
  assign new_n49858_ = ys__n18693 & ~new_n43948_;
  assign new_n49859_ = ~new_n49857_ & ~new_n49858_;
  assign ys__n32795 = ~new_n43951_ & ~new_n49859_;
  assign new_n49861_ = ys__n38104 & new_n43944_;
  assign new_n49862_ = ys__n18696 & ~new_n43948_;
  assign new_n49863_ = ~new_n49861_ & ~new_n49862_;
  assign ys__n32796 = ~new_n43951_ & ~new_n49863_;
  assign new_n49865_ = ys__n38105 & new_n43944_;
  assign new_n49866_ = ys__n18699 & ~new_n43948_;
  assign new_n49867_ = ~new_n49865_ & ~new_n49866_;
  assign ys__n32797 = ~new_n43951_ & ~new_n49867_;
  assign new_n49869_ = ys__n38106 & new_n43944_;
  assign new_n49870_ = ys__n18702 & ~new_n43948_;
  assign new_n49871_ = ~new_n49869_ & ~new_n49870_;
  assign ys__n32798 = ~new_n43951_ & ~new_n49871_;
  assign new_n49873_ = ys__n38107 & new_n43944_;
  assign new_n49874_ = ys__n18705 & ~new_n43948_;
  assign new_n49875_ = ~new_n49873_ & ~new_n49874_;
  assign ys__n32799 = ~new_n43951_ & ~new_n49875_;
  assign new_n49877_ = ys__n38108 & new_n43944_;
  assign new_n49878_ = ys__n18708 & ~new_n43948_;
  assign new_n49879_ = ~new_n49877_ & ~new_n49878_;
  assign ys__n32800 = ~new_n43951_ & ~new_n49879_;
  assign new_n49881_ = ys__n38109 & new_n43944_;
  assign new_n49882_ = ys__n18711 & ~new_n43948_;
  assign new_n49883_ = ~new_n49881_ & ~new_n49882_;
  assign ys__n32801 = ~new_n43951_ & ~new_n49883_;
  assign new_n49885_ = ys__n38110 & new_n43944_;
  assign new_n49886_ = ys__n18714 & ~new_n43948_;
  assign new_n49887_ = ~new_n49885_ & ~new_n49886_;
  assign ys__n32802 = ~new_n43951_ & ~new_n49887_;
  assign new_n49889_ = ys__n38111 & new_n43944_;
  assign new_n49890_ = ys__n18717 & ~new_n43948_;
  assign new_n49891_ = ~new_n49889_ & ~new_n49890_;
  assign ys__n32803 = ~new_n43951_ & ~new_n49891_;
  assign new_n49893_ = ys__n38112 & new_n43944_;
  assign new_n49894_ = ys__n18720 & ~new_n43948_;
  assign new_n49895_ = ~new_n49893_ & ~new_n49894_;
  assign ys__n32804 = ~new_n43951_ & ~new_n49895_;
  assign new_n49897_ = ys__n38113 & new_n43944_;
  assign new_n49898_ = ys__n18723 & ~new_n43948_;
  assign new_n49899_ = ~new_n49897_ & ~new_n49898_;
  assign ys__n32805 = ~new_n43951_ & ~new_n49899_;
  assign new_n49901_ = ys__n38114 & new_n43944_;
  assign new_n49902_ = ys__n18726 & ~new_n43948_;
  assign new_n49903_ = ~new_n49901_ & ~new_n49902_;
  assign ys__n32806 = ~new_n43951_ & ~new_n49903_;
  assign new_n49905_ = ys__n38115 & new_n43944_;
  assign new_n49906_ = ys__n18729 & ~new_n43948_;
  assign new_n49907_ = ~new_n49905_ & ~new_n49906_;
  assign ys__n32807 = ~new_n43951_ & ~new_n49907_;
  assign new_n49909_ = ys__n38116 & new_n43944_;
  assign new_n49910_ = ys__n18732 & ~new_n43948_;
  assign new_n49911_ = ~new_n49909_ & ~new_n49910_;
  assign ys__n32808 = ~new_n43951_ & ~new_n49911_;
  assign new_n49913_ = ys__n38117 & new_n43944_;
  assign new_n49914_ = ys__n18735 & ~new_n43948_;
  assign new_n49915_ = ~new_n49913_ & ~new_n49914_;
  assign ys__n32809 = ~new_n43951_ & ~new_n49915_;
  assign new_n49917_ = ys__n38118 & new_n43944_;
  assign new_n49918_ = ys__n18738 & ~new_n43948_;
  assign new_n49919_ = ~new_n49917_ & ~new_n49918_;
  assign ys__n32810 = ~new_n43951_ & ~new_n49919_;
  assign new_n49921_ = ys__n38119 & new_n43944_;
  assign new_n49922_ = ys__n18741 & ~new_n43948_;
  assign new_n49923_ = ~new_n49921_ & ~new_n49922_;
  assign ys__n32811 = ~new_n43951_ & ~new_n49923_;
  assign new_n49925_ = ys__n38120 & new_n43944_;
  assign new_n49926_ = ys__n18744 & ~new_n43948_;
  assign new_n49927_ = ~new_n49925_ & ~new_n49926_;
  assign ys__n32812 = ~new_n43951_ & ~new_n49927_;
  assign new_n49929_ = ys__n38121 & new_n43944_;
  assign new_n49930_ = ys__n18747 & ~new_n43948_;
  assign new_n49931_ = ~new_n49929_ & ~new_n49930_;
  assign ys__n32813 = ~new_n43951_ & ~new_n49931_;
  assign new_n49933_ = ys__n48146 & new_n43799_;
  assign new_n49934_ = ys__n18654 & ~new_n43803_;
  assign new_n49935_ = ~new_n49933_ & ~new_n49934_;
  assign ys__n32814 = ~new_n43806_ & ~new_n49935_;
  assign new_n49937_ = ys__n48147 & new_n43799_;
  assign new_n49938_ = ys__n18657 & ~new_n43803_;
  assign new_n49939_ = ~new_n49937_ & ~new_n49938_;
  assign ys__n32815 = ~new_n43806_ & ~new_n49939_;
  assign new_n49941_ = ys__n48148 & new_n43799_;
  assign new_n49942_ = ys__n18660 & ~new_n43803_;
  assign new_n49943_ = ~new_n49941_ & ~new_n49942_;
  assign ys__n32816 = ~new_n43806_ & ~new_n49943_;
  assign new_n49945_ = ys__n48149 & new_n43799_;
  assign new_n49946_ = ys__n18663 & ~new_n43803_;
  assign new_n49947_ = ~new_n49945_ & ~new_n49946_;
  assign ys__n32817 = ~new_n43806_ & ~new_n49947_;
  assign new_n49949_ = ys__n38122 & new_n43799_;
  assign new_n49950_ = ys__n18666 & ~new_n43803_;
  assign new_n49951_ = ~new_n49949_ & ~new_n49950_;
  assign ys__n32818 = ~new_n43806_ & ~new_n49951_;
  assign new_n49953_ = ys__n38123 & new_n43799_;
  assign new_n49954_ = ys__n18669 & ~new_n43803_;
  assign new_n49955_ = ~new_n49953_ & ~new_n49954_;
  assign ys__n32819 = ~new_n43806_ & ~new_n49955_;
  assign new_n49957_ = ys__n38124 & new_n43799_;
  assign new_n49958_ = ys__n18672 & ~new_n43803_;
  assign new_n49959_ = ~new_n49957_ & ~new_n49958_;
  assign ys__n32820 = ~new_n43806_ & ~new_n49959_;
  assign new_n49961_ = ys__n38125 & new_n43799_;
  assign new_n49962_ = ys__n18675 & ~new_n43803_;
  assign new_n49963_ = ~new_n49961_ & ~new_n49962_;
  assign ys__n32821 = ~new_n43806_ & ~new_n49963_;
  assign new_n49965_ = ys__n38126 & new_n43799_;
  assign new_n49966_ = ys__n18678 & ~new_n43803_;
  assign new_n49967_ = ~new_n49965_ & ~new_n49966_;
  assign ys__n32822 = ~new_n43806_ & ~new_n49967_;
  assign new_n49969_ = ys__n38127 & new_n43799_;
  assign new_n49970_ = ys__n18681 & ~new_n43803_;
  assign new_n49971_ = ~new_n49969_ & ~new_n49970_;
  assign ys__n32823 = ~new_n43806_ & ~new_n49971_;
  assign new_n49973_ = ys__n38128 & new_n43799_;
  assign new_n49974_ = ys__n18684 & ~new_n43803_;
  assign new_n49975_ = ~new_n49973_ & ~new_n49974_;
  assign ys__n32824 = ~new_n43806_ & ~new_n49975_;
  assign new_n49977_ = ys__n38129 & new_n43799_;
  assign new_n49978_ = ys__n18687 & ~new_n43803_;
  assign new_n49979_ = ~new_n49977_ & ~new_n49978_;
  assign ys__n32825 = ~new_n43806_ & ~new_n49979_;
  assign new_n49981_ = ys__n38130 & new_n43799_;
  assign new_n49982_ = ys__n18690 & ~new_n43803_;
  assign new_n49983_ = ~new_n49981_ & ~new_n49982_;
  assign ys__n32826 = ~new_n43806_ & ~new_n49983_;
  assign new_n49985_ = ys__n38131 & new_n43799_;
  assign new_n49986_ = ys__n18693 & ~new_n43803_;
  assign new_n49987_ = ~new_n49985_ & ~new_n49986_;
  assign ys__n32827 = ~new_n43806_ & ~new_n49987_;
  assign new_n49989_ = ys__n38132 & new_n43799_;
  assign new_n49990_ = ys__n18696 & ~new_n43803_;
  assign new_n49991_ = ~new_n49989_ & ~new_n49990_;
  assign ys__n32828 = ~new_n43806_ & ~new_n49991_;
  assign new_n49993_ = ys__n38133 & new_n43799_;
  assign new_n49994_ = ys__n18699 & ~new_n43803_;
  assign new_n49995_ = ~new_n49993_ & ~new_n49994_;
  assign ys__n32829 = ~new_n43806_ & ~new_n49995_;
  assign new_n49997_ = ys__n38134 & new_n43799_;
  assign new_n49998_ = ys__n18702 & ~new_n43803_;
  assign new_n49999_ = ~new_n49997_ & ~new_n49998_;
  assign ys__n32830 = ~new_n43806_ & ~new_n49999_;
  assign new_n50001_ = ys__n38135 & new_n43799_;
  assign new_n50002_ = ys__n18705 & ~new_n43803_;
  assign new_n50003_ = ~new_n50001_ & ~new_n50002_;
  assign ys__n32831 = ~new_n43806_ & ~new_n50003_;
  assign new_n50005_ = ys__n38136 & new_n43799_;
  assign new_n50006_ = ys__n18708 & ~new_n43803_;
  assign new_n50007_ = ~new_n50005_ & ~new_n50006_;
  assign ys__n32832 = ~new_n43806_ & ~new_n50007_;
  assign new_n50009_ = ys__n38137 & new_n43799_;
  assign new_n50010_ = ys__n18711 & ~new_n43803_;
  assign new_n50011_ = ~new_n50009_ & ~new_n50010_;
  assign ys__n32833 = ~new_n43806_ & ~new_n50011_;
  assign new_n50013_ = ys__n38138 & new_n43799_;
  assign new_n50014_ = ys__n18714 & ~new_n43803_;
  assign new_n50015_ = ~new_n50013_ & ~new_n50014_;
  assign ys__n32834 = ~new_n43806_ & ~new_n50015_;
  assign new_n50017_ = ys__n38139 & new_n43799_;
  assign new_n50018_ = ys__n18717 & ~new_n43803_;
  assign new_n50019_ = ~new_n50017_ & ~new_n50018_;
  assign ys__n32835 = ~new_n43806_ & ~new_n50019_;
  assign new_n50021_ = ys__n38140 & new_n43799_;
  assign new_n50022_ = ys__n18720 & ~new_n43803_;
  assign new_n50023_ = ~new_n50021_ & ~new_n50022_;
  assign ys__n32836 = ~new_n43806_ & ~new_n50023_;
  assign new_n50025_ = ys__n38141 & new_n43799_;
  assign new_n50026_ = ys__n18723 & ~new_n43803_;
  assign new_n50027_ = ~new_n50025_ & ~new_n50026_;
  assign ys__n32837 = ~new_n43806_ & ~new_n50027_;
  assign new_n50029_ = ys__n38142 & new_n43799_;
  assign new_n50030_ = ys__n18726 & ~new_n43803_;
  assign new_n50031_ = ~new_n50029_ & ~new_n50030_;
  assign ys__n32838 = ~new_n43806_ & ~new_n50031_;
  assign new_n50033_ = ys__n38143 & new_n43799_;
  assign new_n50034_ = ys__n18729 & ~new_n43803_;
  assign new_n50035_ = ~new_n50033_ & ~new_n50034_;
  assign ys__n32839 = ~new_n43806_ & ~new_n50035_;
  assign new_n50037_ = ys__n38144 & new_n43799_;
  assign new_n50038_ = ys__n18732 & ~new_n43803_;
  assign new_n50039_ = ~new_n50037_ & ~new_n50038_;
  assign ys__n32840 = ~new_n43806_ & ~new_n50039_;
  assign new_n50041_ = ys__n38145 & new_n43799_;
  assign new_n50042_ = ys__n18735 & ~new_n43803_;
  assign new_n50043_ = ~new_n50041_ & ~new_n50042_;
  assign ys__n32841 = ~new_n43806_ & ~new_n50043_;
  assign new_n50045_ = ys__n38146 & new_n43799_;
  assign new_n50046_ = ys__n18738 & ~new_n43803_;
  assign new_n50047_ = ~new_n50045_ & ~new_n50046_;
  assign ys__n32842 = ~new_n43806_ & ~new_n50047_;
  assign new_n50049_ = ys__n38147 & new_n43799_;
  assign new_n50050_ = ys__n18741 & ~new_n43803_;
  assign new_n50051_ = ~new_n50049_ & ~new_n50050_;
  assign ys__n32843 = ~new_n43806_ & ~new_n50051_;
  assign new_n50053_ = ys__n38148 & new_n43799_;
  assign new_n50054_ = ys__n18744 & ~new_n43803_;
  assign new_n50055_ = ~new_n50053_ & ~new_n50054_;
  assign ys__n32844 = ~new_n43806_ & ~new_n50055_;
  assign new_n50057_ = ys__n38149 & new_n43799_;
  assign new_n50058_ = ys__n18747 & ~new_n43803_;
  assign new_n50059_ = ~new_n50057_ & ~new_n50058_;
  assign ys__n32845 = ~new_n43806_ & ~new_n50059_;
  assign new_n50061_ = ys__n48150 & new_n43654_;
  assign new_n50062_ = ys__n18654 & ~new_n43658_;
  assign new_n50063_ = ~new_n50061_ & ~new_n50062_;
  assign ys__n32846 = ~new_n43661_ & ~new_n50063_;
  assign new_n50065_ = ys__n48151 & new_n43654_;
  assign new_n50066_ = ys__n18657 & ~new_n43658_;
  assign new_n50067_ = ~new_n50065_ & ~new_n50066_;
  assign ys__n32847 = ~new_n43661_ & ~new_n50067_;
  assign new_n50069_ = ys__n48152 & new_n43654_;
  assign new_n50070_ = ys__n18660 & ~new_n43658_;
  assign new_n50071_ = ~new_n50069_ & ~new_n50070_;
  assign ys__n32848 = ~new_n43661_ & ~new_n50071_;
  assign new_n50073_ = ys__n48153 & new_n43654_;
  assign new_n50074_ = ys__n18663 & ~new_n43658_;
  assign new_n50075_ = ~new_n50073_ & ~new_n50074_;
  assign ys__n32849 = ~new_n43661_ & ~new_n50075_;
  assign new_n50077_ = ys__n38150 & new_n43654_;
  assign new_n50078_ = ys__n18666 & ~new_n43658_;
  assign new_n50079_ = ~new_n50077_ & ~new_n50078_;
  assign ys__n32850 = ~new_n43661_ & ~new_n50079_;
  assign new_n50081_ = ys__n38151 & new_n43654_;
  assign new_n50082_ = ys__n18669 & ~new_n43658_;
  assign new_n50083_ = ~new_n50081_ & ~new_n50082_;
  assign ys__n32851 = ~new_n43661_ & ~new_n50083_;
  assign new_n50085_ = ys__n38152 & new_n43654_;
  assign new_n50086_ = ys__n18672 & ~new_n43658_;
  assign new_n50087_ = ~new_n50085_ & ~new_n50086_;
  assign ys__n32852 = ~new_n43661_ & ~new_n50087_;
  assign new_n50089_ = ys__n38153 & new_n43654_;
  assign new_n50090_ = ys__n18675 & ~new_n43658_;
  assign new_n50091_ = ~new_n50089_ & ~new_n50090_;
  assign ys__n32853 = ~new_n43661_ & ~new_n50091_;
  assign new_n50093_ = ys__n38154 & new_n43654_;
  assign new_n50094_ = ys__n18678 & ~new_n43658_;
  assign new_n50095_ = ~new_n50093_ & ~new_n50094_;
  assign ys__n32854 = ~new_n43661_ & ~new_n50095_;
  assign new_n50097_ = ys__n38155 & new_n43654_;
  assign new_n50098_ = ys__n18681 & ~new_n43658_;
  assign new_n50099_ = ~new_n50097_ & ~new_n50098_;
  assign ys__n32855 = ~new_n43661_ & ~new_n50099_;
  assign new_n50101_ = ys__n38156 & new_n43654_;
  assign new_n50102_ = ys__n18684 & ~new_n43658_;
  assign new_n50103_ = ~new_n50101_ & ~new_n50102_;
  assign ys__n32856 = ~new_n43661_ & ~new_n50103_;
  assign new_n50105_ = ys__n38157 & new_n43654_;
  assign new_n50106_ = ys__n18687 & ~new_n43658_;
  assign new_n50107_ = ~new_n50105_ & ~new_n50106_;
  assign ys__n32857 = ~new_n43661_ & ~new_n50107_;
  assign new_n50109_ = ys__n38158 & new_n43654_;
  assign new_n50110_ = ys__n18690 & ~new_n43658_;
  assign new_n50111_ = ~new_n50109_ & ~new_n50110_;
  assign ys__n32858 = ~new_n43661_ & ~new_n50111_;
  assign new_n50113_ = ys__n38159 & new_n43654_;
  assign new_n50114_ = ys__n18693 & ~new_n43658_;
  assign new_n50115_ = ~new_n50113_ & ~new_n50114_;
  assign ys__n32859 = ~new_n43661_ & ~new_n50115_;
  assign new_n50117_ = ys__n38160 & new_n43654_;
  assign new_n50118_ = ys__n18696 & ~new_n43658_;
  assign new_n50119_ = ~new_n50117_ & ~new_n50118_;
  assign ys__n32860 = ~new_n43661_ & ~new_n50119_;
  assign new_n50121_ = ys__n38161 & new_n43654_;
  assign new_n50122_ = ys__n18699 & ~new_n43658_;
  assign new_n50123_ = ~new_n50121_ & ~new_n50122_;
  assign ys__n32861 = ~new_n43661_ & ~new_n50123_;
  assign new_n50125_ = ys__n38162 & new_n43654_;
  assign new_n50126_ = ys__n18702 & ~new_n43658_;
  assign new_n50127_ = ~new_n50125_ & ~new_n50126_;
  assign ys__n32862 = ~new_n43661_ & ~new_n50127_;
  assign new_n50129_ = ys__n38163 & new_n43654_;
  assign new_n50130_ = ys__n18705 & ~new_n43658_;
  assign new_n50131_ = ~new_n50129_ & ~new_n50130_;
  assign ys__n32863 = ~new_n43661_ & ~new_n50131_;
  assign new_n50133_ = ys__n38164 & new_n43654_;
  assign new_n50134_ = ys__n18708 & ~new_n43658_;
  assign new_n50135_ = ~new_n50133_ & ~new_n50134_;
  assign ys__n32864 = ~new_n43661_ & ~new_n50135_;
  assign new_n50137_ = ys__n38165 & new_n43654_;
  assign new_n50138_ = ys__n18711 & ~new_n43658_;
  assign new_n50139_ = ~new_n50137_ & ~new_n50138_;
  assign ys__n32865 = ~new_n43661_ & ~new_n50139_;
  assign new_n50141_ = ys__n38166 & new_n43654_;
  assign new_n50142_ = ys__n18714 & ~new_n43658_;
  assign new_n50143_ = ~new_n50141_ & ~new_n50142_;
  assign ys__n32866 = ~new_n43661_ & ~new_n50143_;
  assign new_n50145_ = ys__n38167 & new_n43654_;
  assign new_n50146_ = ys__n18717 & ~new_n43658_;
  assign new_n50147_ = ~new_n50145_ & ~new_n50146_;
  assign ys__n32867 = ~new_n43661_ & ~new_n50147_;
  assign new_n50149_ = ys__n38168 & new_n43654_;
  assign new_n50150_ = ys__n18720 & ~new_n43658_;
  assign new_n50151_ = ~new_n50149_ & ~new_n50150_;
  assign ys__n32868 = ~new_n43661_ & ~new_n50151_;
  assign new_n50153_ = ys__n38169 & new_n43654_;
  assign new_n50154_ = ys__n18723 & ~new_n43658_;
  assign new_n50155_ = ~new_n50153_ & ~new_n50154_;
  assign ys__n32869 = ~new_n43661_ & ~new_n50155_;
  assign new_n50157_ = ys__n38170 & new_n43654_;
  assign new_n50158_ = ys__n18726 & ~new_n43658_;
  assign new_n50159_ = ~new_n50157_ & ~new_n50158_;
  assign ys__n32870 = ~new_n43661_ & ~new_n50159_;
  assign new_n50161_ = ys__n38171 & new_n43654_;
  assign new_n50162_ = ys__n18729 & ~new_n43658_;
  assign new_n50163_ = ~new_n50161_ & ~new_n50162_;
  assign ys__n32871 = ~new_n43661_ & ~new_n50163_;
  assign new_n50165_ = ys__n38172 & new_n43654_;
  assign new_n50166_ = ys__n18732 & ~new_n43658_;
  assign new_n50167_ = ~new_n50165_ & ~new_n50166_;
  assign ys__n32872 = ~new_n43661_ & ~new_n50167_;
  assign new_n50169_ = ys__n38173 & new_n43654_;
  assign new_n50170_ = ys__n18735 & ~new_n43658_;
  assign new_n50171_ = ~new_n50169_ & ~new_n50170_;
  assign ys__n32873 = ~new_n43661_ & ~new_n50171_;
  assign new_n50173_ = ys__n38174 & new_n43654_;
  assign new_n50174_ = ys__n18738 & ~new_n43658_;
  assign new_n50175_ = ~new_n50173_ & ~new_n50174_;
  assign ys__n32874 = ~new_n43661_ & ~new_n50175_;
  assign new_n50177_ = ys__n38175 & new_n43654_;
  assign new_n50178_ = ys__n18741 & ~new_n43658_;
  assign new_n50179_ = ~new_n50177_ & ~new_n50178_;
  assign ys__n32875 = ~new_n43661_ & ~new_n50179_;
  assign new_n50181_ = ys__n38176 & new_n43654_;
  assign new_n50182_ = ys__n18744 & ~new_n43658_;
  assign new_n50183_ = ~new_n50181_ & ~new_n50182_;
  assign ys__n32876 = ~new_n43661_ & ~new_n50183_;
  assign new_n50185_ = ys__n38177 & new_n43654_;
  assign new_n50186_ = ys__n18747 & ~new_n43658_;
  assign new_n50187_ = ~new_n50185_ & ~new_n50186_;
  assign ys__n32877 = ~new_n43661_ & ~new_n50187_;
  assign new_n50189_ = ys__n37757 & new_n48254_;
  assign new_n50190_ = ys__n18759 & ~new_n48258_;
  assign new_n50191_ = ~new_n50189_ & ~new_n50190_;
  assign ys__n32878 = ~new_n48261_ & ~new_n50191_;
  assign new_n50193_ = ys__n37756 & new_n48387_;
  assign new_n50194_ = ys__n18759 & ~new_n48391_;
  assign new_n50195_ = ~new_n50193_ & ~new_n50194_;
  assign ys__n32879 = ~new_n48394_ & ~new_n50195_;
  assign new_n50197_ = ys__n37755 & new_n48520_;
  assign new_n50198_ = ys__n18759 & ~new_n48524_;
  assign new_n50199_ = ~new_n50197_ & ~new_n50198_;
  assign ys__n32880 = ~new_n48527_ & ~new_n50199_;
  assign new_n50201_ = ys__n37754 & new_n45366_;
  assign new_n50202_ = ys__n18759 & ~new_n45370_;
  assign new_n50203_ = ~new_n50201_ & ~new_n50202_;
  assign ys__n32881 = ~new_n45373_ & ~new_n50203_;
  assign new_n50205_ = ys__n37753 & new_n45221_;
  assign new_n50206_ = ys__n18759 & ~new_n45225_;
  assign new_n50207_ = ~new_n50205_ & ~new_n50206_;
  assign ys__n32882 = ~new_n45228_ & ~new_n50207_;
  assign new_n50209_ = ys__n37752 & new_n45076_;
  assign new_n50210_ = ys__n18759 & ~new_n45080_;
  assign new_n50211_ = ~new_n50209_ & ~new_n50210_;
  assign ys__n32883 = ~new_n45083_ & ~new_n50211_;
  assign new_n50213_ = ys__n37751 & new_n44931_;
  assign new_n50214_ = ys__n18759 & ~new_n44935_;
  assign new_n50215_ = ~new_n50213_ & ~new_n50214_;
  assign ys__n32884 = ~new_n44938_ & ~new_n50215_;
  assign new_n50217_ = ys__n37750 & new_n44786_;
  assign new_n50218_ = ys__n18759 & ~new_n44790_;
  assign new_n50219_ = ~new_n50217_ & ~new_n50218_;
  assign ys__n32885 = ~new_n44793_ & ~new_n50219_;
  assign new_n50221_ = ys__n37749 & new_n44641_;
  assign new_n50222_ = ys__n18759 & ~new_n44645_;
  assign new_n50223_ = ~new_n50221_ & ~new_n50222_;
  assign ys__n32886 = ~new_n44648_ & ~new_n50223_;
  assign new_n50225_ = ys__n37748 & new_n44317_;
  assign new_n50226_ = ys__n18759 & ~new_n44321_;
  assign new_n50227_ = ~new_n50225_ & ~new_n50226_;
  assign ys__n32887 = ~new_n44324_ & ~new_n50227_;
  assign new_n50229_ = ys__n37747 & new_n44462_;
  assign new_n50230_ = ys__n18759 & ~new_n44466_;
  assign new_n50231_ = ~new_n50229_ & ~new_n50230_;
  assign ys__n32888 = ~new_n44469_ & ~new_n50231_;
  assign new_n50233_ = ys__n37746 & new_n44172_;
  assign new_n50234_ = ys__n18759 & ~new_n44176_;
  assign new_n50235_ = ~new_n50233_ & ~new_n50234_;
  assign ys__n32889 = ~new_n44179_ & ~new_n50235_;
  assign new_n50237_ = ys__n37745 & new_n43944_;
  assign new_n50238_ = ys__n18759 & ~new_n43948_;
  assign new_n50239_ = ~new_n50237_ & ~new_n50238_;
  assign ys__n32890 = ~new_n43951_ & ~new_n50239_;
  assign new_n50241_ = ys__n37744 & new_n43799_;
  assign new_n50242_ = ys__n18759 & ~new_n43803_;
  assign new_n50243_ = ~new_n50241_ & ~new_n50242_;
  assign ys__n32891 = ~new_n43806_ & ~new_n50243_;
  assign new_n50245_ = ys__n37743 & new_n43654_;
  assign new_n50246_ = ys__n18759 & ~new_n43658_;
  assign new_n50247_ = ~new_n50245_ & ~new_n50246_;
  assign ys__n32892 = ~new_n43661_ & ~new_n50247_;
  assign new_n50249_ = ys__n48154 & new_n48254_;
  assign new_n50250_ = ys__n47202 & ~new_n48258_;
  assign new_n50251_ = ~new_n50249_ & ~new_n50250_;
  assign ys__n32893 = ~new_n48261_ & ~new_n50251_;
  assign new_n50253_ = ys__n48155 & new_n48254_;
  assign new_n50254_ = ys__n47203 & ~new_n48258_;
  assign new_n50255_ = ~new_n50253_ & ~new_n50254_;
  assign ys__n32894 = ~new_n48261_ & ~new_n50255_;
  assign new_n50257_ = ys__n48156 & new_n48254_;
  assign new_n50258_ = ys__n47204 & ~new_n48258_;
  assign new_n50259_ = ~new_n50257_ & ~new_n50258_;
  assign ys__n32895 = ~new_n48261_ & ~new_n50259_;
  assign new_n50261_ = ys__n48157 & new_n48254_;
  assign new_n50262_ = ys__n47205 & ~new_n48258_;
  assign new_n50263_ = ~new_n50261_ & ~new_n50262_;
  assign ys__n32896 = ~new_n48261_ & ~new_n50263_;
  assign new_n50265_ = ys__n48158 & new_n48254_;
  assign new_n50266_ = ys__n47206 & ~new_n48258_;
  assign new_n50267_ = ~new_n50265_ & ~new_n50266_;
  assign ys__n32897 = ~new_n48261_ & ~new_n50267_;
  assign new_n50269_ = ys__n48159 & new_n48254_;
  assign new_n50270_ = ys__n47207 & ~new_n48258_;
  assign new_n50271_ = ~new_n50269_ & ~new_n50270_;
  assign ys__n32898 = ~new_n48261_ & ~new_n50271_;
  assign new_n50273_ = ys__n48160 & new_n48254_;
  assign new_n50274_ = ys__n47208 & ~new_n48258_;
  assign new_n50275_ = ~new_n50273_ & ~new_n50274_;
  assign ys__n32899 = ~new_n48261_ & ~new_n50275_;
  assign new_n50277_ = ys__n48161 & new_n48254_;
  assign new_n50278_ = ys__n47209 & ~new_n48258_;
  assign new_n50279_ = ~new_n50277_ & ~new_n50278_;
  assign ys__n32900 = ~new_n48261_ & ~new_n50279_;
  assign new_n50281_ = ys__n48162 & new_n48254_;
  assign new_n50282_ = ys__n47210 & ~new_n48258_;
  assign new_n50283_ = ~new_n50281_ & ~new_n50282_;
  assign ys__n32901 = ~new_n48261_ & ~new_n50283_;
  assign new_n50285_ = ys__n48163 & new_n48254_;
  assign new_n50286_ = ys__n47211 & ~new_n48258_;
  assign new_n50287_ = ~new_n50285_ & ~new_n50286_;
  assign ys__n32902 = ~new_n48261_ & ~new_n50287_;
  assign new_n50289_ = ys__n48164 & new_n48254_;
  assign new_n50290_ = ys__n47212 & ~new_n48258_;
  assign new_n50291_ = ~new_n50289_ & ~new_n50290_;
  assign ys__n32903 = ~new_n48261_ & ~new_n50291_;
  assign new_n50293_ = ys__n48165 & new_n48254_;
  assign new_n50294_ = ys__n47213 & ~new_n48258_;
  assign new_n50295_ = ~new_n50293_ & ~new_n50294_;
  assign ys__n32904 = ~new_n48261_ & ~new_n50295_;
  assign new_n50297_ = ys__n48166 & new_n48254_;
  assign new_n50298_ = ys__n47214 & ~new_n48258_;
  assign new_n50299_ = ~new_n50297_ & ~new_n50298_;
  assign ys__n32905 = ~new_n48261_ & ~new_n50299_;
  assign new_n50301_ = ys__n48167 & new_n48254_;
  assign new_n50302_ = ys__n47215 & ~new_n48258_;
  assign new_n50303_ = ~new_n50301_ & ~new_n50302_;
  assign ys__n32906 = ~new_n48261_ & ~new_n50303_;
  assign new_n50305_ = ys__n48168 & new_n48254_;
  assign new_n50306_ = ys__n47216 & ~new_n48258_;
  assign new_n50307_ = ~new_n50305_ & ~new_n50306_;
  assign ys__n32907 = ~new_n48261_ & ~new_n50307_;
  assign new_n50309_ = ys__n48169 & new_n48254_;
  assign new_n50310_ = ys__n47217 & ~new_n48258_;
  assign new_n50311_ = ~new_n50309_ & ~new_n50310_;
  assign ys__n32908 = ~new_n48261_ & ~new_n50311_;
  assign new_n50313_ = ys__n48170 & new_n48254_;
  assign new_n50314_ = ys__n47218 & ~new_n48258_;
  assign new_n50315_ = ~new_n50313_ & ~new_n50314_;
  assign ys__n32909 = ~new_n48261_ & ~new_n50315_;
  assign new_n50317_ = ys__n48171 & new_n48254_;
  assign new_n50318_ = ys__n47219 & ~new_n48258_;
  assign new_n50319_ = ~new_n50317_ & ~new_n50318_;
  assign ys__n32910 = ~new_n48261_ & ~new_n50319_;
  assign new_n50321_ = ys__n48172 & new_n48254_;
  assign new_n50322_ = ys__n47220 & ~new_n48258_;
  assign new_n50323_ = ~new_n50321_ & ~new_n50322_;
  assign ys__n32911 = ~new_n48261_ & ~new_n50323_;
  assign new_n50325_ = ys__n48173 & new_n48254_;
  assign new_n50326_ = ys__n47221 & ~new_n48258_;
  assign new_n50327_ = ~new_n50325_ & ~new_n50326_;
  assign ys__n32912 = ~new_n48261_ & ~new_n50327_;
  assign new_n50329_ = ys__n48174 & new_n48254_;
  assign new_n50330_ = ys__n47222 & ~new_n48258_;
  assign new_n50331_ = ~new_n50329_ & ~new_n50330_;
  assign ys__n32913 = ~new_n48261_ & ~new_n50331_;
  assign new_n50333_ = ys__n48175 & new_n48254_;
  assign new_n50334_ = ys__n47223 & ~new_n48258_;
  assign new_n50335_ = ~new_n50333_ & ~new_n50334_;
  assign ys__n32914 = ~new_n48261_ & ~new_n50335_;
  assign new_n50337_ = ys__n48176 & new_n48254_;
  assign new_n50338_ = ys__n47224 & ~new_n48258_;
  assign new_n50339_ = ~new_n50337_ & ~new_n50338_;
  assign ys__n32915 = ~new_n48261_ & ~new_n50339_;
  assign new_n50341_ = ys__n48177 & new_n48254_;
  assign new_n50342_ = ys__n47225 & ~new_n48258_;
  assign new_n50343_ = ~new_n50341_ & ~new_n50342_;
  assign ys__n32916 = ~new_n48261_ & ~new_n50343_;
  assign new_n50345_ = ys__n48178 & new_n48254_;
  assign new_n50346_ = ys__n47226 & ~new_n48258_;
  assign new_n50347_ = ~new_n50345_ & ~new_n50346_;
  assign ys__n32917 = ~new_n48261_ & ~new_n50347_;
  assign new_n50349_ = ys__n48179 & new_n48254_;
  assign new_n50350_ = ys__n47227 & ~new_n48258_;
  assign new_n50351_ = ~new_n50349_ & ~new_n50350_;
  assign ys__n32918 = ~new_n48261_ & ~new_n50351_;
  assign new_n50353_ = ys__n48180 & new_n48254_;
  assign new_n50354_ = ys__n47228 & ~new_n48258_;
  assign new_n50355_ = ~new_n50353_ & ~new_n50354_;
  assign ys__n32919 = ~new_n48261_ & ~new_n50355_;
  assign new_n50357_ = ys__n48181 & new_n48254_;
  assign new_n50358_ = ys__n47229 & ~new_n48258_;
  assign new_n50359_ = ~new_n50357_ & ~new_n50358_;
  assign ys__n32920 = ~new_n48261_ & ~new_n50359_;
  assign new_n50361_ = ys__n48182 & new_n48254_;
  assign new_n50362_ = ys__n47230 & ~new_n48258_;
  assign new_n50363_ = ~new_n50361_ & ~new_n50362_;
  assign ys__n32921 = ~new_n48261_ & ~new_n50363_;
  assign new_n50365_ = ys__n48183 & new_n48254_;
  assign new_n50366_ = ys__n47231 & ~new_n48258_;
  assign new_n50367_ = ~new_n50365_ & ~new_n50366_;
  assign ys__n32922 = ~new_n48261_ & ~new_n50367_;
  assign new_n50369_ = ys__n48184 & new_n48254_;
  assign new_n50370_ = ys__n47232 & ~new_n48258_;
  assign new_n50371_ = ~new_n50369_ & ~new_n50370_;
  assign ys__n32923 = ~new_n48261_ & ~new_n50371_;
  assign new_n50373_ = ys__n48185 & new_n48254_;
  assign new_n50374_ = ys__n47233 & ~new_n48258_;
  assign new_n50375_ = ~new_n50373_ & ~new_n50374_;
  assign ys__n32924 = ~new_n48261_ & ~new_n50375_;
  assign new_n50377_ = ys__n48186 & new_n48254_;
  assign new_n50378_ = ys__n18762 & ~new_n48258_;
  assign new_n50379_ = ~new_n50377_ & ~new_n50378_;
  assign ys__n32925 = ~new_n48261_ & ~new_n50379_;
  assign new_n50381_ = ys__n48187 & new_n48254_;
  assign new_n50382_ = ys__n18750 & ~new_n48258_;
  assign new_n50383_ = ~new_n50381_ & ~new_n50382_;
  assign ys__n32926 = ~new_n48261_ & ~new_n50383_;
  assign new_n50385_ = ys__n48188 & new_n48254_;
  assign new_n50386_ = ys__n18753 & ~new_n48258_;
  assign new_n50387_ = ~new_n50385_ & ~new_n50386_;
  assign ys__n32927 = ~new_n48261_ & ~new_n50387_;
  assign new_n50389_ = ys__n48189 & new_n48387_;
  assign new_n50390_ = ys__n47202 & ~new_n48391_;
  assign new_n50391_ = ~new_n50389_ & ~new_n50390_;
  assign ys__n32928 = ~new_n48394_ & ~new_n50391_;
  assign new_n50393_ = ys__n48190 & new_n48387_;
  assign new_n50394_ = ys__n47203 & ~new_n48391_;
  assign new_n50395_ = ~new_n50393_ & ~new_n50394_;
  assign ys__n32929 = ~new_n48394_ & ~new_n50395_;
  assign new_n50397_ = ys__n48191 & new_n48387_;
  assign new_n50398_ = ys__n47204 & ~new_n48391_;
  assign new_n50399_ = ~new_n50397_ & ~new_n50398_;
  assign ys__n32930 = ~new_n48394_ & ~new_n50399_;
  assign new_n50401_ = ys__n48192 & new_n48387_;
  assign new_n50402_ = ys__n47205 & ~new_n48391_;
  assign new_n50403_ = ~new_n50401_ & ~new_n50402_;
  assign ys__n32931 = ~new_n48394_ & ~new_n50403_;
  assign new_n50405_ = ys__n48193 & new_n48387_;
  assign new_n50406_ = ys__n47206 & ~new_n48391_;
  assign new_n50407_ = ~new_n50405_ & ~new_n50406_;
  assign ys__n32932 = ~new_n48394_ & ~new_n50407_;
  assign new_n50409_ = ys__n48194 & new_n48387_;
  assign new_n50410_ = ys__n47207 & ~new_n48391_;
  assign new_n50411_ = ~new_n50409_ & ~new_n50410_;
  assign ys__n32933 = ~new_n48394_ & ~new_n50411_;
  assign new_n50413_ = ys__n48195 & new_n48387_;
  assign new_n50414_ = ys__n47208 & ~new_n48391_;
  assign new_n50415_ = ~new_n50413_ & ~new_n50414_;
  assign ys__n32934 = ~new_n48394_ & ~new_n50415_;
  assign new_n50417_ = ys__n48196 & new_n48387_;
  assign new_n50418_ = ys__n47209 & ~new_n48391_;
  assign new_n50419_ = ~new_n50417_ & ~new_n50418_;
  assign ys__n32935 = ~new_n48394_ & ~new_n50419_;
  assign new_n50421_ = ys__n48197 & new_n48387_;
  assign new_n50422_ = ys__n47210 & ~new_n48391_;
  assign new_n50423_ = ~new_n50421_ & ~new_n50422_;
  assign ys__n32936 = ~new_n48394_ & ~new_n50423_;
  assign new_n50425_ = ys__n48198 & new_n48387_;
  assign new_n50426_ = ys__n47211 & ~new_n48391_;
  assign new_n50427_ = ~new_n50425_ & ~new_n50426_;
  assign ys__n32937 = ~new_n48394_ & ~new_n50427_;
  assign new_n50429_ = ys__n48199 & new_n48387_;
  assign new_n50430_ = ys__n47212 & ~new_n48391_;
  assign new_n50431_ = ~new_n50429_ & ~new_n50430_;
  assign ys__n32938 = ~new_n48394_ & ~new_n50431_;
  assign new_n50433_ = ys__n48200 & new_n48387_;
  assign new_n50434_ = ys__n47213 & ~new_n48391_;
  assign new_n50435_ = ~new_n50433_ & ~new_n50434_;
  assign ys__n32939 = ~new_n48394_ & ~new_n50435_;
  assign new_n50437_ = ys__n48201 & new_n48387_;
  assign new_n50438_ = ys__n47214 & ~new_n48391_;
  assign new_n50439_ = ~new_n50437_ & ~new_n50438_;
  assign ys__n32940 = ~new_n48394_ & ~new_n50439_;
  assign new_n50441_ = ys__n48202 & new_n48387_;
  assign new_n50442_ = ys__n47215 & ~new_n48391_;
  assign new_n50443_ = ~new_n50441_ & ~new_n50442_;
  assign ys__n32941 = ~new_n48394_ & ~new_n50443_;
  assign new_n50445_ = ys__n48203 & new_n48387_;
  assign new_n50446_ = ys__n47216 & ~new_n48391_;
  assign new_n50447_ = ~new_n50445_ & ~new_n50446_;
  assign ys__n32942 = ~new_n48394_ & ~new_n50447_;
  assign new_n50449_ = ys__n48204 & new_n48387_;
  assign new_n50450_ = ys__n47217 & ~new_n48391_;
  assign new_n50451_ = ~new_n50449_ & ~new_n50450_;
  assign ys__n32943 = ~new_n48394_ & ~new_n50451_;
  assign new_n50453_ = ys__n48205 & new_n48387_;
  assign new_n50454_ = ys__n47218 & ~new_n48391_;
  assign new_n50455_ = ~new_n50453_ & ~new_n50454_;
  assign ys__n32944 = ~new_n48394_ & ~new_n50455_;
  assign new_n50457_ = ys__n48206 & new_n48387_;
  assign new_n50458_ = ys__n47219 & ~new_n48391_;
  assign new_n50459_ = ~new_n50457_ & ~new_n50458_;
  assign ys__n32945 = ~new_n48394_ & ~new_n50459_;
  assign new_n50461_ = ys__n48207 & new_n48387_;
  assign new_n50462_ = ys__n47220 & ~new_n48391_;
  assign new_n50463_ = ~new_n50461_ & ~new_n50462_;
  assign ys__n32946 = ~new_n48394_ & ~new_n50463_;
  assign new_n50465_ = ys__n48208 & new_n48387_;
  assign new_n50466_ = ys__n47221 & ~new_n48391_;
  assign new_n50467_ = ~new_n50465_ & ~new_n50466_;
  assign ys__n32947 = ~new_n48394_ & ~new_n50467_;
  assign new_n50469_ = ys__n48209 & new_n48387_;
  assign new_n50470_ = ys__n47222 & ~new_n48391_;
  assign new_n50471_ = ~new_n50469_ & ~new_n50470_;
  assign ys__n32948 = ~new_n48394_ & ~new_n50471_;
  assign new_n50473_ = ys__n48210 & new_n48387_;
  assign new_n50474_ = ys__n47223 & ~new_n48391_;
  assign new_n50475_ = ~new_n50473_ & ~new_n50474_;
  assign ys__n32949 = ~new_n48394_ & ~new_n50475_;
  assign new_n50477_ = ys__n48211 & new_n48387_;
  assign new_n50478_ = ys__n47224 & ~new_n48391_;
  assign new_n50479_ = ~new_n50477_ & ~new_n50478_;
  assign ys__n32950 = ~new_n48394_ & ~new_n50479_;
  assign new_n50481_ = ys__n48212 & new_n48387_;
  assign new_n50482_ = ys__n47225 & ~new_n48391_;
  assign new_n50483_ = ~new_n50481_ & ~new_n50482_;
  assign ys__n32951 = ~new_n48394_ & ~new_n50483_;
  assign new_n50485_ = ys__n48213 & new_n48387_;
  assign new_n50486_ = ys__n47226 & ~new_n48391_;
  assign new_n50487_ = ~new_n50485_ & ~new_n50486_;
  assign ys__n32952 = ~new_n48394_ & ~new_n50487_;
  assign new_n50489_ = ys__n48214 & new_n48387_;
  assign new_n50490_ = ys__n47227 & ~new_n48391_;
  assign new_n50491_ = ~new_n50489_ & ~new_n50490_;
  assign ys__n32953 = ~new_n48394_ & ~new_n50491_;
  assign new_n50493_ = ys__n48215 & new_n48387_;
  assign new_n50494_ = ys__n47228 & ~new_n48391_;
  assign new_n50495_ = ~new_n50493_ & ~new_n50494_;
  assign ys__n32954 = ~new_n48394_ & ~new_n50495_;
  assign new_n50497_ = ys__n48216 & new_n48387_;
  assign new_n50498_ = ys__n47229 & ~new_n48391_;
  assign new_n50499_ = ~new_n50497_ & ~new_n50498_;
  assign ys__n32955 = ~new_n48394_ & ~new_n50499_;
  assign new_n50501_ = ys__n48217 & new_n48387_;
  assign new_n50502_ = ys__n47230 & ~new_n48391_;
  assign new_n50503_ = ~new_n50501_ & ~new_n50502_;
  assign ys__n32956 = ~new_n48394_ & ~new_n50503_;
  assign new_n50505_ = ys__n48218 & new_n48387_;
  assign new_n50506_ = ys__n47231 & ~new_n48391_;
  assign new_n50507_ = ~new_n50505_ & ~new_n50506_;
  assign ys__n32957 = ~new_n48394_ & ~new_n50507_;
  assign new_n50509_ = ys__n48219 & new_n48387_;
  assign new_n50510_ = ys__n47232 & ~new_n48391_;
  assign new_n50511_ = ~new_n50509_ & ~new_n50510_;
  assign ys__n32958 = ~new_n48394_ & ~new_n50511_;
  assign new_n50513_ = ys__n48220 & new_n48387_;
  assign new_n50514_ = ys__n47233 & ~new_n48391_;
  assign new_n50515_ = ~new_n50513_ & ~new_n50514_;
  assign ys__n32959 = ~new_n48394_ & ~new_n50515_;
  assign new_n50517_ = ys__n48221 & new_n48387_;
  assign new_n50518_ = ys__n18762 & ~new_n48391_;
  assign new_n50519_ = ~new_n50517_ & ~new_n50518_;
  assign ys__n32960 = ~new_n48394_ & ~new_n50519_;
  assign new_n50521_ = ys__n48222 & new_n48387_;
  assign new_n50522_ = ys__n18750 & ~new_n48391_;
  assign new_n50523_ = ~new_n50521_ & ~new_n50522_;
  assign ys__n32961 = ~new_n48394_ & ~new_n50523_;
  assign new_n50525_ = ys__n48223 & new_n48387_;
  assign new_n50526_ = ys__n18753 & ~new_n48391_;
  assign new_n50527_ = ~new_n50525_ & ~new_n50526_;
  assign ys__n32962 = ~new_n48394_ & ~new_n50527_;
  assign new_n50529_ = ys__n48224 & new_n48520_;
  assign new_n50530_ = ys__n47202 & ~new_n48524_;
  assign new_n50531_ = ~new_n50529_ & ~new_n50530_;
  assign ys__n32963 = ~new_n48527_ & ~new_n50531_;
  assign new_n50533_ = ys__n48225 & new_n48520_;
  assign new_n50534_ = ys__n47203 & ~new_n48524_;
  assign new_n50535_ = ~new_n50533_ & ~new_n50534_;
  assign ys__n32964 = ~new_n48527_ & ~new_n50535_;
  assign new_n50537_ = ys__n48226 & new_n48520_;
  assign new_n50538_ = ys__n47204 & ~new_n48524_;
  assign new_n50539_ = ~new_n50537_ & ~new_n50538_;
  assign ys__n32965 = ~new_n48527_ & ~new_n50539_;
  assign new_n50541_ = ys__n48227 & new_n48520_;
  assign new_n50542_ = ys__n47205 & ~new_n48524_;
  assign new_n50543_ = ~new_n50541_ & ~new_n50542_;
  assign ys__n32966 = ~new_n48527_ & ~new_n50543_;
  assign new_n50545_ = ys__n48228 & new_n48520_;
  assign new_n50546_ = ys__n47206 & ~new_n48524_;
  assign new_n50547_ = ~new_n50545_ & ~new_n50546_;
  assign ys__n32967 = ~new_n48527_ & ~new_n50547_;
  assign new_n50549_ = ys__n48229 & new_n48520_;
  assign new_n50550_ = ys__n47207 & ~new_n48524_;
  assign new_n50551_ = ~new_n50549_ & ~new_n50550_;
  assign ys__n32968 = ~new_n48527_ & ~new_n50551_;
  assign new_n50553_ = ys__n48230 & new_n48520_;
  assign new_n50554_ = ys__n47208 & ~new_n48524_;
  assign new_n50555_ = ~new_n50553_ & ~new_n50554_;
  assign ys__n32969 = ~new_n48527_ & ~new_n50555_;
  assign new_n50557_ = ys__n48231 & new_n48520_;
  assign new_n50558_ = ys__n47209 & ~new_n48524_;
  assign new_n50559_ = ~new_n50557_ & ~new_n50558_;
  assign ys__n32970 = ~new_n48527_ & ~new_n50559_;
  assign new_n50561_ = ys__n48232 & new_n48520_;
  assign new_n50562_ = ys__n47210 & ~new_n48524_;
  assign new_n50563_ = ~new_n50561_ & ~new_n50562_;
  assign ys__n32971 = ~new_n48527_ & ~new_n50563_;
  assign new_n50565_ = ys__n48233 & new_n48520_;
  assign new_n50566_ = ys__n47211 & ~new_n48524_;
  assign new_n50567_ = ~new_n50565_ & ~new_n50566_;
  assign ys__n32972 = ~new_n48527_ & ~new_n50567_;
  assign new_n50569_ = ys__n48234 & new_n48520_;
  assign new_n50570_ = ys__n47212 & ~new_n48524_;
  assign new_n50571_ = ~new_n50569_ & ~new_n50570_;
  assign ys__n32973 = ~new_n48527_ & ~new_n50571_;
  assign new_n50573_ = ys__n48235 & new_n48520_;
  assign new_n50574_ = ys__n47213 & ~new_n48524_;
  assign new_n50575_ = ~new_n50573_ & ~new_n50574_;
  assign ys__n32974 = ~new_n48527_ & ~new_n50575_;
  assign new_n50577_ = ys__n48236 & new_n48520_;
  assign new_n50578_ = ys__n47214 & ~new_n48524_;
  assign new_n50579_ = ~new_n50577_ & ~new_n50578_;
  assign ys__n32975 = ~new_n48527_ & ~new_n50579_;
  assign new_n50581_ = ys__n48237 & new_n48520_;
  assign new_n50582_ = ys__n47215 & ~new_n48524_;
  assign new_n50583_ = ~new_n50581_ & ~new_n50582_;
  assign ys__n32976 = ~new_n48527_ & ~new_n50583_;
  assign new_n50585_ = ys__n48238 & new_n48520_;
  assign new_n50586_ = ys__n47216 & ~new_n48524_;
  assign new_n50587_ = ~new_n50585_ & ~new_n50586_;
  assign ys__n32977 = ~new_n48527_ & ~new_n50587_;
  assign new_n50589_ = ys__n48239 & new_n48520_;
  assign new_n50590_ = ys__n47217 & ~new_n48524_;
  assign new_n50591_ = ~new_n50589_ & ~new_n50590_;
  assign ys__n32978 = ~new_n48527_ & ~new_n50591_;
  assign new_n50593_ = ys__n48240 & new_n48520_;
  assign new_n50594_ = ys__n47218 & ~new_n48524_;
  assign new_n50595_ = ~new_n50593_ & ~new_n50594_;
  assign ys__n32979 = ~new_n48527_ & ~new_n50595_;
  assign new_n50597_ = ys__n48241 & new_n48520_;
  assign new_n50598_ = ys__n47219 & ~new_n48524_;
  assign new_n50599_ = ~new_n50597_ & ~new_n50598_;
  assign ys__n32980 = ~new_n48527_ & ~new_n50599_;
  assign new_n50601_ = ys__n48242 & new_n48520_;
  assign new_n50602_ = ys__n47220 & ~new_n48524_;
  assign new_n50603_ = ~new_n50601_ & ~new_n50602_;
  assign ys__n32981 = ~new_n48527_ & ~new_n50603_;
  assign new_n50605_ = ys__n48243 & new_n48520_;
  assign new_n50606_ = ys__n47221 & ~new_n48524_;
  assign new_n50607_ = ~new_n50605_ & ~new_n50606_;
  assign ys__n32982 = ~new_n48527_ & ~new_n50607_;
  assign new_n50609_ = ys__n48244 & new_n48520_;
  assign new_n50610_ = ys__n47222 & ~new_n48524_;
  assign new_n50611_ = ~new_n50609_ & ~new_n50610_;
  assign ys__n32983 = ~new_n48527_ & ~new_n50611_;
  assign new_n50613_ = ys__n48245 & new_n48520_;
  assign new_n50614_ = ys__n47223 & ~new_n48524_;
  assign new_n50615_ = ~new_n50613_ & ~new_n50614_;
  assign ys__n32984 = ~new_n48527_ & ~new_n50615_;
  assign new_n50617_ = ys__n48246 & new_n48520_;
  assign new_n50618_ = ys__n47224 & ~new_n48524_;
  assign new_n50619_ = ~new_n50617_ & ~new_n50618_;
  assign ys__n32985 = ~new_n48527_ & ~new_n50619_;
  assign new_n50621_ = ys__n48247 & new_n48520_;
  assign new_n50622_ = ys__n47225 & ~new_n48524_;
  assign new_n50623_ = ~new_n50621_ & ~new_n50622_;
  assign ys__n32986 = ~new_n48527_ & ~new_n50623_;
  assign new_n50625_ = ys__n48248 & new_n48520_;
  assign new_n50626_ = ys__n47226 & ~new_n48524_;
  assign new_n50627_ = ~new_n50625_ & ~new_n50626_;
  assign ys__n32987 = ~new_n48527_ & ~new_n50627_;
  assign new_n50629_ = ys__n48249 & new_n48520_;
  assign new_n50630_ = ys__n47227 & ~new_n48524_;
  assign new_n50631_ = ~new_n50629_ & ~new_n50630_;
  assign ys__n32988 = ~new_n48527_ & ~new_n50631_;
  assign new_n50633_ = ys__n48250 & new_n48520_;
  assign new_n50634_ = ys__n47228 & ~new_n48524_;
  assign new_n50635_ = ~new_n50633_ & ~new_n50634_;
  assign ys__n32989 = ~new_n48527_ & ~new_n50635_;
  assign new_n50637_ = ys__n48251 & new_n48520_;
  assign new_n50638_ = ys__n47229 & ~new_n48524_;
  assign new_n50639_ = ~new_n50637_ & ~new_n50638_;
  assign ys__n32990 = ~new_n48527_ & ~new_n50639_;
  assign new_n50641_ = ys__n48252 & new_n48520_;
  assign new_n50642_ = ys__n47230 & ~new_n48524_;
  assign new_n50643_ = ~new_n50641_ & ~new_n50642_;
  assign ys__n32991 = ~new_n48527_ & ~new_n50643_;
  assign new_n50645_ = ys__n48253 & new_n48520_;
  assign new_n50646_ = ys__n47231 & ~new_n48524_;
  assign new_n50647_ = ~new_n50645_ & ~new_n50646_;
  assign ys__n32992 = ~new_n48527_ & ~new_n50647_;
  assign new_n50649_ = ys__n48254 & new_n48520_;
  assign new_n50650_ = ys__n47232 & ~new_n48524_;
  assign new_n50651_ = ~new_n50649_ & ~new_n50650_;
  assign ys__n32993 = ~new_n48527_ & ~new_n50651_;
  assign new_n50653_ = ys__n48255 & new_n48520_;
  assign new_n50654_ = ys__n47233 & ~new_n48524_;
  assign new_n50655_ = ~new_n50653_ & ~new_n50654_;
  assign ys__n32994 = ~new_n48527_ & ~new_n50655_;
  assign new_n50657_ = ys__n48256 & new_n48520_;
  assign new_n50658_ = ys__n18762 & ~new_n48524_;
  assign new_n50659_ = ~new_n50657_ & ~new_n50658_;
  assign ys__n32995 = ~new_n48527_ & ~new_n50659_;
  assign new_n50661_ = ys__n48257 & new_n48520_;
  assign new_n50662_ = ys__n18750 & ~new_n48524_;
  assign new_n50663_ = ~new_n50661_ & ~new_n50662_;
  assign ys__n32996 = ~new_n48527_ & ~new_n50663_;
  assign new_n50665_ = ys__n48258 & new_n48520_;
  assign new_n50666_ = ys__n18753 & ~new_n48524_;
  assign new_n50667_ = ~new_n50665_ & ~new_n50666_;
  assign ys__n32997 = ~new_n48527_ & ~new_n50667_;
  assign ys__n32998 = new_n13477_ & ~new_n13486_;
  assign new_n50670_ = ys__n140 & ~ys__n214;
  assign new_n50671_ = new_n13288_ & new_n50670_;
  assign new_n50672_ = ~new_n13290_ & ~new_n50671_;
  assign new_n50673_ = new_n13287_ & new_n50672_;
  assign new_n50674_ = new_n18038_ & new_n50673_;
  assign new_n50675_ = ~ys__n740 & new_n18038_;
  assign new_n50676_ = new_n13284_ & new_n50675_;
  assign new_n50677_ = ys__n30223 & new_n18038_;
  assign new_n50678_ = new_n13286_ & new_n50677_;
  assign new_n50679_ = ~new_n50676_ & ~new_n50678_;
  assign new_n50680_ = ~ys__n1020 & new_n13563_;
  assign new_n50681_ = new_n18038_ & new_n50680_;
  assign new_n50682_ = new_n13290_ & new_n50681_;
  assign new_n50683_ = new_n50671_ & new_n50675_;
  assign new_n50684_ = ~new_n50682_ & ~new_n50683_;
  assign new_n50685_ = new_n50679_ & new_n50684_;
  assign new_n50686_ = ~new_n50673_ & ~new_n50685_;
  assign ys__n33014 = new_n50674_ | new_n50686_;
  assign new_n50688_ = new_n13264_ & new_n50673_;
  assign new_n50689_ = ~ys__n740 & new_n13264_;
  assign new_n50690_ = new_n13284_ & new_n50689_;
  assign new_n50691_ = ys__n30223 & new_n13264_;
  assign new_n50692_ = new_n13286_ & new_n50691_;
  assign new_n50693_ = ~new_n50690_ & ~new_n50692_;
  assign new_n50694_ = new_n13264_ & new_n50680_;
  assign new_n50695_ = new_n13290_ & new_n50694_;
  assign new_n50696_ = new_n50671_ & new_n50689_;
  assign new_n50697_ = ~new_n50695_ & ~new_n50696_;
  assign new_n50698_ = new_n50693_ & new_n50697_;
  assign new_n50699_ = ~new_n50673_ & ~new_n50698_;
  assign ys__n33015 = new_n50688_ | new_n50699_;
  assign new_n50701_ = new_n13246_ & new_n50673_;
  assign new_n50702_ = ~ys__n740 & new_n13246_;
  assign new_n50703_ = new_n13284_ & new_n50702_;
  assign new_n50704_ = ys__n30223 & new_n13246_;
  assign new_n50705_ = new_n13286_ & new_n50704_;
  assign new_n50706_ = ~new_n50703_ & ~new_n50705_;
  assign new_n50707_ = new_n13246_ & new_n50680_;
  assign new_n50708_ = new_n13290_ & new_n50707_;
  assign new_n50709_ = new_n50671_ & new_n50702_;
  assign new_n50710_ = ~new_n50708_ & ~new_n50709_;
  assign new_n50711_ = new_n50706_ & new_n50710_;
  assign new_n50712_ = ~new_n50673_ & ~new_n50711_;
  assign ys__n33016 = new_n50701_ | new_n50712_;
  assign new_n50714_ = new_n13188_ & new_n50673_;
  assign new_n50715_ = ~ys__n740 & new_n13188_;
  assign new_n50716_ = new_n13284_ & new_n50715_;
  assign new_n50717_ = ys__n30223 & new_n13188_;
  assign new_n50718_ = new_n13286_ & new_n50717_;
  assign new_n50719_ = ~new_n50716_ & ~new_n50718_;
  assign new_n50720_ = new_n13188_ & new_n50680_;
  assign new_n50721_ = new_n13290_ & new_n50720_;
  assign new_n50722_ = new_n50671_ & new_n50715_;
  assign new_n50723_ = ~new_n50721_ & ~new_n50722_;
  assign new_n50724_ = new_n50719_ & new_n50723_;
  assign new_n50725_ = ~new_n50673_ & ~new_n50724_;
  assign ys__n33017 = new_n50714_ | new_n50725_;
  assign new_n50727_ = new_n11739_ & new_n50673_;
  assign new_n50728_ = new_n11739_ & ~ys__n740;
  assign new_n50729_ = new_n13284_ & new_n50728_;
  assign new_n50730_ = new_n11739_ & ys__n30223;
  assign new_n50731_ = new_n13286_ & new_n50730_;
  assign new_n50732_ = ~new_n50729_ & ~new_n50731_;
  assign new_n50733_ = new_n11739_ & new_n50680_;
  assign new_n50734_ = new_n13290_ & new_n50733_;
  assign new_n50735_ = new_n50671_ & new_n50728_;
  assign new_n50736_ = ~new_n50734_ & ~new_n50735_;
  assign new_n50737_ = new_n50732_ & new_n50736_;
  assign new_n50738_ = ~new_n50673_ & ~new_n50737_;
  assign ys__n33018 = new_n50727_ | new_n50738_;
  assign new_n50740_ = new_n45663_ & new_n50673_;
  assign new_n50741_ = ~ys__n740 & new_n45663_;
  assign new_n50742_ = new_n13284_ & new_n50741_;
  assign new_n50743_ = ys__n30223 & new_n45663_;
  assign new_n50744_ = new_n13286_ & new_n50743_;
  assign new_n50745_ = ~new_n50742_ & ~new_n50744_;
  assign new_n50746_ = new_n45663_ & new_n50680_;
  assign new_n50747_ = new_n13290_ & new_n50746_;
  assign new_n50748_ = new_n50671_ & new_n50741_;
  assign new_n50749_ = ~new_n50747_ & ~new_n50748_;
  assign new_n50750_ = new_n50745_ & new_n50749_;
  assign new_n50751_ = ~new_n50673_ & ~new_n50750_;
  assign ys__n33019 = new_n50740_ | new_n50751_;
  assign new_n50753_ = new_n27304_ & new_n50673_;
  assign new_n50754_ = ~ys__n740 & new_n27304_;
  assign new_n50755_ = new_n13284_ & new_n50754_;
  assign new_n50756_ = ys__n30223 & new_n27304_;
  assign new_n50757_ = new_n13286_ & new_n50756_;
  assign new_n50758_ = ~new_n50755_ & ~new_n50757_;
  assign new_n50759_ = new_n27304_ & new_n50680_;
  assign new_n50760_ = new_n13290_ & new_n50759_;
  assign new_n50761_ = new_n50671_ & new_n50754_;
  assign new_n50762_ = ~new_n50760_ & ~new_n50761_;
  assign new_n50763_ = new_n50758_ & new_n50762_;
  assign new_n50764_ = ~new_n50673_ & ~new_n50763_;
  assign ys__n33020 = new_n50753_ | new_n50764_;
  assign new_n50766_ = new_n27315_ & new_n50673_;
  assign new_n50767_ = ~ys__n740 & new_n27315_;
  assign new_n50768_ = new_n13284_ & new_n50767_;
  assign new_n50769_ = ys__n30223 & new_n27315_;
  assign new_n50770_ = new_n13286_ & new_n50769_;
  assign new_n50771_ = ~new_n50768_ & ~new_n50770_;
  assign new_n50772_ = new_n27315_ & new_n50680_;
  assign new_n50773_ = new_n13290_ & new_n50772_;
  assign new_n50774_ = new_n50671_ & new_n50767_;
  assign new_n50775_ = ~new_n50773_ & ~new_n50774_;
  assign new_n50776_ = new_n50771_ & new_n50775_;
  assign new_n50777_ = ~new_n50673_ & ~new_n50776_;
  assign ys__n33021 = new_n50766_ | new_n50777_;
  assign new_n50779_ = new_n27326_ & new_n50673_;
  assign new_n50780_ = ~ys__n740 & new_n27326_;
  assign new_n50781_ = new_n13284_ & new_n50780_;
  assign new_n50782_ = ys__n30223 & new_n27326_;
  assign new_n50783_ = new_n13286_ & new_n50782_;
  assign new_n50784_ = ~new_n50781_ & ~new_n50783_;
  assign new_n50785_ = new_n27326_ & new_n50680_;
  assign new_n50786_ = new_n13290_ & new_n50785_;
  assign new_n50787_ = new_n50671_ & new_n50780_;
  assign new_n50788_ = ~new_n50786_ & ~new_n50787_;
  assign new_n50789_ = new_n50784_ & new_n50788_;
  assign new_n50790_ = ~new_n50673_ & ~new_n50789_;
  assign ys__n33022 = new_n50779_ | new_n50790_;
  assign new_n50792_ = new_n18026_ & new_n50673_;
  assign new_n50793_ = ~ys__n740 & new_n18026_;
  assign new_n50794_ = new_n13284_ & new_n50793_;
  assign new_n50795_ = ys__n30223 & new_n18026_;
  assign new_n50796_ = new_n13286_ & new_n50795_;
  assign new_n50797_ = ~new_n50794_ & ~new_n50796_;
  assign new_n50798_ = new_n18026_ & new_n50680_;
  assign new_n50799_ = new_n13290_ & new_n50798_;
  assign new_n50800_ = new_n50671_ & new_n50793_;
  assign new_n50801_ = ~new_n50799_ & ~new_n50800_;
  assign new_n50802_ = new_n50797_ & new_n50801_;
  assign new_n50803_ = ~new_n50673_ & ~new_n50802_;
  assign ys__n33023 = new_n50792_ | new_n50803_;
  assign new_n50805_ = new_n45674_ & new_n50673_;
  assign new_n50806_ = ~ys__n740 & new_n45674_;
  assign new_n50807_ = new_n13284_ & new_n50806_;
  assign new_n50808_ = ys__n30223 & new_n45674_;
  assign new_n50809_ = new_n13286_ & new_n50808_;
  assign new_n50810_ = ~new_n50807_ & ~new_n50809_;
  assign new_n50811_ = new_n45674_ & new_n50680_;
  assign new_n50812_ = new_n13290_ & new_n50811_;
  assign new_n50813_ = new_n50671_ & new_n50806_;
  assign new_n50814_ = ~new_n50812_ & ~new_n50813_;
  assign new_n50815_ = new_n50810_ & new_n50814_;
  assign new_n50816_ = ~new_n50673_ & ~new_n50815_;
  assign ys__n33024 = new_n50805_ | new_n50816_;
  assign new_n50818_ = new_n45685_ & new_n50673_;
  assign new_n50819_ = ~ys__n740 & new_n45685_;
  assign new_n50820_ = new_n13284_ & new_n50819_;
  assign new_n50821_ = ys__n30223 & new_n45685_;
  assign new_n50822_ = new_n13286_ & new_n50821_;
  assign new_n50823_ = ~new_n50820_ & ~new_n50822_;
  assign new_n50824_ = new_n45685_ & new_n50680_;
  assign new_n50825_ = new_n13290_ & new_n50824_;
  assign new_n50826_ = new_n50671_ & new_n50819_;
  assign new_n50827_ = ~new_n50825_ & ~new_n50826_;
  assign new_n50828_ = new_n50823_ & new_n50827_;
  assign new_n50829_ = ~new_n50673_ & ~new_n50828_;
  assign ys__n33025 = new_n50818_ | new_n50829_;
  assign new_n50831_ = new_n45696_ & new_n50673_;
  assign new_n50832_ = ~ys__n740 & new_n45696_;
  assign new_n50833_ = new_n13284_ & new_n50832_;
  assign new_n50834_ = ys__n30223 & new_n45696_;
  assign new_n50835_ = new_n13286_ & new_n50834_;
  assign new_n50836_ = ~new_n50833_ & ~new_n50835_;
  assign new_n50837_ = new_n45696_ & new_n50680_;
  assign new_n50838_ = new_n13290_ & new_n50837_;
  assign new_n50839_ = new_n50671_ & new_n50832_;
  assign new_n50840_ = ~new_n50838_ & ~new_n50839_;
  assign new_n50841_ = new_n50836_ & new_n50840_;
  assign new_n50842_ = ~new_n50673_ & ~new_n50841_;
  assign ys__n33026 = new_n50831_ | new_n50842_;
  assign new_n50844_ = new_n45707_ & new_n50673_;
  assign new_n50845_ = ~ys__n740 & new_n45707_;
  assign new_n50846_ = new_n13284_ & new_n50845_;
  assign new_n50847_ = ys__n30223 & new_n45707_;
  assign new_n50848_ = new_n13286_ & new_n50847_;
  assign new_n50849_ = ~new_n50846_ & ~new_n50848_;
  assign new_n50850_ = new_n45707_ & new_n50680_;
  assign new_n50851_ = new_n13290_ & new_n50850_;
  assign new_n50852_ = new_n50671_ & new_n50845_;
  assign new_n50853_ = ~new_n50851_ & ~new_n50852_;
  assign new_n50854_ = new_n50849_ & new_n50853_;
  assign new_n50855_ = ~new_n50673_ & ~new_n50854_;
  assign ys__n33027 = new_n50844_ | new_n50855_;
  assign new_n50857_ = new_n45720_ & new_n50673_;
  assign new_n50858_ = ~ys__n740 & new_n45720_;
  assign new_n50859_ = new_n13284_ & new_n50858_;
  assign new_n50860_ = ys__n30223 & new_n45720_;
  assign new_n50861_ = new_n13286_ & new_n50860_;
  assign new_n50862_ = ~new_n50859_ & ~new_n50861_;
  assign new_n50863_ = new_n45720_ & new_n50680_;
  assign new_n50864_ = new_n13290_ & new_n50863_;
  assign new_n50865_ = new_n50671_ & new_n50858_;
  assign new_n50866_ = ~new_n50864_ & ~new_n50865_;
  assign new_n50867_ = new_n50862_ & new_n50866_;
  assign new_n50868_ = ~new_n50673_ & ~new_n50867_;
  assign ys__n33028 = new_n50857_ | new_n50868_;
  assign new_n50870_ = new_n45731_ & new_n50673_;
  assign new_n50871_ = ~ys__n740 & new_n45731_;
  assign new_n50872_ = new_n13284_ & new_n50871_;
  assign new_n50873_ = ys__n30223 & new_n45731_;
  assign new_n50874_ = new_n13286_ & new_n50873_;
  assign new_n50875_ = ~new_n50872_ & ~new_n50874_;
  assign new_n50876_ = new_n45731_ & new_n50680_;
  assign new_n50877_ = new_n13290_ & new_n50876_;
  assign new_n50878_ = new_n50671_ & new_n50871_;
  assign new_n50879_ = ~new_n50877_ & ~new_n50878_;
  assign new_n50880_ = new_n50875_ & new_n50879_;
  assign new_n50881_ = ~new_n50673_ & ~new_n50880_;
  assign ys__n33029 = new_n50870_ | new_n50881_;
  assign new_n50883_ = new_n18041_ & new_n50673_;
  assign new_n50884_ = ~ys__n740 & new_n18041_;
  assign new_n50885_ = new_n13284_ & new_n50884_;
  assign new_n50886_ = ys__n30223 & new_n18041_;
  assign new_n50887_ = new_n13286_ & new_n50886_;
  assign new_n50888_ = ~new_n50885_ & ~new_n50887_;
  assign new_n50889_ = new_n18041_ & new_n50680_;
  assign new_n50890_ = new_n13290_ & new_n50889_;
  assign new_n50891_ = new_n50671_ & new_n50884_;
  assign new_n50892_ = ~new_n50890_ & ~new_n50891_;
  assign new_n50893_ = new_n50888_ & new_n50892_;
  assign new_n50894_ = ~new_n50673_ & ~new_n50893_;
  assign ys__n33030 = new_n50883_ | new_n50894_;
  assign new_n50896_ = new_n13267_ & new_n50673_;
  assign new_n50897_ = ~ys__n740 & new_n13267_;
  assign new_n50898_ = new_n13284_ & new_n50897_;
  assign new_n50899_ = ys__n30223 & new_n13267_;
  assign new_n50900_ = new_n13286_ & new_n50899_;
  assign new_n50901_ = ~new_n50898_ & ~new_n50900_;
  assign new_n50902_ = new_n13267_ & new_n50680_;
  assign new_n50903_ = new_n13290_ & new_n50902_;
  assign new_n50904_ = new_n50671_ & new_n50897_;
  assign new_n50905_ = ~new_n50903_ & ~new_n50904_;
  assign new_n50906_ = new_n50901_ & new_n50905_;
  assign new_n50907_ = ~new_n50673_ & ~new_n50906_;
  assign ys__n33031 = new_n50896_ | new_n50907_;
  assign new_n50909_ = new_n13249_ & new_n50673_;
  assign new_n50910_ = ~ys__n740 & new_n13249_;
  assign new_n50911_ = new_n13284_ & new_n50910_;
  assign new_n50912_ = ys__n30223 & new_n13249_;
  assign new_n50913_ = new_n13286_ & new_n50912_;
  assign new_n50914_ = ~new_n50911_ & ~new_n50913_;
  assign new_n50915_ = new_n13249_ & new_n50680_;
  assign new_n50916_ = new_n13290_ & new_n50915_;
  assign new_n50917_ = new_n50671_ & new_n50910_;
  assign new_n50918_ = ~new_n50916_ & ~new_n50917_;
  assign new_n50919_ = new_n50914_ & new_n50918_;
  assign new_n50920_ = ~new_n50673_ & ~new_n50919_;
  assign ys__n33032 = new_n50909_ | new_n50920_;
  assign new_n50922_ = new_n13191_ & new_n50673_;
  assign new_n50923_ = ~ys__n740 & new_n13191_;
  assign new_n50924_ = new_n13284_ & new_n50923_;
  assign new_n50925_ = ys__n30223 & new_n13191_;
  assign new_n50926_ = new_n13286_ & new_n50925_;
  assign new_n50927_ = ~new_n50924_ & ~new_n50926_;
  assign new_n50928_ = new_n13191_ & new_n50680_;
  assign new_n50929_ = new_n13290_ & new_n50928_;
  assign new_n50930_ = new_n50671_ & new_n50923_;
  assign new_n50931_ = ~new_n50929_ & ~new_n50930_;
  assign new_n50932_ = new_n50927_ & new_n50931_;
  assign new_n50933_ = ~new_n50673_ & ~new_n50932_;
  assign ys__n33033 = new_n50922_ | new_n50933_;
  assign new_n50935_ = new_n11754_ & new_n50673_;
  assign new_n50936_ = new_n11754_ & ~ys__n740;
  assign new_n50937_ = new_n13284_ & new_n50936_;
  assign new_n50938_ = new_n11754_ & ys__n30223;
  assign new_n50939_ = new_n13286_ & new_n50938_;
  assign new_n50940_ = ~new_n50937_ & ~new_n50939_;
  assign new_n50941_ = new_n11754_ & new_n50680_;
  assign new_n50942_ = new_n13290_ & new_n50941_;
  assign new_n50943_ = new_n50671_ & new_n50936_;
  assign new_n50944_ = ~new_n50942_ & ~new_n50943_;
  assign new_n50945_ = new_n50940_ & new_n50944_;
  assign new_n50946_ = ~new_n50673_ & ~new_n50945_;
  assign ys__n33034 = new_n50935_ | new_n50946_;
  assign new_n50948_ = ~ys__n740 & new_n13320_;
  assign new_n50949_ = ~ys__n23850 & new_n13317_;
  assign new_n50950_ = ~new_n50948_ & ~new_n50949_;
  assign new_n50951_ = ~new_n13324_ & ~new_n50950_;
  assign ys__n33035 = new_n13324_ | new_n50951_;
  assign new_n50953_ = ys__n140 & ~ys__n210;
  assign new_n50954_ = new_n13299_ & new_n50953_;
  assign new_n50955_ = ~new_n13301_ & ~new_n50954_;
  assign new_n50956_ = new_n13298_ & new_n50955_;
  assign new_n50957_ = new_n18038_ & new_n50956_;
  assign new_n50958_ = new_n13295_ & new_n50675_;
  assign new_n50959_ = new_n13297_ & new_n50677_;
  assign new_n50960_ = ~new_n50958_ & ~new_n50959_;
  assign new_n50961_ = new_n13301_ & new_n50681_;
  assign new_n50962_ = new_n50675_ & new_n50954_;
  assign new_n50963_ = ~new_n50961_ & ~new_n50962_;
  assign new_n50964_ = new_n50960_ & new_n50963_;
  assign new_n50965_ = ~new_n50956_ & ~new_n50964_;
  assign ys__n33036 = new_n50957_ | new_n50965_;
  assign new_n50967_ = new_n13264_ & new_n50956_;
  assign new_n50968_ = new_n13295_ & new_n50689_;
  assign new_n50969_ = new_n13297_ & new_n50691_;
  assign new_n50970_ = ~new_n50968_ & ~new_n50969_;
  assign new_n50971_ = new_n13301_ & new_n50694_;
  assign new_n50972_ = new_n50689_ & new_n50954_;
  assign new_n50973_ = ~new_n50971_ & ~new_n50972_;
  assign new_n50974_ = new_n50970_ & new_n50973_;
  assign new_n50975_ = ~new_n50956_ & ~new_n50974_;
  assign ys__n33037 = new_n50967_ | new_n50975_;
  assign new_n50977_ = new_n13246_ & new_n50956_;
  assign new_n50978_ = new_n13295_ & new_n50702_;
  assign new_n50979_ = new_n13297_ & new_n50704_;
  assign new_n50980_ = ~new_n50978_ & ~new_n50979_;
  assign new_n50981_ = new_n13301_ & new_n50707_;
  assign new_n50982_ = new_n50702_ & new_n50954_;
  assign new_n50983_ = ~new_n50981_ & ~new_n50982_;
  assign new_n50984_ = new_n50980_ & new_n50983_;
  assign new_n50985_ = ~new_n50956_ & ~new_n50984_;
  assign ys__n33038 = new_n50977_ | new_n50985_;
  assign new_n50987_ = new_n13188_ & new_n50956_;
  assign new_n50988_ = new_n13295_ & new_n50715_;
  assign new_n50989_ = new_n13297_ & new_n50717_;
  assign new_n50990_ = ~new_n50988_ & ~new_n50989_;
  assign new_n50991_ = new_n13301_ & new_n50720_;
  assign new_n50992_ = new_n50715_ & new_n50954_;
  assign new_n50993_ = ~new_n50991_ & ~new_n50992_;
  assign new_n50994_ = new_n50990_ & new_n50993_;
  assign new_n50995_ = ~new_n50956_ & ~new_n50994_;
  assign ys__n33039 = new_n50987_ | new_n50995_;
  assign new_n50997_ = new_n11739_ & new_n50956_;
  assign new_n50998_ = new_n13295_ & new_n50728_;
  assign new_n50999_ = new_n13297_ & new_n50730_;
  assign new_n51000_ = ~new_n50998_ & ~new_n50999_;
  assign new_n51001_ = new_n13301_ & new_n50733_;
  assign new_n51002_ = new_n50728_ & new_n50954_;
  assign new_n51003_ = ~new_n51001_ & ~new_n51002_;
  assign new_n51004_ = new_n51000_ & new_n51003_;
  assign new_n51005_ = ~new_n50956_ & ~new_n51004_;
  assign ys__n33040 = new_n50997_ | new_n51005_;
  assign new_n51007_ = new_n45663_ & new_n50956_;
  assign new_n51008_ = new_n13295_ & new_n50741_;
  assign new_n51009_ = new_n13297_ & new_n50743_;
  assign new_n51010_ = ~new_n51008_ & ~new_n51009_;
  assign new_n51011_ = new_n13301_ & new_n50746_;
  assign new_n51012_ = new_n50741_ & new_n50954_;
  assign new_n51013_ = ~new_n51011_ & ~new_n51012_;
  assign new_n51014_ = new_n51010_ & new_n51013_;
  assign new_n51015_ = ~new_n50956_ & ~new_n51014_;
  assign ys__n33041 = new_n51007_ | new_n51015_;
  assign new_n51017_ = new_n27304_ & new_n50956_;
  assign new_n51018_ = new_n13295_ & new_n50754_;
  assign new_n51019_ = new_n13297_ & new_n50756_;
  assign new_n51020_ = ~new_n51018_ & ~new_n51019_;
  assign new_n51021_ = new_n13301_ & new_n50759_;
  assign new_n51022_ = new_n50754_ & new_n50954_;
  assign new_n51023_ = ~new_n51021_ & ~new_n51022_;
  assign new_n51024_ = new_n51020_ & new_n51023_;
  assign new_n51025_ = ~new_n50956_ & ~new_n51024_;
  assign ys__n33042 = new_n51017_ | new_n51025_;
  assign new_n51027_ = new_n27315_ & new_n50956_;
  assign new_n51028_ = new_n13295_ & new_n50767_;
  assign new_n51029_ = new_n13297_ & new_n50769_;
  assign new_n51030_ = ~new_n51028_ & ~new_n51029_;
  assign new_n51031_ = new_n13301_ & new_n50772_;
  assign new_n51032_ = new_n50767_ & new_n50954_;
  assign new_n51033_ = ~new_n51031_ & ~new_n51032_;
  assign new_n51034_ = new_n51030_ & new_n51033_;
  assign new_n51035_ = ~new_n50956_ & ~new_n51034_;
  assign ys__n33043 = new_n51027_ | new_n51035_;
  assign new_n51037_ = new_n27326_ & new_n50956_;
  assign new_n51038_ = new_n13295_ & new_n50780_;
  assign new_n51039_ = new_n13297_ & new_n50782_;
  assign new_n51040_ = ~new_n51038_ & ~new_n51039_;
  assign new_n51041_ = new_n13301_ & new_n50785_;
  assign new_n51042_ = new_n50780_ & new_n50954_;
  assign new_n51043_ = ~new_n51041_ & ~new_n51042_;
  assign new_n51044_ = new_n51040_ & new_n51043_;
  assign new_n51045_ = ~new_n50956_ & ~new_n51044_;
  assign ys__n33044 = new_n51037_ | new_n51045_;
  assign new_n51047_ = new_n18026_ & new_n50956_;
  assign new_n51048_ = new_n13295_ & new_n50793_;
  assign new_n51049_ = new_n13297_ & new_n50795_;
  assign new_n51050_ = ~new_n51048_ & ~new_n51049_;
  assign new_n51051_ = new_n13301_ & new_n50798_;
  assign new_n51052_ = new_n50793_ & new_n50954_;
  assign new_n51053_ = ~new_n51051_ & ~new_n51052_;
  assign new_n51054_ = new_n51050_ & new_n51053_;
  assign new_n51055_ = ~new_n50956_ & ~new_n51054_;
  assign ys__n33045 = new_n51047_ | new_n51055_;
  assign new_n51057_ = new_n45674_ & new_n50956_;
  assign new_n51058_ = new_n13295_ & new_n50806_;
  assign new_n51059_ = new_n13297_ & new_n50808_;
  assign new_n51060_ = ~new_n51058_ & ~new_n51059_;
  assign new_n51061_ = new_n13301_ & new_n50811_;
  assign new_n51062_ = new_n50806_ & new_n50954_;
  assign new_n51063_ = ~new_n51061_ & ~new_n51062_;
  assign new_n51064_ = new_n51060_ & new_n51063_;
  assign new_n51065_ = ~new_n50956_ & ~new_n51064_;
  assign ys__n33046 = new_n51057_ | new_n51065_;
  assign new_n51067_ = new_n45685_ & new_n50956_;
  assign new_n51068_ = new_n13295_ & new_n50819_;
  assign new_n51069_ = new_n13297_ & new_n50821_;
  assign new_n51070_ = ~new_n51068_ & ~new_n51069_;
  assign new_n51071_ = new_n13301_ & new_n50824_;
  assign new_n51072_ = new_n50819_ & new_n50954_;
  assign new_n51073_ = ~new_n51071_ & ~new_n51072_;
  assign new_n51074_ = new_n51070_ & new_n51073_;
  assign new_n51075_ = ~new_n50956_ & ~new_n51074_;
  assign ys__n33047 = new_n51067_ | new_n51075_;
  assign new_n51077_ = new_n45696_ & new_n50956_;
  assign new_n51078_ = new_n13295_ & new_n50832_;
  assign new_n51079_ = new_n13297_ & new_n50834_;
  assign new_n51080_ = ~new_n51078_ & ~new_n51079_;
  assign new_n51081_ = new_n13301_ & new_n50837_;
  assign new_n51082_ = new_n50832_ & new_n50954_;
  assign new_n51083_ = ~new_n51081_ & ~new_n51082_;
  assign new_n51084_ = new_n51080_ & new_n51083_;
  assign new_n51085_ = ~new_n50956_ & ~new_n51084_;
  assign ys__n33048 = new_n51077_ | new_n51085_;
  assign new_n51087_ = new_n45707_ & new_n50956_;
  assign new_n51088_ = new_n13295_ & new_n50845_;
  assign new_n51089_ = new_n13297_ & new_n50847_;
  assign new_n51090_ = ~new_n51088_ & ~new_n51089_;
  assign new_n51091_ = new_n13301_ & new_n50850_;
  assign new_n51092_ = new_n50845_ & new_n50954_;
  assign new_n51093_ = ~new_n51091_ & ~new_n51092_;
  assign new_n51094_ = new_n51090_ & new_n51093_;
  assign new_n51095_ = ~new_n50956_ & ~new_n51094_;
  assign ys__n33049 = new_n51087_ | new_n51095_;
  assign new_n51097_ = new_n45720_ & new_n50956_;
  assign new_n51098_ = new_n13295_ & new_n50858_;
  assign new_n51099_ = new_n13297_ & new_n50860_;
  assign new_n51100_ = ~new_n51098_ & ~new_n51099_;
  assign new_n51101_ = new_n13301_ & new_n50863_;
  assign new_n51102_ = new_n50858_ & new_n50954_;
  assign new_n51103_ = ~new_n51101_ & ~new_n51102_;
  assign new_n51104_ = new_n51100_ & new_n51103_;
  assign new_n51105_ = ~new_n50956_ & ~new_n51104_;
  assign ys__n33050 = new_n51097_ | new_n51105_;
  assign new_n51107_ = new_n45731_ & new_n50956_;
  assign new_n51108_ = new_n13295_ & new_n50871_;
  assign new_n51109_ = new_n13297_ & new_n50873_;
  assign new_n51110_ = ~new_n51108_ & ~new_n51109_;
  assign new_n51111_ = new_n13301_ & new_n50876_;
  assign new_n51112_ = new_n50871_ & new_n50954_;
  assign new_n51113_ = ~new_n51111_ & ~new_n51112_;
  assign new_n51114_ = new_n51110_ & new_n51113_;
  assign new_n51115_ = ~new_n50956_ & ~new_n51114_;
  assign ys__n33051 = new_n51107_ | new_n51115_;
  assign new_n51117_ = new_n18041_ & new_n50956_;
  assign new_n51118_ = new_n13295_ & new_n50884_;
  assign new_n51119_ = new_n13297_ & new_n50886_;
  assign new_n51120_ = ~new_n51118_ & ~new_n51119_;
  assign new_n51121_ = new_n13301_ & new_n50889_;
  assign new_n51122_ = new_n50884_ & new_n50954_;
  assign new_n51123_ = ~new_n51121_ & ~new_n51122_;
  assign new_n51124_ = new_n51120_ & new_n51123_;
  assign new_n51125_ = ~new_n50956_ & ~new_n51124_;
  assign ys__n33052 = new_n51117_ | new_n51125_;
  assign new_n51127_ = new_n13267_ & new_n50956_;
  assign new_n51128_ = new_n13295_ & new_n50897_;
  assign new_n51129_ = new_n13297_ & new_n50899_;
  assign new_n51130_ = ~new_n51128_ & ~new_n51129_;
  assign new_n51131_ = new_n13301_ & new_n50902_;
  assign new_n51132_ = new_n50897_ & new_n50954_;
  assign new_n51133_ = ~new_n51131_ & ~new_n51132_;
  assign new_n51134_ = new_n51130_ & new_n51133_;
  assign new_n51135_ = ~new_n50956_ & ~new_n51134_;
  assign ys__n33053 = new_n51127_ | new_n51135_;
  assign new_n51137_ = new_n13249_ & new_n50956_;
  assign new_n51138_ = new_n13295_ & new_n50910_;
  assign new_n51139_ = new_n13297_ & new_n50912_;
  assign new_n51140_ = ~new_n51138_ & ~new_n51139_;
  assign new_n51141_ = new_n13301_ & new_n50915_;
  assign new_n51142_ = new_n50910_ & new_n50954_;
  assign new_n51143_ = ~new_n51141_ & ~new_n51142_;
  assign new_n51144_ = new_n51140_ & new_n51143_;
  assign new_n51145_ = ~new_n50956_ & ~new_n51144_;
  assign ys__n33054 = new_n51137_ | new_n51145_;
  assign new_n51147_ = new_n13191_ & new_n50956_;
  assign new_n51148_ = new_n13295_ & new_n50923_;
  assign new_n51149_ = new_n13297_ & new_n50925_;
  assign new_n51150_ = ~new_n51148_ & ~new_n51149_;
  assign new_n51151_ = new_n13301_ & new_n50928_;
  assign new_n51152_ = new_n50923_ & new_n50954_;
  assign new_n51153_ = ~new_n51151_ & ~new_n51152_;
  assign new_n51154_ = new_n51150_ & new_n51153_;
  assign new_n51155_ = ~new_n50956_ & ~new_n51154_;
  assign ys__n33055 = new_n51147_ | new_n51155_;
  assign new_n51157_ = new_n11754_ & new_n50956_;
  assign new_n51158_ = new_n13295_ & new_n50936_;
  assign new_n51159_ = new_n13297_ & new_n50938_;
  assign new_n51160_ = ~new_n51158_ & ~new_n51159_;
  assign new_n51161_ = new_n13301_ & new_n50941_;
  assign new_n51162_ = new_n50936_ & new_n50954_;
  assign new_n51163_ = ~new_n51161_ & ~new_n51162_;
  assign new_n51164_ = new_n51160_ & new_n51163_;
  assign new_n51165_ = ~new_n50956_ & ~new_n51164_;
  assign ys__n33056 = new_n51157_ | new_n51165_;
  assign new_n51167_ = ~ys__n740 & new_n13309_;
  assign new_n51168_ = ~ys__n23850 & new_n13306_;
  assign new_n51169_ = ~new_n51167_ & ~new_n51168_;
  assign new_n51170_ = ~new_n13313_ & ~new_n51169_;
  assign ys__n33058 = new_n13313_ | new_n51170_;
  assign new_n51172_ = ~ys__n138 & ys__n140;
  assign new_n51173_ = new_n13332_ & new_n51172_;
  assign new_n51174_ = ~new_n13334_ & ~new_n51173_;
  assign new_n51175_ = new_n13331_ & new_n51174_;
  assign new_n51176_ = new_n18038_ & new_n51175_;
  assign new_n51177_ = new_n13328_ & new_n50675_;
  assign new_n51178_ = new_n13330_ & new_n50677_;
  assign new_n51179_ = ~new_n51177_ & ~new_n51178_;
  assign new_n51180_ = new_n13334_ & new_n50681_;
  assign new_n51181_ = new_n50675_ & new_n51173_;
  assign new_n51182_ = ~new_n51180_ & ~new_n51181_;
  assign new_n51183_ = new_n51179_ & new_n51182_;
  assign new_n51184_ = ~new_n51175_ & ~new_n51183_;
  assign ys__n33059 = new_n51176_ | new_n51184_;
  assign new_n51186_ = new_n13264_ & new_n51175_;
  assign new_n51187_ = new_n13328_ & new_n50689_;
  assign new_n51188_ = new_n13330_ & new_n50691_;
  assign new_n51189_ = ~new_n51187_ & ~new_n51188_;
  assign new_n51190_ = new_n13334_ & new_n50694_;
  assign new_n51191_ = new_n50689_ & new_n51173_;
  assign new_n51192_ = ~new_n51190_ & ~new_n51191_;
  assign new_n51193_ = new_n51189_ & new_n51192_;
  assign new_n51194_ = ~new_n51175_ & ~new_n51193_;
  assign ys__n33060 = new_n51186_ | new_n51194_;
  assign new_n51196_ = new_n13246_ & new_n51175_;
  assign new_n51197_ = new_n13328_ & new_n50702_;
  assign new_n51198_ = new_n13330_ & new_n50704_;
  assign new_n51199_ = ~new_n51197_ & ~new_n51198_;
  assign new_n51200_ = new_n13334_ & new_n50707_;
  assign new_n51201_ = new_n50702_ & new_n51173_;
  assign new_n51202_ = ~new_n51200_ & ~new_n51201_;
  assign new_n51203_ = new_n51199_ & new_n51202_;
  assign new_n51204_ = ~new_n51175_ & ~new_n51203_;
  assign ys__n33061 = new_n51196_ | new_n51204_;
  assign new_n51206_ = new_n13188_ & new_n51175_;
  assign new_n51207_ = new_n13328_ & new_n50715_;
  assign new_n51208_ = new_n13330_ & new_n50717_;
  assign new_n51209_ = ~new_n51207_ & ~new_n51208_;
  assign new_n51210_ = new_n13334_ & new_n50720_;
  assign new_n51211_ = new_n50715_ & new_n51173_;
  assign new_n51212_ = ~new_n51210_ & ~new_n51211_;
  assign new_n51213_ = new_n51209_ & new_n51212_;
  assign new_n51214_ = ~new_n51175_ & ~new_n51213_;
  assign ys__n33062 = new_n51206_ | new_n51214_;
  assign new_n51216_ = new_n11739_ & new_n51175_;
  assign new_n51217_ = new_n13328_ & new_n50728_;
  assign new_n51218_ = new_n13330_ & new_n50730_;
  assign new_n51219_ = ~new_n51217_ & ~new_n51218_;
  assign new_n51220_ = new_n13334_ & new_n50733_;
  assign new_n51221_ = new_n50728_ & new_n51173_;
  assign new_n51222_ = ~new_n51220_ & ~new_n51221_;
  assign new_n51223_ = new_n51219_ & new_n51222_;
  assign new_n51224_ = ~new_n51175_ & ~new_n51223_;
  assign ys__n33063 = new_n51216_ | new_n51224_;
  assign new_n51226_ = new_n45663_ & new_n51175_;
  assign new_n51227_ = new_n13328_ & new_n50741_;
  assign new_n51228_ = new_n13330_ & new_n50743_;
  assign new_n51229_ = ~new_n51227_ & ~new_n51228_;
  assign new_n51230_ = new_n13334_ & new_n50746_;
  assign new_n51231_ = new_n50741_ & new_n51173_;
  assign new_n51232_ = ~new_n51230_ & ~new_n51231_;
  assign new_n51233_ = new_n51229_ & new_n51232_;
  assign new_n51234_ = ~new_n51175_ & ~new_n51233_;
  assign ys__n33064 = new_n51226_ | new_n51234_;
  assign new_n51236_ = new_n27304_ & new_n51175_;
  assign new_n51237_ = new_n13328_ & new_n50754_;
  assign new_n51238_ = new_n13330_ & new_n50756_;
  assign new_n51239_ = ~new_n51237_ & ~new_n51238_;
  assign new_n51240_ = new_n13334_ & new_n50759_;
  assign new_n51241_ = new_n50754_ & new_n51173_;
  assign new_n51242_ = ~new_n51240_ & ~new_n51241_;
  assign new_n51243_ = new_n51239_ & new_n51242_;
  assign new_n51244_ = ~new_n51175_ & ~new_n51243_;
  assign ys__n33065 = new_n51236_ | new_n51244_;
  assign new_n51246_ = new_n27315_ & new_n51175_;
  assign new_n51247_ = new_n13328_ & new_n50767_;
  assign new_n51248_ = new_n13330_ & new_n50769_;
  assign new_n51249_ = ~new_n51247_ & ~new_n51248_;
  assign new_n51250_ = new_n13334_ & new_n50772_;
  assign new_n51251_ = new_n50767_ & new_n51173_;
  assign new_n51252_ = ~new_n51250_ & ~new_n51251_;
  assign new_n51253_ = new_n51249_ & new_n51252_;
  assign new_n51254_ = ~new_n51175_ & ~new_n51253_;
  assign ys__n33066 = new_n51246_ | new_n51254_;
  assign new_n51256_ = new_n27326_ & new_n51175_;
  assign new_n51257_ = new_n13328_ & new_n50780_;
  assign new_n51258_ = new_n13330_ & new_n50782_;
  assign new_n51259_ = ~new_n51257_ & ~new_n51258_;
  assign new_n51260_ = new_n13334_ & new_n50785_;
  assign new_n51261_ = new_n50780_ & new_n51173_;
  assign new_n51262_ = ~new_n51260_ & ~new_n51261_;
  assign new_n51263_ = new_n51259_ & new_n51262_;
  assign new_n51264_ = ~new_n51175_ & ~new_n51263_;
  assign ys__n33067 = new_n51256_ | new_n51264_;
  assign new_n51266_ = new_n18026_ & new_n51175_;
  assign new_n51267_ = new_n13328_ & new_n50793_;
  assign new_n51268_ = new_n13330_ & new_n50795_;
  assign new_n51269_ = ~new_n51267_ & ~new_n51268_;
  assign new_n51270_ = new_n13334_ & new_n50798_;
  assign new_n51271_ = new_n50793_ & new_n51173_;
  assign new_n51272_ = ~new_n51270_ & ~new_n51271_;
  assign new_n51273_ = new_n51269_ & new_n51272_;
  assign new_n51274_ = ~new_n51175_ & ~new_n51273_;
  assign ys__n33068 = new_n51266_ | new_n51274_;
  assign new_n51276_ = new_n45674_ & new_n51175_;
  assign new_n51277_ = new_n13328_ & new_n50806_;
  assign new_n51278_ = new_n13330_ & new_n50808_;
  assign new_n51279_ = ~new_n51277_ & ~new_n51278_;
  assign new_n51280_ = new_n13334_ & new_n50811_;
  assign new_n51281_ = new_n50806_ & new_n51173_;
  assign new_n51282_ = ~new_n51280_ & ~new_n51281_;
  assign new_n51283_ = new_n51279_ & new_n51282_;
  assign new_n51284_ = ~new_n51175_ & ~new_n51283_;
  assign ys__n33069 = new_n51276_ | new_n51284_;
  assign new_n51286_ = new_n45685_ & new_n51175_;
  assign new_n51287_ = new_n13328_ & new_n50819_;
  assign new_n51288_ = new_n13330_ & new_n50821_;
  assign new_n51289_ = ~new_n51287_ & ~new_n51288_;
  assign new_n51290_ = new_n13334_ & new_n50824_;
  assign new_n51291_ = new_n50819_ & new_n51173_;
  assign new_n51292_ = ~new_n51290_ & ~new_n51291_;
  assign new_n51293_ = new_n51289_ & new_n51292_;
  assign new_n51294_ = ~new_n51175_ & ~new_n51293_;
  assign ys__n33070 = new_n51286_ | new_n51294_;
  assign new_n51296_ = new_n45696_ & new_n51175_;
  assign new_n51297_ = new_n13328_ & new_n50832_;
  assign new_n51298_ = new_n13330_ & new_n50834_;
  assign new_n51299_ = ~new_n51297_ & ~new_n51298_;
  assign new_n51300_ = new_n13334_ & new_n50837_;
  assign new_n51301_ = new_n50832_ & new_n51173_;
  assign new_n51302_ = ~new_n51300_ & ~new_n51301_;
  assign new_n51303_ = new_n51299_ & new_n51302_;
  assign new_n51304_ = ~new_n51175_ & ~new_n51303_;
  assign ys__n33071 = new_n51296_ | new_n51304_;
  assign new_n51306_ = new_n45707_ & new_n51175_;
  assign new_n51307_ = new_n13328_ & new_n50845_;
  assign new_n51308_ = new_n13330_ & new_n50847_;
  assign new_n51309_ = ~new_n51307_ & ~new_n51308_;
  assign new_n51310_ = new_n13334_ & new_n50850_;
  assign new_n51311_ = new_n50845_ & new_n51173_;
  assign new_n51312_ = ~new_n51310_ & ~new_n51311_;
  assign new_n51313_ = new_n51309_ & new_n51312_;
  assign new_n51314_ = ~new_n51175_ & ~new_n51313_;
  assign ys__n33072 = new_n51306_ | new_n51314_;
  assign new_n51316_ = new_n45720_ & new_n51175_;
  assign new_n51317_ = new_n13328_ & new_n50858_;
  assign new_n51318_ = new_n13330_ & new_n50860_;
  assign new_n51319_ = ~new_n51317_ & ~new_n51318_;
  assign new_n51320_ = new_n13334_ & new_n50863_;
  assign new_n51321_ = new_n50858_ & new_n51173_;
  assign new_n51322_ = ~new_n51320_ & ~new_n51321_;
  assign new_n51323_ = new_n51319_ & new_n51322_;
  assign new_n51324_ = ~new_n51175_ & ~new_n51323_;
  assign ys__n33073 = new_n51316_ | new_n51324_;
  assign new_n51326_ = new_n45731_ & new_n51175_;
  assign new_n51327_ = new_n13328_ & new_n50871_;
  assign new_n51328_ = new_n13330_ & new_n50873_;
  assign new_n51329_ = ~new_n51327_ & ~new_n51328_;
  assign new_n51330_ = new_n13334_ & new_n50876_;
  assign new_n51331_ = new_n50871_ & new_n51173_;
  assign new_n51332_ = ~new_n51330_ & ~new_n51331_;
  assign new_n51333_ = new_n51329_ & new_n51332_;
  assign new_n51334_ = ~new_n51175_ & ~new_n51333_;
  assign ys__n33074 = new_n51326_ | new_n51334_;
  assign new_n51336_ = new_n18041_ & new_n51175_;
  assign new_n51337_ = new_n13328_ & new_n50884_;
  assign new_n51338_ = new_n13330_ & new_n50886_;
  assign new_n51339_ = ~new_n51337_ & ~new_n51338_;
  assign new_n51340_ = new_n13334_ & new_n50889_;
  assign new_n51341_ = new_n50884_ & new_n51173_;
  assign new_n51342_ = ~new_n51340_ & ~new_n51341_;
  assign new_n51343_ = new_n51339_ & new_n51342_;
  assign new_n51344_ = ~new_n51175_ & ~new_n51343_;
  assign ys__n33075 = new_n51336_ | new_n51344_;
  assign new_n51346_ = new_n13267_ & new_n51175_;
  assign new_n51347_ = new_n13328_ & new_n50897_;
  assign new_n51348_ = new_n13330_ & new_n50899_;
  assign new_n51349_ = ~new_n51347_ & ~new_n51348_;
  assign new_n51350_ = new_n13334_ & new_n50902_;
  assign new_n51351_ = new_n50897_ & new_n51173_;
  assign new_n51352_ = ~new_n51350_ & ~new_n51351_;
  assign new_n51353_ = new_n51349_ & new_n51352_;
  assign new_n51354_ = ~new_n51175_ & ~new_n51353_;
  assign ys__n33076 = new_n51346_ | new_n51354_;
  assign new_n51356_ = new_n13249_ & new_n51175_;
  assign new_n51357_ = new_n13328_ & new_n50910_;
  assign new_n51358_ = new_n13330_ & new_n50912_;
  assign new_n51359_ = ~new_n51357_ & ~new_n51358_;
  assign new_n51360_ = new_n13334_ & new_n50915_;
  assign new_n51361_ = new_n50910_ & new_n51173_;
  assign new_n51362_ = ~new_n51360_ & ~new_n51361_;
  assign new_n51363_ = new_n51359_ & new_n51362_;
  assign new_n51364_ = ~new_n51175_ & ~new_n51363_;
  assign ys__n33077 = new_n51356_ | new_n51364_;
  assign new_n51366_ = new_n13191_ & new_n51175_;
  assign new_n51367_ = new_n13328_ & new_n50923_;
  assign new_n51368_ = new_n13330_ & new_n50925_;
  assign new_n51369_ = ~new_n51367_ & ~new_n51368_;
  assign new_n51370_ = new_n13334_ & new_n50928_;
  assign new_n51371_ = new_n50923_ & new_n51173_;
  assign new_n51372_ = ~new_n51370_ & ~new_n51371_;
  assign new_n51373_ = new_n51369_ & new_n51372_;
  assign new_n51374_ = ~new_n51175_ & ~new_n51373_;
  assign ys__n33078 = new_n51366_ | new_n51374_;
  assign new_n51376_ = new_n11754_ & new_n51175_;
  assign new_n51377_ = new_n13328_ & new_n50936_;
  assign new_n51378_ = new_n13330_ & new_n50938_;
  assign new_n51379_ = ~new_n51377_ & ~new_n51378_;
  assign new_n51380_ = new_n13334_ & new_n50941_;
  assign new_n51381_ = new_n50936_ & new_n51173_;
  assign new_n51382_ = ~new_n51380_ & ~new_n51381_;
  assign new_n51383_ = new_n51379_ & new_n51382_;
  assign new_n51384_ = ~new_n51175_ & ~new_n51383_;
  assign ys__n33079 = new_n51376_ | new_n51384_;
  assign new_n51386_ = ys__n17803 & new_n13372_;
  assign new_n51387_ = new_n13371_ & ~new_n25394_;
  assign new_n51388_ = ~new_n51386_ & ~new_n51387_;
  assign ys__n33178 = ys__n920 & ~new_n51388_;
  assign new_n51390_ = ys__n17804 & ~ys__n30553;
  assign new_n51391_ = ys__n30553 & ~new_n41063_;
  assign new_n51392_ = ~new_n51390_ & ~new_n51391_;
  assign new_n51393_ = new_n13372_ & ~new_n51392_;
  assign new_n51394_ = new_n13371_ & ~new_n25463_;
  assign new_n51395_ = ~new_n51393_ & ~new_n51394_;
  assign ys__n33179 = ys__n920 & ~new_n51395_;
  assign new_n51397_ = ys__n17806 & ~ys__n30553;
  assign new_n51398_ = ys__n30553 & ~new_n41090_;
  assign new_n51399_ = ~new_n51397_ & ~new_n51398_;
  assign new_n51400_ = new_n13372_ & ~new_n51399_;
  assign new_n51401_ = new_n13371_ & ~new_n25535_;
  assign new_n51402_ = ~new_n51400_ & ~new_n51401_;
  assign ys__n33180 = ys__n920 & ~new_n51402_;
  assign new_n51404_ = ys__n17807 & ~ys__n30553;
  assign new_n51405_ = ys__n30553 & ~new_n41117_;
  assign new_n51406_ = ~new_n51404_ & ~new_n51405_;
  assign new_n51407_ = new_n13372_ & ~new_n51406_;
  assign new_n51408_ = new_n13371_ & ~new_n25610_;
  assign new_n51409_ = ~new_n51407_ & ~new_n51408_;
  assign ys__n33181 = ys__n920 & ~new_n51409_;
  assign new_n51411_ = ys__n17809 & ~ys__n30553;
  assign new_n51412_ = ys__n30553 & ~new_n41142_;
  assign new_n51413_ = ~new_n51411_ & ~new_n51412_;
  assign new_n51414_ = new_n13372_ & ~new_n51413_;
  assign new_n51415_ = new_n13371_ & ~new_n25687_;
  assign new_n51416_ = ~new_n51414_ & ~new_n51415_;
  assign ys__n33182 = ys__n920 & ~new_n51416_;
  assign new_n51418_ = ys__n17810 & ~ys__n30553;
  assign new_n51419_ = ys__n30553 & ~new_n41168_;
  assign new_n51420_ = ~new_n51418_ & ~new_n51419_;
  assign new_n51421_ = new_n13372_ & ~new_n51420_;
  assign new_n51422_ = new_n13371_ & ~new_n25763_;
  assign new_n51423_ = ~new_n51421_ & ~new_n51422_;
  assign ys__n33183 = ys__n920 & ~new_n51423_;
  assign new_n51425_ = ys__n17812 & ~ys__n30553;
  assign new_n51426_ = ys__n30553 & ~new_n41197_;
  assign new_n51427_ = ~new_n51425_ & ~new_n51426_;
  assign new_n51428_ = new_n13372_ & ~new_n51427_;
  assign new_n51429_ = new_n13371_ & ~new_n25843_;
  assign new_n51430_ = ~new_n51428_ & ~new_n51429_;
  assign ys__n33184 = ys__n920 & ~new_n51430_;
  assign new_n51432_ = ys__n17813 & ~ys__n30553;
  assign new_n51433_ = ys__n30553 & ~new_n41226_;
  assign new_n51434_ = ~new_n51432_ & ~new_n51433_;
  assign new_n51435_ = new_n13372_ & ~new_n51434_;
  assign new_n51436_ = new_n13371_ & ~new_n25919_;
  assign new_n51437_ = ~new_n51435_ & ~new_n51436_;
  assign ys__n33185 = ys__n920 & ~new_n51437_;
  assign new_n51439_ = ys__n17815 & ~ys__n30553;
  assign new_n51440_ = ys__n30553 & ~new_n41254_;
  assign new_n51441_ = ~new_n51439_ & ~new_n51440_;
  assign new_n51442_ = new_n13372_ & ~new_n51441_;
  assign new_n51443_ = new_n13371_ & ~new_n26000_;
  assign new_n51444_ = ~new_n51442_ & ~new_n51443_;
  assign ys__n33186 = ys__n920 & ~new_n51444_;
  assign new_n51446_ = ys__n17816 & ~ys__n30553;
  assign new_n51447_ = ys__n30553 & ~new_n41280_;
  assign new_n51448_ = ~new_n51446_ & ~new_n51447_;
  assign new_n51449_ = new_n13372_ & ~new_n51448_;
  assign new_n51450_ = new_n13371_ & ~new_n26076_;
  assign new_n51451_ = ~new_n51449_ & ~new_n51450_;
  assign ys__n33187 = ys__n920 & ~new_n51451_;
  assign new_n51453_ = ys__n17818 & ~ys__n30553;
  assign new_n51454_ = ys__n30553 & ~new_n41309_;
  assign new_n51455_ = ~new_n51453_ & ~new_n51454_;
  assign new_n51456_ = new_n13372_ & ~new_n51455_;
  assign new_n51457_ = new_n13371_ & ~new_n26156_;
  assign new_n51458_ = ~new_n51456_ & ~new_n51457_;
  assign ys__n33188 = ys__n920 & ~new_n51458_;
  assign new_n51460_ = ys__n17819 & ~ys__n30553;
  assign new_n51461_ = ys__n30553 & ~new_n41338_;
  assign new_n51462_ = ~new_n51460_ & ~new_n51461_;
  assign new_n51463_ = new_n13372_ & ~new_n51462_;
  assign new_n51464_ = new_n13371_ & ~new_n26232_;
  assign new_n51465_ = ~new_n51463_ & ~new_n51464_;
  assign ys__n33189 = ys__n920 & ~new_n51465_;
  assign new_n51467_ = ys__n17821 & ~ys__n30553;
  assign new_n51468_ = ys__n30553 & ~new_n41367_;
  assign new_n51469_ = ~new_n51467_ & ~new_n51468_;
  assign new_n51470_ = new_n13372_ & ~new_n51469_;
  assign new_n51471_ = new_n13371_ & ~new_n26316_;
  assign new_n51472_ = ~new_n51470_ & ~new_n51471_;
  assign ys__n33190 = ys__n920 & ~new_n51472_;
  assign new_n51474_ = ys__n17822 & ~ys__n30553;
  assign new_n51475_ = ys__n30553 & ~new_n41396_;
  assign new_n51476_ = ~new_n51474_ & ~new_n51475_;
  assign new_n51477_ = new_n13372_ & ~new_n51476_;
  assign new_n51478_ = new_n13371_ & ~new_n26392_;
  assign new_n51479_ = ~new_n51477_ & ~new_n51478_;
  assign ys__n33191 = ys__n920 & ~new_n51479_;
  assign new_n51481_ = ys__n17824 & ~ys__n30553;
  assign new_n51482_ = ys__n30553 & ~new_n41425_;
  assign new_n51483_ = ~new_n51481_ & ~new_n51482_;
  assign new_n51484_ = new_n13372_ & ~new_n51483_;
  assign new_n51485_ = new_n13371_ & ~new_n26472_;
  assign new_n51486_ = ~new_n51484_ & ~new_n51485_;
  assign ys__n33192 = ys__n920 & ~new_n51486_;
  assign new_n51488_ = ys__n17825 & ~ys__n30553;
  assign new_n51489_ = ys__n30553 & ~new_n41454_;
  assign new_n51490_ = ~new_n51488_ & ~new_n51489_;
  assign new_n51491_ = new_n13372_ & ~new_n51490_;
  assign new_n51492_ = new_n13371_ & ~new_n26546_;
  assign new_n51493_ = ~new_n51491_ & ~new_n51492_;
  assign ys__n33193 = ys__n920 & ~new_n51493_;
  assign new_n51495_ = ys__n17827 & ~ys__n30553;
  assign new_n51496_ = ys__n30553 & ~new_n41482_;
  assign new_n51497_ = ~new_n51495_ & ~new_n51496_;
  assign new_n51498_ = new_n13372_ & ~new_n51497_;
  assign new_n51499_ = new_n13371_ & ~new_n25361_;
  assign new_n51500_ = ~new_n51498_ & ~new_n51499_;
  assign ys__n33194 = ys__n920 & ~new_n51500_;
  assign new_n51502_ = ys__n17828 & ~ys__n30553;
  assign new_n51503_ = ys__n30553 & ~new_n41508_;
  assign new_n51504_ = ~new_n51502_ & ~new_n51503_;
  assign new_n51505_ = new_n13372_ & ~new_n51504_;
  assign new_n51506_ = new_n13371_ & ~new_n25440_;
  assign new_n51507_ = ~new_n51505_ & ~new_n51506_;
  assign ys__n33195 = ys__n920 & ~new_n51507_;
  assign new_n51509_ = ys__n17830 & ~ys__n30553;
  assign new_n51510_ = ys__n30553 & ~new_n41543_;
  assign new_n51511_ = ~new_n51509_ & ~new_n51510_;
  assign new_n51512_ = new_n13372_ & ~new_n51511_;
  assign new_n51513_ = new_n13371_ & ~new_n25512_;
  assign new_n51514_ = ~new_n51512_ & ~new_n51513_;
  assign ys__n33196 = ys__n920 & ~new_n51514_;
  assign new_n51516_ = ys__n17831 & ~ys__n30553;
  assign new_n51517_ = ys__n30553 & ~new_n41578_;
  assign new_n51518_ = ~new_n51516_ & ~new_n51517_;
  assign new_n51519_ = new_n13372_ & ~new_n51518_;
  assign new_n51520_ = new_n13371_ & ~new_n25585_;
  assign new_n51521_ = ~new_n51519_ & ~new_n51520_;
  assign ys__n33197 = ys__n920 & ~new_n51521_;
  assign new_n51523_ = ys__n17833 & ~ys__n30553;
  assign new_n51524_ = ys__n30553 & ~new_n41613_;
  assign new_n51525_ = ~new_n51523_ & ~new_n51524_;
  assign new_n51526_ = new_n13372_ & ~new_n51525_;
  assign new_n51527_ = new_n13371_ & ~new_n25664_;
  assign new_n51528_ = ~new_n51526_ & ~new_n51527_;
  assign ys__n33198 = ys__n920 & ~new_n51528_;
  assign new_n51530_ = ys__n17834 & ~ys__n30553;
  assign new_n51531_ = ys__n30553 & ~new_n41648_;
  assign new_n51532_ = ~new_n51530_ & ~new_n51531_;
  assign new_n51533_ = new_n13372_ & ~new_n51532_;
  assign new_n51534_ = new_n13371_ & ~new_n25737_;
  assign new_n51535_ = ~new_n51533_ & ~new_n51534_;
  assign ys__n33199 = ys__n920 & ~new_n51535_;
  assign new_n51537_ = ys__n17836 & ~ys__n30553;
  assign new_n51538_ = ys__n30553 & ~new_n41686_;
  assign new_n51539_ = ~new_n51537_ & ~new_n51538_;
  assign new_n51540_ = new_n13372_ & ~new_n51539_;
  assign new_n51541_ = new_n13371_ & ~new_n25817_;
  assign new_n51542_ = ~new_n51540_ & ~new_n51541_;
  assign ys__n33200 = ys__n920 & ~new_n51542_;
  assign new_n51544_ = ys__n17837 & ~ys__n30553;
  assign new_n51545_ = ys__n30553 & ~new_n41724_;
  assign new_n51546_ = ~new_n51544_ & ~new_n51545_;
  assign new_n51547_ = new_n13372_ & ~new_n51546_;
  assign new_n51548_ = new_n13371_ & ~new_n25893_;
  assign new_n51549_ = ~new_n51547_ & ~new_n51548_;
  assign ys__n33201 = ys__n920 & ~new_n51549_;
  assign new_n51551_ = ys__n17839 & ~ys__n30553;
  assign new_n51552_ = ys__n30553 & ~new_n41762_;
  assign new_n51553_ = ~new_n51551_ & ~new_n51552_;
  assign new_n51554_ = new_n13372_ & ~new_n51553_;
  assign new_n51555_ = new_n13371_ & ~new_n25977_;
  assign new_n51556_ = ~new_n51554_ & ~new_n51555_;
  assign ys__n33202 = ys__n920 & ~new_n51556_;
  assign new_n51558_ = ys__n17840 & ~ys__n30553;
  assign new_n51559_ = ys__n30553 & ~new_n41797_;
  assign new_n51560_ = ~new_n51558_ & ~new_n51559_;
  assign new_n51561_ = new_n13372_ & ~new_n51560_;
  assign new_n51562_ = new_n13371_ & ~new_n26050_;
  assign new_n51563_ = ~new_n51561_ & ~new_n51562_;
  assign ys__n33203 = ys__n920 & ~new_n51563_;
  assign new_n51565_ = ys__n17842 & ~ys__n30553;
  assign new_n51566_ = ys__n30553 & ~new_n41835_;
  assign new_n51567_ = ~new_n51565_ & ~new_n51566_;
  assign new_n51568_ = new_n13372_ & ~new_n51567_;
  assign new_n51569_ = new_n13371_ & ~new_n26130_;
  assign new_n51570_ = ~new_n51568_ & ~new_n51569_;
  assign ys__n33204 = ys__n920 & ~new_n51570_;
  assign new_n51572_ = ys__n17843 & ~ys__n30553;
  assign new_n51573_ = ys__n30553 & ~new_n41873_;
  assign new_n51574_ = ~new_n51572_ & ~new_n51573_;
  assign new_n51575_ = new_n13372_ & ~new_n51574_;
  assign new_n51576_ = new_n13371_ & ~new_n26206_;
  assign new_n51577_ = ~new_n51575_ & ~new_n51576_;
  assign ys__n33205 = ys__n920 & ~new_n51577_;
  assign new_n51579_ = ys__n17845 & ~ys__n30553;
  assign new_n51580_ = ys__n30553 & ~new_n41911_;
  assign new_n51581_ = ~new_n51579_ & ~new_n51580_;
  assign new_n51582_ = new_n13372_ & ~new_n51581_;
  assign new_n51583_ = new_n13371_ & ~new_n26290_;
  assign new_n51584_ = ~new_n51582_ & ~new_n51583_;
  assign ys__n33206 = ys__n920 & ~new_n51584_;
  assign new_n51586_ = ys__n17846 & ~ys__n30553;
  assign new_n51587_ = ys__n30553 & ~new_n41948_;
  assign new_n51588_ = ~new_n51586_ & ~new_n51587_;
  assign new_n51589_ = new_n13372_ & ~new_n51588_;
  assign new_n51590_ = new_n13371_ & ~new_n26366_;
  assign new_n51591_ = ~new_n51589_ & ~new_n51590_;
  assign ys__n33207 = ys__n920 & ~new_n51591_;
  assign new_n51593_ = ys__n17848 & ~ys__n30553;
  assign new_n51594_ = ys__n30553 & ~new_n41986_;
  assign new_n51595_ = ~new_n51593_ & ~new_n51594_;
  assign new_n51596_ = new_n13372_ & ~new_n51595_;
  assign new_n51597_ = new_n13371_ & ~new_n26446_;
  assign new_n51598_ = ~new_n51596_ & ~new_n51597_;
  assign ys__n33208 = ys__n920 & ~new_n51598_;
  assign new_n51600_ = ys__n17849 & ~ys__n30553;
  assign new_n51601_ = ys__n30553 & ~new_n42023_;
  assign new_n51602_ = ~new_n51600_ & ~new_n51601_;
  assign new_n51603_ = new_n13372_ & ~new_n51602_;
  assign new_n51604_ = new_n13371_ & ~new_n26520_;
  assign new_n51605_ = ~new_n51603_ & ~new_n51604_;
  assign ys__n33209 = ys__n920 & ~new_n51605_;
  assign new_n51607_ = ~ys__n740 & new_n13342_;
  assign new_n51608_ = ~ys__n23850 & new_n13339_;
  assign new_n51609_ = ~new_n51607_ & ~new_n51608_;
  assign new_n51610_ = ~new_n13346_ & ~new_n51609_;
  assign ys__n33211 = new_n13346_ | new_n51610_;
  assign new_n51612_ = new_n12309_ & ~new_n12762_;
  assign ys__n33366 = new_n11954_ & new_n51612_;
  assign ys__n33438 = ~ys__n1084 & ~new_n11979_;
  assign new_n51615_ = ~ys__n30216 & ~ys__n30219;
  assign new_n51616_ = new_n23621_ & new_n51615_;
  assign new_n51617_ = ys__n1106 & ~new_n51616_;
  assign new_n51618_ = ~ys__n24464 & ~ys__n24483;
  assign new_n51619_ = ~ys__n38649 & new_n51618_;
  assign new_n51620_ = ~ys__n1116 & ~ys__n1119;
  assign new_n51621_ = ~ys__n24461 & ~ys__n24463;
  assign new_n51622_ = new_n51620_ & new_n51621_;
  assign new_n51623_ = new_n15125_ & new_n23587_;
  assign new_n51624_ = new_n51622_ & new_n51623_;
  assign new_n51625_ = new_n51619_ & new_n51624_;
  assign ys__n33454 = ~new_n51617_ & new_n51625_;
  assign new_n51627_ = ys__n1153 & ys__n33515;
  assign new_n51628_ = new_n17356_ & new_n51615_;
  assign new_n51629_ = ys__n1151 & ~new_n51628_;
  assign new_n51630_ = ys__n33515 & new_n51629_;
  assign new_n51631_ = new_n24597_ & ~new_n51630_;
  assign ys__n33514 = ~new_n51627_ & new_n51631_;
  assign ys__n34952 = ~ys__n18166 & ~ys__n18165;
  assign ys__n34953 = ~ys__n2651 & ~ys__n18166;
  assign new_n51635_ = ys__n18317 & new_n13407_;
  assign ys__n34962 = new_n13418_ & new_n51635_;
  assign new_n51637_ = ys__n46248 & new_n44610_;
  assign new_n51638_ = ~ys__n46242 & ~ys__n46244;
  assign new_n51639_ = ~ys__n46245 & ~ys__n46247;
  assign new_n51640_ = new_n51638_ & new_n51639_;
  assign ys__n35052 = new_n51637_ | ~new_n51640_;
  assign new_n51642_ = ys__n33081 & ~ys__n33080;
  assign new_n51643_ = ~ys__n33081 & ys__n33080;
  assign ys__n35144 = new_n51642_ | new_n51643_;
  assign new_n51645_ = ~ys__n33081 & ~ys__n33080;
  assign new_n51646_ = ys__n33082 & new_n51645_;
  assign new_n51647_ = ~ys__n33082 & ~new_n51645_;
  assign ys__n35146 = new_n51646_ | new_n51647_;
  assign new_n51649_ = ~ys__n33082 & new_n51645_;
  assign new_n51650_ = ys__n33083 & new_n51649_;
  assign new_n51651_ = ~ys__n33083 & ~new_n51649_;
  assign ys__n35148 = new_n51650_ | new_n51651_;
  assign new_n51653_ = ~ys__n33082 & ~ys__n33083;
  assign new_n51654_ = new_n51645_ & new_n51653_;
  assign new_n51655_ = ys__n33084 & new_n51654_;
  assign new_n51656_ = ~ys__n33084 & ~new_n51654_;
  assign ys__n35150 = new_n51655_ | new_n51656_;
  assign new_n51658_ = ~ys__n33084 & new_n51654_;
  assign new_n51659_ = ys__n33085 & new_n51658_;
  assign new_n51660_ = ~ys__n33085 & ~new_n51658_;
  assign ys__n35152 = new_n51659_ | new_n51660_;
  assign new_n51662_ = ~ys__n33085 & ~ys__n33084;
  assign new_n51663_ = new_n51654_ & new_n51662_;
  assign new_n51664_ = ys__n33086 & new_n51663_;
  assign new_n51665_ = ~ys__n33086 & ~new_n51663_;
  assign ys__n35154 = new_n51664_ | new_n51665_;
  assign new_n51667_ = ~ys__n33086 & new_n51663_;
  assign new_n51668_ = ys__n33087 & new_n51667_;
  assign new_n51669_ = ~ys__n33087 & ~new_n51667_;
  assign ys__n35156 = new_n51668_ | new_n51669_;
  assign new_n51671_ = ~ys__n33087 & ~ys__n33086;
  assign new_n51672_ = new_n51662_ & new_n51671_;
  assign new_n51673_ = new_n51654_ & new_n51672_;
  assign new_n51674_ = ys__n33088 & new_n51673_;
  assign new_n51675_ = ~ys__n33088 & ~new_n51673_;
  assign ys__n35158 = new_n51674_ | new_n51675_;
  assign new_n51677_ = ~ys__n33088 & new_n51673_;
  assign new_n51678_ = ys__n33089 & new_n51677_;
  assign new_n51679_ = ~ys__n33089 & ~new_n51677_;
  assign ys__n35160 = new_n51678_ | new_n51679_;
  assign new_n51681_ = ~ys__n33089 & ~ys__n33088;
  assign new_n51682_ = new_n51673_ & new_n51681_;
  assign new_n51683_ = ys__n33090 & new_n51682_;
  assign new_n51684_ = ~ys__n33090 & ~new_n51682_;
  assign ys__n35162 = new_n51683_ | new_n51684_;
  assign new_n51686_ = ~ys__n33090 & new_n51682_;
  assign new_n51687_ = ys__n33091 & new_n51686_;
  assign new_n51688_ = ~ys__n33091 & ~new_n51686_;
  assign ys__n35164 = new_n51687_ | new_n51688_;
  assign new_n51690_ = ~ys__n33091 & ~ys__n33090;
  assign new_n51691_ = new_n51681_ & new_n51690_;
  assign new_n51692_ = new_n51673_ & new_n51691_;
  assign new_n51693_ = ys__n33092 & new_n51692_;
  assign new_n51694_ = ~ys__n33092 & ~new_n51692_;
  assign ys__n35166 = new_n51693_ | new_n51694_;
  assign new_n51696_ = ~ys__n33092 & new_n51692_;
  assign new_n51697_ = ys__n33093 & new_n51696_;
  assign new_n51698_ = ~ys__n33093 & ~new_n51696_;
  assign ys__n35168 = new_n51697_ | new_n51698_;
  assign new_n51700_ = ~ys__n33093 & ~ys__n33092;
  assign new_n51701_ = new_n51692_ & new_n51700_;
  assign new_n51702_ = ys__n33094 & new_n51701_;
  assign new_n51703_ = ~ys__n33094 & ~new_n51701_;
  assign ys__n35170 = new_n51702_ | new_n51703_;
  assign new_n51705_ = ~ys__n33094 & new_n51701_;
  assign new_n51706_ = ys__n33095 & new_n51705_;
  assign new_n51707_ = ~ys__n33095 & ~new_n51705_;
  assign ys__n35172 = new_n51706_ | new_n51707_;
  assign new_n51709_ = ~ys__n33095 & ~ys__n33094;
  assign new_n51710_ = new_n51700_ & new_n51709_;
  assign new_n51711_ = new_n51691_ & new_n51710_;
  assign new_n51712_ = new_n51673_ & new_n51711_;
  assign new_n51713_ = ys__n33096 & new_n51712_;
  assign new_n51714_ = ~ys__n33096 & ~new_n51712_;
  assign ys__n35174 = new_n51713_ | new_n51714_;
  assign new_n51716_ = ~ys__n33096 & new_n51712_;
  assign new_n51717_ = ys__n33097 & new_n51716_;
  assign new_n51718_ = ~ys__n33097 & ~new_n51716_;
  assign ys__n35176 = new_n51717_ | new_n51718_;
  assign new_n51720_ = ~ys__n33096 & ~ys__n33097;
  assign new_n51721_ = new_n51712_ & new_n51720_;
  assign new_n51722_ = ys__n33098 & new_n51721_;
  assign new_n51723_ = ~ys__n33098 & ~new_n51721_;
  assign ys__n35178 = new_n51722_ | new_n51723_;
  assign new_n51725_ = ~ys__n33098 & new_n51721_;
  assign new_n51726_ = ys__n33099 & new_n51725_;
  assign new_n51727_ = ~ys__n33099 & ~new_n51725_;
  assign ys__n35180 = new_n51726_ | new_n51727_;
  assign new_n51729_ = ~ys__n33098 & ~ys__n33099;
  assign new_n51730_ = new_n51720_ & new_n51729_;
  assign new_n51731_ = new_n51712_ & new_n51730_;
  assign new_n51732_ = ys__n33100 & new_n51731_;
  assign new_n51733_ = ~ys__n33100 & ~new_n51731_;
  assign ys__n35182 = new_n51732_ | new_n51733_;
  assign new_n51735_ = ~ys__n33100 & new_n51731_;
  assign new_n51736_ = ys__n33101 & new_n51735_;
  assign new_n51737_ = ~ys__n33101 & ~new_n51735_;
  assign ys__n35184 = new_n51736_ | new_n51737_;
  assign new_n51739_ = ~ys__n33100 & ~ys__n33101;
  assign new_n51740_ = new_n51731_ & new_n51739_;
  assign new_n51741_ = ys__n33102 & new_n51740_;
  assign new_n51742_ = ~ys__n33102 & ~new_n51740_;
  assign ys__n35186 = new_n51741_ | new_n51742_;
  assign new_n51744_ = ~ys__n33102 & new_n51740_;
  assign new_n51745_ = ys__n33103 & new_n51744_;
  assign new_n51746_ = ~ys__n33103 & ~new_n51744_;
  assign ys__n35188 = new_n51745_ | new_n51746_;
  assign new_n51748_ = ~ys__n33102 & ~ys__n33103;
  assign new_n51749_ = new_n51739_ & new_n51748_;
  assign new_n51750_ = new_n51730_ & new_n51749_;
  assign new_n51751_ = new_n51712_ & new_n51750_;
  assign new_n51752_ = ys__n33104 & new_n51751_;
  assign new_n51753_ = ~ys__n33104 & ~new_n51751_;
  assign ys__n35190 = new_n51752_ | new_n51753_;
  assign new_n51755_ = ~ys__n33104 & new_n51751_;
  assign new_n51756_ = ys__n33105 & new_n51755_;
  assign new_n51757_ = ~ys__n33105 & ~new_n51755_;
  assign ys__n35192 = new_n51756_ | new_n51757_;
  assign new_n51759_ = ~ys__n33104 & ~ys__n33105;
  assign new_n51760_ = new_n51751_ & new_n51759_;
  assign new_n51761_ = ys__n33106 & new_n51760_;
  assign new_n51762_ = ~ys__n33106 & ~new_n51760_;
  assign ys__n35194 = new_n51761_ | new_n51762_;
  assign new_n51764_ = ~ys__n33106 & new_n51760_;
  assign new_n51765_ = ys__n33107 & new_n51764_;
  assign new_n51766_ = ~ys__n33107 & ~new_n51764_;
  assign ys__n35196 = new_n51765_ | new_n51766_;
  assign new_n51768_ = ~ys__n33106 & ~ys__n33107;
  assign new_n51769_ = new_n51759_ & new_n51768_;
  assign new_n51770_ = new_n51751_ & new_n51769_;
  assign new_n51771_ = ys__n33108 & new_n51770_;
  assign new_n51772_ = ~ys__n33108 & ~new_n51770_;
  assign ys__n35198 = new_n51771_ | new_n51772_;
  assign new_n51774_ = ~ys__n33108 & new_n51770_;
  assign new_n51775_ = ys__n33109 & new_n51774_;
  assign new_n51776_ = ~ys__n33109 & ~new_n51774_;
  assign ys__n35200 = new_n51775_ | new_n51776_;
  assign new_n51778_ = ~ys__n33108 & ~ys__n33109;
  assign new_n51779_ = new_n51770_ & new_n51778_;
  assign new_n51780_ = ys__n33110 & new_n51779_;
  assign new_n51781_ = ~ys__n33110 & ~new_n51779_;
  assign ys__n35202 = new_n51780_ | new_n51781_;
  assign new_n51783_ = ~ys__n33110 & new_n51779_;
  assign new_n51784_ = ys__n33111 & new_n51783_;
  assign new_n51785_ = ~ys__n33111 & ~new_n51783_;
  assign ys__n35204 = new_n51784_ | new_n51785_;
  assign new_n51787_ = ~ys__n33110 & ~ys__n33111;
  assign new_n51788_ = new_n51778_ & new_n51787_;
  assign new_n51789_ = new_n51769_ & new_n51788_;
  assign new_n51790_ = new_n51712_ & new_n51789_;
  assign new_n51791_ = new_n51750_ & new_n51790_;
  assign new_n51792_ = ys__n30668 & new_n51791_;
  assign new_n51793_ = ~ys__n30668 & ~new_n51791_;
  assign ys__n35206 = new_n51792_ | new_n51793_;
  assign new_n51795_ = ys__n456 & ~ys__n710;
  assign new_n51796_ = ~ys__n456 & ys__n710;
  assign ys__n35402 = new_n51795_ | new_n51796_;
  assign new_n51798_ = ~ys__n708 & new_n17630_;
  assign new_n51799_ = ys__n708 & ~new_n17630_;
  assign ys__n35404 = new_n51798_ | new_n51799_;
  assign new_n51801_ = ys__n708 & new_n17630_;
  assign new_n51802_ = ~ys__n706 & new_n51801_;
  assign new_n51803_ = ys__n706 & ~new_n51801_;
  assign ys__n35406 = new_n51802_ | new_n51803_;
  assign new_n51805_ = ~ys__n702 & new_n17632_;
  assign new_n51806_ = ys__n702 & ~new_n17632_;
  assign ys__n35408 = new_n51805_ | new_n51806_;
  assign new_n51808_ = ys__n702 & new_n17632_;
  assign new_n51809_ = ~ys__n700 & new_n51808_;
  assign new_n51810_ = ys__n700 & ~new_n51808_;
  assign ys__n35410 = new_n51809_ | new_n51810_;
  assign new_n51812_ = new_n17632_ & new_n17633_;
  assign new_n51813_ = ~ys__n704 & new_n51812_;
  assign new_n51814_ = ys__n704 & ~new_n51812_;
  assign ys__n35412 = new_n51813_ | new_n51814_;
  assign new_n51816_ = ys__n414 & ~ys__n728;
  assign new_n51817_ = ~ys__n414 & ys__n728;
  assign ys__n35706 = new_n51816_ | new_n51817_;
  assign new_n51819_ = ~ys__n726 & new_n17616_;
  assign new_n51820_ = ys__n726 & ~new_n17616_;
  assign ys__n35708 = new_n51819_ | new_n51820_;
  assign new_n51822_ = ys__n726 & new_n17616_;
  assign new_n51823_ = ~ys__n724 & new_n51822_;
  assign new_n51824_ = ys__n724 & ~new_n51822_;
  assign ys__n35710 = new_n51823_ | new_n51824_;
  assign new_n51826_ = ~ys__n720 & new_n17618_;
  assign new_n51827_ = ys__n720 & ~new_n17618_;
  assign ys__n35712 = new_n51826_ | new_n51827_;
  assign new_n51829_ = ys__n720 & new_n17618_;
  assign new_n51830_ = ~ys__n718 & new_n51829_;
  assign new_n51831_ = ys__n718 & ~new_n51829_;
  assign ys__n35714 = new_n51830_ | new_n51831_;
  assign new_n51833_ = new_n17618_ & new_n17619_;
  assign new_n51834_ = ~ys__n722 & new_n51833_;
  assign new_n51835_ = ys__n722 & ~new_n51833_;
  assign ys__n35716 = new_n51834_ | new_n51835_;
  assign new_n51837_ = ys__n3214 & ys__n19159;
  assign new_n51838_ = ~new_n12925_ & ~new_n51837_;
  assign ys__n37687 = new_n12934_ | ~new_n51838_;
  assign ys__n37695 = ~new_n13231_ & new_n13237_;
  assign ys__n37697 = ~new_n13232_ & new_n13237_;
  assign new_n51842_ = ys__n33313 & ~new_n13237_;
  assign new_n51843_ = ys__n3214 & ~new_n51842_;
  assign ys__n37699 = new_n18154_ | new_n51843_;
  assign new_n51845_ = ys__n33311 & ~ys__n33313;
  assign new_n51846_ = ~new_n13237_ & new_n51845_;
  assign new_n51847_ = ys__n18070 & ~new_n51846_;
  assign ys__n37702 = new_n12259_ | new_n51847_;
  assign new_n51849_ = ys__n33309 & ~ys__n33311;
  assign new_n51850_ = ~ys__n33313 & new_n51849_;
  assign new_n51851_ = ~new_n13237_ & new_n51850_;
  assign new_n51852_ = ys__n18071 & ~new_n51851_;
  assign ys__n37707 = new_n12256_ | new_n51852_;
  assign new_n51854_ = ~ys__n844 & ~ys__n37710;
  assign new_n51855_ = ~ys__n37712 & ys__n37713;
  assign ys__n37714 = new_n51854_ & new_n51855_;
  assign ys__n37731 = ys__n24112 & ~ys__n33317;
  assign ys__n37732 = ys__n18380 & ys__n33317;
  assign ys__n37733 = ys__n18383 & ys__n33317;
  assign new_n51860_ = ~ys__n37668 & ys__n37669;
  assign new_n51861_ = ys__n37668 & ~ys__n37669;
  assign new_n51862_ = ~new_n51860_ & ~new_n51861_;
  assign new_n51863_ = ~ys__n18393 & ~new_n51862_;
  assign new_n51864_ = ys__n18393 & ys__n27598;
  assign new_n51865_ = ~new_n51863_ & ~new_n51864_;
  assign ys__n37738 = ys__n33320 & ~new_n51865_;
  assign new_n51867_ = ys__n33318 & ~ys__n33320;
  assign new_n51868_ = ~new_n51865_ & new_n51867_;
  assign ys__n37739 = new_n34730_ | new_n51868_;
  assign new_n51870_ = ~ys__n33318 & ~ys__n33320;
  assign new_n51871_ = ~new_n51865_ & new_n51870_;
  assign new_n51872_ = ys__n18208 & new_n34827_;
  assign ys__n37741 = new_n51871_ | new_n51872_;
  assign new_n51874_ = ys__n812 & ~ys__n3250;
  assign new_n51875_ = ys__n19171 & ys__n18287;
  assign new_n51876_ = ~ys__n18284 & new_n51875_;
  assign new_n51877_ = ys__n18284 & ys__n18763;
  assign new_n51878_ = ~new_n51876_ & ~new_n51877_;
  assign new_n51879_ = ~ys__n18281 & ~new_n51878_;
  assign new_n51880_ = ys__n18281 & ys__n18652;
  assign new_n51881_ = ~new_n51879_ & ~new_n51880_;
  assign new_n51882_ = ~ys__n18278 & ~new_n51881_;
  assign new_n51883_ = ~ys__n18278 & ~new_n51882_;
  assign new_n51884_ = ~ys__n3252 & ~new_n51883_;
  assign new_n51885_ = new_n51874_ & new_n51884_;
  assign new_n51886_ = ys__n804 & ys__n806;
  assign new_n51887_ = ys__n808 & ys__n810;
  assign new_n51888_ = new_n51886_ & new_n51887_;
  assign new_n51889_ = ys__n796 & ys__n798;
  assign new_n51890_ = ys__n800 & ys__n802;
  assign new_n51891_ = new_n51889_ & new_n51890_;
  assign new_n51892_ = new_n51888_ & new_n51891_;
  assign ys__n37742 = new_n51885_ & new_n51892_;
  assign ys__n38180 = ys__n38179 | ys__n18088;
  assign new_n51895_ = ~ys__n240 & new_n34939_;
  assign new_n51896_ = ~new_n34939_ & new_n51895_;
  assign new_n51897_ = ~ys__n1535 & ~new_n51896_;
  assign new_n51898_ = ~ys__n1535 & ~new_n51897_;
  assign new_n51899_ = ys__n28243 & ~ys__n4566;
  assign ys__n38182 = ~new_n51898_ & new_n51899_;
  assign ys__n38184 = ys__n38183 & ~ys__n4566;
  assign ys__n38205 = ~ys__n23627 | ~ys__n738;
  assign new_n51903_ = ys__n45704 & new_n14079_;
  assign new_n51904_ = ys__n45541 & new_n14389_;
  assign new_n51905_ = ~new_n51903_ & ~new_n51904_;
  assign new_n51906_ = ys__n45377 & new_n14700_;
  assign new_n51907_ = ys__n45214 & new_n15010_;
  assign new_n51908_ = ~new_n51906_ & ~new_n51907_;
  assign new_n51909_ = new_n51905_ & new_n51908_;
  assign new_n51910_ = ~new_n15017_ & ~new_n51909_;
  assign new_n51911_ = ~ys__n38282 & ~ys__n38283;
  assign new_n51912_ = ~ys__n38286 & ~ys__n38300;
  assign new_n51913_ = new_n51911_ & new_n51912_;
  assign new_n51914_ = ~new_n51910_ & new_n51913_;
  assign ys__n38207 = ~ys__n4566 & ~new_n51914_;
  assign new_n51916_ = ys__n45771 & ys__n46074;
  assign new_n51917_ = ~ys__n45771 & ~ys__n46074;
  assign new_n51918_ = ~ys__n46116 & ~new_n51917_;
  assign new_n51919_ = ~new_n51916_ & new_n51918_;
  assign new_n51920_ = ys__n45774 & ys__n46076;
  assign new_n51921_ = ~ys__n45774 & ~ys__n46076;
  assign new_n51922_ = ~ys__n46117 & ~new_n51921_;
  assign new_n51923_ = ~new_n51920_ & new_n51922_;
  assign new_n51924_ = ~new_n51919_ & ~new_n51923_;
  assign new_n51925_ = ys__n45777 & ys__n46078;
  assign new_n51926_ = ~ys__n45777 & ~ys__n46078;
  assign new_n51927_ = ~ys__n46118 & ~new_n51926_;
  assign new_n51928_ = ~new_n51925_ & new_n51927_;
  assign new_n51929_ = ys__n45780 & ys__n46080;
  assign new_n51930_ = ~ys__n45780 & ~ys__n46080;
  assign new_n51931_ = ~ys__n46119 & ~new_n51930_;
  assign new_n51932_ = ~new_n51929_ & new_n51931_;
  assign new_n51933_ = ~new_n51928_ & ~new_n51932_;
  assign new_n51934_ = new_n51924_ & new_n51933_;
  assign new_n51935_ = ys__n45759 & ys__n46066;
  assign new_n51936_ = ~ys__n45759 & ~ys__n46066;
  assign new_n51937_ = ~ys__n46112 & ~new_n51936_;
  assign new_n51938_ = ~new_n51935_ & new_n51937_;
  assign new_n51939_ = ys__n45762 & ys__n46068;
  assign new_n51940_ = ~ys__n45762 & ~ys__n46068;
  assign new_n51941_ = ~ys__n46113 & ~new_n51940_;
  assign new_n51942_ = ~new_n51939_ & new_n51941_;
  assign new_n51943_ = ~new_n51938_ & ~new_n51942_;
  assign new_n51944_ = ys__n45765 & ys__n46070;
  assign new_n51945_ = ~ys__n45765 & ~ys__n46070;
  assign new_n51946_ = ~ys__n46114 & ~new_n51945_;
  assign new_n51947_ = ~new_n51944_ & new_n51946_;
  assign new_n51948_ = ys__n45768 & ys__n46072;
  assign new_n51949_ = ~ys__n45768 & ~ys__n46072;
  assign new_n51950_ = ~ys__n46115 & ~new_n51949_;
  assign new_n51951_ = ~new_n51948_ & new_n51950_;
  assign new_n51952_ = ~new_n51947_ & ~new_n51951_;
  assign new_n51953_ = new_n51943_ & new_n51952_;
  assign new_n51954_ = new_n51934_ & new_n51953_;
  assign new_n51955_ = ys__n45801 & ys__n46094;
  assign new_n51956_ = ~ys__n45801 & ~ys__n46094;
  assign new_n51957_ = ~ys__n46126 & ~new_n51956_;
  assign new_n51958_ = ~new_n51955_ & new_n51957_;
  assign new_n51959_ = ys__n45795 & ys__n46090;
  assign new_n51960_ = ~ys__n45795 & ~ys__n46090;
  assign new_n51961_ = ~ys__n46124 & ~new_n51960_;
  assign new_n51962_ = ~new_n51959_ & new_n51961_;
  assign new_n51963_ = ys__n45798 & ys__n46092;
  assign new_n51964_ = ~ys__n45798 & ~ys__n46092;
  assign new_n51965_ = ~ys__n46125 & ~new_n51964_;
  assign new_n51966_ = ~new_n51963_ & new_n51965_;
  assign new_n51967_ = ~new_n51962_ & ~new_n51966_;
  assign new_n51968_ = ~new_n51958_ & new_n51967_;
  assign new_n51969_ = ys__n45783 & ys__n46082;
  assign new_n51970_ = ~ys__n45783 & ~ys__n46082;
  assign new_n51971_ = ~ys__n46120 & ~new_n51970_;
  assign new_n51972_ = ~new_n51969_ & new_n51971_;
  assign new_n51973_ = ys__n45786 & ys__n46084;
  assign new_n51974_ = ~ys__n45786 & ~ys__n46084;
  assign new_n51975_ = ~ys__n46121 & ~new_n51974_;
  assign new_n51976_ = ~new_n51973_ & new_n51975_;
  assign new_n51977_ = ~new_n51972_ & ~new_n51976_;
  assign new_n51978_ = ys__n45789 & ys__n46086;
  assign new_n51979_ = ~ys__n45789 & ~ys__n46086;
  assign new_n51980_ = ~ys__n46122 & ~new_n51979_;
  assign new_n51981_ = ~new_n51978_ & new_n51980_;
  assign new_n51982_ = ys__n45792 & ys__n46088;
  assign new_n51983_ = ~ys__n45792 & ~ys__n46088;
  assign new_n51984_ = ~ys__n46123 & ~new_n51983_;
  assign new_n51985_ = ~new_n51982_ & new_n51984_;
  assign new_n51986_ = ~new_n51981_ & ~new_n51985_;
  assign new_n51987_ = new_n51977_ & new_n51986_;
  assign new_n51988_ = new_n51968_ & new_n51987_;
  assign new_n51989_ = new_n51954_ & new_n51988_;
  assign new_n51990_ = ys__n45723 & ys__n46042;
  assign new_n51991_ = ~ys__n45723 & ~ys__n46042;
  assign new_n51992_ = ~ys__n46100 & ~new_n51991_;
  assign new_n51993_ = ~new_n51990_ & new_n51992_;
  assign new_n51994_ = ys__n45726 & ys__n46044;
  assign new_n51995_ = ~ys__n45726 & ~ys__n46044;
  assign new_n51996_ = ~ys__n46101 & ~new_n51995_;
  assign new_n51997_ = ~new_n51994_ & new_n51996_;
  assign new_n51998_ = ~new_n51993_ & ~new_n51997_;
  assign new_n51999_ = ys__n45729 & ys__n46046;
  assign new_n52000_ = ~ys__n45729 & ~ys__n46046;
  assign new_n52001_ = ~ys__n46102 & ~new_n52000_;
  assign new_n52002_ = ~new_n51999_ & new_n52001_;
  assign new_n52003_ = ys__n45732 & ys__n46048;
  assign new_n52004_ = ~ys__n45732 & ~ys__n46048;
  assign new_n52005_ = ~ys__n46103 & ~new_n52004_;
  assign new_n52006_ = ~new_n52003_ & new_n52005_;
  assign new_n52007_ = ~new_n52002_ & ~new_n52006_;
  assign new_n52008_ = new_n51998_ & new_n52007_;
  assign new_n52009_ = ys__n45711 & ys__n46034;
  assign new_n52010_ = ~ys__n45711 & ~ys__n46034;
  assign new_n52011_ = ~ys__n46096 & ~new_n52010_;
  assign new_n52012_ = ~new_n52009_ & new_n52011_;
  assign new_n52013_ = ys__n45714 & ys__n46036;
  assign new_n52014_ = ~ys__n45714 & ~ys__n46036;
  assign new_n52015_ = ~ys__n46097 & ~new_n52014_;
  assign new_n52016_ = ~new_n52013_ & new_n52015_;
  assign new_n52017_ = ~new_n52012_ & ~new_n52016_;
  assign new_n52018_ = ys__n45717 & ys__n46038;
  assign new_n52019_ = ~ys__n45717 & ~ys__n46038;
  assign new_n52020_ = ~ys__n46098 & ~new_n52019_;
  assign new_n52021_ = ~new_n52018_ & new_n52020_;
  assign new_n52022_ = ys__n45720 & ys__n46040;
  assign new_n52023_ = ~ys__n45720 & ~ys__n46040;
  assign new_n52024_ = ~ys__n46099 & ~new_n52023_;
  assign new_n52025_ = ~new_n52022_ & new_n52024_;
  assign new_n52026_ = ~new_n52021_ & ~new_n52025_;
  assign new_n52027_ = new_n52017_ & new_n52026_;
  assign new_n52028_ = new_n52008_ & new_n52027_;
  assign new_n52029_ = ys__n45747 & ys__n46058;
  assign new_n52030_ = ~ys__n45747 & ~ys__n46058;
  assign new_n52031_ = ~ys__n46108 & ~new_n52030_;
  assign new_n52032_ = ~new_n52029_ & new_n52031_;
  assign new_n52033_ = ys__n45750 & ys__n46060;
  assign new_n52034_ = ~ys__n45750 & ~ys__n46060;
  assign new_n52035_ = ~ys__n46109 & ~new_n52034_;
  assign new_n52036_ = ~new_n52033_ & new_n52035_;
  assign new_n52037_ = ~new_n52032_ & ~new_n52036_;
  assign new_n52038_ = ys__n45753 & ys__n46062;
  assign new_n52039_ = ~ys__n45753 & ~ys__n46062;
  assign new_n52040_ = ~ys__n46110 & ~new_n52039_;
  assign new_n52041_ = ~new_n52038_ & new_n52040_;
  assign new_n52042_ = ys__n45756 & ys__n46064;
  assign new_n52043_ = ~ys__n45756 & ~ys__n46064;
  assign new_n52044_ = ~ys__n46111 & ~new_n52043_;
  assign new_n52045_ = ~new_n52042_ & new_n52044_;
  assign new_n52046_ = ~new_n52041_ & ~new_n52045_;
  assign new_n52047_ = new_n52037_ & new_n52046_;
  assign new_n52048_ = ys__n45735 & ys__n46050;
  assign new_n52049_ = ~ys__n45735 & ~ys__n46050;
  assign new_n52050_ = ~ys__n46104 & ~new_n52049_;
  assign new_n52051_ = ~new_n52048_ & new_n52050_;
  assign new_n52052_ = ys__n45738 & ys__n46052;
  assign new_n52053_ = ~ys__n45738 & ~ys__n46052;
  assign new_n52054_ = ~ys__n46105 & ~new_n52053_;
  assign new_n52055_ = ~new_n52052_ & new_n52054_;
  assign new_n52056_ = ~new_n52051_ & ~new_n52055_;
  assign new_n52057_ = ys__n45741 & ys__n46054;
  assign new_n52058_ = ~ys__n45741 & ~ys__n46054;
  assign new_n52059_ = ~ys__n46106 & ~new_n52058_;
  assign new_n52060_ = ~new_n52057_ & new_n52059_;
  assign new_n52061_ = ys__n45744 & ys__n46056;
  assign new_n52062_ = ~ys__n45744 & ~ys__n46056;
  assign new_n52063_ = ~ys__n46107 & ~new_n52062_;
  assign new_n52064_ = ~new_n52061_ & new_n52063_;
  assign new_n52065_ = ~new_n52060_ & ~new_n52064_;
  assign new_n52066_ = new_n52056_ & new_n52065_;
  assign new_n52067_ = new_n52047_ & new_n52066_;
  assign new_n52068_ = new_n52028_ & new_n52067_;
  assign new_n52069_ = new_n51989_ & new_n52068_;
  assign new_n52070_ = ys__n46128 & new_n52069_;
  assign new_n52071_ = ys__n45771 & ys__n45976;
  assign new_n52072_ = ~ys__n45771 & ~ys__n45976;
  assign new_n52073_ = ~ys__n46018 & ~new_n52072_;
  assign new_n52074_ = ~new_n52071_ & new_n52073_;
  assign new_n52075_ = ys__n45774 & ys__n45978;
  assign new_n52076_ = ~ys__n45774 & ~ys__n45978;
  assign new_n52077_ = ~ys__n46019 & ~new_n52076_;
  assign new_n52078_ = ~new_n52075_ & new_n52077_;
  assign new_n52079_ = ~new_n52074_ & ~new_n52078_;
  assign new_n52080_ = ys__n45777 & ys__n45980;
  assign new_n52081_ = ~ys__n45777 & ~ys__n45980;
  assign new_n52082_ = ~ys__n46020 & ~new_n52081_;
  assign new_n52083_ = ~new_n52080_ & new_n52082_;
  assign new_n52084_ = ys__n45780 & ys__n45982;
  assign new_n52085_ = ~ys__n45780 & ~ys__n45982;
  assign new_n52086_ = ~ys__n46021 & ~new_n52085_;
  assign new_n52087_ = ~new_n52084_ & new_n52086_;
  assign new_n52088_ = ~new_n52083_ & ~new_n52087_;
  assign new_n52089_ = new_n52079_ & new_n52088_;
  assign new_n52090_ = ys__n45759 & ys__n45968;
  assign new_n52091_ = ~ys__n45759 & ~ys__n45968;
  assign new_n52092_ = ~ys__n46014 & ~new_n52091_;
  assign new_n52093_ = ~new_n52090_ & new_n52092_;
  assign new_n52094_ = ys__n45762 & ys__n45970;
  assign new_n52095_ = ~ys__n45762 & ~ys__n45970;
  assign new_n52096_ = ~ys__n46015 & ~new_n52095_;
  assign new_n52097_ = ~new_n52094_ & new_n52096_;
  assign new_n52098_ = ~new_n52093_ & ~new_n52097_;
  assign new_n52099_ = ys__n45765 & ys__n45972;
  assign new_n52100_ = ~ys__n45765 & ~ys__n45972;
  assign new_n52101_ = ~ys__n46016 & ~new_n52100_;
  assign new_n52102_ = ~new_n52099_ & new_n52101_;
  assign new_n52103_ = ys__n45768 & ys__n45974;
  assign new_n52104_ = ~ys__n45768 & ~ys__n45974;
  assign new_n52105_ = ~ys__n46017 & ~new_n52104_;
  assign new_n52106_ = ~new_n52103_ & new_n52105_;
  assign new_n52107_ = ~new_n52102_ & ~new_n52106_;
  assign new_n52108_ = new_n52098_ & new_n52107_;
  assign new_n52109_ = new_n52089_ & new_n52108_;
  assign new_n52110_ = ys__n45801 & ys__n45996;
  assign new_n52111_ = ~ys__n45801 & ~ys__n45996;
  assign new_n52112_ = ~ys__n46028 & ~new_n52111_;
  assign new_n52113_ = ~new_n52110_ & new_n52112_;
  assign new_n52114_ = ys__n45795 & ys__n45992;
  assign new_n52115_ = ~ys__n45795 & ~ys__n45992;
  assign new_n52116_ = ~ys__n46026 & ~new_n52115_;
  assign new_n52117_ = ~new_n52114_ & new_n52116_;
  assign new_n52118_ = ys__n45798 & ys__n45994;
  assign new_n52119_ = ~ys__n45798 & ~ys__n45994;
  assign new_n52120_ = ~ys__n46027 & ~new_n52119_;
  assign new_n52121_ = ~new_n52118_ & new_n52120_;
  assign new_n52122_ = ~new_n52117_ & ~new_n52121_;
  assign new_n52123_ = ~new_n52113_ & new_n52122_;
  assign new_n52124_ = ys__n45783 & ys__n45984;
  assign new_n52125_ = ~ys__n45783 & ~ys__n45984;
  assign new_n52126_ = ~ys__n46022 & ~new_n52125_;
  assign new_n52127_ = ~new_n52124_ & new_n52126_;
  assign new_n52128_ = ys__n45786 & ys__n45986;
  assign new_n52129_ = ~ys__n45786 & ~ys__n45986;
  assign new_n52130_ = ~ys__n46023 & ~new_n52129_;
  assign new_n52131_ = ~new_n52128_ & new_n52130_;
  assign new_n52132_ = ~new_n52127_ & ~new_n52131_;
  assign new_n52133_ = ys__n45789 & ys__n45988;
  assign new_n52134_ = ~ys__n45789 & ~ys__n45988;
  assign new_n52135_ = ~ys__n46024 & ~new_n52134_;
  assign new_n52136_ = ~new_n52133_ & new_n52135_;
  assign new_n52137_ = ys__n45792 & ys__n45990;
  assign new_n52138_ = ~ys__n45792 & ~ys__n45990;
  assign new_n52139_ = ~ys__n46025 & ~new_n52138_;
  assign new_n52140_ = ~new_n52137_ & new_n52139_;
  assign new_n52141_ = ~new_n52136_ & ~new_n52140_;
  assign new_n52142_ = new_n52132_ & new_n52141_;
  assign new_n52143_ = new_n52123_ & new_n52142_;
  assign new_n52144_ = new_n52109_ & new_n52143_;
  assign new_n52145_ = ys__n45723 & ys__n45944;
  assign new_n52146_ = ~ys__n45723 & ~ys__n45944;
  assign new_n52147_ = ~ys__n46002 & ~new_n52146_;
  assign new_n52148_ = ~new_n52145_ & new_n52147_;
  assign new_n52149_ = ys__n45726 & ys__n45946;
  assign new_n52150_ = ~ys__n45726 & ~ys__n45946;
  assign new_n52151_ = ~ys__n46003 & ~new_n52150_;
  assign new_n52152_ = ~new_n52149_ & new_n52151_;
  assign new_n52153_ = ~new_n52148_ & ~new_n52152_;
  assign new_n52154_ = ys__n45729 & ys__n45948;
  assign new_n52155_ = ~ys__n45729 & ~ys__n45948;
  assign new_n52156_ = ~ys__n46004 & ~new_n52155_;
  assign new_n52157_ = ~new_n52154_ & new_n52156_;
  assign new_n52158_ = ys__n45732 & ys__n45950;
  assign new_n52159_ = ~ys__n45732 & ~ys__n45950;
  assign new_n52160_ = ~ys__n46005 & ~new_n52159_;
  assign new_n52161_ = ~new_n52158_ & new_n52160_;
  assign new_n52162_ = ~new_n52157_ & ~new_n52161_;
  assign new_n52163_ = new_n52153_ & new_n52162_;
  assign new_n52164_ = ys__n45711 & ys__n45936;
  assign new_n52165_ = ~ys__n45711 & ~ys__n45936;
  assign new_n52166_ = ~ys__n45998 & ~new_n52165_;
  assign new_n52167_ = ~new_n52164_ & new_n52166_;
  assign new_n52168_ = ys__n45714 & ys__n45938;
  assign new_n52169_ = ~ys__n45714 & ~ys__n45938;
  assign new_n52170_ = ~ys__n45999 & ~new_n52169_;
  assign new_n52171_ = ~new_n52168_ & new_n52170_;
  assign new_n52172_ = ~new_n52167_ & ~new_n52171_;
  assign new_n52173_ = ys__n45717 & ys__n45940;
  assign new_n52174_ = ~ys__n45717 & ~ys__n45940;
  assign new_n52175_ = ~ys__n46000 & ~new_n52174_;
  assign new_n52176_ = ~new_n52173_ & new_n52175_;
  assign new_n52177_ = ys__n45720 & ys__n45942;
  assign new_n52178_ = ~ys__n45720 & ~ys__n45942;
  assign new_n52179_ = ~ys__n46001 & ~new_n52178_;
  assign new_n52180_ = ~new_n52177_ & new_n52179_;
  assign new_n52181_ = ~new_n52176_ & ~new_n52180_;
  assign new_n52182_ = new_n52172_ & new_n52181_;
  assign new_n52183_ = new_n52163_ & new_n52182_;
  assign new_n52184_ = ys__n45747 & ys__n45960;
  assign new_n52185_ = ~ys__n45747 & ~ys__n45960;
  assign new_n52186_ = ~ys__n46010 & ~new_n52185_;
  assign new_n52187_ = ~new_n52184_ & new_n52186_;
  assign new_n52188_ = ys__n45750 & ys__n45962;
  assign new_n52189_ = ~ys__n45750 & ~ys__n45962;
  assign new_n52190_ = ~ys__n46011 & ~new_n52189_;
  assign new_n52191_ = ~new_n52188_ & new_n52190_;
  assign new_n52192_ = ~new_n52187_ & ~new_n52191_;
  assign new_n52193_ = ys__n45753 & ys__n45964;
  assign new_n52194_ = ~ys__n45753 & ~ys__n45964;
  assign new_n52195_ = ~ys__n46012 & ~new_n52194_;
  assign new_n52196_ = ~new_n52193_ & new_n52195_;
  assign new_n52197_ = ys__n45756 & ys__n45966;
  assign new_n52198_ = ~ys__n45756 & ~ys__n45966;
  assign new_n52199_ = ~ys__n46013 & ~new_n52198_;
  assign new_n52200_ = ~new_n52197_ & new_n52199_;
  assign new_n52201_ = ~new_n52196_ & ~new_n52200_;
  assign new_n52202_ = new_n52192_ & new_n52201_;
  assign new_n52203_ = ys__n45735 & ys__n45952;
  assign new_n52204_ = ~ys__n45735 & ~ys__n45952;
  assign new_n52205_ = ~ys__n46006 & ~new_n52204_;
  assign new_n52206_ = ~new_n52203_ & new_n52205_;
  assign new_n52207_ = ys__n45738 & ys__n45954;
  assign new_n52208_ = ~ys__n45738 & ~ys__n45954;
  assign new_n52209_ = ~ys__n46007 & ~new_n52208_;
  assign new_n52210_ = ~new_n52207_ & new_n52209_;
  assign new_n52211_ = ~new_n52206_ & ~new_n52210_;
  assign new_n52212_ = ys__n45741 & ys__n45956;
  assign new_n52213_ = ~ys__n45741 & ~ys__n45956;
  assign new_n52214_ = ~ys__n46008 & ~new_n52213_;
  assign new_n52215_ = ~new_n52212_ & new_n52214_;
  assign new_n52216_ = ys__n45744 & ys__n45958;
  assign new_n52217_ = ~ys__n45744 & ~ys__n45958;
  assign new_n52218_ = ~ys__n46009 & ~new_n52217_;
  assign new_n52219_ = ~new_n52216_ & new_n52218_;
  assign new_n52220_ = ~new_n52215_ & ~new_n52219_;
  assign new_n52221_ = new_n52211_ & new_n52220_;
  assign new_n52222_ = new_n52202_ & new_n52221_;
  assign new_n52223_ = new_n52183_ & new_n52222_;
  assign new_n52224_ = new_n52144_ & new_n52223_;
  assign new_n52225_ = ys__n46031 & new_n52224_;
  assign new_n52226_ = ~new_n52070_ & ~new_n52225_;
  assign new_n52227_ = ys__n45771 & ys__n45878;
  assign new_n52228_ = ~ys__n45771 & ~ys__n45878;
  assign new_n52229_ = ~ys__n45920 & ~new_n52228_;
  assign new_n52230_ = ~new_n52227_ & new_n52229_;
  assign new_n52231_ = ys__n45774 & ys__n45880;
  assign new_n52232_ = ~ys__n45774 & ~ys__n45880;
  assign new_n52233_ = ~ys__n45921 & ~new_n52232_;
  assign new_n52234_ = ~new_n52231_ & new_n52233_;
  assign new_n52235_ = ~new_n52230_ & ~new_n52234_;
  assign new_n52236_ = ys__n45777 & ys__n45882;
  assign new_n52237_ = ~ys__n45777 & ~ys__n45882;
  assign new_n52238_ = ~ys__n45922 & ~new_n52237_;
  assign new_n52239_ = ~new_n52236_ & new_n52238_;
  assign new_n52240_ = ys__n45780 & ys__n45884;
  assign new_n52241_ = ~ys__n45780 & ~ys__n45884;
  assign new_n52242_ = ~ys__n45923 & ~new_n52241_;
  assign new_n52243_ = ~new_n52240_ & new_n52242_;
  assign new_n52244_ = ~new_n52239_ & ~new_n52243_;
  assign new_n52245_ = new_n52235_ & new_n52244_;
  assign new_n52246_ = ys__n45759 & ys__n45870;
  assign new_n52247_ = ~ys__n45759 & ~ys__n45870;
  assign new_n52248_ = ~ys__n45916 & ~new_n52247_;
  assign new_n52249_ = ~new_n52246_ & new_n52248_;
  assign new_n52250_ = ys__n45762 & ys__n45872;
  assign new_n52251_ = ~ys__n45762 & ~ys__n45872;
  assign new_n52252_ = ~ys__n45917 & ~new_n52251_;
  assign new_n52253_ = ~new_n52250_ & new_n52252_;
  assign new_n52254_ = ~new_n52249_ & ~new_n52253_;
  assign new_n52255_ = ys__n45765 & ys__n45874;
  assign new_n52256_ = ~ys__n45765 & ~ys__n45874;
  assign new_n52257_ = ~ys__n45918 & ~new_n52256_;
  assign new_n52258_ = ~new_n52255_ & new_n52257_;
  assign new_n52259_ = ys__n45768 & ys__n45876;
  assign new_n52260_ = ~ys__n45768 & ~ys__n45876;
  assign new_n52261_ = ~ys__n45919 & ~new_n52260_;
  assign new_n52262_ = ~new_n52259_ & new_n52261_;
  assign new_n52263_ = ~new_n52258_ & ~new_n52262_;
  assign new_n52264_ = new_n52254_ & new_n52263_;
  assign new_n52265_ = new_n52245_ & new_n52264_;
  assign new_n52266_ = ys__n45801 & ys__n45898;
  assign new_n52267_ = ~ys__n45801 & ~ys__n45898;
  assign new_n52268_ = ~ys__n45930 & ~new_n52267_;
  assign new_n52269_ = ~new_n52266_ & new_n52268_;
  assign new_n52270_ = ys__n45795 & ys__n45894;
  assign new_n52271_ = ~ys__n45795 & ~ys__n45894;
  assign new_n52272_ = ~ys__n45928 & ~new_n52271_;
  assign new_n52273_ = ~new_n52270_ & new_n52272_;
  assign new_n52274_ = ys__n45798 & ys__n45896;
  assign new_n52275_ = ~ys__n45798 & ~ys__n45896;
  assign new_n52276_ = ~ys__n45929 & ~new_n52275_;
  assign new_n52277_ = ~new_n52274_ & new_n52276_;
  assign new_n52278_ = ~new_n52273_ & ~new_n52277_;
  assign new_n52279_ = ~new_n52269_ & new_n52278_;
  assign new_n52280_ = ys__n45783 & ys__n45886;
  assign new_n52281_ = ~ys__n45783 & ~ys__n45886;
  assign new_n52282_ = ~ys__n45924 & ~new_n52281_;
  assign new_n52283_ = ~new_n52280_ & new_n52282_;
  assign new_n52284_ = ys__n45786 & ys__n45888;
  assign new_n52285_ = ~ys__n45786 & ~ys__n45888;
  assign new_n52286_ = ~ys__n45925 & ~new_n52285_;
  assign new_n52287_ = ~new_n52284_ & new_n52286_;
  assign new_n52288_ = ~new_n52283_ & ~new_n52287_;
  assign new_n52289_ = ys__n45789 & ys__n45890;
  assign new_n52290_ = ~ys__n45789 & ~ys__n45890;
  assign new_n52291_ = ~ys__n45926 & ~new_n52290_;
  assign new_n52292_ = ~new_n52289_ & new_n52291_;
  assign new_n52293_ = ys__n45792 & ys__n45892;
  assign new_n52294_ = ~ys__n45792 & ~ys__n45892;
  assign new_n52295_ = ~ys__n45927 & ~new_n52294_;
  assign new_n52296_ = ~new_n52293_ & new_n52295_;
  assign new_n52297_ = ~new_n52292_ & ~new_n52296_;
  assign new_n52298_ = new_n52288_ & new_n52297_;
  assign new_n52299_ = new_n52279_ & new_n52298_;
  assign new_n52300_ = new_n52265_ & new_n52299_;
  assign new_n52301_ = ys__n45723 & ys__n45846;
  assign new_n52302_ = ~ys__n45723 & ~ys__n45846;
  assign new_n52303_ = ~ys__n45904 & ~new_n52302_;
  assign new_n52304_ = ~new_n52301_ & new_n52303_;
  assign new_n52305_ = ys__n45726 & ys__n45848;
  assign new_n52306_ = ~ys__n45726 & ~ys__n45848;
  assign new_n52307_ = ~ys__n45905 & ~new_n52306_;
  assign new_n52308_ = ~new_n52305_ & new_n52307_;
  assign new_n52309_ = ~new_n52304_ & ~new_n52308_;
  assign new_n52310_ = ys__n45729 & ys__n45850;
  assign new_n52311_ = ~ys__n45729 & ~ys__n45850;
  assign new_n52312_ = ~ys__n45906 & ~new_n52311_;
  assign new_n52313_ = ~new_n52310_ & new_n52312_;
  assign new_n52314_ = ys__n45732 & ys__n45852;
  assign new_n52315_ = ~ys__n45732 & ~ys__n45852;
  assign new_n52316_ = ~ys__n45907 & ~new_n52315_;
  assign new_n52317_ = ~new_n52314_ & new_n52316_;
  assign new_n52318_ = ~new_n52313_ & ~new_n52317_;
  assign new_n52319_ = new_n52309_ & new_n52318_;
  assign new_n52320_ = ys__n45711 & ys__n45838;
  assign new_n52321_ = ~ys__n45711 & ~ys__n45838;
  assign new_n52322_ = ~ys__n45900 & ~new_n52321_;
  assign new_n52323_ = ~new_n52320_ & new_n52322_;
  assign new_n52324_ = ys__n45714 & ys__n45840;
  assign new_n52325_ = ~ys__n45714 & ~ys__n45840;
  assign new_n52326_ = ~ys__n45901 & ~new_n52325_;
  assign new_n52327_ = ~new_n52324_ & new_n52326_;
  assign new_n52328_ = ~new_n52323_ & ~new_n52327_;
  assign new_n52329_ = ys__n45717 & ys__n45842;
  assign new_n52330_ = ~ys__n45717 & ~ys__n45842;
  assign new_n52331_ = ~ys__n45902 & ~new_n52330_;
  assign new_n52332_ = ~new_n52329_ & new_n52331_;
  assign new_n52333_ = ys__n45720 & ys__n45844;
  assign new_n52334_ = ~ys__n45720 & ~ys__n45844;
  assign new_n52335_ = ~ys__n45903 & ~new_n52334_;
  assign new_n52336_ = ~new_n52333_ & new_n52335_;
  assign new_n52337_ = ~new_n52332_ & ~new_n52336_;
  assign new_n52338_ = new_n52328_ & new_n52337_;
  assign new_n52339_ = new_n52319_ & new_n52338_;
  assign new_n52340_ = ys__n45747 & ys__n45862;
  assign new_n52341_ = ~ys__n45747 & ~ys__n45862;
  assign new_n52342_ = ~ys__n45912 & ~new_n52341_;
  assign new_n52343_ = ~new_n52340_ & new_n52342_;
  assign new_n52344_ = ys__n45750 & ys__n45864;
  assign new_n52345_ = ~ys__n45750 & ~ys__n45864;
  assign new_n52346_ = ~ys__n45913 & ~new_n52345_;
  assign new_n52347_ = ~new_n52344_ & new_n52346_;
  assign new_n52348_ = ~new_n52343_ & ~new_n52347_;
  assign new_n52349_ = ys__n45753 & ys__n45866;
  assign new_n52350_ = ~ys__n45753 & ~ys__n45866;
  assign new_n52351_ = ~ys__n45914 & ~new_n52350_;
  assign new_n52352_ = ~new_n52349_ & new_n52351_;
  assign new_n52353_ = ys__n45756 & ys__n45868;
  assign new_n52354_ = ~ys__n45756 & ~ys__n45868;
  assign new_n52355_ = ~ys__n45915 & ~new_n52354_;
  assign new_n52356_ = ~new_n52353_ & new_n52355_;
  assign new_n52357_ = ~new_n52352_ & ~new_n52356_;
  assign new_n52358_ = new_n52348_ & new_n52357_;
  assign new_n52359_ = ys__n45735 & ys__n45854;
  assign new_n52360_ = ~ys__n45735 & ~ys__n45854;
  assign new_n52361_ = ~ys__n45908 & ~new_n52360_;
  assign new_n52362_ = ~new_n52359_ & new_n52361_;
  assign new_n52363_ = ys__n45738 & ys__n45856;
  assign new_n52364_ = ~ys__n45738 & ~ys__n45856;
  assign new_n52365_ = ~ys__n45909 & ~new_n52364_;
  assign new_n52366_ = ~new_n52363_ & new_n52365_;
  assign new_n52367_ = ~new_n52362_ & ~new_n52366_;
  assign new_n52368_ = ys__n45741 & ys__n45858;
  assign new_n52369_ = ~ys__n45741 & ~ys__n45858;
  assign new_n52370_ = ~ys__n45910 & ~new_n52369_;
  assign new_n52371_ = ~new_n52368_ & new_n52370_;
  assign new_n52372_ = ys__n45744 & ys__n45860;
  assign new_n52373_ = ~ys__n45744 & ~ys__n45860;
  assign new_n52374_ = ~ys__n45911 & ~new_n52373_;
  assign new_n52375_ = ~new_n52372_ & new_n52374_;
  assign new_n52376_ = ~new_n52371_ & ~new_n52375_;
  assign new_n52377_ = new_n52367_ & new_n52376_;
  assign new_n52378_ = new_n52358_ & new_n52377_;
  assign new_n52379_ = new_n52339_ & new_n52378_;
  assign new_n52380_ = new_n52300_ & new_n52379_;
  assign new_n52381_ = ys__n45933 & new_n52380_;
  assign new_n52382_ = ys__n45771 & ys__n45772;
  assign new_n52383_ = ~ys__n45771 & ~ys__n45772;
  assign new_n52384_ = ~ys__n45824 & ~new_n52383_;
  assign new_n52385_ = ~new_n52382_ & new_n52384_;
  assign new_n52386_ = ys__n45774 & ys__n45775;
  assign new_n52387_ = ~ys__n45774 & ~ys__n45775;
  assign new_n52388_ = ~ys__n45825 & ~new_n52387_;
  assign new_n52389_ = ~new_n52386_ & new_n52388_;
  assign new_n52390_ = ~new_n52385_ & ~new_n52389_;
  assign new_n52391_ = ys__n45777 & ys__n45778;
  assign new_n52392_ = ~ys__n45777 & ~ys__n45778;
  assign new_n52393_ = ~ys__n45826 & ~new_n52392_;
  assign new_n52394_ = ~new_n52391_ & new_n52393_;
  assign new_n52395_ = ys__n45780 & ys__n45781;
  assign new_n52396_ = ~ys__n45780 & ~ys__n45781;
  assign new_n52397_ = ~ys__n45827 & ~new_n52396_;
  assign new_n52398_ = ~new_n52395_ & new_n52397_;
  assign new_n52399_ = ~new_n52394_ & ~new_n52398_;
  assign new_n52400_ = new_n52390_ & new_n52399_;
  assign new_n52401_ = ys__n45759 & ys__n45760;
  assign new_n52402_ = ~ys__n45759 & ~ys__n45760;
  assign new_n52403_ = ~ys__n45820 & ~new_n52402_;
  assign new_n52404_ = ~new_n52401_ & new_n52403_;
  assign new_n52405_ = ys__n45762 & ys__n45763;
  assign new_n52406_ = ~ys__n45762 & ~ys__n45763;
  assign new_n52407_ = ~ys__n45821 & ~new_n52406_;
  assign new_n52408_ = ~new_n52405_ & new_n52407_;
  assign new_n52409_ = ~new_n52404_ & ~new_n52408_;
  assign new_n52410_ = ys__n45765 & ys__n45766;
  assign new_n52411_ = ~ys__n45765 & ~ys__n45766;
  assign new_n52412_ = ~ys__n45822 & ~new_n52411_;
  assign new_n52413_ = ~new_n52410_ & new_n52412_;
  assign new_n52414_ = ys__n45768 & ys__n45769;
  assign new_n52415_ = ~ys__n45768 & ~ys__n45769;
  assign new_n52416_ = ~ys__n45823 & ~new_n52415_;
  assign new_n52417_ = ~new_n52414_ & new_n52416_;
  assign new_n52418_ = ~new_n52413_ & ~new_n52417_;
  assign new_n52419_ = new_n52409_ & new_n52418_;
  assign new_n52420_ = new_n52400_ & new_n52419_;
  assign new_n52421_ = ys__n45801 & ys__n45802;
  assign new_n52422_ = ~ys__n45801 & ~ys__n45802;
  assign new_n52423_ = ~ys__n45834 & ~new_n52422_;
  assign new_n52424_ = ~new_n52421_ & new_n52423_;
  assign new_n52425_ = ys__n45795 & ys__n45796;
  assign new_n52426_ = ~ys__n45795 & ~ys__n45796;
  assign new_n52427_ = ~ys__n45832 & ~new_n52426_;
  assign new_n52428_ = ~new_n52425_ & new_n52427_;
  assign new_n52429_ = ys__n45798 & ys__n45799;
  assign new_n52430_ = ~ys__n45798 & ~ys__n45799;
  assign new_n52431_ = ~ys__n45833 & ~new_n52430_;
  assign new_n52432_ = ~new_n52429_ & new_n52431_;
  assign new_n52433_ = ~new_n52428_ & ~new_n52432_;
  assign new_n52434_ = ~new_n52424_ & new_n52433_;
  assign new_n52435_ = ys__n45783 & ys__n45784;
  assign new_n52436_ = ~ys__n45783 & ~ys__n45784;
  assign new_n52437_ = ~ys__n45828 & ~new_n52436_;
  assign new_n52438_ = ~new_n52435_ & new_n52437_;
  assign new_n52439_ = ys__n45786 & ys__n45787;
  assign new_n52440_ = ~ys__n45786 & ~ys__n45787;
  assign new_n52441_ = ~ys__n45829 & ~new_n52440_;
  assign new_n52442_ = ~new_n52439_ & new_n52441_;
  assign new_n52443_ = ~new_n52438_ & ~new_n52442_;
  assign new_n52444_ = ys__n45789 & ys__n45790;
  assign new_n52445_ = ~ys__n45789 & ~ys__n45790;
  assign new_n52446_ = ~ys__n45830 & ~new_n52445_;
  assign new_n52447_ = ~new_n52444_ & new_n52446_;
  assign new_n52448_ = ys__n45792 & ys__n45793;
  assign new_n52449_ = ~ys__n45792 & ~ys__n45793;
  assign new_n52450_ = ~ys__n45831 & ~new_n52449_;
  assign new_n52451_ = ~new_n52448_ & new_n52450_;
  assign new_n52452_ = ~new_n52447_ & ~new_n52451_;
  assign new_n52453_ = new_n52443_ & new_n52452_;
  assign new_n52454_ = new_n52434_ & new_n52453_;
  assign new_n52455_ = new_n52420_ & new_n52454_;
  assign new_n52456_ = ys__n45723 & ys__n45724;
  assign new_n52457_ = ~ys__n45723 & ~ys__n45724;
  assign new_n52458_ = ~ys__n45808 & ~new_n52457_;
  assign new_n52459_ = ~new_n52456_ & new_n52458_;
  assign new_n52460_ = ys__n45726 & ys__n45727;
  assign new_n52461_ = ~ys__n45726 & ~ys__n45727;
  assign new_n52462_ = ~ys__n45809 & ~new_n52461_;
  assign new_n52463_ = ~new_n52460_ & new_n52462_;
  assign new_n52464_ = ~new_n52459_ & ~new_n52463_;
  assign new_n52465_ = ys__n45729 & ys__n45730;
  assign new_n52466_ = ~ys__n45729 & ~ys__n45730;
  assign new_n52467_ = ~ys__n45810 & ~new_n52466_;
  assign new_n52468_ = ~new_n52465_ & new_n52467_;
  assign new_n52469_ = ys__n45732 & ys__n45733;
  assign new_n52470_ = ~ys__n45732 & ~ys__n45733;
  assign new_n52471_ = ~ys__n45811 & ~new_n52470_;
  assign new_n52472_ = ~new_n52469_ & new_n52471_;
  assign new_n52473_ = ~new_n52468_ & ~new_n52472_;
  assign new_n52474_ = new_n52464_ & new_n52473_;
  assign new_n52475_ = ys__n45711 & ys__n45712;
  assign new_n52476_ = ~ys__n45711 & ~ys__n45712;
  assign new_n52477_ = ~ys__n45804 & ~new_n52476_;
  assign new_n52478_ = ~new_n52475_ & new_n52477_;
  assign new_n52479_ = ys__n45714 & ys__n45715;
  assign new_n52480_ = ~ys__n45714 & ~ys__n45715;
  assign new_n52481_ = ~ys__n45805 & ~new_n52480_;
  assign new_n52482_ = ~new_n52479_ & new_n52481_;
  assign new_n52483_ = ~new_n52478_ & ~new_n52482_;
  assign new_n52484_ = ys__n45717 & ys__n45718;
  assign new_n52485_ = ~ys__n45717 & ~ys__n45718;
  assign new_n52486_ = ~ys__n45806 & ~new_n52485_;
  assign new_n52487_ = ~new_n52484_ & new_n52486_;
  assign new_n52488_ = ys__n45720 & ys__n45721;
  assign new_n52489_ = ~ys__n45720 & ~ys__n45721;
  assign new_n52490_ = ~ys__n45807 & ~new_n52489_;
  assign new_n52491_ = ~new_n52488_ & new_n52490_;
  assign new_n52492_ = ~new_n52487_ & ~new_n52491_;
  assign new_n52493_ = new_n52483_ & new_n52492_;
  assign new_n52494_ = new_n52474_ & new_n52493_;
  assign new_n52495_ = ys__n45747 & ys__n45748;
  assign new_n52496_ = ~ys__n45747 & ~ys__n45748;
  assign new_n52497_ = ~ys__n45816 & ~new_n52496_;
  assign new_n52498_ = ~new_n52495_ & new_n52497_;
  assign new_n52499_ = ys__n45750 & ys__n45751;
  assign new_n52500_ = ~ys__n45750 & ~ys__n45751;
  assign new_n52501_ = ~ys__n45817 & ~new_n52500_;
  assign new_n52502_ = ~new_n52499_ & new_n52501_;
  assign new_n52503_ = ~new_n52498_ & ~new_n52502_;
  assign new_n52504_ = ys__n45753 & ys__n45754;
  assign new_n52505_ = ~ys__n45753 & ~ys__n45754;
  assign new_n52506_ = ~ys__n45818 & ~new_n52505_;
  assign new_n52507_ = ~new_n52504_ & new_n52506_;
  assign new_n52508_ = ys__n45756 & ys__n45757;
  assign new_n52509_ = ~ys__n45756 & ~ys__n45757;
  assign new_n52510_ = ~ys__n45819 & ~new_n52509_;
  assign new_n52511_ = ~new_n52508_ & new_n52510_;
  assign new_n52512_ = ~new_n52507_ & ~new_n52511_;
  assign new_n52513_ = new_n52503_ & new_n52512_;
  assign new_n52514_ = ys__n45735 & ys__n45736;
  assign new_n52515_ = ~ys__n45735 & ~ys__n45736;
  assign new_n52516_ = ~ys__n45812 & ~new_n52515_;
  assign new_n52517_ = ~new_n52514_ & new_n52516_;
  assign new_n52518_ = ys__n45738 & ys__n45739;
  assign new_n52519_ = ~ys__n45738 & ~ys__n45739;
  assign new_n52520_ = ~ys__n45813 & ~new_n52519_;
  assign new_n52521_ = ~new_n52518_ & new_n52520_;
  assign new_n52522_ = ~new_n52517_ & ~new_n52521_;
  assign new_n52523_ = ys__n45741 & ys__n45742;
  assign new_n52524_ = ~ys__n45741 & ~ys__n45742;
  assign new_n52525_ = ~ys__n45814 & ~new_n52524_;
  assign new_n52526_ = ~new_n52523_ & new_n52525_;
  assign new_n52527_ = ys__n45744 & ys__n45745;
  assign new_n52528_ = ~ys__n45744 & ~ys__n45745;
  assign new_n52529_ = ~ys__n45815 & ~new_n52528_;
  assign new_n52530_ = ~new_n52527_ & new_n52529_;
  assign new_n52531_ = ~new_n52526_ & ~new_n52530_;
  assign new_n52532_ = new_n52522_ & new_n52531_;
  assign new_n52533_ = new_n52513_ & new_n52532_;
  assign new_n52534_ = new_n52494_ & new_n52533_;
  assign new_n52535_ = new_n52455_ & new_n52534_;
  assign new_n52536_ = ys__n45836 & new_n52535_;
  assign new_n52537_ = ~new_n52381_ & ~new_n52536_;
  assign new_n52538_ = new_n52226_ & new_n52537_;
  assign new_n52539_ = ~ys__n30225 & ys__n38910;
  assign new_n52540_ = ~ys__n1020 & new_n52539_;
  assign new_n52541_ = ~ys__n38908 & ~new_n52540_;
  assign new_n52542_ = ~new_n52538_ & ~new_n52541_;
  assign new_n52543_ = ~ys__n38288 & ~new_n52542_;
  assign ys__n38209 = ~ys__n4566 & ~new_n52543_;
  assign new_n52545_ = ys__n46127 & new_n52069_;
  assign new_n52546_ = ys__n46029 & new_n52224_;
  assign new_n52547_ = ~new_n52545_ & ~new_n52546_;
  assign new_n52548_ = ys__n45931 & new_n52380_;
  assign new_n52549_ = ys__n45835 & new_n52535_;
  assign new_n52550_ = ~new_n52548_ & ~new_n52549_;
  assign new_n52551_ = new_n52547_ & new_n52550_;
  assign new_n52552_ = ~new_n52541_ & ~new_n52551_;
  assign new_n52553_ = ~ys__n38290 & ~new_n52552_;
  assign ys__n38211 = ~ys__n4566 & ~new_n52553_;
  assign ys__n38213 = ys__n38212 & ~ys__n4566;
  assign new_n52556_ = ~ys__n18101 & ~ys__n18106;
  assign new_n52557_ = ~ys__n33375 & ys__n38315;
  assign new_n52558_ = new_n52556_ & new_n52557_;
  assign new_n52559_ = ys__n38311 & new_n52558_;
  assign new_n52560_ = ~new_n11954_ & new_n52559_;
  assign new_n52561_ = new_n17588_ & new_n52558_;
  assign new_n52562_ = ys__n23272 & ~ys__n23335;
  assign new_n52563_ = ys__n23332 & new_n52558_;
  assign new_n52564_ = ~new_n52562_ & ~new_n52563_;
  assign new_n52565_ = new_n12314_ & ~new_n52564_;
  assign new_n52566_ = ~new_n52561_ & ~new_n52565_;
  assign new_n52567_ = new_n11954_ & ~new_n52566_;
  assign new_n52568_ = ~new_n52560_ & ~new_n52567_;
  assign ys__n38214 = ~ys__n4566 & ~new_n52568_;
  assign ys__n38216 = ys__n38215 & ~ys__n4566;
  assign ys__n38218 = ys__n38217 & ~ys__n4566;
  assign ys__n38222 = ~ys__n33340 & ys__n478;
  assign new_n52573_ = ys__n22818 & ~ys__n33342;
  assign ys__n38224 = ys__n935 | new_n52573_;
  assign ys__n38246 = ~new_n15018_ & new_n15036_;
  assign ys__n38247 = ~new_n15018_ & new_n15032_;
  assign ys__n38248 = ~new_n15018_ & new_n15030_;
  assign new_n52578_ = new_n15018_ & new_n15048_;
  assign ys__n38250 = new_n15037_ | new_n52578_;
  assign new_n52580_ = new_n15018_ & new_n15047_;
  assign ys__n38252 = new_n15038_ | new_n52580_;
  assign new_n52582_ = ~ys__n33364 & ys__n38237;
  assign new_n52583_ = new_n15018_ & new_n52582_;
  assign new_n52584_ = ~ys__n33350 & ~new_n52583_;
  assign ys__n38263 = ~new_n15085_ & ~new_n52584_;
  assign new_n52586_ = ~ys__n33364 & ys__n38236;
  assign new_n52587_ = new_n15018_ & new_n52586_;
  assign new_n52588_ = ~ys__n33352 & ~new_n52587_;
  assign ys__n38266 = ~new_n15085_ & ~new_n52588_;
  assign ys__n38281 = ys__n738 & ~new_n51911_;
  assign new_n52591_ = ~ys__n38286 & ~new_n51910_;
  assign ys__n38285 = ys__n738 & ~new_n52591_;
  assign ys__n38287 = ys__n738 & ~new_n52543_;
  assign ys__n38289 = ys__n738 & ~new_n52553_;
  assign ys__n38292 = ys__n34959 | ys__n38291;
  assign new_n52596_ = ys__n422 & ys__n432;
  assign new_n52597_ = new_n12716_ & new_n52596_;
  assign new_n52598_ = new_n12821_ & new_n52597_;
  assign new_n52599_ = ~ys__n436 & ~ys__n34959;
  assign new_n52600_ = ys__n38291 & new_n52599_;
  assign new_n52601_ = new_n12741_ & new_n52600_;
  assign ys__n38294 = new_n52598_ & new_n52601_;
  assign new_n52603_ = ~ys__n935 & ~ys__n34959;
  assign ys__n38296 = ~ys__n33366 & ~new_n52603_;
  assign new_n52605_ = new_n17091_ & ~new_n17097_;
  assign new_n52606_ = ~new_n17099_ & ~new_n52605_;
  assign new_n52607_ = ~ys__n28243 & ~new_n52606_;
  assign new_n52608_ = ys__n28243 & ~new_n52607_;
  assign new_n52609_ = ys__n23480 & new_n52607_;
  assign ys__n38303 = new_n52608_ | new_n52609_;
  assign new_n52611_ = ys__n23339 & ~new_n12457_;
  assign new_n52612_ = ~ys__n28243 & new_n12457_;
  assign new_n52613_ = ~new_n52611_ & ~new_n52612_;
  assign new_n52614_ = ~new_n12309_ & ~new_n52613_;
  assign new_n52615_ = ~new_n35685_ & ~new_n52614_;
  assign new_n52616_ = ~new_n12314_ & ~new_n52615_;
  assign new_n52617_ = ys__n23335 & new_n12314_;
  assign new_n52618_ = ~new_n52616_ & ~new_n52617_;
  assign new_n52619_ = new_n11954_ & ~new_n52618_;
  assign new_n52620_ = ys__n23339 & ~new_n11954_;
  assign new_n52621_ = ~new_n52619_ & ~new_n52620_;
  assign ys__n38325 = ~ys__n4566 & ~new_n52621_;
  assign new_n52623_ = new_n12326_ & ~new_n12328_;
  assign new_n52624_ = ~ys__n516 & ~ys__n520;
  assign new_n52625_ = ~ys__n2024 & ~ys__n4478;
  assign new_n52626_ = ~ys__n4480 & new_n52625_;
  assign new_n52627_ = new_n52624_ & new_n52626_;
  assign new_n52628_ = new_n12346_ & new_n52627_;
  assign new_n52629_ = ~new_n52623_ & new_n52628_;
  assign new_n52630_ = new_n12464_ & ~new_n52629_;
  assign new_n52631_ = ~new_n12327_ & new_n12336_;
  assign new_n52632_ = new_n52623_ & new_n52631_;
  assign new_n52633_ = ~ys__n28243 & ~new_n52632_;
  assign new_n52634_ = ~new_n52630_ & new_n52633_;
  assign new_n52635_ = new_n12341_ & ~new_n17097_;
  assign new_n52636_ = new_n12391_ & new_n17094_;
  assign new_n52637_ = new_n17092_ & new_n52636_;
  assign new_n52638_ = ~new_n17096_ & ~new_n52637_;
  assign new_n52639_ = new_n17097_ & ~new_n52638_;
  assign new_n52640_ = new_n12341_ & ~new_n52639_;
  assign new_n52641_ = ~ys__n28243 & ~new_n52640_;
  assign new_n52642_ = ~new_n52635_ & new_n52641_;
  assign new_n52643_ = ~ys__n23730 & new_n17105_;
  assign new_n52644_ = ~ys__n23730 & ~new_n52643_;
  assign new_n52645_ = ys__n28243 & ~new_n52644_;
  assign new_n52646_ = ~new_n52642_ & ~new_n52645_;
  assign ys__n38326 = new_n52634_ | ~new_n52646_;
  assign ys__n38327 = ys__n33359 & ~ys__n4566;
  assign ys__n38328 = ys__n256 & ~ys__n4566;
  assign new_n52650_ = new_n11764_ & new_n11782_;
  assign new_n52651_ = new_n11792_ & new_n12318_;
  assign new_n52652_ = new_n52650_ & new_n52651_;
  assign ys__n38330 = ~ys__n4566 & new_n52652_;
  assign ys__n38331 = ys__n262 & ~ys__n4566;
  assign ys__n38332 = ys__n18105 & ~ys__n4566;
  assign new_n52656_ = new_n12318_ & new_n12337_;
  assign ys__n38334 = ~ys__n4566 & new_n52656_;
  assign new_n52658_ = new_n12318_ & new_n12384_;
  assign new_n52659_ = new_n12394_ & new_n52658_;
  assign ys__n38336 = ~ys__n4566 & new_n52659_;
  assign new_n52661_ = ys__n550 & ~ys__n23730;
  assign new_n52662_ = ys__n28243 & new_n52661_;
  assign new_n52663_ = new_n12337_ & new_n52662_;
  assign ys__n38337 = ~ys__n4566 & new_n52663_;
  assign new_n52665_ = ~ys__n28243 & new_n12334_;
  assign ys__n38339 = ~ys__n4566 & new_n52665_;
  assign new_n52667_ = ~new_n12356_ & ~new_n12363_;
  assign new_n52668_ = ~ys__n28243 & new_n12327_;
  assign new_n52669_ = ~new_n52667_ & new_n52668_;
  assign ys__n38340 = ~ys__n4566 & new_n52669_;
  assign new_n52671_ = ~new_n12351_ & ~new_n12362_;
  assign new_n52672_ = new_n52668_ & ~new_n52671_;
  assign ys__n38341 = ~ys__n4566 & new_n52672_;
  assign new_n52674_ = ~ys__n28243 & new_n12332_;
  assign ys__n38342 = ~ys__n4566 & new_n52674_;
  assign new_n52676_ = ~ys__n28243 & new_n11780_;
  assign new_n52677_ = ~ys__n23730 & new_n11769_;
  assign new_n52678_ = new_n11767_ & new_n52677_;
  assign new_n52679_ = ~ys__n23730 & new_n11780_;
  assign new_n52680_ = ~new_n52678_ & ~new_n52679_;
  assign new_n52681_ = ~new_n11767_ & ~new_n11780_;
  assign new_n52682_ = ys__n28243 & ~new_n52681_;
  assign new_n52683_ = ~new_n52680_ & new_n52682_;
  assign new_n52684_ = ~new_n52676_ & ~new_n52683_;
  assign ys__n38343 = ~ys__n4566 & ~new_n52684_;
  assign new_n52686_ = ~ys__n28243 & new_n11777_;
  assign new_n52687_ = ~ys__n23730 & new_n11771_;
  assign new_n52688_ = new_n11767_ & new_n52687_;
  assign new_n52689_ = ~ys__n23730 & new_n11777_;
  assign new_n52690_ = ~new_n52688_ & ~new_n52689_;
  assign new_n52691_ = ~new_n11767_ & ~new_n11777_;
  assign new_n52692_ = ys__n28243 & ~new_n52691_;
  assign new_n52693_ = ~new_n52690_ & new_n52692_;
  assign new_n52694_ = ~new_n52686_ & ~new_n52693_;
  assign ys__n38344 = ~ys__n4566 & ~new_n52694_;
  assign new_n52696_ = ~ys__n28243 & new_n52639_;
  assign new_n52697_ = ys__n28243 & new_n12384_;
  assign new_n52698_ = new_n12395_ & new_n52697_;
  assign new_n52699_ = ~new_n52696_ & ~new_n52698_;
  assign ys__n38345 = ~ys__n4566 & ~new_n52699_;
  assign ys__n38347 = ys__n38346 & ~ys__n4566;
  assign new_n52702_ = ys__n22648 & ys__n28432;
  assign new_n52703_ = ys__n22650 & ys__n28434;
  assign new_n52704_ = ~new_n52702_ & ~new_n52703_;
  assign new_n52705_ = ys__n22652 & ys__n28436;
  assign new_n52706_ = ys__n22654 & ys__n28438;
  assign new_n52707_ = ~new_n52705_ & ~new_n52706_;
  assign new_n52708_ = new_n52704_ & new_n52707_;
  assign new_n52709_ = ys__n22640 & ys__n28424;
  assign new_n52710_ = ys__n22642 & ys__n28426;
  assign new_n52711_ = ~new_n52709_ & ~new_n52710_;
  assign new_n52712_ = ys__n22644 & ys__n28428;
  assign new_n52713_ = ys__n22646 & ys__n28430;
  assign new_n52714_ = ~new_n52712_ & ~new_n52713_;
  assign new_n52715_ = new_n52711_ & new_n52714_;
  assign new_n52716_ = new_n52708_ & new_n52715_;
  assign new_n52717_ = ~ys__n33370 & ~ys__n33389;
  assign new_n52718_ = ys__n38427 & new_n52717_;
  assign new_n52719_ = ~new_n52716_ & new_n52718_;
  assign new_n52720_ = ~ys__n4566 & new_n52719_;
  assign ys__n38349 = ~ys__n18120 & new_n52720_;
  assign new_n52722_ = ~ys__n38420 & new_n45794_;
  assign new_n52723_ = ~new_n45790_ & new_n52722_;
  assign new_n52724_ = new_n45788_ & new_n52723_;
  assign ys__n38351 = ~ys__n4566 & ~new_n52724_;
  assign new_n52726_ = ~ys__n28243 & new_n12298_;
  assign ys__n38352 = ~ys__n4566 & new_n52726_;
  assign new_n52728_ = ys__n748 & ys__n750;
  assign new_n52729_ = new_n11796_ & new_n52728_;
  assign new_n52730_ = ys__n742 & ~ys__n744;
  assign new_n52731_ = new_n11778_ & new_n52730_;
  assign new_n52732_ = new_n52728_ & new_n52731_;
  assign new_n52733_ = ~new_n12328_ & ~new_n52732_;
  assign new_n52734_ = ~new_n52729_ & new_n52733_;
  assign ys__n38353 = new_n38358_ & ~new_n52734_;
  assign new_n52736_ = new_n11784_ & new_n52728_;
  assign new_n52737_ = new_n11782_ & new_n52730_;
  assign new_n52738_ = new_n52728_ & new_n52737_;
  assign new_n52739_ = ~new_n12325_ & ~new_n52738_;
  assign new_n52740_ = ~new_n52736_ & new_n52739_;
  assign ys__n38354 = new_n38358_ & ~new_n52740_;
  assign new_n52742_ = new_n11802_ & new_n52728_;
  assign new_n52743_ = new_n11801_ & new_n52730_;
  assign new_n52744_ = new_n52728_ & new_n52743_;
  assign new_n52745_ = ~new_n12324_ & ~new_n52744_;
  assign new_n52746_ = ~new_n52742_ & new_n52745_;
  assign ys__n38355 = new_n38358_ & ~new_n52746_;
  assign new_n52748_ = new_n11763_ & new_n52730_;
  assign new_n52749_ = new_n11766_ & new_n52748_;
  assign new_n52750_ = ~ys__n530 & ys__n752;
  assign new_n52751_ = new_n12393_ & new_n52750_;
  assign new_n52752_ = ys__n526 & ~ys__n528;
  assign new_n52753_ = new_n12392_ & new_n52750_;
  assign new_n52754_ = new_n52752_ & new_n52753_;
  assign new_n52755_ = ~new_n52751_ & ~new_n52754_;
  assign new_n52756_ = new_n17097_ & ~new_n52755_;
  assign new_n52757_ = ~new_n52749_ & ~new_n52756_;
  assign new_n52758_ = ~new_n17097_ & ~new_n52749_;
  assign new_n52759_ = ~ys__n28243 & ~new_n52758_;
  assign new_n52760_ = ~ys__n4566 & new_n52759_;
  assign ys__n38356 = ~new_n52757_ & new_n52760_;
  assign new_n52762_ = ~ys__n28243 & new_n12299_;
  assign new_n52763_ = new_n17092_ & new_n17093_;
  assign new_n52764_ = new_n52762_ & new_n52763_;
  assign new_n52765_ = new_n17097_ & new_n52764_;
  assign new_n52766_ = ~ys__n522 & ys__n524;
  assign new_n52767_ = new_n17093_ & new_n52766_;
  assign new_n52768_ = ~ys__n530 & ys__n28243;
  assign new_n52769_ = new_n52767_ & new_n52768_;
  assign new_n52770_ = new_n12384_ & new_n52769_;
  assign new_n52771_ = ~new_n52765_ & ~new_n52770_;
  assign ys__n38357 = ~ys__n4566 & ~new_n52771_;
  assign new_n52773_ = new_n12391_ & new_n17092_;
  assign new_n52774_ = new_n52762_ & new_n52773_;
  assign new_n52775_ = new_n17097_ & new_n52774_;
  assign ys__n38359 = ~ys__n4566 & new_n52775_;
  assign new_n52777_ = new_n12392_ & new_n17093_;
  assign new_n52778_ = new_n17092_ & new_n52777_;
  assign new_n52779_ = new_n12299_ & new_n52750_;
  assign new_n52780_ = ys__n530 & ys__n752;
  assign new_n52781_ = ~new_n12303_ & ~new_n52780_;
  assign new_n52782_ = ~new_n52779_ & new_n52781_;
  assign new_n52783_ = ~new_n52778_ & new_n52782_;
  assign new_n52784_ = new_n17092_ & new_n52767_;
  assign new_n52785_ = ys__n522 & ~ys__n530;
  assign new_n52786_ = ~ys__n524 & ys__n526;
  assign new_n52787_ = ~ys__n752 & new_n52786_;
  assign new_n52788_ = new_n52785_ & new_n52787_;
  assign new_n52789_ = ~new_n52784_ & ~new_n52788_;
  assign new_n52790_ = ys__n524 & ys__n526;
  assign new_n52791_ = ~ys__n752 & new_n52790_;
  assign new_n52792_ = new_n52785_ & new_n52791_;
  assign new_n52793_ = ~ys__n524 & ~ys__n526;
  assign new_n52794_ = ys__n752 & new_n52793_;
  assign new_n52795_ = new_n52785_ & new_n52794_;
  assign new_n52796_ = ~new_n52792_ & ~new_n52795_;
  assign new_n52797_ = new_n52789_ & new_n52796_;
  assign new_n52798_ = new_n52783_ & new_n52797_;
  assign new_n52799_ = new_n17097_ & ~new_n52798_;
  assign new_n52800_ = ys__n744 & ys__n746;
  assign new_n52801_ = ys__n742 & ys__n750;
  assign new_n52802_ = new_n52800_ & new_n52801_;
  assign new_n52803_ = ys__n748 & new_n52802_;
  assign new_n52804_ = new_n11765_ & new_n52728_;
  assign new_n52805_ = new_n12338_ & new_n52728_;
  assign new_n52806_ = ~new_n52804_ & ~new_n52805_;
  assign new_n52807_ = ~new_n52803_ & new_n52806_;
  assign new_n52808_ = ~ys__n742 & ys__n748;
  assign new_n52809_ = ~ys__n750 & new_n52808_;
  assign new_n52810_ = new_n52800_ & new_n52809_;
  assign new_n52811_ = new_n11792_ & new_n52737_;
  assign new_n52812_ = ~new_n52810_ & ~new_n52811_;
  assign new_n52813_ = new_n11791_ & new_n52728_;
  assign new_n52814_ = new_n52728_ & new_n52748_;
  assign new_n52815_ = ~new_n52813_ & ~new_n52814_;
  assign new_n52816_ = new_n52812_ & new_n52815_;
  assign new_n52817_ = new_n11775_ & new_n12297_;
  assign new_n52818_ = new_n12297_ & new_n52730_;
  assign new_n52819_ = ~new_n52817_ & ~new_n52818_;
  assign new_n52820_ = new_n11764_ & new_n11792_;
  assign new_n52821_ = new_n11775_ & new_n52728_;
  assign new_n52822_ = ~new_n52820_ & ~new_n52821_;
  assign new_n52823_ = new_n52819_ & new_n52822_;
  assign new_n52824_ = ~ys__n748 & new_n52802_;
  assign new_n52825_ = ~new_n11804_ & ~new_n52824_;
  assign new_n52826_ = new_n52823_ & new_n52825_;
  assign new_n52827_ = new_n52816_ & new_n52826_;
  assign new_n52828_ = new_n52807_ & new_n52827_;
  assign new_n52829_ = new_n12301_ & new_n52780_;
  assign new_n52830_ = new_n11765_ & new_n12297_;
  assign new_n52831_ = ~new_n52829_ & new_n52830_;
  assign new_n52832_ = new_n12303_ & new_n52636_;
  assign new_n52833_ = new_n12298_ & new_n52832_;
  assign new_n52834_ = ~new_n52831_ & ~new_n52833_;
  assign new_n52835_ = new_n52828_ & new_n52834_;
  assign new_n52836_ = ~new_n52799_ & new_n52835_;
  assign new_n52837_ = ~new_n12298_ & ~new_n17097_;
  assign new_n52838_ = ~new_n52830_ & new_n52837_;
  assign new_n52839_ = new_n52828_ & new_n52838_;
  assign new_n52840_ = ~ys__n28243 & ~new_n52839_;
  assign new_n52841_ = ~new_n52836_ & new_n52840_;
  assign new_n52842_ = new_n11764_ & new_n11801_;
  assign new_n52843_ = new_n11766_ & new_n52842_;
  assign new_n52844_ = ~new_n12334_ & ~new_n52843_;
  assign new_n52845_ = new_n11792_ & new_n12333_;
  assign new_n52846_ = new_n11792_ & new_n52842_;
  assign new_n52847_ = ~new_n52845_ & ~new_n52846_;
  assign new_n52848_ = new_n52844_ & new_n52847_;
  assign new_n52849_ = ~new_n11767_ & ~new_n12332_;
  assign new_n52850_ = new_n11765_ & new_n11792_;
  assign new_n52851_ = ~new_n12384_ & ~new_n52749_;
  assign new_n52852_ = ~new_n52850_ & new_n52851_;
  assign new_n52853_ = new_n52849_ & new_n52852_;
  assign new_n52854_ = new_n52848_ & new_n52853_;
  assign new_n52855_ = ys__n47659 & new_n12384_;
  assign new_n52856_ = ys__n530 & new_n52749_;
  assign new_n52857_ = ~new_n12391_ & ~new_n52752_;
  assign new_n52858_ = new_n52850_ & ~new_n52857_;
  assign new_n52859_ = ~new_n52856_ & ~new_n52858_;
  assign new_n52860_ = ~new_n52855_ & new_n52859_;
  assign new_n52861_ = ys__n550 & new_n11770_;
  assign new_n52862_ = ~ys__n518 & ys__n548;
  assign new_n52863_ = ys__n550 & new_n52862_;
  assign new_n52864_ = ~new_n52861_ & ~new_n52863_;
  assign new_n52865_ = new_n11767_ & ~new_n52864_;
  assign new_n52866_ = new_n12332_ & new_n17093_;
  assign new_n52867_ = ~new_n52865_ & ~new_n52866_;
  assign new_n52868_ = new_n52848_ & new_n52867_;
  assign new_n52869_ = new_n52860_ & new_n52868_;
  assign new_n52870_ = ys__n28243 & ~new_n52869_;
  assign new_n52871_ = ~new_n52854_ & new_n52870_;
  assign new_n52872_ = ~new_n52841_ & ~new_n52871_;
  assign ys__n38360 = ~ys__n4566 & ~new_n52872_;
  assign ys__n38362 = ys__n38361 & ~ys__n4566;
  assign new_n52875_ = ys__n520 & new_n52780_;
  assign new_n52876_ = new_n52636_ & new_n52875_;
  assign new_n52877_ = new_n52726_ & new_n52876_;
  assign ys__n38364 = ~ys__n4566 & new_n52877_;
  assign new_n52879_ = ~ys__n512 & ~ys__n520;
  assign new_n52880_ = ~ys__n632 & new_n52879_;
  assign new_n52881_ = new_n12344_ & new_n52880_;
  assign new_n52882_ = ys__n23705 & ~ys__n28243;
  assign new_n52883_ = new_n12298_ & new_n52882_;
  assign new_n52884_ = new_n52881_ & new_n52883_;
  assign ys__n38365 = ~ys__n4566 & new_n52884_;
  assign new_n52886_ = ys__n23706 & ~ys__n28243;
  assign new_n52887_ = new_n12298_ & new_n52886_;
  assign new_n52888_ = new_n52881_ & new_n52887_;
  assign ys__n38366 = ~ys__n4566 & new_n52888_;
  assign new_n52890_ = ys__n23707 & ~ys__n28243;
  assign new_n52891_ = new_n12298_ & new_n52890_;
  assign new_n52892_ = new_n52881_ & new_n52891_;
  assign ys__n38367 = ~ys__n4566 & new_n52892_;
  assign new_n52894_ = ys__n23708 & ~ys__n28243;
  assign new_n52895_ = new_n12298_ & new_n52894_;
  assign new_n52896_ = new_n52881_ & new_n52895_;
  assign ys__n38368 = ~ys__n4566 & new_n52896_;
  assign new_n52898_ = ys__n23709 & ~ys__n28243;
  assign new_n52899_ = new_n12298_ & new_n52898_;
  assign new_n52900_ = new_n52881_ & new_n52899_;
  assign ys__n38369 = ~ys__n4566 & new_n52900_;
  assign new_n52902_ = ys__n23710 & ~ys__n28243;
  assign new_n52903_ = new_n12298_ & new_n52902_;
  assign new_n52904_ = new_n52881_ & new_n52903_;
  assign ys__n38370 = ~ys__n4566 & new_n52904_;
  assign new_n52906_ = ys__n23711 & ~ys__n28243;
  assign new_n52907_ = new_n12298_ & new_n52906_;
  assign new_n52908_ = new_n52881_ & new_n52907_;
  assign ys__n38371 = ~ys__n4566 & new_n52908_;
  assign new_n52910_ = ys__n23712 & ~ys__n28243;
  assign new_n52911_ = new_n12298_ & new_n52910_;
  assign new_n52912_ = new_n52881_ & new_n52911_;
  assign ys__n38372 = ~ys__n4566 & new_n52912_;
  assign new_n52914_ = ys__n23713 & ~ys__n28243;
  assign new_n52915_ = new_n12298_ & new_n52914_;
  assign new_n52916_ = new_n52881_ & new_n52915_;
  assign ys__n38373 = ~ys__n4566 & new_n52916_;
  assign new_n52918_ = ys__n23714 & ~ys__n28243;
  assign new_n52919_ = new_n12298_ & new_n52918_;
  assign new_n52920_ = new_n52881_ & new_n52919_;
  assign ys__n38374 = ~ys__n4566 & new_n52920_;
  assign new_n52922_ = ys__n23715 & ~ys__n28243;
  assign new_n52923_ = new_n12298_ & new_n52922_;
  assign new_n52924_ = new_n52881_ & new_n52923_;
  assign ys__n38375 = ~ys__n4566 & new_n52924_;
  assign ys__n38377 = ys__n38376 & ~ys__n4566;
  assign ys__n38379 = ys__n38378 & ~ys__n4566;
  assign ys__n38381 = ys__n38380 & ~ys__n4566;
  assign ys__n38383 = ys__n38382 & ~ys__n4566;
  assign ys__n38385 = ys__n38384 & ~ys__n4566;
  assign ys__n38387 = ys__n38386 & ~ys__n4566;
  assign new_n52932_ = ys__n632 & new_n52879_;
  assign new_n52933_ = new_n12344_ & new_n52932_;
  assign new_n52934_ = ys__n634 & ys__n636;
  assign new_n52935_ = ~ys__n638 & ~ys__n640;
  assign new_n52936_ = ~ys__n642 & ~ys__n28243;
  assign new_n52937_ = new_n52935_ & new_n52936_;
  assign new_n52938_ = new_n52934_ & new_n52937_;
  assign new_n52939_ = new_n12298_ & new_n52938_;
  assign new_n52940_ = new_n52933_ & new_n52939_;
  assign ys__n38388 = ~ys__n4566 & new_n52940_;
  assign new_n52942_ = ~ys__n638 & ys__n640;
  assign new_n52943_ = new_n52934_ & new_n52936_;
  assign new_n52944_ = new_n52942_ & new_n52943_;
  assign new_n52945_ = new_n12298_ & new_n52944_;
  assign new_n52946_ = new_n52933_ & new_n52945_;
  assign ys__n38389 = ~ys__n4566 & new_n52946_;
  assign new_n52948_ = ~ys__n634 & ys__n636;
  assign new_n52949_ = new_n12699_ & new_n52948_;
  assign new_n52950_ = new_n52935_ & new_n52949_;
  assign new_n52951_ = new_n12298_ & new_n52950_;
  assign new_n52952_ = new_n52933_ & new_n52951_;
  assign ys__n38390 = ~ys__n4566 & new_n52952_;
  assign new_n52954_ = ~ys__n634 & ~ys__n636;
  assign new_n52955_ = new_n12699_ & new_n52935_;
  assign new_n52956_ = new_n52954_ & new_n52955_;
  assign new_n52957_ = new_n12298_ & new_n52956_;
  assign new_n52958_ = new_n52933_ & new_n52957_;
  assign ys__n38391 = ~ys__n4566 & new_n52958_;
  assign new_n52960_ = new_n12699_ & new_n52942_;
  assign new_n52961_ = new_n52954_ & new_n52960_;
  assign new_n52962_ = new_n12298_ & new_n52961_;
  assign new_n52963_ = new_n52933_ & new_n52962_;
  assign ys__n38392 = ~ys__n4566 & new_n52963_;
  assign new_n52965_ = ys__n640 & ys__n642;
  assign new_n52966_ = new_n12600_ & new_n52965_;
  assign new_n52967_ = new_n52934_ & new_n52966_;
  assign new_n52968_ = new_n12298_ & new_n52967_;
  assign new_n52969_ = new_n52933_ & new_n52968_;
  assign ys__n38393 = ~ys__n4566 & new_n52969_;
  assign new_n52971_ = ~ys__n4458 & ~ys__n4461;
  assign new_n52972_ = ~ys__n4465 & new_n52971_;
  assign new_n52973_ = ~ys__n4454 & ~ys__n4455;
  assign new_n52974_ = new_n35223_ & new_n52973_;
  assign new_n52975_ = new_n35099_ & new_n35261_;
  assign new_n52976_ = new_n52974_ & new_n52975_;
  assign new_n52977_ = new_n52972_ & new_n52976_;
  assign ys__n38394 = ~ys__n4566 & ~new_n52977_;
  assign new_n52979_ = ~ys__n28243 & new_n12344_;
  assign new_n52980_ = new_n12350_ & new_n52979_;
  assign new_n52981_ = new_n12393_ & new_n52980_;
  assign new_n52982_ = ~ys__n516 & ~ys__n550;
  assign new_n52983_ = new_n11770_ & new_n52982_;
  assign new_n52984_ = new_n12304_ & new_n52983_;
  assign new_n52985_ = ~ys__n640 & ~ys__n642;
  assign new_n52986_ = ~ys__n736 & ~ys__n4488;
  assign new_n52987_ = new_n52985_ & new_n52986_;
  assign new_n52988_ = ~ys__n632 & ~ys__n634;
  assign new_n52989_ = ~ys__n636 & ~ys__n638;
  assign new_n52990_ = new_n52988_ & new_n52989_;
  assign new_n52991_ = new_n52987_ & new_n52990_;
  assign new_n52992_ = new_n52984_ & new_n52991_;
  assign new_n52993_ = new_n12298_ & new_n52992_;
  assign new_n52994_ = new_n52981_ & new_n52993_;
  assign ys__n38396 = ~ys__n4566 & new_n52994_;
  assign new_n52996_ = ~ys__n28243 & new_n52829_;
  assign new_n52997_ = new_n52830_ & new_n52996_;
  assign new_n52998_ = ~ys__n23730 & new_n52768_;
  assign new_n52999_ = new_n52777_ & new_n52998_;
  assign new_n53000_ = new_n12384_ & new_n52999_;
  assign new_n53001_ = ~new_n52997_ & ~new_n53000_;
  assign ys__n38397 = ~ys__n4566 & ~new_n53001_;
  assign new_n53003_ = new_n19558_ & ~new_n21909_;
  assign new_n53004_ = ~new_n19558_ & new_n21909_;
  assign new_n53005_ = ~new_n53003_ & ~new_n53004_;
  assign new_n53006_ = ys__n38418 & ~ys__n4566;
  assign ys__n38417 = ~new_n53005_ & new_n53006_;
  assign new_n53008_ = new_n12124_ & new_n12137_;
  assign new_n53009_ = ys__n23717 & ys__n33403;
  assign new_n53010_ = ~new_n53008_ & new_n53009_;
  assign new_n53011_ = new_n12140_ & new_n53010_;
  assign new_n53012_ = ~ys__n935 & ~ys__n38473;
  assign new_n53013_ = ys__n33403 & new_n12127_;
  assign new_n53014_ = new_n53012_ & ~new_n53013_;
  assign new_n53015_ = ~new_n12124_ & ~new_n53014_;
  assign new_n53016_ = ys__n738 & new_n53015_;
  assign new_n53017_ = ys__n935 & ~new_n12124_;
  assign new_n53018_ = new_n13717_ & new_n53017_;
  assign new_n53019_ = ~new_n53016_ & ~new_n53018_;
  assign new_n53020_ = ~new_n53011_ & new_n53019_;
  assign new_n53021_ = ~new_n45599_ & ~new_n53020_;
  assign new_n53022_ = ~new_n13689_ & ~new_n13763_;
  assign new_n53023_ = ~new_n42890_ & ~new_n42905_;
  assign new_n53024_ = new_n13763_ & ~new_n53023_;
  assign new_n53025_ = ~new_n53022_ & ~new_n53024_;
  assign new_n53026_ = ~ys__n33396 & ~ys__n33398;
  assign new_n53027_ = ys__n33403 & new_n53026_;
  assign new_n53028_ = ~ys__n4566 & new_n53027_;
  assign new_n53029_ = new_n12140_ & new_n53028_;
  assign new_n53030_ = ~new_n53025_ & new_n53029_;
  assign new_n53031_ = new_n53012_ & ~new_n53028_;
  assign new_n53032_ = ys__n738 & ~new_n53031_;
  assign new_n53033_ = ~new_n53025_ & new_n53032_;
  assign new_n53034_ = ys__n935 & new_n13689_;
  assign new_n53035_ = ys__n935 & ~new_n53034_;
  assign new_n53036_ = new_n13717_ & new_n53035_;
  assign new_n53037_ = ~new_n53033_ & ~new_n53036_;
  assign new_n53038_ = ~new_n53030_ & new_n53037_;
  assign new_n53039_ = ~new_n45599_ & ~new_n53038_;
  assign new_n53040_ = ~new_n53021_ & ~new_n53039_;
  assign ys__n38456 = ys__n30863 & ~new_n53040_;
  assign new_n53042_ = ~ys__n626 & ys__n664;
  assign new_n53043_ = new_n23014_ & new_n53042_;
  assign new_n53044_ = ~ys__n662 & ~ys__n668;
  assign new_n53045_ = new_n23013_ & new_n53044_;
  assign new_n53046_ = new_n53042_ & new_n53045_;
  assign new_n53047_ = ys__n662 & ~ys__n668;
  assign new_n53048_ = new_n23013_ & new_n53042_;
  assign new_n53049_ = new_n53047_ & new_n53048_;
  assign new_n53050_ = ~new_n53046_ & ~new_n53049_;
  assign new_n53051_ = ~new_n53043_ & new_n53050_;
  assign ys__n38508 = ys__n33414 & ~new_n53051_;
  assign new_n53053_ = new_n22986_ & new_n53044_;
  assign new_n53054_ = new_n53042_ & new_n53053_;
  assign new_n53055_ = ys__n660 & ~ys__n666;
  assign new_n53056_ = new_n53042_ & new_n53044_;
  assign new_n53057_ = new_n53055_ & new_n53056_;
  assign new_n53058_ = ~new_n53054_ & ~new_n53057_;
  assign new_n53059_ = new_n22987_ & new_n53042_;
  assign new_n53060_ = new_n22986_ & new_n53042_;
  assign new_n53061_ = new_n53047_ & new_n53060_;
  assign new_n53062_ = new_n53042_ & new_n53047_;
  assign new_n53063_ = new_n53055_ & new_n53062_;
  assign new_n53064_ = ~new_n53061_ & ~new_n53063_;
  assign new_n53065_ = ~new_n53059_ & new_n53064_;
  assign new_n53066_ = new_n53058_ & new_n53065_;
  assign ys__n38509 = ys__n33414 & ~new_n53066_;
  assign ys__n38510 = ys__n846 | ~new_n23752_;
  assign ys__n38515 = ~ys__n18120 & new_n23194_;
  assign new_n53070_ = ~ys__n33431 & ys__n38553;
  assign new_n53071_ = ~ys__n24131 & ~new_n53070_;
  assign ys__n38518 = ~ys__n1036 & ~new_n53071_;
  assign new_n53073_ = ys__n24145 & ys__n38518;
  assign ys__n38520 = ~ys__n24145 | new_n53073_;
  assign new_n53075_ = ~ys__n4185 & new_n23148_;
  assign ys__n38523 = ys__n38522 | new_n53075_;
  assign ys__n38525 = ys__n1029 | ys__n1036;
  assign new_n53078_ = ys__n33442 & ~ys__n18120;
  assign ys__n38552 = new_n23521_ & ~new_n53078_;
  assign new_n53080_ = ~ys__n24228 & ~new_n53070_;
  assign ys__n38555 = ~ys__n1076 & ~new_n53080_;
  assign new_n53082_ = ys__n24236 & ys__n38555;
  assign ys__n38563 = ~ys__n24236 | new_n53082_;
  assign new_n53084_ = ys__n33491 & ys__n33497;
  assign new_n53085_ = ~ys__n33495 & ~new_n53084_;
  assign new_n53086_ = ~ys__n4566 & new_n53085_;
  assign ys__n38615 = ys__n24271 & new_n53086_;
  assign new_n53088_ = ~ys__n33451 & ys__n38620;
  assign new_n53089_ = ~ys__n33499 & ~new_n53088_;
  assign ys__n38623 = ~ys__n1094 & ~new_n53089_;
  assign ys__n38650 = ~ys__n33455 & ys__n33454;
  assign new_n53092_ = ~ys__n33457 & ys__n24268;
  assign new_n53093_ = ys__n24502 & new_n53092_;
  assign ys__n38662 = ys__n24255 | new_n53093_;
  assign new_n53095_ = ~ys__n24447 & ~ys__n24541;
  assign new_n53096_ = ~ys__n24502 & new_n53095_;
  assign new_n53097_ = new_n17716_ & ys__n38623;
  assign new_n53098_ = ~ys__n4566 & new_n53097_;
  assign new_n53099_ = ~ys__n24259 & new_n53098_;
  assign new_n53100_ = ~ys__n24262 & new_n53099_;
  assign new_n53101_ = ys__n24502 & new_n53100_;
  assign ys__n38668 = new_n53096_ | new_n53101_;
  assign ys__n38669 = ys__n38662 | ys__n38668;
  assign new_n53104_ = ys__n18214 & ~ys__n18216;
  assign ys__n38672 = ys__n18218 & new_n53104_;
  assign new_n53106_ = ys__n1511 & ys__n30216;
  assign ys__n38674 = ~ys__n4566 & new_n53106_;
  assign new_n53108_ = ys__n1110 & ys__n33488;
  assign ys__n38689 = new_n24561_ | new_n53108_;
  assign new_n53110_ = ys__n33552 & new_n13606_;
  assign new_n53111_ = ~new_n24498_ & ~new_n53110_;
  assign new_n53112_ = ~ys__n33491 & ~new_n53111_;
  assign new_n53113_ = ~ys__n33491 & ys__n33552;
  assign new_n53114_ = new_n13606_ & ~new_n53113_;
  assign new_n53115_ = ~new_n23601_ & new_n53114_;
  assign new_n53116_ = ~new_n53112_ & ~new_n53115_;
  assign new_n53117_ = ~ys__n4566 & new_n23581_;
  assign new_n53118_ = ~new_n53116_ & new_n53117_;
  assign ys__n38742 = ~ys__n4696 & new_n53118_;
  assign new_n53120_ = ys__n1106 & new_n13606_;
  assign new_n53121_ = ~new_n53113_ & new_n53120_;
  assign new_n53122_ = new_n17716_ & new_n53121_;
  assign new_n53123_ = ~new_n23601_ & new_n53122_;
  assign new_n53124_ = new_n23580_ & new_n53123_;
  assign new_n53125_ = ~ys__n4566 & new_n53124_;
  assign ys__n38768 = ~ys__n4696 & new_n53125_;
  assign ys__n38795 = ys__n33515 & ys__n33514;
  assign new_n53128_ = ~ys__n24581 & ~ys__n24604;
  assign new_n53129_ = new_n17742_ & new_n53128_;
  assign ys__n38799 = ys__n18136 | new_n53129_;
  assign ys__n38884 = ~ys__n29117 & ys__n38883;
  assign ys__n38886 = ~ys__n29117 & ys__n38885;
  assign new_n53133_ = ys__n48 & ~ys__n50;
  assign new_n53134_ = ys__n52 & new_n53133_;
  assign new_n53135_ = ys__n56 & ys__n58;
  assign new_n53136_ = ys__n60 & ys__n62;
  assign new_n53137_ = new_n53135_ & new_n53136_;
  assign new_n53138_ = ys__n48 & ys__n50;
  assign new_n53139_ = ys__n52 & ys__n54;
  assign new_n53140_ = new_n53138_ & new_n53139_;
  assign new_n53141_ = new_n53137_ & new_n53140_;
  assign ys__n38887 = new_n53134_ | new_n53141_;
  assign ys__n38900 = ~ys__n33558 & ys__n740;
  assign new_n53144_ = ys__n30214 & ~ys__n3039;
  assign ys__n38912 = ys__n23850 | new_n53144_;
  assign ys__n38913 = ys__n30217 & ~ys__n4566;
  assign new_n53147_ = ys__n30216 & ~ys__n740;
  assign new_n53148_ = ys__n30217 & ys__n740;
  assign new_n53149_ = ~new_n53147_ & ~new_n53148_;
  assign ys__n38914 = ~ys__n4566 & ~new_n53149_;
  assign new_n53151_ = ys__n30219 & ~ys__n740;
  assign new_n53152_ = ys__n30220 & ys__n740;
  assign new_n53153_ = ~new_n53151_ & ~new_n53152_;
  assign ys__n38915 = ~ys__n4566 & ~new_n53153_;
  assign new_n53155_ = ys__n30225 & ~ys__n30223;
  assign ys__n38917 = ys__n1020 | new_n53155_;
  assign new_n53157_ = ys__n28438 & ~ys__n33574;
  assign new_n53158_ = ys__n28434 & ~ys__n33570;
  assign new_n53159_ = ys__n28436 & ~ys__n33572;
  assign new_n53160_ = ~new_n53158_ & ~new_n53159_;
  assign new_n53161_ = ~new_n53157_ & new_n53160_;
  assign new_n53162_ = ys__n28428 & ~ys__n33564;
  assign new_n53163_ = ~ys__n38277 & ~new_n53162_;
  assign new_n53164_ = ys__n28430 & ~ys__n33566;
  assign new_n53165_ = ys__n28432 & ~ys__n33568;
  assign new_n53166_ = ~new_n53164_ & ~new_n53165_;
  assign new_n53167_ = new_n53163_ & new_n53166_;
  assign ys__n38923 = ~new_n53161_ | ~new_n53167_;
  assign new_n53169_ = ~ys__n33576 & ys__n38927;
  assign new_n53170_ = ys__n38928 & ys__n38929;
  assign ys__n38925 = new_n53169_ & new_n53170_;
  assign ys__n38930 = ~ys__n398 & ~new_n15136_;
  assign new_n53173_ = ys__n196 & ys__n198;
  assign new_n53174_ = ~ys__n2830 & new_n53173_;
  assign new_n53175_ = ys__n196 & ys__n2830;
  assign new_n53176_ = ~ys__n196 & ~ys__n2830;
  assign new_n53177_ = ~new_n53175_ & ~new_n53176_;
  assign new_n53178_ = ~new_n53174_ & new_n53177_;
  assign new_n53179_ = ~ys__n196 & new_n42060_;
  assign new_n53180_ = ys__n196 & ~ys__n198;
  assign new_n53181_ = ~ys__n2830 & new_n53180_;
  assign new_n53182_ = ~ys__n196 & new_n53175_;
  assign new_n53183_ = ~new_n53181_ & ~new_n53182_;
  assign new_n53184_ = ~new_n53179_ & new_n53183_;
  assign new_n53185_ = new_n53178_ & new_n53184_;
  assign new_n53186_ = ys__n48259 & new_n53181_;
  assign new_n53187_ = ys__n48259 & new_n53175_;
  assign ys__n44968 = ys__n352 & ys__n27855;
  assign new_n53189_ = new_n53176_ & ys__n44968;
  assign new_n53190_ = ~new_n53187_ & ~new_n53189_;
  assign new_n53191_ = ~new_n53186_ & new_n53190_;
  assign new_n53192_ = new_n53179_ & ys__n44968;
  assign new_n53193_ = ys__n48259 & new_n53174_;
  assign ys__n44952 = ys__n352 & ys__n28015;
  assign new_n53195_ = new_n53182_ & ys__n44952;
  assign new_n53196_ = ~new_n53193_ & ~new_n53195_;
  assign new_n53197_ = ~new_n53192_ & new_n53196_;
  assign new_n53198_ = new_n53191_ & new_n53197_;
  assign new_n53199_ = ~new_n53185_ & ~new_n53198_;
  assign new_n53200_ = ys__n48275 & new_n53174_;
  assign new_n53201_ = ~new_n53185_ & new_n53200_;
  assign new_n53202_ = new_n53199_ & ~new_n53201_;
  assign new_n53203_ = new_n53199_ & ~new_n53202_;
  assign new_n53204_ = ys__n48260 & new_n53181_;
  assign new_n53205_ = ys__n48260 & new_n53175_;
  assign ys__n44969 = ys__n352 & ys__n27857;
  assign new_n53207_ = new_n53176_ & ys__n44969;
  assign new_n53208_ = ~new_n53205_ & ~new_n53207_;
  assign new_n53209_ = ~new_n53204_ & new_n53208_;
  assign new_n53210_ = new_n53179_ & ys__n44969;
  assign new_n53211_ = ys__n48260 & new_n53174_;
  assign ys__n44953 = ys__n352 & ys__n28016;
  assign new_n53213_ = new_n53182_ & ys__n44953;
  assign new_n53214_ = ~new_n53211_ & ~new_n53213_;
  assign new_n53215_ = ~new_n53210_ & new_n53214_;
  assign new_n53216_ = new_n53209_ & new_n53215_;
  assign new_n53217_ = ~new_n53185_ & ~new_n53216_;
  assign new_n53218_ = ~new_n53203_ & ~new_n53217_;
  assign new_n53219_ = ys__n48261 & new_n53181_;
  assign new_n53220_ = ys__n48261 & new_n53175_;
  assign ys__n44970 = ys__n352 & ys__n27859;
  assign new_n53222_ = new_n53176_ & ys__n44970;
  assign new_n53223_ = ~new_n53220_ & ~new_n53222_;
  assign new_n53224_ = ~new_n53219_ & new_n53223_;
  assign new_n53225_ = new_n53179_ & ys__n44970;
  assign new_n53226_ = ys__n48261 & new_n53174_;
  assign ys__n44954 = ys__n352 & ys__n28017;
  assign new_n53228_ = new_n53182_ & ys__n44954;
  assign new_n53229_ = ~new_n53226_ & ~new_n53228_;
  assign new_n53230_ = ~new_n53225_ & new_n53229_;
  assign new_n53231_ = new_n53224_ & new_n53230_;
  assign new_n53232_ = ~new_n53185_ & ~new_n53231_;
  assign new_n53233_ = new_n53218_ & ~new_n53232_;
  assign new_n53234_ = ~new_n53199_ & ~new_n53201_;
  assign new_n53235_ = new_n53217_ & new_n53234_;
  assign new_n53236_ = new_n53217_ & ~new_n53235_;
  assign new_n53237_ = new_n53232_ & ~new_n53236_;
  assign new_n53238_ = ~new_n53233_ & ~new_n53237_;
  assign new_n53239_ = ys__n162 & ~ys__n346;
  assign new_n53240_ = new_n13473_ & new_n53239_;
  assign new_n53241_ = ys__n352 & new_n42806_;
  assign new_n53242_ = new_n53240_ & new_n53241_;
  assign new_n53243_ = ys__n352 & new_n42813_;
  assign new_n53244_ = new_n53240_ & new_n53243_;
  assign new_n53245_ = ~new_n53242_ & ~new_n53244_;
  assign new_n53246_ = new_n13732_ & new_n53240_;
  assign new_n53247_ = new_n13478_ & new_n13730_;
  assign new_n53248_ = ys__n352 & new_n53240_;
  assign new_n53249_ = new_n53247_ & new_n53248_;
  assign new_n53250_ = ~new_n53246_ & ~new_n53249_;
  assign new_n53251_ = new_n53245_ & new_n53250_;
  assign new_n53252_ = new_n42811_ & new_n42824_;
  assign new_n53253_ = new_n13738_ & new_n42815_;
  assign new_n53254_ = new_n53252_ & new_n53253_;
  assign new_n53255_ = ~ys__n196 & ys__n948;
  assign ys__n44836 = ~new_n53254_ & new_n53255_;
  assign new_n53257_ = ys__n1817 & ys__n44836;
  assign new_n53258_ = new_n53251_ & ~new_n53257_;
  assign new_n53259_ = ys__n948 & ~new_n53258_;
  assign new_n53260_ = ys__n196 & ys__n44833;
  assign new_n53261_ = ~new_n53259_ & ~new_n53260_;
  assign new_n53262_ = new_n53238_ & ~new_n53261_;
  assign new_n53263_ = ~new_n53238_ & new_n53261_;
  assign ys__n39395 = new_n53262_ | new_n53263_;
  assign new_n53265_ = new_n53199_ & new_n53201_;
  assign new_n53266_ = ~new_n53217_ & new_n53265_;
  assign new_n53267_ = ~new_n53235_ & ~new_n53266_;
  assign new_n53268_ = ~new_n53232_ & ~new_n53267_;
  assign new_n53269_ = ~new_n53199_ & new_n53201_;
  assign new_n53270_ = ~new_n53199_ & ~new_n53269_;
  assign new_n53271_ = new_n53217_ & ~new_n53270_;
  assign new_n53272_ = ~new_n53218_ & ~new_n53271_;
  assign new_n53273_ = new_n53232_ & ~new_n53272_;
  assign new_n53274_ = ~new_n53268_ & ~new_n53273_;
  assign new_n53275_ = ~new_n53261_ & new_n53274_;
  assign new_n53276_ = new_n53261_ & ~new_n53274_;
  assign ys__n39396 = new_n53275_ | new_n53276_;
  assign new_n53278_ = ~new_n53217_ & new_n53234_;
  assign new_n53279_ = ~new_n53202_ & ~new_n53269_;
  assign new_n53280_ = new_n53217_ & ~new_n53279_;
  assign new_n53281_ = ~new_n53278_ & ~new_n53280_;
  assign new_n53282_ = ~new_n53232_ & ~new_n53281_;
  assign new_n53283_ = ~new_n53234_ & ~new_n53265_;
  assign new_n53284_ = ~new_n53217_ & ~new_n53283_;
  assign new_n53285_ = ~new_n53203_ & new_n53217_;
  assign new_n53286_ = ~new_n53284_ & ~new_n53285_;
  assign new_n53287_ = new_n53232_ & ~new_n53286_;
  assign new_n53288_ = ~new_n53282_ & ~new_n53287_;
  assign new_n53289_ = ~new_n53261_ & new_n53288_;
  assign new_n53290_ = new_n53261_ & ~new_n53288_;
  assign ys__n39397 = new_n53289_ | new_n53290_;
  assign new_n53292_ = new_n53217_ & ~new_n53232_;
  assign new_n53293_ = new_n53265_ & new_n53292_;
  assign new_n53294_ = ~new_n53217_ & ~new_n53270_;
  assign new_n53295_ = ~new_n53217_ & ~new_n53294_;
  assign new_n53296_ = new_n53232_ & ~new_n53295_;
  assign new_n53297_ = ~new_n53293_ & ~new_n53296_;
  assign new_n53298_ = ~new_n53261_ & new_n53297_;
  assign new_n53299_ = new_n53261_ & ~new_n53297_;
  assign ys__n39398 = new_n53298_ | new_n53299_;
  assign new_n53301_ = ys__n48262 & new_n53181_;
  assign new_n53302_ = ys__n48262 & new_n53175_;
  assign ys__n44971 = ys__n352 & ys__n27861;
  assign new_n53304_ = new_n53176_ & ys__n44971;
  assign new_n53305_ = ~new_n53302_ & ~new_n53304_;
  assign new_n53306_ = ~new_n53301_ & new_n53305_;
  assign new_n53307_ = new_n53179_ & ys__n44971;
  assign new_n53308_ = ys__n48262 & new_n53174_;
  assign ys__n44955 = ys__n352 & ys__n28018;
  assign new_n53310_ = new_n53182_ & ys__n44955;
  assign new_n53311_ = ~new_n53308_ & ~new_n53310_;
  assign new_n53312_ = ~new_n53307_ & new_n53311_;
  assign new_n53313_ = new_n53306_ & new_n53312_;
  assign new_n53314_ = ~new_n53185_ & ~new_n53313_;
  assign new_n53315_ = ~new_n53232_ & new_n53314_;
  assign new_n53316_ = new_n53314_ & ~new_n53315_;
  assign new_n53317_ = ys__n48263 & new_n53181_;
  assign new_n53318_ = ys__n48263 & new_n53175_;
  assign ys__n44972 = ys__n352 & ys__n27863;
  assign new_n53320_ = new_n53176_ & ys__n44972;
  assign new_n53321_ = ~new_n53318_ & ~new_n53320_;
  assign new_n53322_ = ~new_n53317_ & new_n53321_;
  assign new_n53323_ = new_n53179_ & ys__n44972;
  assign new_n53324_ = ys__n48263 & new_n53174_;
  assign ys__n44956 = ys__n352 & ys__n28019;
  assign new_n53326_ = new_n53182_ & ys__n44956;
  assign new_n53327_ = ~new_n53324_ & ~new_n53326_;
  assign new_n53328_ = ~new_n53323_ & new_n53327_;
  assign new_n53329_ = new_n53322_ & new_n53328_;
  assign new_n53330_ = ~new_n53185_ & ~new_n53329_;
  assign new_n53331_ = ~new_n53316_ & ~new_n53330_;
  assign new_n53332_ = ys__n48264 & new_n53181_;
  assign new_n53333_ = ys__n48264 & new_n53175_;
  assign ys__n44973 = ys__n352 & ys__n27865;
  assign new_n53335_ = new_n53176_ & ys__n44973;
  assign new_n53336_ = ~new_n53333_ & ~new_n53335_;
  assign new_n53337_ = ~new_n53332_ & new_n53336_;
  assign new_n53338_ = new_n53179_ & ys__n44973;
  assign new_n53339_ = ys__n48264 & new_n53174_;
  assign ys__n44957 = ys__n352 & ys__n28020;
  assign new_n53341_ = new_n53182_ & ys__n44957;
  assign new_n53342_ = ~new_n53339_ & ~new_n53341_;
  assign new_n53343_ = ~new_n53338_ & new_n53342_;
  assign new_n53344_ = new_n53337_ & new_n53343_;
  assign new_n53345_ = ~new_n53185_ & ~new_n53344_;
  assign new_n53346_ = new_n53331_ & ~new_n53345_;
  assign new_n53347_ = ~new_n53232_ & ~new_n53314_;
  assign new_n53348_ = new_n53330_ & new_n53347_;
  assign new_n53349_ = new_n53330_ & ~new_n53348_;
  assign new_n53350_ = new_n53345_ & ~new_n53349_;
  assign new_n53351_ = ~new_n53346_ & ~new_n53350_;
  assign new_n53352_ = ~new_n53261_ & new_n53351_;
  assign new_n53353_ = new_n53261_ & ~new_n53351_;
  assign ys__n39399 = new_n53352_ | new_n53353_;
  assign new_n53355_ = new_n53232_ & new_n53314_;
  assign new_n53356_ = ~new_n53330_ & new_n53355_;
  assign new_n53357_ = ~new_n53348_ & ~new_n53356_;
  assign new_n53358_ = ~new_n53345_ & ~new_n53357_;
  assign new_n53359_ = new_n53232_ & ~new_n53314_;
  assign new_n53360_ = ~new_n53314_ & ~new_n53359_;
  assign new_n53361_ = new_n53330_ & ~new_n53360_;
  assign new_n53362_ = ~new_n53331_ & ~new_n53361_;
  assign new_n53363_ = new_n53345_ & ~new_n53362_;
  assign new_n53364_ = ~new_n53358_ & ~new_n53363_;
  assign new_n53365_ = ~new_n53261_ & new_n53364_;
  assign new_n53366_ = new_n53261_ & ~new_n53364_;
  assign ys__n39400 = new_n53365_ | new_n53366_;
  assign new_n53368_ = ~new_n53330_ & new_n53347_;
  assign new_n53369_ = ~new_n53315_ & ~new_n53359_;
  assign new_n53370_ = new_n53330_ & ~new_n53369_;
  assign new_n53371_ = ~new_n53368_ & ~new_n53370_;
  assign new_n53372_ = ~new_n53345_ & ~new_n53371_;
  assign new_n53373_ = ~new_n53347_ & ~new_n53355_;
  assign new_n53374_ = ~new_n53330_ & ~new_n53373_;
  assign new_n53375_ = ~new_n53316_ & new_n53330_;
  assign new_n53376_ = ~new_n53374_ & ~new_n53375_;
  assign new_n53377_ = new_n53345_ & ~new_n53376_;
  assign new_n53378_ = ~new_n53372_ & ~new_n53377_;
  assign new_n53379_ = ~new_n53261_ & new_n53378_;
  assign new_n53380_ = new_n53261_ & ~new_n53378_;
  assign ys__n39401 = new_n53379_ | new_n53380_;
  assign new_n53382_ = new_n53330_ & ~new_n53345_;
  assign new_n53383_ = new_n53355_ & new_n53382_;
  assign new_n53384_ = ~new_n53330_ & ~new_n53360_;
  assign new_n53385_ = ~new_n53330_ & ~new_n53384_;
  assign new_n53386_ = new_n53345_ & ~new_n53385_;
  assign new_n53387_ = ~new_n53383_ & ~new_n53386_;
  assign new_n53388_ = ~new_n53261_ & new_n53387_;
  assign new_n53389_ = new_n53261_ & ~new_n53387_;
  assign ys__n39402 = new_n53388_ | new_n53389_;
  assign new_n53391_ = ys__n48265 & new_n53181_;
  assign new_n53392_ = ys__n48265 & new_n53175_;
  assign ys__n44974 = ys__n352 & ys__n27867;
  assign new_n53394_ = new_n53176_ & ys__n44974;
  assign new_n53395_ = ~new_n53392_ & ~new_n53394_;
  assign new_n53396_ = ~new_n53391_ & new_n53395_;
  assign new_n53397_ = new_n53179_ & ys__n44974;
  assign new_n53398_ = ys__n48265 & new_n53174_;
  assign ys__n44958 = ys__n352 & ys__n28021;
  assign new_n53400_ = new_n53182_ & ys__n44958;
  assign new_n53401_ = ~new_n53398_ & ~new_n53400_;
  assign new_n53402_ = ~new_n53397_ & new_n53401_;
  assign new_n53403_ = new_n53396_ & new_n53402_;
  assign new_n53404_ = ~new_n53185_ & ~new_n53403_;
  assign new_n53405_ = ~new_n53345_ & new_n53404_;
  assign new_n53406_ = new_n53404_ & ~new_n53405_;
  assign new_n53407_ = ys__n48266 & new_n53181_;
  assign new_n53408_ = ys__n48266 & new_n53175_;
  assign ys__n44975 = ys__n352 & ys__n27869;
  assign new_n53410_ = new_n53176_ & ys__n44975;
  assign new_n53411_ = ~new_n53408_ & ~new_n53410_;
  assign new_n53412_ = ~new_n53407_ & new_n53411_;
  assign new_n53413_ = new_n53179_ & ys__n44975;
  assign new_n53414_ = ys__n48266 & new_n53174_;
  assign ys__n44959 = ys__n352 & ys__n28022;
  assign new_n53416_ = new_n53182_ & ys__n44959;
  assign new_n53417_ = ~new_n53414_ & ~new_n53416_;
  assign new_n53418_ = ~new_n53413_ & new_n53417_;
  assign new_n53419_ = new_n53412_ & new_n53418_;
  assign new_n53420_ = ~new_n53185_ & ~new_n53419_;
  assign new_n53421_ = ~new_n53406_ & ~new_n53420_;
  assign new_n53422_ = ys__n48267 & new_n53181_;
  assign new_n53423_ = ys__n48267 & new_n53175_;
  assign ys__n44976 = ys__n352 & ys__n27871;
  assign new_n53425_ = new_n53176_ & ys__n44976;
  assign new_n53426_ = ~new_n53423_ & ~new_n53425_;
  assign new_n53427_ = ~new_n53422_ & new_n53426_;
  assign new_n53428_ = new_n53179_ & ys__n44976;
  assign new_n53429_ = ys__n48267 & new_n53174_;
  assign ys__n44960 = ys__n352 & ys__n28023;
  assign new_n53431_ = new_n53182_ & ys__n44960;
  assign new_n53432_ = ~new_n53429_ & ~new_n53431_;
  assign new_n53433_ = ~new_n53428_ & new_n53432_;
  assign new_n53434_ = new_n53427_ & new_n53433_;
  assign new_n53435_ = ~new_n53185_ & ~new_n53434_;
  assign new_n53436_ = new_n53421_ & ~new_n53435_;
  assign new_n53437_ = ~new_n53345_ & ~new_n53404_;
  assign new_n53438_ = new_n53420_ & new_n53437_;
  assign new_n53439_ = new_n53420_ & ~new_n53438_;
  assign new_n53440_ = new_n53435_ & ~new_n53439_;
  assign new_n53441_ = ~new_n53436_ & ~new_n53440_;
  assign new_n53442_ = ~new_n53261_ & new_n53441_;
  assign new_n53443_ = new_n53261_ & ~new_n53441_;
  assign ys__n39403 = new_n53442_ | new_n53443_;
  assign new_n53445_ = new_n53345_ & new_n53404_;
  assign new_n53446_ = ~new_n53420_ & new_n53445_;
  assign new_n53447_ = ~new_n53438_ & ~new_n53446_;
  assign new_n53448_ = ~new_n53435_ & ~new_n53447_;
  assign new_n53449_ = new_n53345_ & ~new_n53404_;
  assign new_n53450_ = ~new_n53404_ & ~new_n53449_;
  assign new_n53451_ = new_n53420_ & ~new_n53450_;
  assign new_n53452_ = ~new_n53421_ & ~new_n53451_;
  assign new_n53453_ = new_n53435_ & ~new_n53452_;
  assign new_n53454_ = ~new_n53448_ & ~new_n53453_;
  assign new_n53455_ = ~new_n53261_ & new_n53454_;
  assign new_n53456_ = new_n53261_ & ~new_n53454_;
  assign ys__n39404 = new_n53455_ | new_n53456_;
  assign new_n53458_ = ~new_n53420_ & new_n53437_;
  assign new_n53459_ = ~new_n53405_ & ~new_n53449_;
  assign new_n53460_ = new_n53420_ & ~new_n53459_;
  assign new_n53461_ = ~new_n53458_ & ~new_n53460_;
  assign new_n53462_ = ~new_n53435_ & ~new_n53461_;
  assign new_n53463_ = ~new_n53437_ & ~new_n53445_;
  assign new_n53464_ = ~new_n53420_ & ~new_n53463_;
  assign new_n53465_ = ~new_n53406_ & new_n53420_;
  assign new_n53466_ = ~new_n53464_ & ~new_n53465_;
  assign new_n53467_ = new_n53435_ & ~new_n53466_;
  assign new_n53468_ = ~new_n53462_ & ~new_n53467_;
  assign new_n53469_ = ~new_n53261_ & new_n53468_;
  assign new_n53470_ = new_n53261_ & ~new_n53468_;
  assign ys__n39405 = new_n53469_ | new_n53470_;
  assign new_n53472_ = new_n53420_ & ~new_n53435_;
  assign new_n53473_ = new_n53445_ & new_n53472_;
  assign new_n53474_ = ~new_n53420_ & ~new_n53450_;
  assign new_n53475_ = ~new_n53420_ & ~new_n53474_;
  assign new_n53476_ = new_n53435_ & ~new_n53475_;
  assign new_n53477_ = ~new_n53473_ & ~new_n53476_;
  assign new_n53478_ = ~new_n53261_ & new_n53477_;
  assign new_n53479_ = new_n53261_ & ~new_n53477_;
  assign ys__n39406 = new_n53478_ | new_n53479_;
  assign new_n53481_ = ys__n48268 & new_n53181_;
  assign new_n53482_ = ys__n48268 & new_n53175_;
  assign ys__n44977 = ys__n352 & ys__n27873;
  assign new_n53484_ = new_n53176_ & ys__n44977;
  assign new_n53485_ = ~new_n53482_ & ~new_n53484_;
  assign new_n53486_ = ~new_n53481_ & new_n53485_;
  assign new_n53487_ = new_n53179_ & ys__n44977;
  assign new_n53488_ = ys__n48268 & new_n53174_;
  assign ys__n44961 = ys__n352 & ys__n28024;
  assign new_n53490_ = new_n53182_ & ys__n44961;
  assign new_n53491_ = ~new_n53488_ & ~new_n53490_;
  assign new_n53492_ = ~new_n53487_ & new_n53491_;
  assign new_n53493_ = new_n53486_ & new_n53492_;
  assign new_n53494_ = ~new_n53185_ & ~new_n53493_;
  assign new_n53495_ = ~new_n53435_ & new_n53494_;
  assign new_n53496_ = new_n53494_ & ~new_n53495_;
  assign new_n53497_ = ys__n48269 & new_n53181_;
  assign new_n53498_ = ys__n48269 & new_n53175_;
  assign ys__n44978 = ys__n352 & ys__n27875;
  assign new_n53500_ = new_n53176_ & ys__n44978;
  assign new_n53501_ = ~new_n53498_ & ~new_n53500_;
  assign new_n53502_ = ~new_n53497_ & new_n53501_;
  assign new_n53503_ = new_n53179_ & ys__n44978;
  assign new_n53504_ = ys__n48269 & new_n53174_;
  assign ys__n44962 = ys__n352 & ys__n28025;
  assign new_n53506_ = new_n53182_ & ys__n44962;
  assign new_n53507_ = ~new_n53504_ & ~new_n53506_;
  assign new_n53508_ = ~new_n53503_ & new_n53507_;
  assign new_n53509_ = new_n53502_ & new_n53508_;
  assign new_n53510_ = ~new_n53185_ & ~new_n53509_;
  assign new_n53511_ = ~new_n53496_ & ~new_n53510_;
  assign new_n53512_ = ys__n48270 & new_n53181_;
  assign new_n53513_ = ys__n48270 & new_n53175_;
  assign ys__n44979 = ys__n352 & ys__n27877;
  assign new_n53515_ = new_n53176_ & ys__n44979;
  assign new_n53516_ = ~new_n53513_ & ~new_n53515_;
  assign new_n53517_ = ~new_n53512_ & new_n53516_;
  assign new_n53518_ = new_n53179_ & ys__n44979;
  assign new_n53519_ = ys__n48270 & new_n53174_;
  assign ys__n44963 = ys__n352 & ys__n28026;
  assign new_n53521_ = new_n53182_ & ys__n44963;
  assign new_n53522_ = ~new_n53519_ & ~new_n53521_;
  assign new_n53523_ = ~new_n53518_ & new_n53522_;
  assign new_n53524_ = new_n53517_ & new_n53523_;
  assign new_n53525_ = ~new_n53185_ & ~new_n53524_;
  assign new_n53526_ = new_n53511_ & ~new_n53525_;
  assign new_n53527_ = ~new_n53435_ & ~new_n53494_;
  assign new_n53528_ = new_n53510_ & new_n53527_;
  assign new_n53529_ = new_n53510_ & ~new_n53528_;
  assign new_n53530_ = new_n53525_ & ~new_n53529_;
  assign new_n53531_ = ~new_n53526_ & ~new_n53530_;
  assign new_n53532_ = ~new_n53261_ & new_n53531_;
  assign new_n53533_ = new_n53261_ & ~new_n53531_;
  assign ys__n39407 = new_n53532_ | new_n53533_;
  assign new_n53535_ = new_n53435_ & new_n53494_;
  assign new_n53536_ = ~new_n53510_ & new_n53535_;
  assign new_n53537_ = ~new_n53528_ & ~new_n53536_;
  assign new_n53538_ = ~new_n53525_ & ~new_n53537_;
  assign new_n53539_ = new_n53435_ & ~new_n53494_;
  assign new_n53540_ = ~new_n53494_ & ~new_n53539_;
  assign new_n53541_ = new_n53510_ & ~new_n53540_;
  assign new_n53542_ = ~new_n53511_ & ~new_n53541_;
  assign new_n53543_ = new_n53525_ & ~new_n53542_;
  assign new_n53544_ = ~new_n53538_ & ~new_n53543_;
  assign new_n53545_ = ~new_n53261_ & new_n53544_;
  assign new_n53546_ = new_n53261_ & ~new_n53544_;
  assign ys__n39408 = new_n53545_ | new_n53546_;
  assign new_n53548_ = ~new_n53510_ & new_n53527_;
  assign new_n53549_ = ~new_n53495_ & ~new_n53539_;
  assign new_n53550_ = new_n53510_ & ~new_n53549_;
  assign new_n53551_ = ~new_n53548_ & ~new_n53550_;
  assign new_n53552_ = ~new_n53525_ & ~new_n53551_;
  assign new_n53553_ = ~new_n53527_ & ~new_n53535_;
  assign new_n53554_ = ~new_n53510_ & ~new_n53553_;
  assign new_n53555_ = ~new_n53496_ & new_n53510_;
  assign new_n53556_ = ~new_n53554_ & ~new_n53555_;
  assign new_n53557_ = new_n53525_ & ~new_n53556_;
  assign new_n53558_ = ~new_n53552_ & ~new_n53557_;
  assign new_n53559_ = ~new_n53261_ & new_n53558_;
  assign new_n53560_ = new_n53261_ & ~new_n53558_;
  assign ys__n39409 = new_n53559_ | new_n53560_;
  assign new_n53562_ = new_n53510_ & ~new_n53525_;
  assign new_n53563_ = new_n53535_ & new_n53562_;
  assign new_n53564_ = ~new_n53510_ & ~new_n53540_;
  assign new_n53565_ = ~new_n53510_ & ~new_n53564_;
  assign new_n53566_ = new_n53525_ & ~new_n53565_;
  assign new_n53567_ = ~new_n53563_ & ~new_n53566_;
  assign new_n53568_ = ~new_n53261_ & new_n53567_;
  assign new_n53569_ = new_n53261_ & ~new_n53567_;
  assign ys__n39410 = new_n53568_ | new_n53569_;
  assign new_n53571_ = ys__n48271 & new_n53181_;
  assign new_n53572_ = ys__n48271 & new_n53175_;
  assign ys__n44980 = ys__n352 & ys__n27879;
  assign new_n53574_ = new_n53176_ & ys__n44980;
  assign new_n53575_ = ~new_n53572_ & ~new_n53574_;
  assign new_n53576_ = ~new_n53571_ & new_n53575_;
  assign new_n53577_ = new_n53179_ & ys__n44980;
  assign new_n53578_ = ys__n48271 & new_n53174_;
  assign ys__n44964 = ys__n352 & ys__n28027;
  assign new_n53580_ = new_n53182_ & ys__n44964;
  assign new_n53581_ = ~new_n53578_ & ~new_n53580_;
  assign new_n53582_ = ~new_n53577_ & new_n53581_;
  assign new_n53583_ = new_n53576_ & new_n53582_;
  assign new_n53584_ = ~new_n53185_ & ~new_n53583_;
  assign new_n53585_ = ~new_n53525_ & new_n53584_;
  assign new_n53586_ = new_n53584_ & ~new_n53585_;
  assign new_n53587_ = ys__n48272 & new_n53181_;
  assign new_n53588_ = ys__n48272 & new_n53175_;
  assign ys__n44981 = ys__n352 & ys__n27881;
  assign new_n53590_ = new_n53176_ & ys__n44981;
  assign new_n53591_ = ~new_n53588_ & ~new_n53590_;
  assign new_n53592_ = ~new_n53587_ & new_n53591_;
  assign new_n53593_ = new_n53179_ & ys__n44981;
  assign new_n53594_ = ys__n48272 & new_n53174_;
  assign ys__n44965 = ys__n352 & ys__n28028;
  assign new_n53596_ = new_n53182_ & ys__n44965;
  assign new_n53597_ = ~new_n53594_ & ~new_n53596_;
  assign new_n53598_ = ~new_n53593_ & new_n53597_;
  assign new_n53599_ = new_n53592_ & new_n53598_;
  assign new_n53600_ = ~new_n53185_ & ~new_n53599_;
  assign new_n53601_ = ~new_n53586_ & ~new_n53600_;
  assign new_n53602_ = ys__n48273 & new_n53181_;
  assign new_n53603_ = ys__n48273 & new_n53175_;
  assign ys__n44982 = ys__n352 & ys__n27883;
  assign new_n53605_ = new_n53176_ & ys__n44982;
  assign new_n53606_ = ~new_n53603_ & ~new_n53605_;
  assign new_n53607_ = ~new_n53602_ & new_n53606_;
  assign new_n53608_ = new_n53179_ & ys__n44982;
  assign new_n53609_ = ys__n48273 & new_n53174_;
  assign ys__n44966 = ys__n352 & ys__n28029;
  assign new_n53611_ = new_n53182_ & ys__n44966;
  assign new_n53612_ = ~new_n53609_ & ~new_n53611_;
  assign new_n53613_ = ~new_n53608_ & new_n53612_;
  assign new_n53614_ = new_n53607_ & new_n53613_;
  assign new_n53615_ = ~new_n53185_ & ~new_n53614_;
  assign new_n53616_ = new_n53601_ & ~new_n53615_;
  assign new_n53617_ = ~new_n53525_ & ~new_n53584_;
  assign new_n53618_ = new_n53600_ & new_n53617_;
  assign new_n53619_ = new_n53600_ & ~new_n53618_;
  assign new_n53620_ = new_n53615_ & ~new_n53619_;
  assign new_n53621_ = ~new_n53616_ & ~new_n53620_;
  assign new_n53622_ = ~new_n53261_ & new_n53621_;
  assign new_n53623_ = new_n53261_ & ~new_n53621_;
  assign ys__n39411 = new_n53622_ | new_n53623_;
  assign new_n53625_ = new_n53525_ & new_n53584_;
  assign new_n53626_ = ~new_n53600_ & new_n53625_;
  assign new_n53627_ = ~new_n53618_ & ~new_n53626_;
  assign new_n53628_ = ~new_n53615_ & ~new_n53627_;
  assign new_n53629_ = new_n53525_ & ~new_n53584_;
  assign new_n53630_ = ~new_n53584_ & ~new_n53629_;
  assign new_n53631_ = new_n53600_ & ~new_n53630_;
  assign new_n53632_ = ~new_n53601_ & ~new_n53631_;
  assign new_n53633_ = new_n53615_ & ~new_n53632_;
  assign new_n53634_ = ~new_n53628_ & ~new_n53633_;
  assign new_n53635_ = ~new_n53261_ & new_n53634_;
  assign new_n53636_ = new_n53261_ & ~new_n53634_;
  assign ys__n39412 = new_n53635_ | new_n53636_;
  assign new_n53638_ = ~new_n53600_ & new_n53617_;
  assign new_n53639_ = ~new_n53585_ & ~new_n53629_;
  assign new_n53640_ = new_n53600_ & ~new_n53639_;
  assign new_n53641_ = ~new_n53638_ & ~new_n53640_;
  assign new_n53642_ = ~new_n53615_ & ~new_n53641_;
  assign new_n53643_ = ~new_n53617_ & ~new_n53625_;
  assign new_n53644_ = ~new_n53600_ & ~new_n53643_;
  assign new_n53645_ = ~new_n53586_ & new_n53600_;
  assign new_n53646_ = ~new_n53644_ & ~new_n53645_;
  assign new_n53647_ = new_n53615_ & ~new_n53646_;
  assign new_n53648_ = ~new_n53642_ & ~new_n53647_;
  assign new_n53649_ = ~new_n53261_ & new_n53648_;
  assign new_n53650_ = new_n53261_ & ~new_n53648_;
  assign ys__n39413 = new_n53649_ | new_n53650_;
  assign new_n53652_ = new_n53600_ & ~new_n53615_;
  assign new_n53653_ = new_n53625_ & new_n53652_;
  assign new_n53654_ = ~new_n53600_ & ~new_n53630_;
  assign new_n53655_ = ~new_n53600_ & ~new_n53654_;
  assign new_n53656_ = new_n53615_ & ~new_n53655_;
  assign new_n53657_ = ~new_n53653_ & ~new_n53656_;
  assign new_n53658_ = ~new_n53261_ & new_n53657_;
  assign new_n53659_ = new_n53261_ & ~new_n53657_;
  assign ys__n39414 = new_n53658_ | new_n53659_;
  assign ys__n44983 = ys__n352 & ys__n27885;
  assign new_n53662_ = new_n53176_ & ys__n44983;
  assign new_n53663_ = ys__n48274 & new_n53181_;
  assign new_n53664_ = ys__n48274 & new_n53174_;
  assign new_n53665_ = ~new_n53663_ & ~new_n53664_;
  assign new_n53666_ = ~new_n53662_ & new_n53665_;
  assign new_n53667_ = ~new_n53185_ & ~new_n53666_;
  assign new_n53668_ = new_n53179_ & ys__n44983;
  assign ys__n44967 = ys__n352 & ys__n28030;
  assign new_n53670_ = new_n53182_ & ys__n44967;
  assign new_n53671_ = ys__n48274 & new_n53175_;
  assign new_n53672_ = ~new_n53662_ & ~new_n53671_;
  assign new_n53673_ = ~new_n53670_ & new_n53672_;
  assign new_n53674_ = ~new_n53668_ & new_n53673_;
  assign new_n53675_ = new_n53665_ & new_n53674_;
  assign new_n53676_ = ~new_n53185_ & ~new_n53675_;
  assign new_n53677_ = ~new_n53615_ & new_n53676_;
  assign new_n53678_ = new_n53676_ & ~new_n53677_;
  assign new_n53679_ = ~new_n53667_ & ~new_n53678_;
  assign new_n53680_ = ~new_n53667_ & new_n53679_;
  assign new_n53681_ = ~new_n53615_ & ~new_n53676_;
  assign new_n53682_ = new_n53667_ & new_n53681_;
  assign new_n53683_ = new_n53667_ & ~new_n53682_;
  assign new_n53684_ = new_n53667_ & ~new_n53683_;
  assign new_n53685_ = ~new_n53680_ & ~new_n53684_;
  assign new_n53686_ = ~new_n53261_ & new_n53685_;
  assign new_n53687_ = new_n53261_ & ~new_n53685_;
  assign ys__n39415 = new_n53686_ | new_n53687_;
  assign new_n53689_ = new_n53615_ & new_n53676_;
  assign new_n53690_ = ~new_n53667_ & new_n53689_;
  assign new_n53691_ = ~new_n53682_ & ~new_n53690_;
  assign new_n53692_ = ~new_n53667_ & ~new_n53691_;
  assign new_n53693_ = new_n53615_ & ~new_n53676_;
  assign new_n53694_ = ~new_n53676_ & ~new_n53693_;
  assign new_n53695_ = new_n53667_ & ~new_n53694_;
  assign new_n53696_ = ~new_n53679_ & ~new_n53695_;
  assign new_n53697_ = new_n53667_ & ~new_n53696_;
  assign new_n53698_ = ~new_n53692_ & ~new_n53697_;
  assign new_n53699_ = ~new_n53261_ & new_n53698_;
  assign new_n53700_ = new_n53261_ & ~new_n53698_;
  assign ys__n39416 = new_n53699_ | new_n53700_;
  assign new_n53702_ = ~new_n53667_ & new_n53681_;
  assign new_n53703_ = ~new_n53677_ & ~new_n53693_;
  assign new_n53704_ = new_n53667_ & ~new_n53703_;
  assign new_n53705_ = ~new_n53702_ & ~new_n53704_;
  assign new_n53706_ = ~new_n53667_ & ~new_n53705_;
  assign new_n53707_ = ~new_n53681_ & ~new_n53689_;
  assign new_n53708_ = ~new_n53667_ & ~new_n53707_;
  assign new_n53709_ = new_n53667_ & ~new_n53678_;
  assign new_n53710_ = ~new_n53708_ & ~new_n53709_;
  assign new_n53711_ = new_n53667_ & ~new_n53710_;
  assign new_n53712_ = ~new_n53706_ & ~new_n53711_;
  assign new_n53713_ = ~new_n53261_ & new_n53712_;
  assign new_n53714_ = new_n53261_ & ~new_n53712_;
  assign ys__n39417 = new_n53713_ | new_n53714_;
  assign new_n53716_ = ~new_n53667_ & ~new_n53694_;
  assign new_n53717_ = ~new_n53667_ & ~new_n53716_;
  assign new_n53718_ = new_n53667_ & ~new_n53717_;
  assign new_n53719_ = ~new_n53261_ & ~new_n53718_;
  assign new_n53720_ = new_n53261_ & new_n53718_;
  assign ys__n39418 = new_n53719_ | new_n53720_;
  assign new_n53722_ = ys__n33634 & ys__n33636;
  assign new_n53723_ = ys__n33632 & new_n53722_;
  assign new_n53724_ = ys__n39718 & new_n53723_;
  assign new_n53725_ = ys__n33632 & ys__n33636;
  assign new_n53726_ = ys__n33638 & new_n53725_;
  assign new_n53727_ = ys__n24741 & new_n53726_;
  assign new_n53728_ = ~new_n53724_ & ~new_n53727_;
  assign new_n53729_ = ~ys__n33632 & ~ys__n33634;
  assign new_n53730_ = ~ys__n33638 & new_n53729_;
  assign new_n53731_ = ys__n33683 & new_n53730_;
  assign new_n53732_ = ys__n33632 & ys__n33634;
  assign new_n53733_ = ys__n33638 & new_n53732_;
  assign new_n53734_ = ~ys__n33683 & new_n53733_;
  assign new_n53735_ = ~new_n53731_ & ~new_n53734_;
  assign new_n53736_ = new_n53728_ & new_n53735_;
  assign new_n53737_ = ~ys__n33634 & ~ys__n33636;
  assign new_n53738_ = ~ys__n33638 & new_n53737_;
  assign new_n53739_ = ys__n24747 & new_n53738_;
  assign new_n53740_ = ~ys__n33632 & new_n53737_;
  assign new_n53741_ = ys__n24744 & new_n53740_;
  assign new_n53742_ = ~new_n53739_ & ~new_n53741_;
  assign new_n53743_ = ~ys__n33632 & ~ys__n33636;
  assign new_n53744_ = ~ys__n33638 & new_n53743_;
  assign new_n53745_ = ys__n24741 & new_n53744_;
  assign new_n53746_ = ys__n33638 & new_n53722_;
  assign new_n53747_ = ys__n39720 & new_n53746_;
  assign new_n53748_ = ~new_n53745_ & ~new_n53747_;
  assign new_n53749_ = new_n53742_ & new_n53748_;
  assign ys__n40052 = ~new_n53736_ | ~new_n53749_;
  assign ys__n42129 = new_n26586_ & new_n26624_;
  assign new_n53752_ = ys__n33658 & ys__n33660;
  assign new_n53753_ = ys__n33662 & new_n53752_;
  assign new_n53754_ = ys__n33656 & ys__n33660;
  assign new_n53755_ = ys__n33662 & new_n53754_;
  assign new_n53756_ = ys__n33656 & new_n53752_;
  assign new_n53757_ = ~new_n53755_ & ~new_n53756_;
  assign new_n53758_ = ~new_n53753_ & new_n53757_;
  assign new_n53759_ = ys__n39520 & ~new_n53758_;
  assign new_n53760_ = ~ys__n33658 & ~ys__n33660;
  assign new_n53761_ = ~ys__n33662 & new_n53760_;
  assign new_n53762_ = ~ys__n33656 & ~ys__n33660;
  assign new_n53763_ = ~ys__n33662 & new_n53762_;
  assign new_n53764_ = ~ys__n33656 & new_n53760_;
  assign new_n53765_ = ~new_n53763_ & ~new_n53764_;
  assign new_n53766_ = ~new_n53761_ & new_n53765_;
  assign new_n53767_ = ys__n39518 & ~new_n53766_;
  assign new_n53768_ = ~ys__n33656 & ~ys__n33658;
  assign new_n53769_ = ~ys__n33662 & new_n53768_;
  assign new_n53770_ = ys__n33747 & new_n53769_;
  assign new_n53771_ = ys__n33656 & ys__n33658;
  assign new_n53772_ = ys__n33662 & new_n53771_;
  assign new_n53773_ = ~ys__n33747 & new_n53772_;
  assign new_n53774_ = ~new_n53770_ & ~new_n53773_;
  assign new_n53775_ = ~new_n53767_ & new_n53774_;
  assign new_n53776_ = ~new_n53759_ & new_n53775_;
  assign new_n53777_ = ys__n33666 & ys__n33668;
  assign new_n53778_ = ys__n33670 & new_n53777_;
  assign new_n53779_ = ys__n33664 & ys__n33668;
  assign new_n53780_ = ys__n33670 & new_n53779_;
  assign new_n53781_ = ys__n33664 & new_n53777_;
  assign new_n53782_ = ~new_n53780_ & ~new_n53781_;
  assign new_n53783_ = ~new_n53778_ & new_n53782_;
  assign new_n53784_ = ys__n39520 & ~new_n53783_;
  assign new_n53785_ = ~ys__n33666 & ~ys__n33668;
  assign new_n53786_ = ~ys__n33670 & new_n53785_;
  assign new_n53787_ = ~ys__n33664 & ~ys__n33668;
  assign new_n53788_ = ~ys__n33670 & new_n53787_;
  assign new_n53789_ = ~ys__n33664 & new_n53785_;
  assign new_n53790_ = ~new_n53788_ & ~new_n53789_;
  assign new_n53791_ = ~new_n53786_ & new_n53790_;
  assign new_n53792_ = ys__n39518 & ~new_n53791_;
  assign new_n53793_ = ~ys__n33664 & ~ys__n33666;
  assign new_n53794_ = ~ys__n33670 & new_n53793_;
  assign new_n53795_ = ys__n33747 & new_n53794_;
  assign new_n53796_ = ys__n33664 & ys__n33666;
  assign new_n53797_ = ys__n33670 & new_n53796_;
  assign new_n53798_ = ~ys__n33747 & new_n53797_;
  assign new_n53799_ = ~new_n53795_ & ~new_n53798_;
  assign new_n53800_ = ~new_n53792_ & new_n53799_;
  assign new_n53801_ = ~new_n53784_ & new_n53800_;
  assign new_n53802_ = ~ys__n33672 & ~ys__n33676;
  assign new_n53803_ = ~ys__n33678 & new_n53802_;
  assign new_n53804_ = ~ys__n33674 & ~ys__n33676;
  assign new_n53805_ = ~ys__n33678 & new_n53804_;
  assign new_n53806_ = ~ys__n33672 & new_n53804_;
  assign new_n53807_ = ~new_n53805_ & ~new_n53806_;
  assign new_n53808_ = ~new_n53803_ & new_n53807_;
  assign new_n53809_ = ys__n39518 & ~new_n53808_;
  assign new_n53810_ = ys__n33672 & ys__n33676;
  assign new_n53811_ = ys__n33678 & new_n53810_;
  assign new_n53812_ = ys__n33674 & ys__n33676;
  assign new_n53813_ = ys__n33678 & new_n53812_;
  assign new_n53814_ = ys__n33672 & new_n53812_;
  assign new_n53815_ = ~new_n53813_ & ~new_n53814_;
  assign new_n53816_ = ~new_n53811_ & new_n53815_;
  assign new_n53817_ = ys__n39520 & ~new_n53816_;
  assign new_n53818_ = ~new_n53809_ & ~new_n53817_;
  assign new_n53819_ = ~new_n53801_ & ~new_n53818_;
  assign new_n53820_ = ~new_n53776_ & new_n53819_;
  assign new_n53821_ = new_n53801_ & new_n53818_;
  assign new_n53822_ = ~new_n53776_ & new_n53821_;
  assign new_n53823_ = ~new_n53820_ & ~new_n53822_;
  assign new_n53824_ = ~new_n53801_ & new_n53818_;
  assign new_n53825_ = new_n53776_ & new_n53824_;
  assign new_n53826_ = new_n53801_ & ~new_n53818_;
  assign new_n53827_ = new_n53776_ & new_n53826_;
  assign new_n53828_ = ~new_n53825_ & ~new_n53827_;
  assign new_n53829_ = new_n53823_ & new_n53828_;
  assign new_n53830_ = ys__n33642 & ys__n33644;
  assign new_n53831_ = ys__n33646 & new_n53830_;
  assign new_n53832_ = ys__n33640 & ys__n33644;
  assign new_n53833_ = ys__n33646 & new_n53832_;
  assign new_n53834_ = ys__n33640 & new_n53830_;
  assign new_n53835_ = ~new_n53833_ & ~new_n53834_;
  assign new_n53836_ = ~new_n53831_ & new_n53835_;
  assign new_n53837_ = ys__n39520 & ~new_n53836_;
  assign new_n53838_ = ~ys__n33642 & ~ys__n33644;
  assign new_n53839_ = ~ys__n33646 & new_n53838_;
  assign new_n53840_ = ~ys__n33640 & ~ys__n33644;
  assign new_n53841_ = ~ys__n33646 & new_n53840_;
  assign new_n53842_ = ~ys__n33640 & new_n53838_;
  assign new_n53843_ = ~new_n53841_ & ~new_n53842_;
  assign new_n53844_ = ~new_n53839_ & new_n53843_;
  assign new_n53845_ = ys__n39518 & ~new_n53844_;
  assign new_n53846_ = ~ys__n33640 & ~ys__n33642;
  assign new_n53847_ = ~ys__n33646 & new_n53846_;
  assign new_n53848_ = ys__n33747 & new_n53847_;
  assign new_n53849_ = ys__n33640 & ys__n33642;
  assign new_n53850_ = ys__n33646 & new_n53849_;
  assign new_n53851_ = ~ys__n33747 & new_n53850_;
  assign new_n53852_ = ~new_n53848_ & ~new_n53851_;
  assign new_n53853_ = ~new_n53845_ & new_n53852_;
  assign new_n53854_ = ~new_n53837_ & new_n53853_;
  assign new_n53855_ = ~new_n53723_ & ~new_n53746_;
  assign new_n53856_ = ~new_n53726_ & new_n53855_;
  assign new_n53857_ = ys__n39520 & ~new_n53856_;
  assign new_n53858_ = ~new_n53738_ & ~new_n53740_;
  assign new_n53859_ = ~new_n53744_ & new_n53858_;
  assign new_n53860_ = ys__n39518 & ~new_n53859_;
  assign new_n53861_ = ys__n33747 & new_n53730_;
  assign new_n53862_ = ~ys__n33747 & new_n53733_;
  assign new_n53863_ = ~new_n53861_ & ~new_n53862_;
  assign new_n53864_ = ~new_n53860_ & new_n53863_;
  assign new_n53865_ = ~new_n53857_ & new_n53864_;
  assign new_n53866_ = ~new_n53854_ & ~new_n53865_;
  assign new_n53867_ = ys__n33650 & ys__n33652;
  assign new_n53868_ = ys__n33654 & new_n53867_;
  assign new_n53869_ = ys__n33648 & ys__n33652;
  assign new_n53870_ = ys__n33654 & new_n53869_;
  assign new_n53871_ = ys__n33648 & new_n53867_;
  assign new_n53872_ = ~new_n53870_ & ~new_n53871_;
  assign new_n53873_ = ~new_n53868_ & new_n53872_;
  assign new_n53874_ = ys__n39520 & ~new_n53873_;
  assign new_n53875_ = ~ys__n33650 & ~ys__n33652;
  assign new_n53876_ = ~ys__n33654 & new_n53875_;
  assign new_n53877_ = ~ys__n33648 & ~ys__n33652;
  assign new_n53878_ = ~ys__n33654 & new_n53877_;
  assign new_n53879_ = ~ys__n33648 & new_n53875_;
  assign new_n53880_ = ~new_n53878_ & ~new_n53879_;
  assign new_n53881_ = ~new_n53876_ & new_n53880_;
  assign new_n53882_ = ys__n39518 & ~new_n53881_;
  assign new_n53883_ = ~ys__n33648 & ~ys__n33650;
  assign new_n53884_ = ~ys__n33654 & new_n53883_;
  assign new_n53885_ = ys__n33747 & new_n53884_;
  assign new_n53886_ = ys__n33648 & ys__n33650;
  assign new_n53887_ = ys__n33654 & new_n53886_;
  assign new_n53888_ = ~ys__n33747 & new_n53887_;
  assign new_n53889_ = ~new_n53885_ & ~new_n53888_;
  assign new_n53890_ = ~new_n53882_ & new_n53889_;
  assign new_n53891_ = ~new_n53874_ & new_n53890_;
  assign new_n53892_ = ~new_n53854_ & ~new_n53891_;
  assign new_n53893_ = ~new_n53865_ & ~new_n53891_;
  assign new_n53894_ = ~new_n53892_ & ~new_n53893_;
  assign new_n53895_ = ~new_n53866_ & new_n53894_;
  assign new_n53896_ = ys__n39518 & new_n53805_;
  assign new_n53897_ = ys__n39520 & new_n53813_;
  assign new_n53898_ = ~new_n53896_ & ~new_n53897_;
  assign new_n53899_ = ys__n39518 & new_n53806_;
  assign new_n53900_ = ys__n39520 & new_n53814_;
  assign new_n53901_ = ~new_n53899_ & ~new_n53900_;
  assign new_n53902_ = new_n53898_ & new_n53901_;
  assign new_n53903_ = ~new_n53776_ & ~new_n53902_;
  assign new_n53904_ = ~new_n53776_ & ~new_n53801_;
  assign new_n53905_ = ~new_n53801_ & ~new_n53902_;
  assign new_n53906_ = ~new_n53904_ & ~new_n53905_;
  assign new_n53907_ = ~new_n53903_ & new_n53906_;
  assign new_n53908_ = ~new_n53895_ & ~new_n53907_;
  assign new_n53909_ = ~new_n53829_ & new_n53908_;
  assign new_n53910_ = ~new_n53895_ & new_n53907_;
  assign new_n53911_ = new_n53829_ & new_n53910_;
  assign new_n53912_ = ~new_n53909_ & ~new_n53911_;
  assign new_n53913_ = new_n53895_ & new_n53907_;
  assign new_n53914_ = ~new_n53829_ & new_n53913_;
  assign new_n53915_ = new_n53895_ & ~new_n53907_;
  assign new_n53916_ = new_n53829_ & new_n53915_;
  assign new_n53917_ = ~new_n53914_ & ~new_n53916_;
  assign new_n53918_ = new_n53912_ & new_n53917_;
  assign new_n53919_ = ~new_n53776_ & new_n53905_;
  assign new_n53920_ = new_n53801_ & new_n53902_;
  assign new_n53921_ = ~new_n53776_ & new_n53920_;
  assign new_n53922_ = ~new_n53919_ & ~new_n53921_;
  assign new_n53923_ = ~new_n53801_ & new_n53902_;
  assign new_n53924_ = new_n53776_ & new_n53923_;
  assign new_n53925_ = new_n53801_ & ~new_n53902_;
  assign new_n53926_ = new_n53776_ & new_n53925_;
  assign new_n53927_ = ~new_n53924_ & ~new_n53926_;
  assign new_n53928_ = new_n53922_ & new_n53927_;
  assign new_n53929_ = ~new_n53895_ & ~new_n53928_;
  assign new_n53930_ = ys__n24834 & new_n53806_;
  assign new_n53931_ = ~new_n53896_ & ~new_n53930_;
  assign new_n53932_ = ys__n39778 & new_n53814_;
  assign new_n53933_ = ~new_n53897_ & ~new_n53932_;
  assign new_n53934_ = new_n53931_ & new_n53933_;
  assign new_n53935_ = ~new_n53801_ & ~new_n53934_;
  assign new_n53936_ = ~new_n53776_ & ~new_n53934_;
  assign new_n53937_ = ~new_n53935_ & ~new_n53936_;
  assign new_n53938_ = ~new_n53904_ & new_n53937_;
  assign new_n53939_ = ~new_n53928_ & ~new_n53938_;
  assign new_n53940_ = ~new_n53895_ & ~new_n53938_;
  assign new_n53941_ = ~new_n53939_ & ~new_n53940_;
  assign new_n53942_ = ~new_n53929_ & new_n53941_;
  assign new_n53943_ = ~new_n53865_ & new_n53892_;
  assign new_n53944_ = new_n53854_ & new_n53891_;
  assign new_n53945_ = ~new_n53865_ & new_n53944_;
  assign new_n53946_ = ~new_n53943_ & ~new_n53945_;
  assign new_n53947_ = ~new_n53854_ & new_n53891_;
  assign new_n53948_ = new_n53865_ & new_n53947_;
  assign new_n53949_ = new_n53854_ & ~new_n53891_;
  assign new_n53950_ = new_n53865_ & new_n53949_;
  assign new_n53951_ = ~new_n53948_ & ~new_n53950_;
  assign new_n53952_ = new_n53946_ & new_n53951_;
  assign new_n53953_ = ~new_n53942_ & ~new_n53952_;
  assign new_n53954_ = ~new_n53918_ & new_n53953_;
  assign new_n53955_ = new_n53942_ & ~new_n53952_;
  assign new_n53956_ = new_n53918_ & new_n53955_;
  assign new_n53957_ = ~new_n53954_ & ~new_n53956_;
  assign new_n53958_ = new_n53942_ & new_n53952_;
  assign new_n53959_ = ~new_n53918_ & new_n53958_;
  assign new_n53960_ = ~new_n53942_ & new_n53952_;
  assign new_n53961_ = new_n53918_ & new_n53960_;
  assign new_n53962_ = ~new_n53959_ & ~new_n53961_;
  assign ys__n42153 = ~new_n53957_ | ~new_n53962_;
  assign new_n53964_ = ~new_n53895_ & new_n53939_;
  assign new_n53965_ = new_n53895_ & ~new_n53938_;
  assign new_n53966_ = new_n53928_ & new_n53965_;
  assign new_n53967_ = ~new_n53895_ & new_n53938_;
  assign new_n53968_ = new_n53928_ & new_n53967_;
  assign new_n53969_ = new_n53895_ & new_n53938_;
  assign new_n53970_ = ~new_n53928_ & new_n53969_;
  assign new_n53971_ = ~new_n53968_ & ~new_n53970_;
  assign new_n53972_ = ~new_n53966_ & new_n53971_;
  assign new_n53973_ = ~new_n53964_ & new_n53972_;
  assign new_n53974_ = ~new_n53952_ & ~new_n53973_;
  assign new_n53975_ = ~new_n53776_ & new_n53935_;
  assign new_n53976_ = new_n53801_ & new_n53934_;
  assign new_n53977_ = ~new_n53776_ & new_n53976_;
  assign new_n53978_ = ~new_n53975_ & ~new_n53977_;
  assign new_n53979_ = ~new_n53801_ & new_n53934_;
  assign new_n53980_ = new_n53776_ & new_n53979_;
  assign new_n53981_ = new_n53801_ & ~new_n53934_;
  assign new_n53982_ = new_n53776_ & new_n53981_;
  assign new_n53983_ = ~new_n53980_ & ~new_n53982_;
  assign new_n53984_ = new_n53978_ & new_n53983_;
  assign new_n53985_ = ~new_n53895_ & ~new_n53984_;
  assign new_n53986_ = ys__n39518 & new_n53788_;
  assign new_n53987_ = ys__n39520 & new_n53778_;
  assign new_n53988_ = ~new_n53986_ & ~new_n53987_;
  assign new_n53989_ = ys__n39520 & new_n53781_;
  assign new_n53990_ = ys__n39520 & new_n53780_;
  assign new_n53991_ = ~new_n53989_ & ~new_n53990_;
  assign new_n53992_ = new_n53988_ & new_n53991_;
  assign new_n53993_ = ys__n39518 & new_n53786_;
  assign new_n53994_ = ys__n39518 & new_n53789_;
  assign new_n53995_ = ~new_n53993_ & ~new_n53994_;
  assign new_n53996_ = new_n53799_ & new_n53995_;
  assign new_n53997_ = new_n53992_ & new_n53996_;
  assign new_n53998_ = ~new_n53776_ & ~new_n53997_;
  assign new_n53999_ = ys__n24834 & new_n53805_;
  assign new_n54000_ = ys__n24831 & new_n53806_;
  assign new_n54001_ = ~new_n53999_ & ~new_n54000_;
  assign new_n54002_ = ys__n39778 & new_n53813_;
  assign new_n54003_ = ys__n39776 & new_n53814_;
  assign new_n54004_ = ~new_n54002_ & ~new_n54003_;
  assign new_n54005_ = new_n54001_ & new_n54004_;
  assign new_n54006_ = ~new_n53997_ & ~new_n54005_;
  assign new_n54007_ = ~new_n53776_ & ~new_n54005_;
  assign new_n54008_ = ~new_n54006_ & ~new_n54007_;
  assign new_n54009_ = ~new_n53998_ & new_n54008_;
  assign new_n54010_ = ~new_n53984_ & ~new_n54009_;
  assign new_n54011_ = ~new_n53895_ & ~new_n54009_;
  assign new_n54012_ = ~new_n54010_ & ~new_n54011_;
  assign new_n54013_ = ~new_n53985_ & new_n54012_;
  assign new_n54014_ = ~new_n53973_ & ~new_n54013_;
  assign new_n54015_ = ~new_n53952_ & ~new_n54013_;
  assign new_n54016_ = ~new_n54014_ & ~new_n54015_;
  assign ys__n42189 = new_n53974_ | ~new_n54016_;
  assign new_n54018_ = ~new_n53952_ & new_n54014_;
  assign new_n54019_ = new_n53952_ & ~new_n54013_;
  assign new_n54020_ = new_n53973_ & new_n54019_;
  assign new_n54021_ = ~new_n53952_ & new_n54013_;
  assign new_n54022_ = new_n53973_ & new_n54021_;
  assign new_n54023_ = new_n53952_ & new_n54013_;
  assign new_n54024_ = ~new_n53973_ & new_n54023_;
  assign new_n54025_ = ~new_n54022_ & ~new_n54024_;
  assign new_n54026_ = ~new_n54020_ & new_n54025_;
  assign ys__n42194 = new_n54018_ | ~new_n54026_;
  assign new_n54028_ = ~new_n53895_ & new_n54010_;
  assign new_n54029_ = new_n53895_ & ~new_n54009_;
  assign new_n54030_ = new_n53984_ & new_n54029_;
  assign new_n54031_ = ~new_n53895_ & new_n54009_;
  assign new_n54032_ = new_n53984_ & new_n54031_;
  assign new_n54033_ = new_n53895_ & new_n54009_;
  assign new_n54034_ = ~new_n53984_ & new_n54033_;
  assign new_n54035_ = ~new_n54032_ & ~new_n54034_;
  assign new_n54036_ = ~new_n54030_ & new_n54035_;
  assign new_n54037_ = ~new_n54028_ & new_n54036_;
  assign new_n54038_ = ~new_n53952_ & ~new_n54037_;
  assign new_n54039_ = ~new_n53776_ & new_n54006_;
  assign new_n54040_ = new_n53997_ & new_n54005_;
  assign new_n54041_ = ~new_n53776_ & new_n54040_;
  assign new_n54042_ = ~new_n54039_ & ~new_n54041_;
  assign new_n54043_ = ~new_n53997_ & new_n54005_;
  assign new_n54044_ = new_n53776_ & new_n54043_;
  assign new_n54045_ = new_n53997_ & ~new_n54005_;
  assign new_n54046_ = new_n53776_ & new_n54045_;
  assign new_n54047_ = ~new_n54044_ & ~new_n54046_;
  assign new_n54048_ = new_n54042_ & new_n54047_;
  assign new_n54049_ = ~new_n53895_ & ~new_n54048_;
  assign new_n54050_ = ys__n24834 & new_n53788_;
  assign new_n54051_ = ys__n39778 & new_n53780_;
  assign new_n54052_ = ~new_n54050_ & ~new_n54051_;
  assign new_n54053_ = ys__n33745 & new_n53794_;
  assign new_n54054_ = ~ys__n33745 & new_n53797_;
  assign new_n54055_ = ~new_n54053_ & ~new_n54054_;
  assign new_n54056_ = new_n54052_ & new_n54055_;
  assign new_n54057_ = ~new_n53987_ & ~new_n53989_;
  assign new_n54058_ = new_n53995_ & new_n54057_;
  assign new_n54059_ = new_n54056_ & new_n54058_;
  assign new_n54060_ = ~new_n53776_ & ~new_n54059_;
  assign new_n54061_ = ys__n24831 & new_n53805_;
  assign new_n54062_ = ys__n24828 & new_n53806_;
  assign new_n54063_ = ~new_n54061_ & ~new_n54062_;
  assign new_n54064_ = ys__n39776 & new_n53813_;
  assign new_n54065_ = ys__n39774 & new_n53814_;
  assign new_n54066_ = ~new_n54064_ & ~new_n54065_;
  assign new_n54067_ = new_n54063_ & new_n54066_;
  assign new_n54068_ = ~new_n54059_ & ~new_n54067_;
  assign new_n54069_ = ~new_n53776_ & ~new_n54067_;
  assign new_n54070_ = ~new_n54068_ & ~new_n54069_;
  assign new_n54071_ = ~new_n54060_ & new_n54070_;
  assign new_n54072_ = ~new_n54048_ & ~new_n54071_;
  assign new_n54073_ = ~new_n53895_ & ~new_n54071_;
  assign new_n54074_ = ~new_n54072_ & ~new_n54073_;
  assign new_n54075_ = ~new_n54049_ & new_n54074_;
  assign new_n54076_ = ~new_n54037_ & ~new_n54075_;
  assign new_n54077_ = ~new_n53952_ & ~new_n54075_;
  assign new_n54078_ = ~new_n54076_ & ~new_n54077_;
  assign ys__n42229 = new_n54038_ | ~new_n54078_;
  assign new_n54080_ = ~new_n53952_ & new_n54076_;
  assign new_n54081_ = new_n53952_ & ~new_n54075_;
  assign new_n54082_ = new_n54037_ & new_n54081_;
  assign new_n54083_ = ~new_n53952_ & new_n54075_;
  assign new_n54084_ = new_n54037_ & new_n54083_;
  assign new_n54085_ = new_n53952_ & new_n54075_;
  assign new_n54086_ = ~new_n54037_ & new_n54085_;
  assign new_n54087_ = ~new_n54084_ & ~new_n54086_;
  assign new_n54088_ = ~new_n54082_ & new_n54087_;
  assign ys__n42234 = new_n54080_ | ~new_n54088_;
  assign new_n54090_ = ~new_n53895_ & new_n54072_;
  assign new_n54091_ = ~new_n53895_ & new_n54071_;
  assign new_n54092_ = new_n54048_ & new_n54091_;
  assign new_n54093_ = ~new_n54090_ & ~new_n54092_;
  assign new_n54094_ = new_n53895_ & new_n54071_;
  assign new_n54095_ = ~new_n54048_ & new_n54094_;
  assign new_n54096_ = new_n53895_ & ~new_n54071_;
  assign new_n54097_ = new_n54048_ & new_n54096_;
  assign new_n54098_ = ~new_n54095_ & ~new_n54097_;
  assign new_n54099_ = new_n54093_ & new_n54098_;
  assign new_n54100_ = ~new_n53952_ & ~new_n54099_;
  assign new_n54101_ = ~new_n53776_ & new_n54068_;
  assign new_n54102_ = new_n54059_ & new_n54067_;
  assign new_n54103_ = ~new_n53776_ & new_n54102_;
  assign new_n54104_ = ~new_n54101_ & ~new_n54103_;
  assign new_n54105_ = ~new_n54059_ & new_n54067_;
  assign new_n54106_ = new_n53776_ & new_n54105_;
  assign new_n54107_ = new_n54059_ & ~new_n54067_;
  assign new_n54108_ = new_n53776_ & new_n54107_;
  assign new_n54109_ = ~new_n54106_ & ~new_n54108_;
  assign new_n54110_ = new_n54104_ & new_n54109_;
  assign new_n54111_ = ~new_n53895_ & ~new_n54110_;
  assign new_n54112_ = ys__n39778 & new_n53781_;
  assign new_n54113_ = ys__n39776 & new_n53780_;
  assign new_n54114_ = ~new_n54112_ & ~new_n54113_;
  assign new_n54115_ = ys__n33743 & new_n53794_;
  assign new_n54116_ = ~ys__n33743 & new_n53797_;
  assign new_n54117_ = ~new_n54115_ & ~new_n54116_;
  assign new_n54118_ = new_n54114_ & new_n54117_;
  assign new_n54119_ = ~new_n53987_ & ~new_n53993_;
  assign new_n54120_ = ys__n24834 & new_n53789_;
  assign new_n54121_ = ys__n24831 & new_n53788_;
  assign new_n54122_ = ~new_n54120_ & ~new_n54121_;
  assign new_n54123_ = new_n54119_ & new_n54122_;
  assign new_n54124_ = new_n54118_ & new_n54123_;
  assign new_n54125_ = ~new_n53776_ & ~new_n54124_;
  assign new_n54126_ = ys__n24828 & new_n53805_;
  assign new_n54127_ = ys__n24825 & new_n53806_;
  assign new_n54128_ = ~new_n54126_ & ~new_n54127_;
  assign new_n54129_ = ys__n39774 & new_n53813_;
  assign new_n54130_ = ys__n39772 & new_n53814_;
  assign new_n54131_ = ~new_n54129_ & ~new_n54130_;
  assign new_n54132_ = new_n54128_ & new_n54131_;
  assign new_n54133_ = ~new_n54124_ & ~new_n54132_;
  assign new_n54134_ = ~new_n53776_ & ~new_n54132_;
  assign new_n54135_ = ~new_n54133_ & ~new_n54134_;
  assign new_n54136_ = ~new_n54125_ & new_n54135_;
  assign new_n54137_ = ~new_n54110_ & ~new_n54136_;
  assign new_n54138_ = ~new_n53895_ & ~new_n54136_;
  assign new_n54139_ = ~new_n54137_ & ~new_n54138_;
  assign new_n54140_ = ~new_n54111_ & new_n54139_;
  assign new_n54141_ = ~new_n54099_ & ~new_n54140_;
  assign new_n54142_ = ~new_n53952_ & ~new_n54140_;
  assign new_n54143_ = ~new_n54141_ & ~new_n54142_;
  assign ys__n42270 = new_n54100_ | ~new_n54143_;
  assign new_n54145_ = ~new_n53952_ & new_n54141_;
  assign new_n54146_ = new_n53952_ & ~new_n54140_;
  assign new_n54147_ = new_n54099_ & new_n54146_;
  assign new_n54148_ = ~new_n53952_ & new_n54140_;
  assign new_n54149_ = new_n54099_ & new_n54148_;
  assign new_n54150_ = new_n53952_ & new_n54140_;
  assign new_n54151_ = ~new_n54099_ & new_n54150_;
  assign new_n54152_ = ~new_n54149_ & ~new_n54151_;
  assign new_n54153_ = ~new_n54147_ & new_n54152_;
  assign ys__n42275 = new_n54145_ | ~new_n54153_;
  assign new_n54155_ = ~new_n53895_ & new_n54137_;
  assign new_n54156_ = ~new_n53895_ & new_n54136_;
  assign new_n54157_ = new_n54110_ & new_n54156_;
  assign new_n54158_ = ~new_n54155_ & ~new_n54157_;
  assign new_n54159_ = new_n53895_ & new_n54136_;
  assign new_n54160_ = ~new_n54110_ & new_n54159_;
  assign new_n54161_ = new_n53895_ & ~new_n54136_;
  assign new_n54162_ = new_n54110_ & new_n54161_;
  assign new_n54163_ = ~new_n54160_ & ~new_n54162_;
  assign new_n54164_ = new_n54158_ & new_n54163_;
  assign new_n54165_ = ~new_n53952_ & ~new_n54164_;
  assign new_n54166_ = ~new_n53776_ & new_n54133_;
  assign new_n54167_ = new_n54124_ & new_n54132_;
  assign new_n54168_ = ~new_n53776_ & new_n54167_;
  assign new_n54169_ = ~new_n54166_ & ~new_n54168_;
  assign new_n54170_ = ~new_n54124_ & new_n54132_;
  assign new_n54171_ = new_n53776_ & new_n54170_;
  assign new_n54172_ = new_n54124_ & ~new_n54132_;
  assign new_n54173_ = new_n53776_ & new_n54172_;
  assign new_n54174_ = ~new_n54171_ & ~new_n54173_;
  assign new_n54175_ = new_n54169_ & new_n54174_;
  assign new_n54176_ = ~new_n53895_ & ~new_n54175_;
  assign new_n54177_ = ys__n39776 & new_n53781_;
  assign new_n54178_ = ys__n39774 & new_n53780_;
  assign new_n54179_ = ~new_n54177_ & ~new_n54178_;
  assign new_n54180_ = ys__n33741 & new_n53794_;
  assign new_n54181_ = ~ys__n33741 & new_n53797_;
  assign new_n54182_ = ~new_n54180_ & ~new_n54181_;
  assign new_n54183_ = new_n54179_ & new_n54182_;
  assign new_n54184_ = ys__n24834 & new_n53786_;
  assign new_n54185_ = ys__n24831 & new_n53789_;
  assign new_n54186_ = ~new_n54184_ & ~new_n54185_;
  assign new_n54187_ = ys__n24828 & new_n53788_;
  assign new_n54188_ = ys__n39778 & new_n53778_;
  assign new_n54189_ = ~new_n54187_ & ~new_n54188_;
  assign new_n54190_ = new_n54186_ & new_n54189_;
  assign new_n54191_ = new_n54183_ & new_n54190_;
  assign new_n54192_ = ys__n39518 & new_n53763_;
  assign new_n54193_ = ys__n39520 & new_n53753_;
  assign new_n54194_ = ~new_n54192_ & ~new_n54193_;
  assign new_n54195_ = ys__n39520 & new_n53756_;
  assign new_n54196_ = ys__n39520 & new_n53755_;
  assign new_n54197_ = ~new_n54195_ & ~new_n54196_;
  assign new_n54198_ = new_n54194_ & new_n54197_;
  assign new_n54199_ = ys__n39518 & new_n53761_;
  assign new_n54200_ = ys__n39518 & new_n53764_;
  assign new_n54201_ = ~new_n54199_ & ~new_n54200_;
  assign new_n54202_ = new_n53774_ & new_n54201_;
  assign new_n54203_ = new_n54198_ & new_n54202_;
  assign new_n54204_ = ~new_n54191_ & ~new_n54203_;
  assign new_n54205_ = ys__n24825 & new_n53805_;
  assign new_n54206_ = ys__n24822 & new_n53806_;
  assign new_n54207_ = ~new_n54205_ & ~new_n54206_;
  assign new_n54208_ = ys__n39772 & new_n53813_;
  assign new_n54209_ = ys__n39770 & new_n53814_;
  assign new_n54210_ = ~new_n54208_ & ~new_n54209_;
  assign new_n54211_ = new_n54207_ & new_n54210_;
  assign new_n54212_ = ~new_n54191_ & ~new_n54211_;
  assign new_n54213_ = ~new_n54203_ & ~new_n54211_;
  assign new_n54214_ = ~new_n54212_ & ~new_n54213_;
  assign new_n54215_ = ~new_n54204_ & new_n54214_;
  assign new_n54216_ = ~new_n54175_ & ~new_n54215_;
  assign new_n54217_ = ~new_n53895_ & ~new_n54215_;
  assign new_n54218_ = ~new_n54216_ & ~new_n54217_;
  assign new_n54219_ = ~new_n54176_ & new_n54218_;
  assign new_n54220_ = ~new_n54164_ & ~new_n54219_;
  assign new_n54221_ = ~new_n53952_ & ~new_n54219_;
  assign new_n54222_ = ~new_n54220_ & ~new_n54221_;
  assign ys__n42311 = new_n54165_ | ~new_n54222_;
  assign new_n54224_ = ~new_n53952_ & new_n54220_;
  assign new_n54225_ = new_n53952_ & ~new_n54219_;
  assign new_n54226_ = new_n54164_ & new_n54225_;
  assign new_n54227_ = ~new_n53952_ & new_n54219_;
  assign new_n54228_ = new_n54164_ & new_n54227_;
  assign new_n54229_ = new_n53952_ & new_n54219_;
  assign new_n54230_ = ~new_n54164_ & new_n54229_;
  assign new_n54231_ = ~new_n54228_ & ~new_n54230_;
  assign new_n54232_ = ~new_n54226_ & new_n54231_;
  assign ys__n42316 = new_n54224_ | ~new_n54232_;
  assign new_n54234_ = ~new_n53895_ & new_n54216_;
  assign new_n54235_ = ~new_n53895_ & new_n54215_;
  assign new_n54236_ = new_n54175_ & new_n54235_;
  assign new_n54237_ = ~new_n54234_ & ~new_n54236_;
  assign new_n54238_ = new_n53895_ & new_n54215_;
  assign new_n54239_ = ~new_n54175_ & new_n54238_;
  assign new_n54240_ = new_n53895_ & ~new_n54215_;
  assign new_n54241_ = new_n54175_ & new_n54240_;
  assign new_n54242_ = ~new_n54239_ & ~new_n54241_;
  assign new_n54243_ = new_n54237_ & new_n54242_;
  assign new_n54244_ = ~new_n53952_ & ~new_n54243_;
  assign new_n54245_ = ~new_n54203_ & new_n54212_;
  assign new_n54246_ = new_n54191_ & new_n54211_;
  assign new_n54247_ = ~new_n54203_ & new_n54246_;
  assign new_n54248_ = ~new_n54245_ & ~new_n54247_;
  assign new_n54249_ = ~new_n54191_ & new_n54211_;
  assign new_n54250_ = new_n54203_ & new_n54249_;
  assign new_n54251_ = new_n54191_ & ~new_n54211_;
  assign new_n54252_ = new_n54203_ & new_n54251_;
  assign new_n54253_ = ~new_n54250_ & ~new_n54252_;
  assign new_n54254_ = new_n54248_ & new_n54253_;
  assign new_n54255_ = ~new_n53895_ & ~new_n54254_;
  assign new_n54256_ = ys__n39774 & new_n53781_;
  assign new_n54257_ = ys__n39772 & new_n53780_;
  assign new_n54258_ = ~new_n54256_ & ~new_n54257_;
  assign new_n54259_ = ys__n33739 & new_n53794_;
  assign new_n54260_ = ~ys__n33739 & new_n53797_;
  assign new_n54261_ = ~new_n54259_ & ~new_n54260_;
  assign new_n54262_ = new_n54258_ & new_n54261_;
  assign new_n54263_ = ys__n24831 & new_n53786_;
  assign new_n54264_ = ys__n24828 & new_n53789_;
  assign new_n54265_ = ~new_n54263_ & ~new_n54264_;
  assign new_n54266_ = ys__n24825 & new_n53788_;
  assign new_n54267_ = ys__n39776 & new_n53778_;
  assign new_n54268_ = ~new_n54266_ & ~new_n54267_;
  assign new_n54269_ = new_n54265_ & new_n54268_;
  assign new_n54270_ = new_n54262_ & new_n54269_;
  assign new_n54271_ = ys__n24834 & new_n53763_;
  assign new_n54272_ = ys__n39778 & new_n53755_;
  assign new_n54273_ = ~new_n54271_ & ~new_n54272_;
  assign new_n54274_ = ys__n33745 & new_n53769_;
  assign new_n54275_ = ~ys__n33745 & new_n53772_;
  assign new_n54276_ = ~new_n54274_ & ~new_n54275_;
  assign new_n54277_ = new_n54273_ & new_n54276_;
  assign new_n54278_ = ~new_n54193_ & ~new_n54195_;
  assign new_n54279_ = new_n54201_ & new_n54278_;
  assign new_n54280_ = new_n54277_ & new_n54279_;
  assign new_n54281_ = ~new_n54270_ & ~new_n54280_;
  assign new_n54282_ = ys__n24822 & new_n53805_;
  assign new_n54283_ = ys__n24819 & new_n53806_;
  assign new_n54284_ = ~new_n54282_ & ~new_n54283_;
  assign new_n54285_ = ys__n39770 & new_n53813_;
  assign new_n54286_ = ys__n39768 & new_n53814_;
  assign new_n54287_ = ~new_n54285_ & ~new_n54286_;
  assign new_n54288_ = new_n54284_ & new_n54287_;
  assign new_n54289_ = ~new_n54270_ & ~new_n54288_;
  assign new_n54290_ = ~new_n54280_ & ~new_n54288_;
  assign new_n54291_ = ~new_n54289_ & ~new_n54290_;
  assign new_n54292_ = ~new_n54281_ & new_n54291_;
  assign new_n54293_ = ~new_n54254_ & ~new_n54292_;
  assign new_n54294_ = ~new_n53895_ & ~new_n54292_;
  assign new_n54295_ = ~new_n54293_ & ~new_n54294_;
  assign new_n54296_ = ~new_n54255_ & new_n54295_;
  assign new_n54297_ = ~new_n54243_ & ~new_n54296_;
  assign new_n54298_ = ~new_n53952_ & ~new_n54296_;
  assign new_n54299_ = ~new_n54297_ & ~new_n54298_;
  assign ys__n42352 = new_n54244_ | ~new_n54299_;
  assign new_n54301_ = ~new_n53952_ & new_n54297_;
  assign new_n54302_ = new_n53952_ & ~new_n54296_;
  assign new_n54303_ = new_n54243_ & new_n54302_;
  assign new_n54304_ = ~new_n53952_ & new_n54296_;
  assign new_n54305_ = new_n54243_ & new_n54304_;
  assign new_n54306_ = new_n53952_ & new_n54296_;
  assign new_n54307_ = ~new_n54243_ & new_n54306_;
  assign new_n54308_ = ~new_n54305_ & ~new_n54307_;
  assign new_n54309_ = ~new_n54303_ & new_n54308_;
  assign ys__n42357 = new_n54301_ | ~new_n54309_;
  assign new_n54311_ = ~new_n53895_ & new_n54293_;
  assign new_n54312_ = ~new_n53895_ & new_n54292_;
  assign new_n54313_ = new_n54254_ & new_n54312_;
  assign new_n54314_ = ~new_n54311_ & ~new_n54313_;
  assign new_n54315_ = new_n53895_ & new_n54292_;
  assign new_n54316_ = ~new_n54254_ & new_n54315_;
  assign new_n54317_ = new_n53895_ & ~new_n54292_;
  assign new_n54318_ = new_n54254_ & new_n54317_;
  assign new_n54319_ = ~new_n54316_ & ~new_n54318_;
  assign new_n54320_ = new_n54314_ & new_n54319_;
  assign new_n54321_ = ~new_n53952_ & ~new_n54320_;
  assign new_n54322_ = ~new_n54280_ & new_n54289_;
  assign new_n54323_ = new_n54270_ & new_n54288_;
  assign new_n54324_ = ~new_n54280_ & new_n54323_;
  assign new_n54325_ = ~new_n54322_ & ~new_n54324_;
  assign new_n54326_ = ~new_n54270_ & new_n54288_;
  assign new_n54327_ = new_n54280_ & new_n54326_;
  assign new_n54328_ = new_n54270_ & ~new_n54288_;
  assign new_n54329_ = new_n54280_ & new_n54328_;
  assign new_n54330_ = ~new_n54327_ & ~new_n54329_;
  assign new_n54331_ = new_n54325_ & new_n54330_;
  assign new_n54332_ = ~new_n53895_ & ~new_n54331_;
  assign new_n54333_ = ys__n39772 & new_n53781_;
  assign new_n54334_ = ys__n39770 & new_n53780_;
  assign new_n54335_ = ~new_n54333_ & ~new_n54334_;
  assign new_n54336_ = ys__n33737 & new_n53794_;
  assign new_n54337_ = ~ys__n33737 & new_n53797_;
  assign new_n54338_ = ~new_n54336_ & ~new_n54337_;
  assign new_n54339_ = new_n54335_ & new_n54338_;
  assign new_n54340_ = ys__n24828 & new_n53786_;
  assign new_n54341_ = ys__n24825 & new_n53789_;
  assign new_n54342_ = ~new_n54340_ & ~new_n54341_;
  assign new_n54343_ = ys__n24822 & new_n53788_;
  assign new_n54344_ = ys__n39774 & new_n53778_;
  assign new_n54345_ = ~new_n54343_ & ~new_n54344_;
  assign new_n54346_ = new_n54342_ & new_n54345_;
  assign new_n54347_ = new_n54339_ & new_n54346_;
  assign new_n54348_ = ys__n39778 & new_n53756_;
  assign new_n54349_ = ys__n39776 & new_n53755_;
  assign new_n54350_ = ~new_n54348_ & ~new_n54349_;
  assign new_n54351_ = ys__n33743 & new_n53769_;
  assign new_n54352_ = ~ys__n33743 & new_n53772_;
  assign new_n54353_ = ~new_n54351_ & ~new_n54352_;
  assign new_n54354_ = new_n54350_ & new_n54353_;
  assign new_n54355_ = ~new_n54193_ & ~new_n54199_;
  assign new_n54356_ = ys__n24834 & new_n53764_;
  assign new_n54357_ = ys__n24831 & new_n53763_;
  assign new_n54358_ = ~new_n54356_ & ~new_n54357_;
  assign new_n54359_ = new_n54355_ & new_n54358_;
  assign new_n54360_ = new_n54354_ & new_n54359_;
  assign new_n54361_ = ~new_n54347_ & ~new_n54360_;
  assign new_n54362_ = ys__n24819 & new_n53805_;
  assign new_n54363_ = ys__n24816 & new_n53806_;
  assign new_n54364_ = ~new_n54362_ & ~new_n54363_;
  assign new_n54365_ = ys__n39768 & new_n53813_;
  assign new_n54366_ = ys__n39766 & new_n53814_;
  assign new_n54367_ = ~new_n54365_ & ~new_n54366_;
  assign new_n54368_ = new_n54364_ & new_n54367_;
  assign new_n54369_ = ~new_n54347_ & ~new_n54368_;
  assign new_n54370_ = ~new_n54360_ & ~new_n54368_;
  assign new_n54371_ = ~new_n54369_ & ~new_n54370_;
  assign new_n54372_ = ~new_n54361_ & new_n54371_;
  assign new_n54373_ = ~new_n54331_ & ~new_n54372_;
  assign new_n54374_ = ~new_n53895_ & ~new_n54372_;
  assign new_n54375_ = ~new_n54373_ & ~new_n54374_;
  assign new_n54376_ = ~new_n54332_ & new_n54375_;
  assign new_n54377_ = ~new_n54320_ & ~new_n54376_;
  assign new_n54378_ = ~new_n53952_ & ~new_n54376_;
  assign new_n54379_ = ~new_n54377_ & ~new_n54378_;
  assign ys__n42393 = new_n54321_ | ~new_n54379_;
  assign new_n54381_ = ~new_n53952_ & new_n54377_;
  assign new_n54382_ = new_n53952_ & ~new_n54376_;
  assign new_n54383_ = new_n54320_ & new_n54382_;
  assign new_n54384_ = ~new_n53952_ & new_n54376_;
  assign new_n54385_ = new_n54320_ & new_n54384_;
  assign new_n54386_ = new_n53952_ & new_n54376_;
  assign new_n54387_ = ~new_n54320_ & new_n54386_;
  assign new_n54388_ = ~new_n54385_ & ~new_n54387_;
  assign new_n54389_ = ~new_n54383_ & new_n54388_;
  assign ys__n42398 = new_n54381_ | ~new_n54389_;
  assign new_n54391_ = ~new_n53895_ & new_n54373_;
  assign new_n54392_ = ~new_n53895_ & new_n54372_;
  assign new_n54393_ = new_n54331_ & new_n54392_;
  assign new_n54394_ = ~new_n54391_ & ~new_n54393_;
  assign new_n54395_ = new_n53895_ & new_n54372_;
  assign new_n54396_ = ~new_n54331_ & new_n54395_;
  assign new_n54397_ = new_n53895_ & ~new_n54372_;
  assign new_n54398_ = new_n54331_ & new_n54397_;
  assign new_n54399_ = ~new_n54396_ & ~new_n54398_;
  assign new_n54400_ = new_n54394_ & new_n54399_;
  assign new_n54401_ = ~new_n53952_ & ~new_n54400_;
  assign new_n54402_ = ~new_n54360_ & new_n54369_;
  assign new_n54403_ = new_n54347_ & new_n54368_;
  assign new_n54404_ = ~new_n54360_ & new_n54403_;
  assign new_n54405_ = ~new_n54402_ & ~new_n54404_;
  assign new_n54406_ = ~new_n54347_ & new_n54368_;
  assign new_n54407_ = new_n54360_ & new_n54406_;
  assign new_n54408_ = new_n54347_ & ~new_n54368_;
  assign new_n54409_ = new_n54360_ & new_n54408_;
  assign new_n54410_ = ~new_n54407_ & ~new_n54409_;
  assign new_n54411_ = new_n54405_ & new_n54410_;
  assign new_n54412_ = ys__n39518 & new_n53878_;
  assign new_n54413_ = ys__n39520 & new_n53868_;
  assign new_n54414_ = ~new_n54412_ & ~new_n54413_;
  assign new_n54415_ = ys__n39520 & new_n53871_;
  assign new_n54416_ = ys__n39520 & new_n53870_;
  assign new_n54417_ = ~new_n54415_ & ~new_n54416_;
  assign new_n54418_ = new_n54414_ & new_n54417_;
  assign new_n54419_ = ys__n39518 & new_n53876_;
  assign new_n54420_ = ys__n39518 & new_n53879_;
  assign new_n54421_ = ~new_n54419_ & ~new_n54420_;
  assign new_n54422_ = new_n53889_ & new_n54421_;
  assign new_n54423_ = new_n54418_ & new_n54422_;
  assign new_n54424_ = ~new_n53865_ & ~new_n54423_;
  assign new_n54425_ = ~new_n53854_ & ~new_n54423_;
  assign new_n54426_ = ~new_n53866_ & ~new_n54425_;
  assign new_n54427_ = ~new_n54424_ & new_n54426_;
  assign new_n54428_ = ~new_n54411_ & ~new_n54427_;
  assign new_n54429_ = ys__n39770 & new_n53781_;
  assign new_n54430_ = ys__n39768 & new_n53780_;
  assign new_n54431_ = ~new_n54429_ & ~new_n54430_;
  assign new_n54432_ = ys__n33735 & new_n53794_;
  assign new_n54433_ = ~ys__n33735 & new_n53797_;
  assign new_n54434_ = ~new_n54432_ & ~new_n54433_;
  assign new_n54435_ = new_n54431_ & new_n54434_;
  assign new_n54436_ = ys__n24825 & new_n53786_;
  assign new_n54437_ = ys__n24822 & new_n53789_;
  assign new_n54438_ = ~new_n54436_ & ~new_n54437_;
  assign new_n54439_ = ys__n24819 & new_n53788_;
  assign new_n54440_ = ys__n39772 & new_n53778_;
  assign new_n54441_ = ~new_n54439_ & ~new_n54440_;
  assign new_n54442_ = new_n54438_ & new_n54441_;
  assign new_n54443_ = new_n54435_ & new_n54442_;
  assign new_n54444_ = ys__n39776 & new_n53756_;
  assign new_n54445_ = ys__n39774 & new_n53755_;
  assign new_n54446_ = ~new_n54444_ & ~new_n54445_;
  assign new_n54447_ = ys__n33741 & new_n53769_;
  assign new_n54448_ = ~ys__n33741 & new_n53772_;
  assign new_n54449_ = ~new_n54447_ & ~new_n54448_;
  assign new_n54450_ = new_n54446_ & new_n54449_;
  assign new_n54451_ = ys__n24834 & new_n53761_;
  assign new_n54452_ = ys__n24831 & new_n53764_;
  assign new_n54453_ = ~new_n54451_ & ~new_n54452_;
  assign new_n54454_ = ys__n24828 & new_n53763_;
  assign new_n54455_ = ys__n39778 & new_n53753_;
  assign new_n54456_ = ~new_n54454_ & ~new_n54455_;
  assign new_n54457_ = new_n54453_ & new_n54456_;
  assign new_n54458_ = new_n54450_ & new_n54457_;
  assign new_n54459_ = ~new_n54443_ & ~new_n54458_;
  assign new_n54460_ = ys__n24816 & new_n53805_;
  assign new_n54461_ = ys__n24813 & new_n53806_;
  assign new_n54462_ = ~new_n54460_ & ~new_n54461_;
  assign new_n54463_ = ys__n39766 & new_n53813_;
  assign new_n54464_ = ys__n39764 & new_n53814_;
  assign new_n54465_ = ~new_n54463_ & ~new_n54464_;
  assign new_n54466_ = new_n54462_ & new_n54465_;
  assign new_n54467_ = ~new_n54443_ & ~new_n54466_;
  assign new_n54468_ = ~new_n54458_ & ~new_n54466_;
  assign new_n54469_ = ~new_n54467_ & ~new_n54468_;
  assign new_n54470_ = ~new_n54459_ & new_n54469_;
  assign new_n54471_ = ~new_n54411_ & ~new_n54470_;
  assign new_n54472_ = ~new_n54427_ & ~new_n54470_;
  assign new_n54473_ = ~new_n54471_ & ~new_n54472_;
  assign new_n54474_ = ~new_n54428_ & new_n54473_;
  assign new_n54475_ = ~new_n54400_ & ~new_n54474_;
  assign new_n54476_ = ~new_n53952_ & ~new_n54474_;
  assign new_n54477_ = ~new_n54475_ & ~new_n54476_;
  assign ys__n42434 = new_n54401_ | ~new_n54477_;
  assign new_n54479_ = ~new_n53952_ & new_n54475_;
  assign new_n54480_ = new_n53952_ & ~new_n54474_;
  assign new_n54481_ = new_n54400_ & new_n54480_;
  assign new_n54482_ = ~new_n53952_ & new_n54474_;
  assign new_n54483_ = new_n54400_ & new_n54482_;
  assign new_n54484_ = new_n53952_ & new_n54474_;
  assign new_n54485_ = ~new_n54400_ & new_n54484_;
  assign new_n54486_ = ~new_n54483_ & ~new_n54485_;
  assign new_n54487_ = ~new_n54481_ & new_n54486_;
  assign ys__n42439 = new_n54479_ | ~new_n54487_;
  assign new_n54489_ = ~new_n54427_ & new_n54471_;
  assign new_n54490_ = new_n54411_ & new_n54470_;
  assign new_n54491_ = ~new_n54427_ & new_n54490_;
  assign new_n54492_ = ~new_n54489_ & ~new_n54491_;
  assign new_n54493_ = ~new_n54411_ & new_n54470_;
  assign new_n54494_ = new_n54427_ & new_n54493_;
  assign new_n54495_ = new_n54411_ & ~new_n54470_;
  assign new_n54496_ = new_n54427_ & new_n54495_;
  assign new_n54497_ = ~new_n54494_ & ~new_n54496_;
  assign new_n54498_ = new_n54492_ & new_n54497_;
  assign new_n54499_ = ~new_n53952_ & ~new_n54498_;
  assign new_n54500_ = ~new_n54458_ & new_n54467_;
  assign new_n54501_ = new_n54443_ & new_n54466_;
  assign new_n54502_ = ~new_n54458_ & new_n54501_;
  assign new_n54503_ = ~new_n54500_ & ~new_n54502_;
  assign new_n54504_ = ~new_n54443_ & new_n54466_;
  assign new_n54505_ = new_n54458_ & new_n54504_;
  assign new_n54506_ = new_n54443_ & ~new_n54466_;
  assign new_n54507_ = new_n54458_ & new_n54506_;
  assign new_n54508_ = ~new_n54505_ & ~new_n54507_;
  assign new_n54509_ = new_n54503_ & new_n54508_;
  assign new_n54510_ = ys__n24834 & new_n53878_;
  assign new_n54511_ = ys__n39778 & new_n53870_;
  assign new_n54512_ = ~new_n54510_ & ~new_n54511_;
  assign new_n54513_ = ys__n33745 & new_n53884_;
  assign new_n54514_ = ~ys__n33745 & new_n53887_;
  assign new_n54515_ = ~new_n54513_ & ~new_n54514_;
  assign new_n54516_ = new_n54512_ & new_n54515_;
  assign new_n54517_ = ~new_n54413_ & ~new_n54415_;
  assign new_n54518_ = new_n54421_ & new_n54517_;
  assign new_n54519_ = new_n54516_ & new_n54518_;
  assign new_n54520_ = ~new_n53865_ & ~new_n54519_;
  assign new_n54521_ = ~new_n53854_ & ~new_n54519_;
  assign new_n54522_ = ~new_n53866_ & ~new_n54521_;
  assign new_n54523_ = ~new_n54520_ & new_n54522_;
  assign new_n54524_ = ~new_n54509_ & ~new_n54523_;
  assign new_n54525_ = ys__n39768 & new_n53781_;
  assign new_n54526_ = ys__n39766 & new_n53780_;
  assign new_n54527_ = ~new_n54525_ & ~new_n54526_;
  assign new_n54528_ = ys__n33733 & new_n53794_;
  assign new_n54529_ = ~ys__n33733 & new_n53797_;
  assign new_n54530_ = ~new_n54528_ & ~new_n54529_;
  assign new_n54531_ = new_n54527_ & new_n54530_;
  assign new_n54532_ = ys__n24822 & new_n53786_;
  assign new_n54533_ = ys__n24819 & new_n53789_;
  assign new_n54534_ = ~new_n54532_ & ~new_n54533_;
  assign new_n54535_ = ys__n24816 & new_n53788_;
  assign new_n54536_ = ys__n39770 & new_n53778_;
  assign new_n54537_ = ~new_n54535_ & ~new_n54536_;
  assign new_n54538_ = new_n54534_ & new_n54537_;
  assign new_n54539_ = new_n54531_ & new_n54538_;
  assign new_n54540_ = ys__n39774 & new_n53756_;
  assign new_n54541_ = ys__n39772 & new_n53755_;
  assign new_n54542_ = ~new_n54540_ & ~new_n54541_;
  assign new_n54543_ = ys__n33739 & new_n53769_;
  assign new_n54544_ = ~ys__n33739 & new_n53772_;
  assign new_n54545_ = ~new_n54543_ & ~new_n54544_;
  assign new_n54546_ = new_n54542_ & new_n54545_;
  assign new_n54547_ = ys__n24831 & new_n53761_;
  assign new_n54548_ = ys__n24828 & new_n53764_;
  assign new_n54549_ = ~new_n54547_ & ~new_n54548_;
  assign new_n54550_ = ys__n24825 & new_n53763_;
  assign new_n54551_ = ys__n39776 & new_n53753_;
  assign new_n54552_ = ~new_n54550_ & ~new_n54551_;
  assign new_n54553_ = new_n54549_ & new_n54552_;
  assign new_n54554_ = new_n54546_ & new_n54553_;
  assign new_n54555_ = ~new_n54539_ & ~new_n54554_;
  assign new_n54556_ = ys__n24813 & new_n53805_;
  assign new_n54557_ = ys__n24810 & new_n53806_;
  assign new_n54558_ = ~new_n54556_ & ~new_n54557_;
  assign new_n54559_ = ys__n39764 & new_n53813_;
  assign new_n54560_ = ys__n39762 & new_n53814_;
  assign new_n54561_ = ~new_n54559_ & ~new_n54560_;
  assign new_n54562_ = new_n54558_ & new_n54561_;
  assign new_n54563_ = ~new_n54539_ & ~new_n54562_;
  assign new_n54564_ = ~new_n54554_ & ~new_n54562_;
  assign new_n54565_ = ~new_n54563_ & ~new_n54564_;
  assign new_n54566_ = ~new_n54555_ & new_n54565_;
  assign new_n54567_ = ~new_n54509_ & ~new_n54566_;
  assign new_n54568_ = ~new_n54523_ & ~new_n54566_;
  assign new_n54569_ = ~new_n54567_ & ~new_n54568_;
  assign new_n54570_ = ~new_n54524_ & new_n54569_;
  assign new_n54571_ = ~new_n54498_ & ~new_n54570_;
  assign new_n54572_ = ~new_n53952_ & ~new_n54570_;
  assign new_n54573_ = ~new_n54571_ & ~new_n54572_;
  assign ys__n42488 = new_n54499_ | ~new_n54573_;
  assign new_n54575_ = ~new_n53952_ & new_n54571_;
  assign new_n54576_ = new_n53952_ & ~new_n54570_;
  assign new_n54577_ = new_n54498_ & new_n54576_;
  assign new_n54578_ = ~new_n53952_ & new_n54570_;
  assign new_n54579_ = new_n54498_ & new_n54578_;
  assign new_n54580_ = new_n53952_ & new_n54570_;
  assign new_n54581_ = ~new_n54498_ & new_n54580_;
  assign new_n54582_ = ~new_n54579_ & ~new_n54581_;
  assign new_n54583_ = ~new_n54577_ & new_n54582_;
  assign ys__n42493 = new_n54575_ | ~new_n54583_;
  assign new_n54585_ = ~new_n54523_ & new_n54567_;
  assign new_n54586_ = new_n54509_ & new_n54566_;
  assign new_n54587_ = ~new_n54523_ & new_n54586_;
  assign new_n54588_ = ~new_n54585_ & ~new_n54587_;
  assign new_n54589_ = ~new_n54509_ & new_n54566_;
  assign new_n54590_ = new_n54523_ & new_n54589_;
  assign new_n54591_ = new_n54509_ & ~new_n54566_;
  assign new_n54592_ = new_n54523_ & new_n54591_;
  assign new_n54593_ = ~new_n54590_ & ~new_n54592_;
  assign new_n54594_ = new_n54588_ & new_n54593_;
  assign new_n54595_ = ~new_n53865_ & new_n54425_;
  assign new_n54596_ = new_n53854_ & new_n54423_;
  assign new_n54597_ = ~new_n53865_ & new_n54596_;
  assign new_n54598_ = ~new_n54595_ & ~new_n54597_;
  assign new_n54599_ = ~new_n53854_ & new_n54423_;
  assign new_n54600_ = new_n53865_ & new_n54599_;
  assign new_n54601_ = new_n53854_ & ~new_n54423_;
  assign new_n54602_ = new_n53865_ & new_n54601_;
  assign new_n54603_ = ~new_n54600_ & ~new_n54602_;
  assign new_n54604_ = new_n54598_ & new_n54603_;
  assign new_n54605_ = ~new_n54594_ & ~new_n54604_;
  assign new_n54606_ = ~new_n54554_ & new_n54563_;
  assign new_n54607_ = new_n54539_ & new_n54562_;
  assign new_n54608_ = ~new_n54554_ & new_n54607_;
  assign new_n54609_ = ~new_n54606_ & ~new_n54608_;
  assign new_n54610_ = ~new_n54539_ & new_n54562_;
  assign new_n54611_ = new_n54554_ & new_n54610_;
  assign new_n54612_ = new_n54539_ & ~new_n54562_;
  assign new_n54613_ = new_n54554_ & new_n54612_;
  assign new_n54614_ = ~new_n54611_ & ~new_n54613_;
  assign new_n54615_ = new_n54609_ & new_n54614_;
  assign new_n54616_ = ys__n39778 & new_n53871_;
  assign new_n54617_ = ys__n39776 & new_n53870_;
  assign new_n54618_ = ~new_n54616_ & ~new_n54617_;
  assign new_n54619_ = ys__n33743 & new_n53884_;
  assign new_n54620_ = ~ys__n33743 & new_n53887_;
  assign new_n54621_ = ~new_n54619_ & ~new_n54620_;
  assign new_n54622_ = new_n54618_ & new_n54621_;
  assign new_n54623_ = ~new_n54413_ & ~new_n54419_;
  assign new_n54624_ = ys__n24834 & new_n53879_;
  assign new_n54625_ = ys__n24831 & new_n53878_;
  assign new_n54626_ = ~new_n54624_ & ~new_n54625_;
  assign new_n54627_ = new_n54623_ & new_n54626_;
  assign new_n54628_ = new_n54622_ & new_n54627_;
  assign new_n54629_ = ~new_n53865_ & ~new_n54628_;
  assign new_n54630_ = ~new_n53854_ & ~new_n54628_;
  assign new_n54631_ = ~new_n53866_ & ~new_n54630_;
  assign new_n54632_ = ~new_n54629_ & new_n54631_;
  assign new_n54633_ = ~new_n54615_ & ~new_n54632_;
  assign new_n54634_ = ys__n39766 & new_n53781_;
  assign new_n54635_ = ys__n39764 & new_n53780_;
  assign new_n54636_ = ~new_n54634_ & ~new_n54635_;
  assign new_n54637_ = ys__n33731 & new_n53794_;
  assign new_n54638_ = ~ys__n33731 & new_n53797_;
  assign new_n54639_ = ~new_n54637_ & ~new_n54638_;
  assign new_n54640_ = new_n54636_ & new_n54639_;
  assign new_n54641_ = ys__n24819 & new_n53786_;
  assign new_n54642_ = ys__n24816 & new_n53789_;
  assign new_n54643_ = ~new_n54641_ & ~new_n54642_;
  assign new_n54644_ = ys__n24813 & new_n53788_;
  assign new_n54645_ = ys__n39768 & new_n53778_;
  assign new_n54646_ = ~new_n54644_ & ~new_n54645_;
  assign new_n54647_ = new_n54643_ & new_n54646_;
  assign new_n54648_ = new_n54640_ & new_n54647_;
  assign new_n54649_ = ys__n39772 & new_n53756_;
  assign new_n54650_ = ys__n39770 & new_n53755_;
  assign new_n54651_ = ~new_n54649_ & ~new_n54650_;
  assign new_n54652_ = ys__n33737 & new_n53769_;
  assign new_n54653_ = ~ys__n33737 & new_n53772_;
  assign new_n54654_ = ~new_n54652_ & ~new_n54653_;
  assign new_n54655_ = new_n54651_ & new_n54654_;
  assign new_n54656_ = ys__n24828 & new_n53761_;
  assign new_n54657_ = ys__n24825 & new_n53764_;
  assign new_n54658_ = ~new_n54656_ & ~new_n54657_;
  assign new_n54659_ = ys__n24822 & new_n53763_;
  assign new_n54660_ = ys__n39774 & new_n53753_;
  assign new_n54661_ = ~new_n54659_ & ~new_n54660_;
  assign new_n54662_ = new_n54658_ & new_n54661_;
  assign new_n54663_ = new_n54655_ & new_n54662_;
  assign new_n54664_ = ~new_n54648_ & ~new_n54663_;
  assign new_n54665_ = ys__n24810 & new_n53805_;
  assign new_n54666_ = ys__n24807 & new_n53806_;
  assign new_n54667_ = ~new_n54665_ & ~new_n54666_;
  assign new_n54668_ = ys__n39762 & new_n53813_;
  assign new_n54669_ = ys__n39760 & new_n53814_;
  assign new_n54670_ = ~new_n54668_ & ~new_n54669_;
  assign new_n54671_ = new_n54667_ & new_n54670_;
  assign new_n54672_ = ~new_n54648_ & ~new_n54671_;
  assign new_n54673_ = ~new_n54663_ & ~new_n54671_;
  assign new_n54674_ = ~new_n54672_ & ~new_n54673_;
  assign new_n54675_ = ~new_n54664_ & new_n54674_;
  assign new_n54676_ = ~new_n54615_ & ~new_n54675_;
  assign new_n54677_ = ~new_n54632_ & ~new_n54675_;
  assign new_n54678_ = ~new_n54676_ & ~new_n54677_;
  assign new_n54679_ = ~new_n54633_ & new_n54678_;
  assign new_n54680_ = ~new_n54594_ & ~new_n54679_;
  assign new_n54681_ = ~new_n54604_ & ~new_n54679_;
  assign new_n54682_ = ~new_n54680_ & ~new_n54681_;
  assign ys__n42541 = new_n54605_ | ~new_n54682_;
  assign new_n54684_ = ~new_n54604_ & new_n54680_;
  assign new_n54685_ = new_n54604_ & ~new_n54679_;
  assign new_n54686_ = new_n54594_ & new_n54685_;
  assign new_n54687_ = ~new_n54604_ & new_n54679_;
  assign new_n54688_ = new_n54594_ & new_n54687_;
  assign new_n54689_ = new_n54604_ & new_n54679_;
  assign new_n54690_ = ~new_n54594_ & new_n54689_;
  assign new_n54691_ = ~new_n54688_ & ~new_n54690_;
  assign new_n54692_ = ~new_n54686_ & new_n54691_;
  assign ys__n42546 = new_n54684_ | ~new_n54692_;
  assign new_n54694_ = ~new_n54632_ & new_n54676_;
  assign new_n54695_ = new_n54615_ & new_n54675_;
  assign new_n54696_ = ~new_n54632_ & new_n54695_;
  assign new_n54697_ = ~new_n54694_ & ~new_n54696_;
  assign new_n54698_ = ~new_n54615_ & new_n54675_;
  assign new_n54699_ = new_n54632_ & new_n54698_;
  assign new_n54700_ = new_n54615_ & ~new_n54675_;
  assign new_n54701_ = new_n54632_ & new_n54700_;
  assign new_n54702_ = ~new_n54699_ & ~new_n54701_;
  assign new_n54703_ = new_n54697_ & new_n54702_;
  assign new_n54704_ = ~new_n53865_ & new_n54521_;
  assign new_n54705_ = new_n53854_ & new_n54519_;
  assign new_n54706_ = ~new_n53865_ & new_n54705_;
  assign new_n54707_ = ~new_n54704_ & ~new_n54706_;
  assign new_n54708_ = ~new_n53854_ & new_n54519_;
  assign new_n54709_ = new_n53865_ & new_n54708_;
  assign new_n54710_ = new_n53854_ & ~new_n54519_;
  assign new_n54711_ = new_n53865_ & new_n54710_;
  assign new_n54712_ = ~new_n54709_ & ~new_n54711_;
  assign new_n54713_ = new_n54707_ & new_n54712_;
  assign new_n54714_ = ~new_n54703_ & ~new_n54713_;
  assign new_n54715_ = ~new_n54663_ & new_n54672_;
  assign new_n54716_ = new_n54648_ & new_n54671_;
  assign new_n54717_ = ~new_n54663_ & new_n54716_;
  assign new_n54718_ = ~new_n54715_ & ~new_n54717_;
  assign new_n54719_ = ~new_n54648_ & new_n54671_;
  assign new_n54720_ = new_n54663_ & new_n54719_;
  assign new_n54721_ = new_n54648_ & ~new_n54671_;
  assign new_n54722_ = new_n54663_ & new_n54721_;
  assign new_n54723_ = ~new_n54720_ & ~new_n54722_;
  assign new_n54724_ = new_n54718_ & new_n54723_;
  assign new_n54725_ = ys__n39518 & new_n53841_;
  assign new_n54726_ = ys__n39520 & new_n53831_;
  assign new_n54727_ = ~new_n54725_ & ~new_n54726_;
  assign new_n54728_ = ys__n39520 & new_n53834_;
  assign new_n54729_ = ys__n39520 & new_n53833_;
  assign new_n54730_ = ~new_n54728_ & ~new_n54729_;
  assign new_n54731_ = new_n54727_ & new_n54730_;
  assign new_n54732_ = ys__n39518 & new_n53839_;
  assign new_n54733_ = ys__n39518 & new_n53842_;
  assign new_n54734_ = ~new_n54732_ & ~new_n54733_;
  assign new_n54735_ = new_n53852_ & new_n54734_;
  assign new_n54736_ = new_n54731_ & new_n54735_;
  assign new_n54737_ = ~new_n53865_ & ~new_n54736_;
  assign new_n54738_ = ys__n39776 & new_n53871_;
  assign new_n54739_ = ys__n39774 & new_n53870_;
  assign new_n54740_ = ~new_n54738_ & ~new_n54739_;
  assign new_n54741_ = ys__n33741 & new_n53884_;
  assign new_n54742_ = ~ys__n33741 & new_n53887_;
  assign new_n54743_ = ~new_n54741_ & ~new_n54742_;
  assign new_n54744_ = new_n54740_ & new_n54743_;
  assign new_n54745_ = ys__n24834 & new_n53876_;
  assign new_n54746_ = ys__n24831 & new_n53879_;
  assign new_n54747_ = ~new_n54745_ & ~new_n54746_;
  assign new_n54748_ = ys__n24828 & new_n53878_;
  assign new_n54749_ = ys__n39778 & new_n53868_;
  assign new_n54750_ = ~new_n54748_ & ~new_n54749_;
  assign new_n54751_ = new_n54747_ & new_n54750_;
  assign new_n54752_ = new_n54744_ & new_n54751_;
  assign new_n54753_ = ~new_n54736_ & ~new_n54752_;
  assign new_n54754_ = ~new_n53865_ & ~new_n54752_;
  assign new_n54755_ = ~new_n54753_ & ~new_n54754_;
  assign new_n54756_ = ~new_n54737_ & new_n54755_;
  assign new_n54757_ = ~new_n54724_ & ~new_n54756_;
  assign new_n54758_ = ys__n39764 & new_n53781_;
  assign new_n54759_ = ys__n39762 & new_n53780_;
  assign new_n54760_ = ~new_n54758_ & ~new_n54759_;
  assign new_n54761_ = ys__n33729 & new_n53794_;
  assign new_n54762_ = ~ys__n33729 & new_n53797_;
  assign new_n54763_ = ~new_n54761_ & ~new_n54762_;
  assign new_n54764_ = new_n54760_ & new_n54763_;
  assign new_n54765_ = ys__n24816 & new_n53786_;
  assign new_n54766_ = ys__n24813 & new_n53789_;
  assign new_n54767_ = ~new_n54765_ & ~new_n54766_;
  assign new_n54768_ = ys__n24810 & new_n53788_;
  assign new_n54769_ = ys__n39766 & new_n53778_;
  assign new_n54770_ = ~new_n54768_ & ~new_n54769_;
  assign new_n54771_ = new_n54767_ & new_n54770_;
  assign new_n54772_ = new_n54764_ & new_n54771_;
  assign new_n54773_ = ys__n39770 & new_n53756_;
  assign new_n54774_ = ys__n39768 & new_n53755_;
  assign new_n54775_ = ~new_n54773_ & ~new_n54774_;
  assign new_n54776_ = ys__n33735 & new_n53769_;
  assign new_n54777_ = ~ys__n33735 & new_n53772_;
  assign new_n54778_ = ~new_n54776_ & ~new_n54777_;
  assign new_n54779_ = new_n54775_ & new_n54778_;
  assign new_n54780_ = ys__n24825 & new_n53761_;
  assign new_n54781_ = ys__n24822 & new_n53764_;
  assign new_n54782_ = ~new_n54780_ & ~new_n54781_;
  assign new_n54783_ = ys__n24819 & new_n53763_;
  assign new_n54784_ = ys__n39772 & new_n53753_;
  assign new_n54785_ = ~new_n54783_ & ~new_n54784_;
  assign new_n54786_ = new_n54782_ & new_n54785_;
  assign new_n54787_ = new_n54779_ & new_n54786_;
  assign new_n54788_ = ~new_n54772_ & ~new_n54787_;
  assign new_n54789_ = ys__n24807 & new_n53805_;
  assign new_n54790_ = ys__n24804 & new_n53806_;
  assign new_n54791_ = ~new_n54789_ & ~new_n54790_;
  assign new_n54792_ = ys__n39760 & new_n53813_;
  assign new_n54793_ = ys__n39758 & new_n53814_;
  assign new_n54794_ = ~new_n54792_ & ~new_n54793_;
  assign new_n54795_ = new_n54791_ & new_n54794_;
  assign new_n54796_ = ~new_n54772_ & ~new_n54795_;
  assign new_n54797_ = ~new_n54787_ & ~new_n54795_;
  assign new_n54798_ = ~new_n54796_ & ~new_n54797_;
  assign new_n54799_ = ~new_n54788_ & new_n54798_;
  assign new_n54800_ = ~new_n54724_ & ~new_n54799_;
  assign new_n54801_ = ~new_n54756_ & ~new_n54799_;
  assign new_n54802_ = ~new_n54800_ & ~new_n54801_;
  assign new_n54803_ = ~new_n54757_ & new_n54802_;
  assign new_n54804_ = ~new_n54703_ & ~new_n54803_;
  assign new_n54805_ = ~new_n54713_ & ~new_n54803_;
  assign new_n54806_ = ~new_n54804_ & ~new_n54805_;
  assign ys__n42594 = new_n54714_ | ~new_n54806_;
  assign new_n54808_ = ~new_n54713_ & new_n54804_;
  assign new_n54809_ = new_n54713_ & ~new_n54803_;
  assign new_n54810_ = new_n54703_ & new_n54809_;
  assign new_n54811_ = ~new_n54713_ & new_n54803_;
  assign new_n54812_ = new_n54703_ & new_n54811_;
  assign new_n54813_ = new_n54713_ & new_n54803_;
  assign new_n54814_ = ~new_n54703_ & new_n54813_;
  assign new_n54815_ = ~new_n54812_ & ~new_n54814_;
  assign new_n54816_ = ~new_n54810_ & new_n54815_;
  assign ys__n42599 = new_n54808_ | ~new_n54816_;
  assign new_n54818_ = ~new_n54756_ & new_n54800_;
  assign new_n54819_ = new_n54724_ & new_n54799_;
  assign new_n54820_ = ~new_n54756_ & new_n54819_;
  assign new_n54821_ = ~new_n54818_ & ~new_n54820_;
  assign new_n54822_ = ~new_n54724_ & new_n54799_;
  assign new_n54823_ = new_n54756_ & new_n54822_;
  assign new_n54824_ = new_n54724_ & ~new_n54799_;
  assign new_n54825_ = new_n54756_ & new_n54824_;
  assign new_n54826_ = ~new_n54823_ & ~new_n54825_;
  assign new_n54827_ = new_n54821_ & new_n54826_;
  assign new_n54828_ = ~new_n53865_ & new_n54630_;
  assign new_n54829_ = new_n53854_ & new_n54628_;
  assign new_n54830_ = ~new_n53865_ & new_n54829_;
  assign new_n54831_ = ~new_n54828_ & ~new_n54830_;
  assign new_n54832_ = ~new_n53854_ & new_n54628_;
  assign new_n54833_ = new_n53865_ & new_n54832_;
  assign new_n54834_ = new_n53854_ & ~new_n54628_;
  assign new_n54835_ = new_n53865_ & new_n54834_;
  assign new_n54836_ = ~new_n54833_ & ~new_n54835_;
  assign new_n54837_ = new_n54831_ & new_n54836_;
  assign new_n54838_ = ~new_n54827_ & ~new_n54837_;
  assign new_n54839_ = ~new_n54787_ & new_n54796_;
  assign new_n54840_ = new_n54772_ & new_n54795_;
  assign new_n54841_ = ~new_n54787_ & new_n54840_;
  assign new_n54842_ = ~new_n54839_ & ~new_n54841_;
  assign new_n54843_ = ~new_n54772_ & new_n54795_;
  assign new_n54844_ = new_n54787_ & new_n54843_;
  assign new_n54845_ = new_n54772_ & ~new_n54795_;
  assign new_n54846_ = new_n54787_ & new_n54845_;
  assign new_n54847_ = ~new_n54844_ & ~new_n54846_;
  assign new_n54848_ = new_n54842_ & new_n54847_;
  assign new_n54849_ = ys__n24834 & new_n53841_;
  assign new_n54850_ = ys__n39778 & new_n53833_;
  assign new_n54851_ = ~new_n54849_ & ~new_n54850_;
  assign new_n54852_ = ys__n33745 & new_n53847_;
  assign new_n54853_ = ~ys__n33745 & new_n53850_;
  assign new_n54854_ = ~new_n54852_ & ~new_n54853_;
  assign new_n54855_ = new_n54851_ & new_n54854_;
  assign new_n54856_ = ~new_n54726_ & ~new_n54728_;
  assign new_n54857_ = new_n54734_ & new_n54856_;
  assign new_n54858_ = new_n54855_ & new_n54857_;
  assign new_n54859_ = ~new_n53865_ & ~new_n54858_;
  assign new_n54860_ = ys__n39774 & new_n53871_;
  assign new_n54861_ = ys__n39772 & new_n53870_;
  assign new_n54862_ = ~new_n54860_ & ~new_n54861_;
  assign new_n54863_ = ys__n33739 & new_n53884_;
  assign new_n54864_ = ~ys__n33739 & new_n53887_;
  assign new_n54865_ = ~new_n54863_ & ~new_n54864_;
  assign new_n54866_ = new_n54862_ & new_n54865_;
  assign new_n54867_ = ys__n24831 & new_n53876_;
  assign new_n54868_ = ys__n24828 & new_n53879_;
  assign new_n54869_ = ~new_n54867_ & ~new_n54868_;
  assign new_n54870_ = ys__n24825 & new_n53878_;
  assign new_n54871_ = ys__n39776 & new_n53868_;
  assign new_n54872_ = ~new_n54870_ & ~new_n54871_;
  assign new_n54873_ = new_n54869_ & new_n54872_;
  assign new_n54874_ = new_n54866_ & new_n54873_;
  assign new_n54875_ = ~new_n54858_ & ~new_n54874_;
  assign new_n54876_ = ~new_n53865_ & ~new_n54874_;
  assign new_n54877_ = ~new_n54875_ & ~new_n54876_;
  assign new_n54878_ = ~new_n54859_ & new_n54877_;
  assign new_n54879_ = ~new_n54848_ & ~new_n54878_;
  assign new_n54880_ = ys__n39762 & new_n53781_;
  assign new_n54881_ = ys__n39760 & new_n53780_;
  assign new_n54882_ = ~new_n54880_ & ~new_n54881_;
  assign new_n54883_ = ys__n33727 & new_n53794_;
  assign new_n54884_ = ~ys__n33727 & new_n53797_;
  assign new_n54885_ = ~new_n54883_ & ~new_n54884_;
  assign new_n54886_ = new_n54882_ & new_n54885_;
  assign new_n54887_ = ys__n24813 & new_n53786_;
  assign new_n54888_ = ys__n24810 & new_n53789_;
  assign new_n54889_ = ~new_n54887_ & ~new_n54888_;
  assign new_n54890_ = ys__n24807 & new_n53788_;
  assign new_n54891_ = ys__n39764 & new_n53778_;
  assign new_n54892_ = ~new_n54890_ & ~new_n54891_;
  assign new_n54893_ = new_n54889_ & new_n54892_;
  assign new_n54894_ = new_n54886_ & new_n54893_;
  assign new_n54895_ = ys__n39768 & new_n53756_;
  assign new_n54896_ = ys__n39766 & new_n53755_;
  assign new_n54897_ = ~new_n54895_ & ~new_n54896_;
  assign new_n54898_ = ys__n33733 & new_n53769_;
  assign new_n54899_ = ~ys__n33733 & new_n53772_;
  assign new_n54900_ = ~new_n54898_ & ~new_n54899_;
  assign new_n54901_ = new_n54897_ & new_n54900_;
  assign new_n54902_ = ys__n24822 & new_n53761_;
  assign new_n54903_ = ys__n24819 & new_n53764_;
  assign new_n54904_ = ~new_n54902_ & ~new_n54903_;
  assign new_n54905_ = ys__n24816 & new_n53763_;
  assign new_n54906_ = ys__n39770 & new_n53753_;
  assign new_n54907_ = ~new_n54905_ & ~new_n54906_;
  assign new_n54908_ = new_n54904_ & new_n54907_;
  assign new_n54909_ = new_n54901_ & new_n54908_;
  assign new_n54910_ = ~new_n54894_ & ~new_n54909_;
  assign new_n54911_ = ys__n24804 & new_n53805_;
  assign new_n54912_ = ys__n24801 & new_n53806_;
  assign new_n54913_ = ~new_n54911_ & ~new_n54912_;
  assign new_n54914_ = ys__n39758 & new_n53813_;
  assign new_n54915_ = ys__n39756 & new_n53814_;
  assign new_n54916_ = ~new_n54914_ & ~new_n54915_;
  assign new_n54917_ = new_n54913_ & new_n54916_;
  assign new_n54918_ = ~new_n54894_ & ~new_n54917_;
  assign new_n54919_ = ~new_n54909_ & ~new_n54917_;
  assign new_n54920_ = ~new_n54918_ & ~new_n54919_;
  assign new_n54921_ = ~new_n54910_ & new_n54920_;
  assign new_n54922_ = ~new_n54848_ & ~new_n54921_;
  assign new_n54923_ = ~new_n54878_ & ~new_n54921_;
  assign new_n54924_ = ~new_n54922_ & ~new_n54923_;
  assign new_n54925_ = ~new_n54879_ & new_n54924_;
  assign new_n54926_ = ~new_n54827_ & ~new_n54925_;
  assign new_n54927_ = ~new_n54837_ & ~new_n54925_;
  assign new_n54928_ = ~new_n54926_ & ~new_n54927_;
  assign ys__n42647 = new_n54838_ | ~new_n54928_;
  assign new_n54930_ = ~new_n54837_ & new_n54926_;
  assign new_n54931_ = new_n54837_ & ~new_n54925_;
  assign new_n54932_ = new_n54827_ & new_n54931_;
  assign new_n54933_ = ~new_n54837_ & new_n54925_;
  assign new_n54934_ = new_n54827_ & new_n54933_;
  assign new_n54935_ = new_n54837_ & new_n54925_;
  assign new_n54936_ = ~new_n54827_ & new_n54935_;
  assign new_n54937_ = ~new_n54934_ & ~new_n54936_;
  assign new_n54938_ = ~new_n54932_ & new_n54937_;
  assign ys__n42652 = new_n54930_ | ~new_n54938_;
  assign new_n54940_ = ~new_n54878_ & new_n54922_;
  assign new_n54941_ = new_n54848_ & new_n54921_;
  assign new_n54942_ = ~new_n54878_ & new_n54941_;
  assign new_n54943_ = ~new_n54940_ & ~new_n54942_;
  assign new_n54944_ = ~new_n54848_ & new_n54921_;
  assign new_n54945_ = new_n54878_ & new_n54944_;
  assign new_n54946_ = new_n54848_ & ~new_n54921_;
  assign new_n54947_ = new_n54878_ & new_n54946_;
  assign new_n54948_ = ~new_n54945_ & ~new_n54947_;
  assign new_n54949_ = new_n54943_ & new_n54948_;
  assign new_n54950_ = ~new_n53865_ & new_n54753_;
  assign new_n54951_ = new_n54736_ & new_n54752_;
  assign new_n54952_ = ~new_n53865_ & new_n54951_;
  assign new_n54953_ = ~new_n54950_ & ~new_n54952_;
  assign new_n54954_ = ~new_n54736_ & new_n54752_;
  assign new_n54955_ = new_n53865_ & new_n54954_;
  assign new_n54956_ = new_n54736_ & ~new_n54752_;
  assign new_n54957_ = new_n53865_ & new_n54956_;
  assign new_n54958_ = ~new_n54955_ & ~new_n54957_;
  assign new_n54959_ = new_n54953_ & new_n54958_;
  assign new_n54960_ = ~new_n54949_ & ~new_n54959_;
  assign new_n54961_ = ~new_n54909_ & new_n54918_;
  assign new_n54962_ = new_n54894_ & new_n54917_;
  assign new_n54963_ = ~new_n54909_ & new_n54962_;
  assign new_n54964_ = ~new_n54961_ & ~new_n54963_;
  assign new_n54965_ = ~new_n54894_ & new_n54917_;
  assign new_n54966_ = new_n54909_ & new_n54965_;
  assign new_n54967_ = new_n54894_ & ~new_n54917_;
  assign new_n54968_ = new_n54909_ & new_n54967_;
  assign new_n54969_ = ~new_n54966_ & ~new_n54968_;
  assign new_n54970_ = new_n54964_ & new_n54969_;
  assign new_n54971_ = ys__n39778 & new_n53834_;
  assign new_n54972_ = ys__n39776 & new_n53833_;
  assign new_n54973_ = ~new_n54971_ & ~new_n54972_;
  assign new_n54974_ = ys__n33743 & new_n53847_;
  assign new_n54975_ = ~ys__n33743 & new_n53850_;
  assign new_n54976_ = ~new_n54974_ & ~new_n54975_;
  assign new_n54977_ = new_n54973_ & new_n54976_;
  assign new_n54978_ = ~new_n54726_ & ~new_n54732_;
  assign new_n54979_ = ys__n24834 & new_n53842_;
  assign new_n54980_ = ys__n24831 & new_n53841_;
  assign new_n54981_ = ~new_n54979_ & ~new_n54980_;
  assign new_n54982_ = new_n54978_ & new_n54981_;
  assign new_n54983_ = new_n54977_ & new_n54982_;
  assign new_n54984_ = ~new_n53865_ & ~new_n54983_;
  assign new_n54985_ = ys__n39772 & new_n53871_;
  assign new_n54986_ = ys__n39770 & new_n53870_;
  assign new_n54987_ = ~new_n54985_ & ~new_n54986_;
  assign new_n54988_ = ys__n33737 & new_n53884_;
  assign new_n54989_ = ~ys__n33737 & new_n53887_;
  assign new_n54990_ = ~new_n54988_ & ~new_n54989_;
  assign new_n54991_ = new_n54987_ & new_n54990_;
  assign new_n54992_ = ys__n24828 & new_n53876_;
  assign new_n54993_ = ys__n24825 & new_n53879_;
  assign new_n54994_ = ~new_n54992_ & ~new_n54993_;
  assign new_n54995_ = ys__n24822 & new_n53878_;
  assign new_n54996_ = ys__n39774 & new_n53868_;
  assign new_n54997_ = ~new_n54995_ & ~new_n54996_;
  assign new_n54998_ = new_n54994_ & new_n54997_;
  assign new_n54999_ = new_n54991_ & new_n54998_;
  assign new_n55000_ = ~new_n54983_ & ~new_n54999_;
  assign new_n55001_ = ~new_n53865_ & ~new_n54999_;
  assign new_n55002_ = ~new_n55000_ & ~new_n55001_;
  assign new_n55003_ = ~new_n54984_ & new_n55002_;
  assign new_n55004_ = ~new_n54970_ & ~new_n55003_;
  assign new_n55005_ = ys__n39760 & new_n53781_;
  assign new_n55006_ = ys__n39758 & new_n53780_;
  assign new_n55007_ = ~new_n55005_ & ~new_n55006_;
  assign new_n55008_ = ys__n33725 & new_n53794_;
  assign new_n55009_ = ~ys__n33725 & new_n53797_;
  assign new_n55010_ = ~new_n55008_ & ~new_n55009_;
  assign new_n55011_ = new_n55007_ & new_n55010_;
  assign new_n55012_ = ys__n24810 & new_n53786_;
  assign new_n55013_ = ys__n24807 & new_n53789_;
  assign new_n55014_ = ~new_n55012_ & ~new_n55013_;
  assign new_n55015_ = ys__n24804 & new_n53788_;
  assign new_n55016_ = ys__n39762 & new_n53778_;
  assign new_n55017_ = ~new_n55015_ & ~new_n55016_;
  assign new_n55018_ = new_n55014_ & new_n55017_;
  assign new_n55019_ = new_n55011_ & new_n55018_;
  assign new_n55020_ = ys__n39766 & new_n53756_;
  assign new_n55021_ = ys__n39764 & new_n53755_;
  assign new_n55022_ = ~new_n55020_ & ~new_n55021_;
  assign new_n55023_ = ys__n33731 & new_n53769_;
  assign new_n55024_ = ~ys__n33731 & new_n53772_;
  assign new_n55025_ = ~new_n55023_ & ~new_n55024_;
  assign new_n55026_ = new_n55022_ & new_n55025_;
  assign new_n55027_ = ys__n24819 & new_n53761_;
  assign new_n55028_ = ys__n24816 & new_n53764_;
  assign new_n55029_ = ~new_n55027_ & ~new_n55028_;
  assign new_n55030_ = ys__n24813 & new_n53763_;
  assign new_n55031_ = ys__n39768 & new_n53753_;
  assign new_n55032_ = ~new_n55030_ & ~new_n55031_;
  assign new_n55033_ = new_n55029_ & new_n55032_;
  assign new_n55034_ = new_n55026_ & new_n55033_;
  assign new_n55035_ = ~new_n55019_ & ~new_n55034_;
  assign new_n55036_ = ys__n24801 & new_n53805_;
  assign new_n55037_ = ys__n24798 & new_n53806_;
  assign new_n55038_ = ~new_n55036_ & ~new_n55037_;
  assign new_n55039_ = ys__n39756 & new_n53813_;
  assign new_n55040_ = ys__n39754 & new_n53814_;
  assign new_n55041_ = ~new_n55039_ & ~new_n55040_;
  assign new_n55042_ = new_n55038_ & new_n55041_;
  assign new_n55043_ = ~new_n55019_ & ~new_n55042_;
  assign new_n55044_ = ~new_n55034_ & ~new_n55042_;
  assign new_n55045_ = ~new_n55043_ & ~new_n55044_;
  assign new_n55046_ = ~new_n55035_ & new_n55045_;
  assign new_n55047_ = ~new_n54970_ & ~new_n55046_;
  assign new_n55048_ = ~new_n55003_ & ~new_n55046_;
  assign new_n55049_ = ~new_n55047_ & ~new_n55048_;
  assign new_n55050_ = ~new_n55004_ & new_n55049_;
  assign new_n55051_ = ~new_n54949_ & ~new_n55050_;
  assign new_n55052_ = ~new_n54959_ & ~new_n55050_;
  assign new_n55053_ = ~new_n55051_ & ~new_n55052_;
  assign ys__n42701 = new_n54960_ | ~new_n55053_;
  assign new_n55055_ = ~new_n54959_ & new_n55051_;
  assign new_n55056_ = new_n54959_ & ~new_n55050_;
  assign new_n55057_ = new_n54949_ & new_n55056_;
  assign new_n55058_ = ~new_n54959_ & new_n55050_;
  assign new_n55059_ = new_n54949_ & new_n55058_;
  assign new_n55060_ = new_n54959_ & new_n55050_;
  assign new_n55061_ = ~new_n54949_ & new_n55060_;
  assign new_n55062_ = ~new_n55059_ & ~new_n55061_;
  assign new_n55063_ = ~new_n55057_ & new_n55062_;
  assign ys__n42706 = new_n55055_ | ~new_n55063_;
  assign new_n55065_ = ~new_n55003_ & new_n55047_;
  assign new_n55066_ = new_n54970_ & new_n55046_;
  assign new_n55067_ = ~new_n55003_ & new_n55066_;
  assign new_n55068_ = ~new_n55065_ & ~new_n55067_;
  assign new_n55069_ = ~new_n54970_ & new_n55046_;
  assign new_n55070_ = new_n55003_ & new_n55069_;
  assign new_n55071_ = new_n54970_ & ~new_n55046_;
  assign new_n55072_ = new_n55003_ & new_n55071_;
  assign new_n55073_ = ~new_n55070_ & ~new_n55072_;
  assign new_n55074_ = new_n55068_ & new_n55073_;
  assign new_n55075_ = ~new_n53865_ & new_n54875_;
  assign new_n55076_ = new_n54858_ & new_n54874_;
  assign new_n55077_ = ~new_n53865_ & new_n55076_;
  assign new_n55078_ = ~new_n55075_ & ~new_n55077_;
  assign new_n55079_ = ~new_n54858_ & new_n54874_;
  assign new_n55080_ = new_n53865_ & new_n55079_;
  assign new_n55081_ = new_n54858_ & ~new_n54874_;
  assign new_n55082_ = new_n53865_ & new_n55081_;
  assign new_n55083_ = ~new_n55080_ & ~new_n55082_;
  assign new_n55084_ = new_n55078_ & new_n55083_;
  assign new_n55085_ = ~new_n55074_ & ~new_n55084_;
  assign new_n55086_ = ~new_n55034_ & new_n55043_;
  assign new_n55087_ = new_n55019_ & new_n55042_;
  assign new_n55088_ = ~new_n55034_ & new_n55087_;
  assign new_n55089_ = ~new_n55086_ & ~new_n55088_;
  assign new_n55090_ = ~new_n55019_ & new_n55042_;
  assign new_n55091_ = new_n55034_ & new_n55090_;
  assign new_n55092_ = new_n55019_ & ~new_n55042_;
  assign new_n55093_ = new_n55034_ & new_n55092_;
  assign new_n55094_ = ~new_n55091_ & ~new_n55093_;
  assign new_n55095_ = new_n55089_ & new_n55094_;
  assign new_n55096_ = ys__n39776 & new_n53834_;
  assign new_n55097_ = ys__n39774 & new_n53833_;
  assign new_n55098_ = ~new_n55096_ & ~new_n55097_;
  assign new_n55099_ = ys__n33741 & new_n53847_;
  assign new_n55100_ = ~ys__n33741 & new_n53850_;
  assign new_n55101_ = ~new_n55099_ & ~new_n55100_;
  assign new_n55102_ = new_n55098_ & new_n55101_;
  assign new_n55103_ = ys__n24834 & new_n53839_;
  assign new_n55104_ = ys__n24831 & new_n53842_;
  assign new_n55105_ = ~new_n55103_ & ~new_n55104_;
  assign new_n55106_ = ys__n24828 & new_n53841_;
  assign new_n55107_ = ys__n39778 & new_n53831_;
  assign new_n55108_ = ~new_n55106_ & ~new_n55107_;
  assign new_n55109_ = new_n55105_ & new_n55108_;
  assign new_n55110_ = new_n55102_ & new_n55109_;
  assign new_n55111_ = ys__n39518 & new_n53744_;
  assign new_n55112_ = ys__n39520 & new_n53746_;
  assign new_n55113_ = ~new_n55111_ & ~new_n55112_;
  assign new_n55114_ = ys__n39520 & new_n53723_;
  assign new_n55115_ = ys__n39520 & new_n53726_;
  assign new_n55116_ = ~new_n55114_ & ~new_n55115_;
  assign new_n55117_ = new_n55113_ & new_n55116_;
  assign new_n55118_ = ys__n39518 & new_n53738_;
  assign new_n55119_ = ys__n39518 & new_n53740_;
  assign new_n55120_ = ~new_n55118_ & ~new_n55119_;
  assign new_n55121_ = new_n53863_ & new_n55120_;
  assign new_n55122_ = new_n55117_ & new_n55121_;
  assign new_n55123_ = ~new_n55110_ & ~new_n55122_;
  assign new_n55124_ = ys__n39770 & new_n53871_;
  assign new_n55125_ = ys__n39768 & new_n53870_;
  assign new_n55126_ = ~new_n55124_ & ~new_n55125_;
  assign new_n55127_ = ys__n33735 & new_n53884_;
  assign new_n55128_ = ~ys__n33735 & new_n53887_;
  assign new_n55129_ = ~new_n55127_ & ~new_n55128_;
  assign new_n55130_ = new_n55126_ & new_n55129_;
  assign new_n55131_ = ys__n24825 & new_n53876_;
  assign new_n55132_ = ys__n24822 & new_n53879_;
  assign new_n55133_ = ~new_n55131_ & ~new_n55132_;
  assign new_n55134_ = ys__n24819 & new_n53878_;
  assign new_n55135_ = ys__n39772 & new_n53868_;
  assign new_n55136_ = ~new_n55134_ & ~new_n55135_;
  assign new_n55137_ = new_n55133_ & new_n55136_;
  assign new_n55138_ = new_n55130_ & new_n55137_;
  assign new_n55139_ = ~new_n55110_ & ~new_n55138_;
  assign new_n55140_ = ~new_n55122_ & ~new_n55138_;
  assign new_n55141_ = ~new_n55139_ & ~new_n55140_;
  assign new_n55142_ = ~new_n55123_ & new_n55141_;
  assign new_n55143_ = ~new_n55095_ & ~new_n55142_;
  assign new_n55144_ = ys__n39758 & new_n53781_;
  assign new_n55145_ = ys__n39756 & new_n53780_;
  assign new_n55146_ = ~new_n55144_ & ~new_n55145_;
  assign new_n55147_ = ys__n33723 & new_n53794_;
  assign new_n55148_ = ~ys__n33723 & new_n53797_;
  assign new_n55149_ = ~new_n55147_ & ~new_n55148_;
  assign new_n55150_ = new_n55146_ & new_n55149_;
  assign new_n55151_ = ys__n24807 & new_n53786_;
  assign new_n55152_ = ys__n24804 & new_n53789_;
  assign new_n55153_ = ~new_n55151_ & ~new_n55152_;
  assign new_n55154_ = ys__n24801 & new_n53788_;
  assign new_n55155_ = ys__n39760 & new_n53778_;
  assign new_n55156_ = ~new_n55154_ & ~new_n55155_;
  assign new_n55157_ = new_n55153_ & new_n55156_;
  assign new_n55158_ = new_n55150_ & new_n55157_;
  assign new_n55159_ = ys__n39764 & new_n53756_;
  assign new_n55160_ = ys__n39762 & new_n53755_;
  assign new_n55161_ = ~new_n55159_ & ~new_n55160_;
  assign new_n55162_ = ys__n33729 & new_n53769_;
  assign new_n55163_ = ~ys__n33729 & new_n53772_;
  assign new_n55164_ = ~new_n55162_ & ~new_n55163_;
  assign new_n55165_ = new_n55161_ & new_n55164_;
  assign new_n55166_ = ys__n24816 & new_n53761_;
  assign new_n55167_ = ys__n24813 & new_n53764_;
  assign new_n55168_ = ~new_n55166_ & ~new_n55167_;
  assign new_n55169_ = ys__n24810 & new_n53763_;
  assign new_n55170_ = ys__n39766 & new_n53753_;
  assign new_n55171_ = ~new_n55169_ & ~new_n55170_;
  assign new_n55172_ = new_n55168_ & new_n55171_;
  assign new_n55173_ = new_n55165_ & new_n55172_;
  assign new_n55174_ = ~new_n55158_ & ~new_n55173_;
  assign new_n55175_ = ys__n24798 & new_n53805_;
  assign new_n55176_ = ys__n24795 & new_n53806_;
  assign new_n55177_ = ~new_n55175_ & ~new_n55176_;
  assign new_n55178_ = ys__n39754 & new_n53813_;
  assign new_n55179_ = ys__n39752 & new_n53814_;
  assign new_n55180_ = ~new_n55178_ & ~new_n55179_;
  assign new_n55181_ = new_n55177_ & new_n55180_;
  assign new_n55182_ = ~new_n55158_ & ~new_n55181_;
  assign new_n55183_ = ~new_n55173_ & ~new_n55181_;
  assign new_n55184_ = ~new_n55182_ & ~new_n55183_;
  assign new_n55185_ = ~new_n55174_ & new_n55184_;
  assign new_n55186_ = ~new_n55095_ & ~new_n55185_;
  assign new_n55187_ = ~new_n55142_ & ~new_n55185_;
  assign new_n55188_ = ~new_n55186_ & ~new_n55187_;
  assign new_n55189_ = ~new_n55143_ & new_n55188_;
  assign new_n55190_ = ~new_n55074_ & ~new_n55189_;
  assign new_n55191_ = ~new_n55084_ & ~new_n55189_;
  assign new_n55192_ = ~new_n55190_ & ~new_n55191_;
  assign ys__n42755 = new_n55085_ | ~new_n55192_;
  assign new_n55194_ = ~new_n55084_ & new_n55190_;
  assign new_n55195_ = new_n55084_ & ~new_n55189_;
  assign new_n55196_ = new_n55074_ & new_n55195_;
  assign new_n55197_ = ~new_n55084_ & new_n55189_;
  assign new_n55198_ = new_n55074_ & new_n55197_;
  assign new_n55199_ = new_n55084_ & new_n55189_;
  assign new_n55200_ = ~new_n55074_ & new_n55199_;
  assign new_n55201_ = ~new_n55198_ & ~new_n55200_;
  assign new_n55202_ = ~new_n55196_ & new_n55201_;
  assign ys__n42760 = new_n55194_ | ~new_n55202_;
  assign new_n55204_ = ~new_n55142_ & new_n55186_;
  assign new_n55205_ = new_n55142_ & ~new_n55185_;
  assign new_n55206_ = new_n55095_ & new_n55205_;
  assign new_n55207_ = ~new_n55142_ & new_n55185_;
  assign new_n55208_ = new_n55095_ & new_n55207_;
  assign new_n55209_ = new_n55142_ & new_n55185_;
  assign new_n55210_ = ~new_n55095_ & new_n55209_;
  assign new_n55211_ = ~new_n55208_ & ~new_n55210_;
  assign new_n55212_ = ~new_n55206_ & new_n55211_;
  assign new_n55213_ = ~new_n55204_ & new_n55212_;
  assign new_n55214_ = ~new_n53865_ & new_n55000_;
  assign new_n55215_ = new_n54983_ & new_n54999_;
  assign new_n55216_ = ~new_n53865_ & new_n55215_;
  assign new_n55217_ = ~new_n55214_ & ~new_n55216_;
  assign new_n55218_ = ~new_n54983_ & new_n54999_;
  assign new_n55219_ = new_n53865_ & new_n55218_;
  assign new_n55220_ = new_n54983_ & ~new_n54999_;
  assign new_n55221_ = new_n53865_ & new_n55220_;
  assign new_n55222_ = ~new_n55219_ & ~new_n55221_;
  assign new_n55223_ = new_n55217_ & new_n55222_;
  assign new_n55224_ = ~new_n55213_ & ~new_n55223_;
  assign new_n55225_ = ~new_n55173_ & new_n55182_;
  assign new_n55226_ = new_n55158_ & new_n55181_;
  assign new_n55227_ = ~new_n55173_ & new_n55226_;
  assign new_n55228_ = ~new_n55225_ & ~new_n55227_;
  assign new_n55229_ = ~new_n55158_ & new_n55181_;
  assign new_n55230_ = new_n55173_ & new_n55229_;
  assign new_n55231_ = new_n55158_ & ~new_n55181_;
  assign new_n55232_ = new_n55173_ & new_n55231_;
  assign new_n55233_ = ~new_n55230_ & ~new_n55232_;
  assign new_n55234_ = new_n55228_ & new_n55233_;
  assign new_n55235_ = ys__n39774 & new_n53834_;
  assign new_n55236_ = ys__n39772 & new_n53833_;
  assign new_n55237_ = ~new_n55235_ & ~new_n55236_;
  assign new_n55238_ = ys__n33739 & new_n53847_;
  assign new_n55239_ = ~ys__n33739 & new_n53850_;
  assign new_n55240_ = ~new_n55238_ & ~new_n55239_;
  assign new_n55241_ = new_n55237_ & new_n55240_;
  assign new_n55242_ = ys__n24831 & new_n53839_;
  assign new_n55243_ = ys__n24828 & new_n53842_;
  assign new_n55244_ = ~new_n55242_ & ~new_n55243_;
  assign new_n55245_ = ys__n24825 & new_n53841_;
  assign new_n55246_ = ys__n39776 & new_n53831_;
  assign new_n55247_ = ~new_n55245_ & ~new_n55246_;
  assign new_n55248_ = new_n55244_ & new_n55247_;
  assign new_n55249_ = new_n55241_ & new_n55248_;
  assign new_n55250_ = ys__n24834 & new_n53744_;
  assign new_n55251_ = ys__n39778 & new_n53726_;
  assign new_n55252_ = ~new_n55250_ & ~new_n55251_;
  assign new_n55253_ = ys__n33745 & new_n53730_;
  assign new_n55254_ = ~ys__n33745 & new_n53733_;
  assign new_n55255_ = ~new_n55253_ & ~new_n55254_;
  assign new_n55256_ = new_n55252_ & new_n55255_;
  assign new_n55257_ = ~new_n55112_ & ~new_n55114_;
  assign new_n55258_ = new_n55120_ & new_n55257_;
  assign new_n55259_ = new_n55256_ & new_n55258_;
  assign new_n55260_ = ~new_n55249_ & ~new_n55259_;
  assign new_n55261_ = ys__n39768 & new_n53871_;
  assign new_n55262_ = ys__n39766 & new_n53870_;
  assign new_n55263_ = ~new_n55261_ & ~new_n55262_;
  assign new_n55264_ = ys__n33733 & new_n53884_;
  assign new_n55265_ = ~ys__n33733 & new_n53887_;
  assign new_n55266_ = ~new_n55264_ & ~new_n55265_;
  assign new_n55267_ = new_n55263_ & new_n55266_;
  assign new_n55268_ = ys__n24822 & new_n53876_;
  assign new_n55269_ = ys__n24819 & new_n53879_;
  assign new_n55270_ = ~new_n55268_ & ~new_n55269_;
  assign new_n55271_ = ys__n24816 & new_n53878_;
  assign new_n55272_ = ys__n39770 & new_n53868_;
  assign new_n55273_ = ~new_n55271_ & ~new_n55272_;
  assign new_n55274_ = new_n55270_ & new_n55273_;
  assign new_n55275_ = new_n55267_ & new_n55274_;
  assign new_n55276_ = ~new_n55249_ & ~new_n55275_;
  assign new_n55277_ = ~new_n55259_ & ~new_n55275_;
  assign new_n55278_ = ~new_n55276_ & ~new_n55277_;
  assign new_n55279_ = ~new_n55260_ & new_n55278_;
  assign new_n55280_ = ~new_n55234_ & ~new_n55279_;
  assign new_n55281_ = ys__n39756 & new_n53781_;
  assign new_n55282_ = ys__n39754 & new_n53780_;
  assign new_n55283_ = ~new_n55281_ & ~new_n55282_;
  assign new_n55284_ = ys__n33721 & new_n53794_;
  assign new_n55285_ = ~ys__n33721 & new_n53797_;
  assign new_n55286_ = ~new_n55284_ & ~new_n55285_;
  assign new_n55287_ = new_n55283_ & new_n55286_;
  assign new_n55288_ = ys__n24804 & new_n53786_;
  assign new_n55289_ = ys__n24801 & new_n53789_;
  assign new_n55290_ = ~new_n55288_ & ~new_n55289_;
  assign new_n55291_ = ys__n24798 & new_n53788_;
  assign new_n55292_ = ys__n39758 & new_n53778_;
  assign new_n55293_ = ~new_n55291_ & ~new_n55292_;
  assign new_n55294_ = new_n55290_ & new_n55293_;
  assign new_n55295_ = new_n55287_ & new_n55294_;
  assign new_n55296_ = ys__n39762 & new_n53756_;
  assign new_n55297_ = ys__n39760 & new_n53755_;
  assign new_n55298_ = ~new_n55296_ & ~new_n55297_;
  assign new_n55299_ = ys__n33727 & new_n53769_;
  assign new_n55300_ = ~ys__n33727 & new_n53772_;
  assign new_n55301_ = ~new_n55299_ & ~new_n55300_;
  assign new_n55302_ = new_n55298_ & new_n55301_;
  assign new_n55303_ = ys__n24813 & new_n53761_;
  assign new_n55304_ = ys__n24810 & new_n53764_;
  assign new_n55305_ = ~new_n55303_ & ~new_n55304_;
  assign new_n55306_ = ys__n24807 & new_n53763_;
  assign new_n55307_ = ys__n39764 & new_n53753_;
  assign new_n55308_ = ~new_n55306_ & ~new_n55307_;
  assign new_n55309_ = new_n55305_ & new_n55308_;
  assign new_n55310_ = new_n55302_ & new_n55309_;
  assign new_n55311_ = ~new_n55295_ & ~new_n55310_;
  assign new_n55312_ = ys__n24795 & new_n53805_;
  assign new_n55313_ = ys__n24792 & new_n53806_;
  assign new_n55314_ = ~new_n55312_ & ~new_n55313_;
  assign new_n55315_ = ys__n39752 & new_n53813_;
  assign new_n55316_ = ys__n39750 & new_n53814_;
  assign new_n55317_ = ~new_n55315_ & ~new_n55316_;
  assign new_n55318_ = new_n55314_ & new_n55317_;
  assign new_n55319_ = ~new_n55295_ & ~new_n55318_;
  assign new_n55320_ = ~new_n55310_ & ~new_n55318_;
  assign new_n55321_ = ~new_n55319_ & ~new_n55320_;
  assign new_n55322_ = ~new_n55311_ & new_n55321_;
  assign new_n55323_ = ~new_n55234_ & ~new_n55322_;
  assign new_n55324_ = ~new_n55279_ & ~new_n55322_;
  assign new_n55325_ = ~new_n55323_ & ~new_n55324_;
  assign new_n55326_ = ~new_n55280_ & new_n55325_;
  assign new_n55327_ = ~new_n55213_ & ~new_n55326_;
  assign new_n55328_ = ~new_n55223_ & ~new_n55326_;
  assign new_n55329_ = ~new_n55327_ & ~new_n55328_;
  assign ys__n42809 = new_n55224_ | ~new_n55329_;
  assign new_n55331_ = ~new_n55223_ & new_n55327_;
  assign new_n55332_ = new_n55223_ & ~new_n55326_;
  assign new_n55333_ = new_n55213_ & new_n55332_;
  assign new_n55334_ = ~new_n55223_ & new_n55326_;
  assign new_n55335_ = new_n55213_ & new_n55334_;
  assign new_n55336_ = new_n55223_ & new_n55326_;
  assign new_n55337_ = ~new_n55213_ & new_n55336_;
  assign new_n55338_ = ~new_n55335_ & ~new_n55337_;
  assign new_n55339_ = ~new_n55333_ & new_n55338_;
  assign ys__n42814 = new_n55331_ | ~new_n55339_;
  assign new_n55341_ = ~new_n55279_ & new_n55323_;
  assign new_n55342_ = new_n55279_ & ~new_n55322_;
  assign new_n55343_ = new_n55234_ & new_n55342_;
  assign new_n55344_ = ~new_n55279_ & new_n55322_;
  assign new_n55345_ = new_n55234_ & new_n55344_;
  assign new_n55346_ = new_n55279_ & new_n55322_;
  assign new_n55347_ = ~new_n55234_ & new_n55346_;
  assign new_n55348_ = ~new_n55345_ & ~new_n55347_;
  assign new_n55349_ = ~new_n55343_ & new_n55348_;
  assign new_n55350_ = ~new_n55341_ & new_n55349_;
  assign new_n55351_ = ~new_n55122_ & new_n55139_;
  assign new_n55352_ = new_n55110_ & new_n55138_;
  assign new_n55353_ = ~new_n55122_ & new_n55352_;
  assign new_n55354_ = ~new_n55351_ & ~new_n55353_;
  assign new_n55355_ = ~new_n55110_ & new_n55138_;
  assign new_n55356_ = new_n55122_ & new_n55355_;
  assign new_n55357_ = new_n55110_ & ~new_n55138_;
  assign new_n55358_ = new_n55122_ & new_n55357_;
  assign new_n55359_ = ~new_n55356_ & ~new_n55358_;
  assign new_n55360_ = new_n55354_ & new_n55359_;
  assign new_n55361_ = ~new_n55350_ & ~new_n55360_;
  assign new_n55362_ = ~new_n55310_ & new_n55319_;
  assign new_n55363_ = new_n55295_ & new_n55318_;
  assign new_n55364_ = ~new_n55310_ & new_n55363_;
  assign new_n55365_ = ~new_n55362_ & ~new_n55364_;
  assign new_n55366_ = ~new_n55295_ & new_n55318_;
  assign new_n55367_ = new_n55310_ & new_n55366_;
  assign new_n55368_ = new_n55295_ & ~new_n55318_;
  assign new_n55369_ = new_n55310_ & new_n55368_;
  assign new_n55370_ = ~new_n55367_ & ~new_n55369_;
  assign new_n55371_ = new_n55365_ & new_n55370_;
  assign new_n55372_ = ys__n39772 & new_n53834_;
  assign new_n55373_ = ys__n39770 & new_n53833_;
  assign new_n55374_ = ~new_n55372_ & ~new_n55373_;
  assign new_n55375_ = ys__n33737 & new_n53847_;
  assign new_n55376_ = ~ys__n33737 & new_n53850_;
  assign new_n55377_ = ~new_n55375_ & ~new_n55376_;
  assign new_n55378_ = new_n55374_ & new_n55377_;
  assign new_n55379_ = ys__n24828 & new_n53839_;
  assign new_n55380_ = ys__n24825 & new_n53842_;
  assign new_n55381_ = ~new_n55379_ & ~new_n55380_;
  assign new_n55382_ = ys__n24822 & new_n53841_;
  assign new_n55383_ = ys__n39774 & new_n53831_;
  assign new_n55384_ = ~new_n55382_ & ~new_n55383_;
  assign new_n55385_ = new_n55381_ & new_n55384_;
  assign new_n55386_ = new_n55378_ & new_n55385_;
  assign new_n55387_ = ys__n39778 & new_n53723_;
  assign new_n55388_ = ys__n39776 & new_n53726_;
  assign new_n55389_ = ~new_n55387_ & ~new_n55388_;
  assign new_n55390_ = ys__n33743 & new_n53730_;
  assign new_n55391_ = ~ys__n33743 & new_n53733_;
  assign new_n55392_ = ~new_n55390_ & ~new_n55391_;
  assign new_n55393_ = new_n55389_ & new_n55392_;
  assign new_n55394_ = ~new_n55112_ & ~new_n55118_;
  assign new_n55395_ = ys__n24834 & new_n53740_;
  assign new_n55396_ = ys__n24831 & new_n53744_;
  assign new_n55397_ = ~new_n55395_ & ~new_n55396_;
  assign new_n55398_ = new_n55394_ & new_n55397_;
  assign new_n55399_ = new_n55393_ & new_n55398_;
  assign new_n55400_ = ~new_n55386_ & ~new_n55399_;
  assign new_n55401_ = ys__n39766 & new_n53871_;
  assign new_n55402_ = ys__n39764 & new_n53870_;
  assign new_n55403_ = ~new_n55401_ & ~new_n55402_;
  assign new_n55404_ = ys__n33731 & new_n53884_;
  assign new_n55405_ = ~ys__n33731 & new_n53887_;
  assign new_n55406_ = ~new_n55404_ & ~new_n55405_;
  assign new_n55407_ = new_n55403_ & new_n55406_;
  assign new_n55408_ = ys__n24819 & new_n53876_;
  assign new_n55409_ = ys__n24816 & new_n53879_;
  assign new_n55410_ = ~new_n55408_ & ~new_n55409_;
  assign new_n55411_ = ys__n24813 & new_n53878_;
  assign new_n55412_ = ys__n39768 & new_n53868_;
  assign new_n55413_ = ~new_n55411_ & ~new_n55412_;
  assign new_n55414_ = new_n55410_ & new_n55413_;
  assign new_n55415_ = new_n55407_ & new_n55414_;
  assign new_n55416_ = ~new_n55386_ & ~new_n55415_;
  assign new_n55417_ = ~new_n55399_ & ~new_n55415_;
  assign new_n55418_ = ~new_n55416_ & ~new_n55417_;
  assign new_n55419_ = ~new_n55400_ & new_n55418_;
  assign new_n55420_ = ~new_n55371_ & ~new_n55419_;
  assign new_n55421_ = ys__n39754 & new_n53781_;
  assign new_n55422_ = ys__n39752 & new_n53780_;
  assign new_n55423_ = ~new_n55421_ & ~new_n55422_;
  assign new_n55424_ = ys__n33719 & new_n53794_;
  assign new_n55425_ = ~ys__n33719 & new_n53797_;
  assign new_n55426_ = ~new_n55424_ & ~new_n55425_;
  assign new_n55427_ = new_n55423_ & new_n55426_;
  assign new_n55428_ = ys__n24801 & new_n53786_;
  assign new_n55429_ = ys__n24798 & new_n53789_;
  assign new_n55430_ = ~new_n55428_ & ~new_n55429_;
  assign new_n55431_ = ys__n24795 & new_n53788_;
  assign new_n55432_ = ys__n39756 & new_n53778_;
  assign new_n55433_ = ~new_n55431_ & ~new_n55432_;
  assign new_n55434_ = new_n55430_ & new_n55433_;
  assign new_n55435_ = new_n55427_ & new_n55434_;
  assign new_n55436_ = ys__n39760 & new_n53756_;
  assign new_n55437_ = ys__n39758 & new_n53755_;
  assign new_n55438_ = ~new_n55436_ & ~new_n55437_;
  assign new_n55439_ = ys__n33725 & new_n53769_;
  assign new_n55440_ = ~ys__n33725 & new_n53772_;
  assign new_n55441_ = ~new_n55439_ & ~new_n55440_;
  assign new_n55442_ = new_n55438_ & new_n55441_;
  assign new_n55443_ = ys__n24810 & new_n53761_;
  assign new_n55444_ = ys__n24807 & new_n53764_;
  assign new_n55445_ = ~new_n55443_ & ~new_n55444_;
  assign new_n55446_ = ys__n24804 & new_n53763_;
  assign new_n55447_ = ys__n39762 & new_n53753_;
  assign new_n55448_ = ~new_n55446_ & ~new_n55447_;
  assign new_n55449_ = new_n55445_ & new_n55448_;
  assign new_n55450_ = new_n55442_ & new_n55449_;
  assign new_n55451_ = ~new_n55435_ & ~new_n55450_;
  assign new_n55452_ = ys__n24792 & new_n53805_;
  assign new_n55453_ = ys__n24789 & new_n53806_;
  assign new_n55454_ = ~new_n55452_ & ~new_n55453_;
  assign new_n55455_ = ys__n39750 & new_n53813_;
  assign new_n55456_ = ys__n39748 & new_n53814_;
  assign new_n55457_ = ~new_n55455_ & ~new_n55456_;
  assign new_n55458_ = new_n55454_ & new_n55457_;
  assign new_n55459_ = ~new_n55435_ & ~new_n55458_;
  assign new_n55460_ = ~new_n55450_ & ~new_n55458_;
  assign new_n55461_ = ~new_n55459_ & ~new_n55460_;
  assign new_n55462_ = ~new_n55451_ & new_n55461_;
  assign new_n55463_ = ~new_n55371_ & ~new_n55462_;
  assign new_n55464_ = ~new_n55419_ & ~new_n55462_;
  assign new_n55465_ = ~new_n55463_ & ~new_n55464_;
  assign new_n55466_ = ~new_n55420_ & new_n55465_;
  assign new_n55467_ = ~new_n55350_ & ~new_n55466_;
  assign new_n55468_ = ~new_n55360_ & ~new_n55466_;
  assign new_n55469_ = ~new_n55467_ & ~new_n55468_;
  assign ys__n42863 = new_n55361_ | ~new_n55469_;
  assign new_n55471_ = ~new_n55360_ & new_n55467_;
  assign new_n55472_ = new_n55360_ & ~new_n55466_;
  assign new_n55473_ = new_n55350_ & new_n55472_;
  assign new_n55474_ = ~new_n55360_ & new_n55466_;
  assign new_n55475_ = new_n55350_ & new_n55474_;
  assign new_n55476_ = new_n55360_ & new_n55466_;
  assign new_n55477_ = ~new_n55350_ & new_n55476_;
  assign new_n55478_ = ~new_n55475_ & ~new_n55477_;
  assign new_n55479_ = ~new_n55473_ & new_n55478_;
  assign ys__n42868 = new_n55471_ | ~new_n55479_;
  assign new_n55481_ = ~new_n55419_ & new_n55463_;
  assign new_n55482_ = new_n55419_ & ~new_n55462_;
  assign new_n55483_ = new_n55371_ & new_n55482_;
  assign new_n55484_ = ~new_n55419_ & new_n55462_;
  assign new_n55485_ = new_n55371_ & new_n55484_;
  assign new_n55486_ = new_n55419_ & new_n55462_;
  assign new_n55487_ = ~new_n55371_ & new_n55486_;
  assign new_n55488_ = ~new_n55485_ & ~new_n55487_;
  assign new_n55489_ = ~new_n55483_ & new_n55488_;
  assign new_n55490_ = ~new_n55481_ & new_n55489_;
  assign new_n55491_ = ~new_n55259_ & new_n55276_;
  assign new_n55492_ = new_n55249_ & new_n55275_;
  assign new_n55493_ = ~new_n55259_ & new_n55492_;
  assign new_n55494_ = ~new_n55491_ & ~new_n55493_;
  assign new_n55495_ = ~new_n55249_ & new_n55275_;
  assign new_n55496_ = new_n55259_ & new_n55495_;
  assign new_n55497_ = new_n55249_ & ~new_n55275_;
  assign new_n55498_ = new_n55259_ & new_n55497_;
  assign new_n55499_ = ~new_n55496_ & ~new_n55498_;
  assign new_n55500_ = new_n55494_ & new_n55499_;
  assign new_n55501_ = ~new_n55490_ & ~new_n55500_;
  assign new_n55502_ = ~new_n55450_ & new_n55459_;
  assign new_n55503_ = new_n55435_ & new_n55458_;
  assign new_n55504_ = ~new_n55450_ & new_n55503_;
  assign new_n55505_ = ~new_n55502_ & ~new_n55504_;
  assign new_n55506_ = ~new_n55435_ & new_n55458_;
  assign new_n55507_ = new_n55450_ & new_n55506_;
  assign new_n55508_ = new_n55435_ & ~new_n55458_;
  assign new_n55509_ = new_n55450_ & new_n55508_;
  assign new_n55510_ = ~new_n55507_ & ~new_n55509_;
  assign new_n55511_ = new_n55505_ & new_n55510_;
  assign new_n55512_ = ys__n39770 & new_n53834_;
  assign new_n55513_ = ys__n39768 & new_n53833_;
  assign new_n55514_ = ~new_n55512_ & ~new_n55513_;
  assign new_n55515_ = ys__n33735 & new_n53847_;
  assign new_n55516_ = ~ys__n33735 & new_n53850_;
  assign new_n55517_ = ~new_n55515_ & ~new_n55516_;
  assign new_n55518_ = new_n55514_ & new_n55517_;
  assign new_n55519_ = ys__n24825 & new_n53839_;
  assign new_n55520_ = ys__n24822 & new_n53842_;
  assign new_n55521_ = ~new_n55519_ & ~new_n55520_;
  assign new_n55522_ = ys__n24819 & new_n53841_;
  assign new_n55523_ = ys__n39772 & new_n53831_;
  assign new_n55524_ = ~new_n55522_ & ~new_n55523_;
  assign new_n55525_ = new_n55521_ & new_n55524_;
  assign new_n55526_ = new_n55518_ & new_n55525_;
  assign new_n55527_ = ys__n39776 & new_n53723_;
  assign new_n55528_ = ys__n39774 & new_n53726_;
  assign new_n55529_ = ~new_n55527_ & ~new_n55528_;
  assign new_n55530_ = ys__n33741 & new_n53730_;
  assign new_n55531_ = ~ys__n33741 & new_n53733_;
  assign new_n55532_ = ~new_n55530_ & ~new_n55531_;
  assign new_n55533_ = new_n55529_ & new_n55532_;
  assign new_n55534_ = ys__n24834 & new_n53738_;
  assign new_n55535_ = ys__n24831 & new_n53740_;
  assign new_n55536_ = ~new_n55534_ & ~new_n55535_;
  assign new_n55537_ = ys__n24828 & new_n53744_;
  assign new_n55538_ = ys__n39778 & new_n53746_;
  assign new_n55539_ = ~new_n55537_ & ~new_n55538_;
  assign new_n55540_ = new_n55536_ & new_n55539_;
  assign new_n55541_ = new_n55533_ & new_n55540_;
  assign new_n55542_ = ~new_n55526_ & ~new_n55541_;
  assign new_n55543_ = ys__n39764 & new_n53871_;
  assign new_n55544_ = ys__n39762 & new_n53870_;
  assign new_n55545_ = ~new_n55543_ & ~new_n55544_;
  assign new_n55546_ = ys__n33729 & new_n53884_;
  assign new_n55547_ = ~ys__n33729 & new_n53887_;
  assign new_n55548_ = ~new_n55546_ & ~new_n55547_;
  assign new_n55549_ = new_n55545_ & new_n55548_;
  assign new_n55550_ = ys__n24816 & new_n53876_;
  assign new_n55551_ = ys__n24813 & new_n53879_;
  assign new_n55552_ = ~new_n55550_ & ~new_n55551_;
  assign new_n55553_ = ys__n24810 & new_n53878_;
  assign new_n55554_ = ys__n39766 & new_n53868_;
  assign new_n55555_ = ~new_n55553_ & ~new_n55554_;
  assign new_n55556_ = new_n55552_ & new_n55555_;
  assign new_n55557_ = new_n55549_ & new_n55556_;
  assign new_n55558_ = ~new_n55526_ & ~new_n55557_;
  assign new_n55559_ = ~new_n55541_ & ~new_n55557_;
  assign new_n55560_ = ~new_n55558_ & ~new_n55559_;
  assign new_n55561_ = ~new_n55542_ & new_n55560_;
  assign new_n55562_ = ~new_n55511_ & ~new_n55561_;
  assign new_n55563_ = ys__n39752 & new_n53781_;
  assign new_n55564_ = ys__n39750 & new_n53780_;
  assign new_n55565_ = ~new_n55563_ & ~new_n55564_;
  assign new_n55566_ = ys__n33717 & new_n53794_;
  assign new_n55567_ = ~ys__n33717 & new_n53797_;
  assign new_n55568_ = ~new_n55566_ & ~new_n55567_;
  assign new_n55569_ = new_n55565_ & new_n55568_;
  assign new_n55570_ = ys__n24798 & new_n53786_;
  assign new_n55571_ = ys__n24795 & new_n53789_;
  assign new_n55572_ = ~new_n55570_ & ~new_n55571_;
  assign new_n55573_ = ys__n24792 & new_n53788_;
  assign new_n55574_ = ys__n39754 & new_n53778_;
  assign new_n55575_ = ~new_n55573_ & ~new_n55574_;
  assign new_n55576_ = new_n55572_ & new_n55575_;
  assign new_n55577_ = new_n55569_ & new_n55576_;
  assign new_n55578_ = ys__n39758 & new_n53756_;
  assign new_n55579_ = ys__n39756 & new_n53755_;
  assign new_n55580_ = ~new_n55578_ & ~new_n55579_;
  assign new_n55581_ = ys__n33723 & new_n53769_;
  assign new_n55582_ = ~ys__n33723 & new_n53772_;
  assign new_n55583_ = ~new_n55581_ & ~new_n55582_;
  assign new_n55584_ = new_n55580_ & new_n55583_;
  assign new_n55585_ = ys__n24807 & new_n53761_;
  assign new_n55586_ = ys__n24804 & new_n53764_;
  assign new_n55587_ = ~new_n55585_ & ~new_n55586_;
  assign new_n55588_ = ys__n24801 & new_n53763_;
  assign new_n55589_ = ys__n39760 & new_n53753_;
  assign new_n55590_ = ~new_n55588_ & ~new_n55589_;
  assign new_n55591_ = new_n55587_ & new_n55590_;
  assign new_n55592_ = new_n55584_ & new_n55591_;
  assign new_n55593_ = ~new_n55577_ & ~new_n55592_;
  assign new_n55594_ = ys__n24789 & new_n53805_;
  assign new_n55595_ = ys__n24786 & new_n53806_;
  assign new_n55596_ = ~new_n55594_ & ~new_n55595_;
  assign new_n55597_ = ys__n39748 & new_n53813_;
  assign new_n55598_ = ys__n39746 & new_n53814_;
  assign new_n55599_ = ~new_n55597_ & ~new_n55598_;
  assign new_n55600_ = new_n55596_ & new_n55599_;
  assign new_n55601_ = ~new_n55577_ & ~new_n55600_;
  assign new_n55602_ = ~new_n55592_ & ~new_n55600_;
  assign new_n55603_ = ~new_n55601_ & ~new_n55602_;
  assign new_n55604_ = ~new_n55593_ & new_n55603_;
  assign new_n55605_ = ~new_n55511_ & ~new_n55604_;
  assign new_n55606_ = ~new_n55561_ & ~new_n55604_;
  assign new_n55607_ = ~new_n55605_ & ~new_n55606_;
  assign new_n55608_ = ~new_n55562_ & new_n55607_;
  assign new_n55609_ = ~new_n55490_ & ~new_n55608_;
  assign new_n55610_ = ~new_n55500_ & ~new_n55608_;
  assign new_n55611_ = ~new_n55609_ & ~new_n55610_;
  assign ys__n42917 = new_n55501_ | ~new_n55611_;
  assign new_n55613_ = ~new_n55500_ & new_n55609_;
  assign new_n55614_ = new_n55500_ & ~new_n55608_;
  assign new_n55615_ = new_n55490_ & new_n55614_;
  assign new_n55616_ = ~new_n55500_ & new_n55608_;
  assign new_n55617_ = new_n55490_ & new_n55616_;
  assign new_n55618_ = new_n55500_ & new_n55608_;
  assign new_n55619_ = ~new_n55490_ & new_n55618_;
  assign new_n55620_ = ~new_n55617_ & ~new_n55619_;
  assign new_n55621_ = ~new_n55615_ & new_n55620_;
  assign ys__n42922 = new_n55613_ | ~new_n55621_;
  assign new_n55623_ = ~new_n55561_ & new_n55605_;
  assign new_n55624_ = new_n55561_ & ~new_n55604_;
  assign new_n55625_ = new_n55511_ & new_n55624_;
  assign new_n55626_ = ~new_n55561_ & new_n55604_;
  assign new_n55627_ = new_n55511_ & new_n55626_;
  assign new_n55628_ = new_n55561_ & new_n55604_;
  assign new_n55629_ = ~new_n55511_ & new_n55628_;
  assign new_n55630_ = ~new_n55627_ & ~new_n55629_;
  assign new_n55631_ = ~new_n55625_ & new_n55630_;
  assign new_n55632_ = ~new_n55623_ & new_n55631_;
  assign new_n55633_ = ~new_n55399_ & new_n55416_;
  assign new_n55634_ = new_n55386_ & new_n55415_;
  assign new_n55635_ = ~new_n55399_ & new_n55634_;
  assign new_n55636_ = ~new_n55633_ & ~new_n55635_;
  assign new_n55637_ = ~new_n55386_ & new_n55415_;
  assign new_n55638_ = new_n55399_ & new_n55637_;
  assign new_n55639_ = new_n55386_ & ~new_n55415_;
  assign new_n55640_ = new_n55399_ & new_n55639_;
  assign new_n55641_ = ~new_n55638_ & ~new_n55640_;
  assign new_n55642_ = new_n55636_ & new_n55641_;
  assign new_n55643_ = ~new_n55632_ & ~new_n55642_;
  assign new_n55644_ = ~new_n55592_ & new_n55601_;
  assign new_n55645_ = new_n55577_ & new_n55600_;
  assign new_n55646_ = ~new_n55592_ & new_n55645_;
  assign new_n55647_ = ~new_n55644_ & ~new_n55646_;
  assign new_n55648_ = ~new_n55577_ & new_n55600_;
  assign new_n55649_ = new_n55592_ & new_n55648_;
  assign new_n55650_ = new_n55577_ & ~new_n55600_;
  assign new_n55651_ = new_n55592_ & new_n55650_;
  assign new_n55652_ = ~new_n55649_ & ~new_n55651_;
  assign new_n55653_ = new_n55647_ & new_n55652_;
  assign new_n55654_ = ys__n39768 & new_n53834_;
  assign new_n55655_ = ys__n39766 & new_n53833_;
  assign new_n55656_ = ~new_n55654_ & ~new_n55655_;
  assign new_n55657_ = ys__n33733 & new_n53847_;
  assign new_n55658_ = ~ys__n33733 & new_n53850_;
  assign new_n55659_ = ~new_n55657_ & ~new_n55658_;
  assign new_n55660_ = new_n55656_ & new_n55659_;
  assign new_n55661_ = ys__n24822 & new_n53839_;
  assign new_n55662_ = ys__n24819 & new_n53842_;
  assign new_n55663_ = ~new_n55661_ & ~new_n55662_;
  assign new_n55664_ = ys__n24816 & new_n53841_;
  assign new_n55665_ = ys__n39770 & new_n53831_;
  assign new_n55666_ = ~new_n55664_ & ~new_n55665_;
  assign new_n55667_ = new_n55663_ & new_n55666_;
  assign new_n55668_ = new_n55660_ & new_n55667_;
  assign new_n55669_ = ys__n39774 & new_n53723_;
  assign new_n55670_ = ys__n39772 & new_n53726_;
  assign new_n55671_ = ~new_n55669_ & ~new_n55670_;
  assign new_n55672_ = ys__n33739 & new_n53730_;
  assign new_n55673_ = ~ys__n33739 & new_n53733_;
  assign new_n55674_ = ~new_n55672_ & ~new_n55673_;
  assign new_n55675_ = new_n55671_ & new_n55674_;
  assign new_n55676_ = ys__n24831 & new_n53738_;
  assign new_n55677_ = ys__n24828 & new_n53740_;
  assign new_n55678_ = ~new_n55676_ & ~new_n55677_;
  assign new_n55679_ = ys__n24825 & new_n53744_;
  assign new_n55680_ = ys__n39776 & new_n53746_;
  assign new_n55681_ = ~new_n55679_ & ~new_n55680_;
  assign new_n55682_ = new_n55678_ & new_n55681_;
  assign new_n55683_ = new_n55675_ & new_n55682_;
  assign new_n55684_ = ~new_n55668_ & ~new_n55683_;
  assign new_n55685_ = ys__n39762 & new_n53871_;
  assign new_n55686_ = ys__n39760 & new_n53870_;
  assign new_n55687_ = ~new_n55685_ & ~new_n55686_;
  assign new_n55688_ = ys__n33727 & new_n53884_;
  assign new_n55689_ = ~ys__n33727 & new_n53887_;
  assign new_n55690_ = ~new_n55688_ & ~new_n55689_;
  assign new_n55691_ = new_n55687_ & new_n55690_;
  assign new_n55692_ = ys__n24813 & new_n53876_;
  assign new_n55693_ = ys__n24810 & new_n53879_;
  assign new_n55694_ = ~new_n55692_ & ~new_n55693_;
  assign new_n55695_ = ys__n24807 & new_n53878_;
  assign new_n55696_ = ys__n39764 & new_n53868_;
  assign new_n55697_ = ~new_n55695_ & ~new_n55696_;
  assign new_n55698_ = new_n55694_ & new_n55697_;
  assign new_n55699_ = new_n55691_ & new_n55698_;
  assign new_n55700_ = ~new_n55668_ & ~new_n55699_;
  assign new_n55701_ = ~new_n55683_ & ~new_n55699_;
  assign new_n55702_ = ~new_n55700_ & ~new_n55701_;
  assign new_n55703_ = ~new_n55684_ & new_n55702_;
  assign new_n55704_ = ~new_n55653_ & ~new_n55703_;
  assign new_n55705_ = ys__n39750 & new_n53781_;
  assign new_n55706_ = ys__n39748 & new_n53780_;
  assign new_n55707_ = ~new_n55705_ & ~new_n55706_;
  assign new_n55708_ = ys__n33715 & new_n53794_;
  assign new_n55709_ = ~ys__n33715 & new_n53797_;
  assign new_n55710_ = ~new_n55708_ & ~new_n55709_;
  assign new_n55711_ = new_n55707_ & new_n55710_;
  assign new_n55712_ = ys__n24795 & new_n53786_;
  assign new_n55713_ = ys__n24792 & new_n53789_;
  assign new_n55714_ = ~new_n55712_ & ~new_n55713_;
  assign new_n55715_ = ys__n24789 & new_n53788_;
  assign new_n55716_ = ys__n39752 & new_n53778_;
  assign new_n55717_ = ~new_n55715_ & ~new_n55716_;
  assign new_n55718_ = new_n55714_ & new_n55717_;
  assign new_n55719_ = new_n55711_ & new_n55718_;
  assign new_n55720_ = ys__n39756 & new_n53756_;
  assign new_n55721_ = ys__n39754 & new_n53755_;
  assign new_n55722_ = ~new_n55720_ & ~new_n55721_;
  assign new_n55723_ = ys__n33721 & new_n53769_;
  assign new_n55724_ = ~ys__n33721 & new_n53772_;
  assign new_n55725_ = ~new_n55723_ & ~new_n55724_;
  assign new_n55726_ = new_n55722_ & new_n55725_;
  assign new_n55727_ = ys__n24804 & new_n53761_;
  assign new_n55728_ = ys__n24801 & new_n53764_;
  assign new_n55729_ = ~new_n55727_ & ~new_n55728_;
  assign new_n55730_ = ys__n24798 & new_n53763_;
  assign new_n55731_ = ys__n39758 & new_n53753_;
  assign new_n55732_ = ~new_n55730_ & ~new_n55731_;
  assign new_n55733_ = new_n55729_ & new_n55732_;
  assign new_n55734_ = new_n55726_ & new_n55733_;
  assign new_n55735_ = ~new_n55719_ & ~new_n55734_;
  assign new_n55736_ = ys__n24786 & new_n53805_;
  assign new_n55737_ = ys__n24783 & new_n53806_;
  assign new_n55738_ = ~new_n55736_ & ~new_n55737_;
  assign new_n55739_ = ys__n39746 & new_n53813_;
  assign new_n55740_ = ys__n39744 & new_n53814_;
  assign new_n55741_ = ~new_n55739_ & ~new_n55740_;
  assign new_n55742_ = new_n55738_ & new_n55741_;
  assign new_n55743_ = ~new_n55719_ & ~new_n55742_;
  assign new_n55744_ = ~new_n55734_ & ~new_n55742_;
  assign new_n55745_ = ~new_n55743_ & ~new_n55744_;
  assign new_n55746_ = ~new_n55735_ & new_n55745_;
  assign new_n55747_ = ~new_n55653_ & ~new_n55746_;
  assign new_n55748_ = ~new_n55703_ & ~new_n55746_;
  assign new_n55749_ = ~new_n55747_ & ~new_n55748_;
  assign new_n55750_ = ~new_n55704_ & new_n55749_;
  assign new_n55751_ = ~new_n55632_ & ~new_n55750_;
  assign new_n55752_ = ~new_n55642_ & ~new_n55750_;
  assign new_n55753_ = ~new_n55751_ & ~new_n55752_;
  assign ys__n42971 = new_n55643_ | ~new_n55753_;
  assign new_n55755_ = ~new_n55642_ & new_n55751_;
  assign new_n55756_ = new_n55642_ & ~new_n55750_;
  assign new_n55757_ = new_n55632_ & new_n55756_;
  assign new_n55758_ = ~new_n55642_ & new_n55750_;
  assign new_n55759_ = new_n55632_ & new_n55758_;
  assign new_n55760_ = new_n55642_ & new_n55750_;
  assign new_n55761_ = ~new_n55632_ & new_n55760_;
  assign new_n55762_ = ~new_n55759_ & ~new_n55761_;
  assign new_n55763_ = ~new_n55757_ & new_n55762_;
  assign ys__n42976 = new_n55755_ | ~new_n55763_;
  assign new_n55765_ = ~new_n55703_ & new_n55747_;
  assign new_n55766_ = new_n55703_ & ~new_n55746_;
  assign new_n55767_ = new_n55653_ & new_n55766_;
  assign new_n55768_ = ~new_n55703_ & new_n55746_;
  assign new_n55769_ = new_n55653_ & new_n55768_;
  assign new_n55770_ = new_n55703_ & new_n55746_;
  assign new_n55771_ = ~new_n55653_ & new_n55770_;
  assign new_n55772_ = ~new_n55769_ & ~new_n55771_;
  assign new_n55773_ = ~new_n55767_ & new_n55772_;
  assign new_n55774_ = ~new_n55765_ & new_n55773_;
  assign new_n55775_ = ~new_n55541_ & new_n55558_;
  assign new_n55776_ = new_n55526_ & new_n55557_;
  assign new_n55777_ = ~new_n55541_ & new_n55776_;
  assign new_n55778_ = ~new_n55775_ & ~new_n55777_;
  assign new_n55779_ = ~new_n55526_ & new_n55557_;
  assign new_n55780_ = new_n55541_ & new_n55779_;
  assign new_n55781_ = new_n55526_ & ~new_n55557_;
  assign new_n55782_ = new_n55541_ & new_n55781_;
  assign new_n55783_ = ~new_n55780_ & ~new_n55782_;
  assign new_n55784_ = new_n55778_ & new_n55783_;
  assign new_n55785_ = ~new_n55774_ & ~new_n55784_;
  assign new_n55786_ = ~new_n55734_ & new_n55743_;
  assign new_n55787_ = new_n55719_ & new_n55742_;
  assign new_n55788_ = ~new_n55734_ & new_n55787_;
  assign new_n55789_ = ~new_n55786_ & ~new_n55788_;
  assign new_n55790_ = ~new_n55719_ & new_n55742_;
  assign new_n55791_ = new_n55734_ & new_n55790_;
  assign new_n55792_ = new_n55719_ & ~new_n55742_;
  assign new_n55793_ = new_n55734_ & new_n55792_;
  assign new_n55794_ = ~new_n55791_ & ~new_n55793_;
  assign new_n55795_ = new_n55789_ & new_n55794_;
  assign new_n55796_ = ys__n39766 & new_n53834_;
  assign new_n55797_ = ys__n39764 & new_n53833_;
  assign new_n55798_ = ~new_n55796_ & ~new_n55797_;
  assign new_n55799_ = ys__n33731 & new_n53847_;
  assign new_n55800_ = ~ys__n33731 & new_n53850_;
  assign new_n55801_ = ~new_n55799_ & ~new_n55800_;
  assign new_n55802_ = new_n55798_ & new_n55801_;
  assign new_n55803_ = ys__n24819 & new_n53839_;
  assign new_n55804_ = ys__n24816 & new_n53842_;
  assign new_n55805_ = ~new_n55803_ & ~new_n55804_;
  assign new_n55806_ = ys__n24813 & new_n53841_;
  assign new_n55807_ = ys__n39768 & new_n53831_;
  assign new_n55808_ = ~new_n55806_ & ~new_n55807_;
  assign new_n55809_ = new_n55805_ & new_n55808_;
  assign new_n55810_ = new_n55802_ & new_n55809_;
  assign new_n55811_ = ys__n39772 & new_n53723_;
  assign new_n55812_ = ys__n39770 & new_n53726_;
  assign new_n55813_ = ~new_n55811_ & ~new_n55812_;
  assign new_n55814_ = ys__n33737 & new_n53730_;
  assign new_n55815_ = ~ys__n33737 & new_n53733_;
  assign new_n55816_ = ~new_n55814_ & ~new_n55815_;
  assign new_n55817_ = new_n55813_ & new_n55816_;
  assign new_n55818_ = ys__n24828 & new_n53738_;
  assign new_n55819_ = ys__n24825 & new_n53740_;
  assign new_n55820_ = ~new_n55818_ & ~new_n55819_;
  assign new_n55821_ = ys__n24822 & new_n53744_;
  assign new_n55822_ = ys__n39774 & new_n53746_;
  assign new_n55823_ = ~new_n55821_ & ~new_n55822_;
  assign new_n55824_ = new_n55820_ & new_n55823_;
  assign new_n55825_ = new_n55817_ & new_n55824_;
  assign new_n55826_ = ~new_n55810_ & ~new_n55825_;
  assign new_n55827_ = ys__n39760 & new_n53871_;
  assign new_n55828_ = ys__n39758 & new_n53870_;
  assign new_n55829_ = ~new_n55827_ & ~new_n55828_;
  assign new_n55830_ = ys__n33725 & new_n53884_;
  assign new_n55831_ = ~ys__n33725 & new_n53887_;
  assign new_n55832_ = ~new_n55830_ & ~new_n55831_;
  assign new_n55833_ = new_n55829_ & new_n55832_;
  assign new_n55834_ = ys__n24810 & new_n53876_;
  assign new_n55835_ = ys__n24807 & new_n53879_;
  assign new_n55836_ = ~new_n55834_ & ~new_n55835_;
  assign new_n55837_ = ys__n24804 & new_n53878_;
  assign new_n55838_ = ys__n39762 & new_n53868_;
  assign new_n55839_ = ~new_n55837_ & ~new_n55838_;
  assign new_n55840_ = new_n55836_ & new_n55839_;
  assign new_n55841_ = new_n55833_ & new_n55840_;
  assign new_n55842_ = ~new_n55810_ & ~new_n55841_;
  assign new_n55843_ = ~new_n55825_ & ~new_n55841_;
  assign new_n55844_ = ~new_n55842_ & ~new_n55843_;
  assign new_n55845_ = ~new_n55826_ & new_n55844_;
  assign new_n55846_ = ~new_n55795_ & ~new_n55845_;
  assign new_n55847_ = ys__n39748 & new_n53781_;
  assign new_n55848_ = ys__n39746 & new_n53780_;
  assign new_n55849_ = ~new_n55847_ & ~new_n55848_;
  assign new_n55850_ = ys__n33713 & new_n53794_;
  assign new_n55851_ = ~ys__n33713 & new_n53797_;
  assign new_n55852_ = ~new_n55850_ & ~new_n55851_;
  assign new_n55853_ = new_n55849_ & new_n55852_;
  assign new_n55854_ = ys__n24792 & new_n53786_;
  assign new_n55855_ = ys__n24789 & new_n53789_;
  assign new_n55856_ = ~new_n55854_ & ~new_n55855_;
  assign new_n55857_ = ys__n24786 & new_n53788_;
  assign new_n55858_ = ys__n39750 & new_n53778_;
  assign new_n55859_ = ~new_n55857_ & ~new_n55858_;
  assign new_n55860_ = new_n55856_ & new_n55859_;
  assign new_n55861_ = new_n55853_ & new_n55860_;
  assign new_n55862_ = ys__n39754 & new_n53756_;
  assign new_n55863_ = ys__n39752 & new_n53755_;
  assign new_n55864_ = ~new_n55862_ & ~new_n55863_;
  assign new_n55865_ = ys__n33719 & new_n53769_;
  assign new_n55866_ = ~ys__n33719 & new_n53772_;
  assign new_n55867_ = ~new_n55865_ & ~new_n55866_;
  assign new_n55868_ = new_n55864_ & new_n55867_;
  assign new_n55869_ = ys__n24801 & new_n53761_;
  assign new_n55870_ = ys__n24798 & new_n53764_;
  assign new_n55871_ = ~new_n55869_ & ~new_n55870_;
  assign new_n55872_ = ys__n24795 & new_n53763_;
  assign new_n55873_ = ys__n39756 & new_n53753_;
  assign new_n55874_ = ~new_n55872_ & ~new_n55873_;
  assign new_n55875_ = new_n55871_ & new_n55874_;
  assign new_n55876_ = new_n55868_ & new_n55875_;
  assign new_n55877_ = ~new_n55861_ & ~new_n55876_;
  assign new_n55878_ = ys__n24783 & new_n53805_;
  assign new_n55879_ = ys__n24780 & new_n53806_;
  assign new_n55880_ = ~new_n55878_ & ~new_n55879_;
  assign new_n55881_ = ys__n39744 & new_n53813_;
  assign new_n55882_ = ys__n39742 & new_n53814_;
  assign new_n55883_ = ~new_n55881_ & ~new_n55882_;
  assign new_n55884_ = new_n55880_ & new_n55883_;
  assign new_n55885_ = ~new_n55861_ & ~new_n55884_;
  assign new_n55886_ = ~new_n55876_ & ~new_n55884_;
  assign new_n55887_ = ~new_n55885_ & ~new_n55886_;
  assign new_n55888_ = ~new_n55877_ & new_n55887_;
  assign new_n55889_ = ~new_n55795_ & ~new_n55888_;
  assign new_n55890_ = ~new_n55845_ & ~new_n55888_;
  assign new_n55891_ = ~new_n55889_ & ~new_n55890_;
  assign new_n55892_ = ~new_n55846_ & new_n55891_;
  assign new_n55893_ = ~new_n55774_ & ~new_n55892_;
  assign new_n55894_ = ~new_n55784_ & ~new_n55892_;
  assign new_n55895_ = ~new_n55893_ & ~new_n55894_;
  assign ys__n43025 = new_n55785_ | ~new_n55895_;
  assign new_n55897_ = ~new_n55784_ & new_n55893_;
  assign new_n55898_ = new_n55784_ & ~new_n55892_;
  assign new_n55899_ = new_n55774_ & new_n55898_;
  assign new_n55900_ = ~new_n55784_ & new_n55892_;
  assign new_n55901_ = new_n55774_ & new_n55900_;
  assign new_n55902_ = new_n55784_ & new_n55892_;
  assign new_n55903_ = ~new_n55774_ & new_n55902_;
  assign new_n55904_ = ~new_n55901_ & ~new_n55903_;
  assign new_n55905_ = ~new_n55899_ & new_n55904_;
  assign ys__n43030 = new_n55897_ | ~new_n55905_;
  assign new_n55907_ = ~new_n55845_ & new_n55889_;
  assign new_n55908_ = new_n55845_ & ~new_n55888_;
  assign new_n55909_ = new_n55795_ & new_n55908_;
  assign new_n55910_ = ~new_n55845_ & new_n55888_;
  assign new_n55911_ = new_n55795_ & new_n55910_;
  assign new_n55912_ = new_n55845_ & new_n55888_;
  assign new_n55913_ = ~new_n55795_ & new_n55912_;
  assign new_n55914_ = ~new_n55911_ & ~new_n55913_;
  assign new_n55915_ = ~new_n55909_ & new_n55914_;
  assign new_n55916_ = ~new_n55907_ & new_n55915_;
  assign new_n55917_ = ~new_n55683_ & new_n55700_;
  assign new_n55918_ = new_n55668_ & new_n55699_;
  assign new_n55919_ = ~new_n55683_ & new_n55918_;
  assign new_n55920_ = ~new_n55917_ & ~new_n55919_;
  assign new_n55921_ = ~new_n55668_ & new_n55699_;
  assign new_n55922_ = new_n55683_ & new_n55921_;
  assign new_n55923_ = new_n55668_ & ~new_n55699_;
  assign new_n55924_ = new_n55683_ & new_n55923_;
  assign new_n55925_ = ~new_n55922_ & ~new_n55924_;
  assign new_n55926_ = new_n55920_ & new_n55925_;
  assign new_n55927_ = ~new_n55916_ & ~new_n55926_;
  assign new_n55928_ = ~new_n55876_ & new_n55885_;
  assign new_n55929_ = new_n55861_ & new_n55884_;
  assign new_n55930_ = ~new_n55876_ & new_n55929_;
  assign new_n55931_ = ~new_n55928_ & ~new_n55930_;
  assign new_n55932_ = ~new_n55861_ & new_n55884_;
  assign new_n55933_ = new_n55876_ & new_n55932_;
  assign new_n55934_ = new_n55861_ & ~new_n55884_;
  assign new_n55935_ = new_n55876_ & new_n55934_;
  assign new_n55936_ = ~new_n55933_ & ~new_n55935_;
  assign new_n55937_ = new_n55931_ & new_n55936_;
  assign new_n55938_ = ys__n39764 & new_n53834_;
  assign new_n55939_ = ys__n39762 & new_n53833_;
  assign new_n55940_ = ~new_n55938_ & ~new_n55939_;
  assign new_n55941_ = ys__n33729 & new_n53847_;
  assign new_n55942_ = ~ys__n33729 & new_n53850_;
  assign new_n55943_ = ~new_n55941_ & ~new_n55942_;
  assign new_n55944_ = new_n55940_ & new_n55943_;
  assign new_n55945_ = ys__n24816 & new_n53839_;
  assign new_n55946_ = ys__n24813 & new_n53842_;
  assign new_n55947_ = ~new_n55945_ & ~new_n55946_;
  assign new_n55948_ = ys__n24810 & new_n53841_;
  assign new_n55949_ = ys__n39766 & new_n53831_;
  assign new_n55950_ = ~new_n55948_ & ~new_n55949_;
  assign new_n55951_ = new_n55947_ & new_n55950_;
  assign new_n55952_ = new_n55944_ & new_n55951_;
  assign new_n55953_ = ys__n39770 & new_n53723_;
  assign new_n55954_ = ys__n39768 & new_n53726_;
  assign new_n55955_ = ~new_n55953_ & ~new_n55954_;
  assign new_n55956_ = ys__n33735 & new_n53730_;
  assign new_n55957_ = ~ys__n33735 & new_n53733_;
  assign new_n55958_ = ~new_n55956_ & ~new_n55957_;
  assign new_n55959_ = new_n55955_ & new_n55958_;
  assign new_n55960_ = ys__n24825 & new_n53738_;
  assign new_n55961_ = ys__n24822 & new_n53740_;
  assign new_n55962_ = ~new_n55960_ & ~new_n55961_;
  assign new_n55963_ = ys__n24819 & new_n53744_;
  assign new_n55964_ = ys__n39772 & new_n53746_;
  assign new_n55965_ = ~new_n55963_ & ~new_n55964_;
  assign new_n55966_ = new_n55962_ & new_n55965_;
  assign new_n55967_ = new_n55959_ & new_n55966_;
  assign new_n55968_ = ~new_n55952_ & ~new_n55967_;
  assign new_n55969_ = ys__n39758 & new_n53871_;
  assign new_n55970_ = ys__n39756 & new_n53870_;
  assign new_n55971_ = ~new_n55969_ & ~new_n55970_;
  assign new_n55972_ = ys__n33723 & new_n53884_;
  assign new_n55973_ = ~ys__n33723 & new_n53887_;
  assign new_n55974_ = ~new_n55972_ & ~new_n55973_;
  assign new_n55975_ = new_n55971_ & new_n55974_;
  assign new_n55976_ = ys__n24807 & new_n53876_;
  assign new_n55977_ = ys__n24804 & new_n53879_;
  assign new_n55978_ = ~new_n55976_ & ~new_n55977_;
  assign new_n55979_ = ys__n24801 & new_n53878_;
  assign new_n55980_ = ys__n39760 & new_n53868_;
  assign new_n55981_ = ~new_n55979_ & ~new_n55980_;
  assign new_n55982_ = new_n55978_ & new_n55981_;
  assign new_n55983_ = new_n55975_ & new_n55982_;
  assign new_n55984_ = ~new_n55952_ & ~new_n55983_;
  assign new_n55985_ = ~new_n55967_ & ~new_n55983_;
  assign new_n55986_ = ~new_n55984_ & ~new_n55985_;
  assign new_n55987_ = ~new_n55968_ & new_n55986_;
  assign new_n55988_ = ~new_n55937_ & ~new_n55987_;
  assign new_n55989_ = ys__n39746 & new_n53781_;
  assign new_n55990_ = ys__n39744 & new_n53780_;
  assign new_n55991_ = ~new_n55989_ & ~new_n55990_;
  assign new_n55992_ = ys__n33711 & new_n53794_;
  assign new_n55993_ = ~ys__n33711 & new_n53797_;
  assign new_n55994_ = ~new_n55992_ & ~new_n55993_;
  assign new_n55995_ = new_n55991_ & new_n55994_;
  assign new_n55996_ = ys__n24789 & new_n53786_;
  assign new_n55997_ = ys__n24786 & new_n53789_;
  assign new_n55998_ = ~new_n55996_ & ~new_n55997_;
  assign new_n55999_ = ys__n24783 & new_n53788_;
  assign new_n56000_ = ys__n39748 & new_n53778_;
  assign new_n56001_ = ~new_n55999_ & ~new_n56000_;
  assign new_n56002_ = new_n55998_ & new_n56001_;
  assign new_n56003_ = new_n55995_ & new_n56002_;
  assign new_n56004_ = ys__n39752 & new_n53756_;
  assign new_n56005_ = ys__n39750 & new_n53755_;
  assign new_n56006_ = ~new_n56004_ & ~new_n56005_;
  assign new_n56007_ = ys__n33717 & new_n53769_;
  assign new_n56008_ = ~ys__n33717 & new_n53772_;
  assign new_n56009_ = ~new_n56007_ & ~new_n56008_;
  assign new_n56010_ = new_n56006_ & new_n56009_;
  assign new_n56011_ = ys__n24798 & new_n53761_;
  assign new_n56012_ = ys__n24795 & new_n53764_;
  assign new_n56013_ = ~new_n56011_ & ~new_n56012_;
  assign new_n56014_ = ys__n24792 & new_n53763_;
  assign new_n56015_ = ys__n39754 & new_n53753_;
  assign new_n56016_ = ~new_n56014_ & ~new_n56015_;
  assign new_n56017_ = new_n56013_ & new_n56016_;
  assign new_n56018_ = new_n56010_ & new_n56017_;
  assign new_n56019_ = ~new_n56003_ & ~new_n56018_;
  assign new_n56020_ = ys__n24780 & new_n53805_;
  assign new_n56021_ = ys__n24777 & new_n53806_;
  assign new_n56022_ = ~new_n56020_ & ~new_n56021_;
  assign new_n56023_ = ys__n39742 & new_n53813_;
  assign new_n56024_ = ys__n39740 & new_n53814_;
  assign new_n56025_ = ~new_n56023_ & ~new_n56024_;
  assign new_n56026_ = new_n56022_ & new_n56025_;
  assign new_n56027_ = ~new_n56003_ & ~new_n56026_;
  assign new_n56028_ = ~new_n56018_ & ~new_n56026_;
  assign new_n56029_ = ~new_n56027_ & ~new_n56028_;
  assign new_n56030_ = ~new_n56019_ & new_n56029_;
  assign new_n56031_ = ~new_n55937_ & ~new_n56030_;
  assign new_n56032_ = ~new_n55987_ & ~new_n56030_;
  assign new_n56033_ = ~new_n56031_ & ~new_n56032_;
  assign new_n56034_ = ~new_n55988_ & new_n56033_;
  assign new_n56035_ = ~new_n55916_ & ~new_n56034_;
  assign new_n56036_ = ~new_n55926_ & ~new_n56034_;
  assign new_n56037_ = ~new_n56035_ & ~new_n56036_;
  assign ys__n43079 = new_n55927_ | ~new_n56037_;
  assign new_n56039_ = ~new_n55926_ & new_n56035_;
  assign new_n56040_ = new_n55926_ & ~new_n56034_;
  assign new_n56041_ = new_n55916_ & new_n56040_;
  assign new_n56042_ = ~new_n55926_ & new_n56034_;
  assign new_n56043_ = new_n55916_ & new_n56042_;
  assign new_n56044_ = new_n55926_ & new_n56034_;
  assign new_n56045_ = ~new_n55916_ & new_n56044_;
  assign new_n56046_ = ~new_n56043_ & ~new_n56045_;
  assign new_n56047_ = ~new_n56041_ & new_n56046_;
  assign ys__n43084 = new_n56039_ | ~new_n56047_;
  assign new_n56049_ = ~new_n55987_ & new_n56031_;
  assign new_n56050_ = new_n55987_ & ~new_n56030_;
  assign new_n56051_ = new_n55937_ & new_n56050_;
  assign new_n56052_ = ~new_n55987_ & new_n56030_;
  assign new_n56053_ = new_n55937_ & new_n56052_;
  assign new_n56054_ = new_n55987_ & new_n56030_;
  assign new_n56055_ = ~new_n55937_ & new_n56054_;
  assign new_n56056_ = ~new_n56053_ & ~new_n56055_;
  assign new_n56057_ = ~new_n56051_ & new_n56056_;
  assign new_n56058_ = ~new_n56049_ & new_n56057_;
  assign new_n56059_ = ~new_n55825_ & new_n55842_;
  assign new_n56060_ = new_n55810_ & new_n55841_;
  assign new_n56061_ = ~new_n55825_ & new_n56060_;
  assign new_n56062_ = ~new_n56059_ & ~new_n56061_;
  assign new_n56063_ = ~new_n55810_ & new_n55841_;
  assign new_n56064_ = new_n55825_ & new_n56063_;
  assign new_n56065_ = new_n55810_ & ~new_n55841_;
  assign new_n56066_ = new_n55825_ & new_n56065_;
  assign new_n56067_ = ~new_n56064_ & ~new_n56066_;
  assign new_n56068_ = new_n56062_ & new_n56067_;
  assign new_n56069_ = ~new_n56058_ & ~new_n56068_;
  assign new_n56070_ = ~new_n56018_ & new_n56027_;
  assign new_n56071_ = new_n56003_ & new_n56026_;
  assign new_n56072_ = ~new_n56018_ & new_n56071_;
  assign new_n56073_ = ~new_n56070_ & ~new_n56072_;
  assign new_n56074_ = ~new_n56003_ & new_n56026_;
  assign new_n56075_ = new_n56018_ & new_n56074_;
  assign new_n56076_ = new_n56003_ & ~new_n56026_;
  assign new_n56077_ = new_n56018_ & new_n56076_;
  assign new_n56078_ = ~new_n56075_ & ~new_n56077_;
  assign new_n56079_ = new_n56073_ & new_n56078_;
  assign new_n56080_ = ys__n39762 & new_n53834_;
  assign new_n56081_ = ys__n39760 & new_n53833_;
  assign new_n56082_ = ~new_n56080_ & ~new_n56081_;
  assign new_n56083_ = ys__n33727 & new_n53847_;
  assign new_n56084_ = ~ys__n33727 & new_n53850_;
  assign new_n56085_ = ~new_n56083_ & ~new_n56084_;
  assign new_n56086_ = new_n56082_ & new_n56085_;
  assign new_n56087_ = ys__n24813 & new_n53839_;
  assign new_n56088_ = ys__n24810 & new_n53842_;
  assign new_n56089_ = ~new_n56087_ & ~new_n56088_;
  assign new_n56090_ = ys__n24807 & new_n53841_;
  assign new_n56091_ = ys__n39764 & new_n53831_;
  assign new_n56092_ = ~new_n56090_ & ~new_n56091_;
  assign new_n56093_ = new_n56089_ & new_n56092_;
  assign new_n56094_ = new_n56086_ & new_n56093_;
  assign new_n56095_ = ys__n39768 & new_n53723_;
  assign new_n56096_ = ys__n39766 & new_n53726_;
  assign new_n56097_ = ~new_n56095_ & ~new_n56096_;
  assign new_n56098_ = ys__n33733 & new_n53730_;
  assign new_n56099_ = ~ys__n33733 & new_n53733_;
  assign new_n56100_ = ~new_n56098_ & ~new_n56099_;
  assign new_n56101_ = new_n56097_ & new_n56100_;
  assign new_n56102_ = ys__n24822 & new_n53738_;
  assign new_n56103_ = ys__n24819 & new_n53740_;
  assign new_n56104_ = ~new_n56102_ & ~new_n56103_;
  assign new_n56105_ = ys__n24816 & new_n53744_;
  assign new_n56106_ = ys__n39770 & new_n53746_;
  assign new_n56107_ = ~new_n56105_ & ~new_n56106_;
  assign new_n56108_ = new_n56104_ & new_n56107_;
  assign new_n56109_ = new_n56101_ & new_n56108_;
  assign new_n56110_ = ~new_n56094_ & ~new_n56109_;
  assign new_n56111_ = ys__n39756 & new_n53871_;
  assign new_n56112_ = ys__n39754 & new_n53870_;
  assign new_n56113_ = ~new_n56111_ & ~new_n56112_;
  assign new_n56114_ = ys__n33721 & new_n53884_;
  assign new_n56115_ = ~ys__n33721 & new_n53887_;
  assign new_n56116_ = ~new_n56114_ & ~new_n56115_;
  assign new_n56117_ = new_n56113_ & new_n56116_;
  assign new_n56118_ = ys__n24804 & new_n53876_;
  assign new_n56119_ = ys__n24801 & new_n53879_;
  assign new_n56120_ = ~new_n56118_ & ~new_n56119_;
  assign new_n56121_ = ys__n24798 & new_n53878_;
  assign new_n56122_ = ys__n39758 & new_n53868_;
  assign new_n56123_ = ~new_n56121_ & ~new_n56122_;
  assign new_n56124_ = new_n56120_ & new_n56123_;
  assign new_n56125_ = new_n56117_ & new_n56124_;
  assign new_n56126_ = ~new_n56094_ & ~new_n56125_;
  assign new_n56127_ = ~new_n56109_ & ~new_n56125_;
  assign new_n56128_ = ~new_n56126_ & ~new_n56127_;
  assign new_n56129_ = ~new_n56110_ & new_n56128_;
  assign new_n56130_ = ~new_n56079_ & ~new_n56129_;
  assign new_n56131_ = ys__n39744 & new_n53781_;
  assign new_n56132_ = ys__n39742 & new_n53780_;
  assign new_n56133_ = ~new_n56131_ & ~new_n56132_;
  assign new_n56134_ = ys__n33709 & new_n53794_;
  assign new_n56135_ = ~ys__n33709 & new_n53797_;
  assign new_n56136_ = ~new_n56134_ & ~new_n56135_;
  assign new_n56137_ = new_n56133_ & new_n56136_;
  assign new_n56138_ = ys__n24786 & new_n53786_;
  assign new_n56139_ = ys__n24783 & new_n53789_;
  assign new_n56140_ = ~new_n56138_ & ~new_n56139_;
  assign new_n56141_ = ys__n24780 & new_n53788_;
  assign new_n56142_ = ys__n39746 & new_n53778_;
  assign new_n56143_ = ~new_n56141_ & ~new_n56142_;
  assign new_n56144_ = new_n56140_ & new_n56143_;
  assign new_n56145_ = new_n56137_ & new_n56144_;
  assign new_n56146_ = ys__n39750 & new_n53756_;
  assign new_n56147_ = ys__n39748 & new_n53755_;
  assign new_n56148_ = ~new_n56146_ & ~new_n56147_;
  assign new_n56149_ = ys__n33715 & new_n53769_;
  assign new_n56150_ = ~ys__n33715 & new_n53772_;
  assign new_n56151_ = ~new_n56149_ & ~new_n56150_;
  assign new_n56152_ = new_n56148_ & new_n56151_;
  assign new_n56153_ = ys__n24795 & new_n53761_;
  assign new_n56154_ = ys__n24792 & new_n53764_;
  assign new_n56155_ = ~new_n56153_ & ~new_n56154_;
  assign new_n56156_ = ys__n24789 & new_n53763_;
  assign new_n56157_ = ys__n39752 & new_n53753_;
  assign new_n56158_ = ~new_n56156_ & ~new_n56157_;
  assign new_n56159_ = new_n56155_ & new_n56158_;
  assign new_n56160_ = new_n56152_ & new_n56159_;
  assign new_n56161_ = ~new_n56145_ & ~new_n56160_;
  assign new_n56162_ = ys__n24777 & new_n53805_;
  assign new_n56163_ = ys__n24774 & new_n53806_;
  assign new_n56164_ = ~new_n56162_ & ~new_n56163_;
  assign new_n56165_ = ys__n39740 & new_n53813_;
  assign new_n56166_ = ys__n39738 & new_n53814_;
  assign new_n56167_ = ~new_n56165_ & ~new_n56166_;
  assign new_n56168_ = new_n56164_ & new_n56167_;
  assign new_n56169_ = ~new_n56145_ & ~new_n56168_;
  assign new_n56170_ = ~new_n56160_ & ~new_n56168_;
  assign new_n56171_ = ~new_n56169_ & ~new_n56170_;
  assign new_n56172_ = ~new_n56161_ & new_n56171_;
  assign new_n56173_ = ~new_n56079_ & ~new_n56172_;
  assign new_n56174_ = ~new_n56129_ & ~new_n56172_;
  assign new_n56175_ = ~new_n56173_ & ~new_n56174_;
  assign new_n56176_ = ~new_n56130_ & new_n56175_;
  assign new_n56177_ = ~new_n56058_ & ~new_n56176_;
  assign new_n56178_ = ~new_n56068_ & ~new_n56176_;
  assign new_n56179_ = ~new_n56177_ & ~new_n56178_;
  assign ys__n43133 = new_n56069_ | ~new_n56179_;
  assign new_n56181_ = ~new_n56068_ & new_n56177_;
  assign new_n56182_ = new_n56068_ & ~new_n56176_;
  assign new_n56183_ = new_n56058_ & new_n56182_;
  assign new_n56184_ = ~new_n56068_ & new_n56176_;
  assign new_n56185_ = new_n56058_ & new_n56184_;
  assign new_n56186_ = new_n56068_ & new_n56176_;
  assign new_n56187_ = ~new_n56058_ & new_n56186_;
  assign new_n56188_ = ~new_n56185_ & ~new_n56187_;
  assign new_n56189_ = ~new_n56183_ & new_n56188_;
  assign ys__n43138 = new_n56181_ | ~new_n56189_;
  assign new_n56191_ = ~new_n56129_ & new_n56173_;
  assign new_n56192_ = new_n56129_ & ~new_n56172_;
  assign new_n56193_ = new_n56079_ & new_n56192_;
  assign new_n56194_ = ~new_n56129_ & new_n56172_;
  assign new_n56195_ = new_n56079_ & new_n56194_;
  assign new_n56196_ = new_n56129_ & new_n56172_;
  assign new_n56197_ = ~new_n56079_ & new_n56196_;
  assign new_n56198_ = ~new_n56195_ & ~new_n56197_;
  assign new_n56199_ = ~new_n56193_ & new_n56198_;
  assign new_n56200_ = ~new_n56191_ & new_n56199_;
  assign new_n56201_ = ~new_n55967_ & new_n55984_;
  assign new_n56202_ = new_n55952_ & new_n55983_;
  assign new_n56203_ = ~new_n55967_ & new_n56202_;
  assign new_n56204_ = ~new_n56201_ & ~new_n56203_;
  assign new_n56205_ = ~new_n55952_ & new_n55983_;
  assign new_n56206_ = new_n55967_ & new_n56205_;
  assign new_n56207_ = new_n55952_ & ~new_n55983_;
  assign new_n56208_ = new_n55967_ & new_n56207_;
  assign new_n56209_ = ~new_n56206_ & ~new_n56208_;
  assign new_n56210_ = new_n56204_ & new_n56209_;
  assign new_n56211_ = ~new_n56200_ & ~new_n56210_;
  assign new_n56212_ = ~new_n56160_ & new_n56169_;
  assign new_n56213_ = new_n56145_ & new_n56168_;
  assign new_n56214_ = ~new_n56160_ & new_n56213_;
  assign new_n56215_ = ~new_n56212_ & ~new_n56214_;
  assign new_n56216_ = ~new_n56145_ & new_n56168_;
  assign new_n56217_ = new_n56160_ & new_n56216_;
  assign new_n56218_ = new_n56145_ & ~new_n56168_;
  assign new_n56219_ = new_n56160_ & new_n56218_;
  assign new_n56220_ = ~new_n56217_ & ~new_n56219_;
  assign new_n56221_ = new_n56215_ & new_n56220_;
  assign new_n56222_ = ys__n39760 & new_n53834_;
  assign new_n56223_ = ys__n39758 & new_n53833_;
  assign new_n56224_ = ~new_n56222_ & ~new_n56223_;
  assign new_n56225_ = ys__n33725 & new_n53847_;
  assign new_n56226_ = ~ys__n33725 & new_n53850_;
  assign new_n56227_ = ~new_n56225_ & ~new_n56226_;
  assign new_n56228_ = new_n56224_ & new_n56227_;
  assign new_n56229_ = ys__n24810 & new_n53839_;
  assign new_n56230_ = ys__n24807 & new_n53842_;
  assign new_n56231_ = ~new_n56229_ & ~new_n56230_;
  assign new_n56232_ = ys__n24804 & new_n53841_;
  assign new_n56233_ = ys__n39762 & new_n53831_;
  assign new_n56234_ = ~new_n56232_ & ~new_n56233_;
  assign new_n56235_ = new_n56231_ & new_n56234_;
  assign new_n56236_ = new_n56228_ & new_n56235_;
  assign new_n56237_ = ys__n39766 & new_n53723_;
  assign new_n56238_ = ys__n39764 & new_n53726_;
  assign new_n56239_ = ~new_n56237_ & ~new_n56238_;
  assign new_n56240_ = ys__n33731 & new_n53730_;
  assign new_n56241_ = ~ys__n33731 & new_n53733_;
  assign new_n56242_ = ~new_n56240_ & ~new_n56241_;
  assign new_n56243_ = new_n56239_ & new_n56242_;
  assign new_n56244_ = ys__n24819 & new_n53738_;
  assign new_n56245_ = ys__n24816 & new_n53740_;
  assign new_n56246_ = ~new_n56244_ & ~new_n56245_;
  assign new_n56247_ = ys__n24813 & new_n53744_;
  assign new_n56248_ = ys__n39768 & new_n53746_;
  assign new_n56249_ = ~new_n56247_ & ~new_n56248_;
  assign new_n56250_ = new_n56246_ & new_n56249_;
  assign new_n56251_ = new_n56243_ & new_n56250_;
  assign new_n56252_ = ~new_n56236_ & ~new_n56251_;
  assign new_n56253_ = ys__n39754 & new_n53871_;
  assign new_n56254_ = ys__n39752 & new_n53870_;
  assign new_n56255_ = ~new_n56253_ & ~new_n56254_;
  assign new_n56256_ = ys__n33719 & new_n53884_;
  assign new_n56257_ = ~ys__n33719 & new_n53887_;
  assign new_n56258_ = ~new_n56256_ & ~new_n56257_;
  assign new_n56259_ = new_n56255_ & new_n56258_;
  assign new_n56260_ = ys__n24801 & new_n53876_;
  assign new_n56261_ = ys__n24798 & new_n53879_;
  assign new_n56262_ = ~new_n56260_ & ~new_n56261_;
  assign new_n56263_ = ys__n24795 & new_n53878_;
  assign new_n56264_ = ys__n39756 & new_n53868_;
  assign new_n56265_ = ~new_n56263_ & ~new_n56264_;
  assign new_n56266_ = new_n56262_ & new_n56265_;
  assign new_n56267_ = new_n56259_ & new_n56266_;
  assign new_n56268_ = ~new_n56236_ & ~new_n56267_;
  assign new_n56269_ = ~new_n56251_ & ~new_n56267_;
  assign new_n56270_ = ~new_n56268_ & ~new_n56269_;
  assign new_n56271_ = ~new_n56252_ & new_n56270_;
  assign new_n56272_ = ~new_n56221_ & ~new_n56271_;
  assign new_n56273_ = ys__n39742 & new_n53781_;
  assign new_n56274_ = ys__n39740 & new_n53780_;
  assign new_n56275_ = ~new_n56273_ & ~new_n56274_;
  assign new_n56276_ = ys__n33707 & new_n53794_;
  assign new_n56277_ = ~ys__n33707 & new_n53797_;
  assign new_n56278_ = ~new_n56276_ & ~new_n56277_;
  assign new_n56279_ = new_n56275_ & new_n56278_;
  assign new_n56280_ = ys__n24783 & new_n53786_;
  assign new_n56281_ = ys__n24780 & new_n53789_;
  assign new_n56282_ = ~new_n56280_ & ~new_n56281_;
  assign new_n56283_ = ys__n24777 & new_n53788_;
  assign new_n56284_ = ys__n39744 & new_n53778_;
  assign new_n56285_ = ~new_n56283_ & ~new_n56284_;
  assign new_n56286_ = new_n56282_ & new_n56285_;
  assign new_n56287_ = new_n56279_ & new_n56286_;
  assign new_n56288_ = ys__n39748 & new_n53756_;
  assign new_n56289_ = ys__n39746 & new_n53755_;
  assign new_n56290_ = ~new_n56288_ & ~new_n56289_;
  assign new_n56291_ = ys__n33713 & new_n53769_;
  assign new_n56292_ = ~ys__n33713 & new_n53772_;
  assign new_n56293_ = ~new_n56291_ & ~new_n56292_;
  assign new_n56294_ = new_n56290_ & new_n56293_;
  assign new_n56295_ = ys__n24792 & new_n53761_;
  assign new_n56296_ = ys__n24789 & new_n53764_;
  assign new_n56297_ = ~new_n56295_ & ~new_n56296_;
  assign new_n56298_ = ys__n24786 & new_n53763_;
  assign new_n56299_ = ys__n39750 & new_n53753_;
  assign new_n56300_ = ~new_n56298_ & ~new_n56299_;
  assign new_n56301_ = new_n56297_ & new_n56300_;
  assign new_n56302_ = new_n56294_ & new_n56301_;
  assign new_n56303_ = ~new_n56287_ & ~new_n56302_;
  assign new_n56304_ = ys__n24774 & new_n53805_;
  assign new_n56305_ = ys__n24771 & new_n53806_;
  assign new_n56306_ = ~new_n56304_ & ~new_n56305_;
  assign new_n56307_ = ys__n39738 & new_n53813_;
  assign new_n56308_ = ys__n39736 & new_n53814_;
  assign new_n56309_ = ~new_n56307_ & ~new_n56308_;
  assign new_n56310_ = new_n56306_ & new_n56309_;
  assign new_n56311_ = ~new_n56287_ & ~new_n56310_;
  assign new_n56312_ = ~new_n56302_ & ~new_n56310_;
  assign new_n56313_ = ~new_n56311_ & ~new_n56312_;
  assign new_n56314_ = ~new_n56303_ & new_n56313_;
  assign new_n56315_ = ~new_n56221_ & ~new_n56314_;
  assign new_n56316_ = ~new_n56271_ & ~new_n56314_;
  assign new_n56317_ = ~new_n56315_ & ~new_n56316_;
  assign new_n56318_ = ~new_n56272_ & new_n56317_;
  assign new_n56319_ = ~new_n56200_ & ~new_n56318_;
  assign new_n56320_ = ~new_n56210_ & ~new_n56318_;
  assign new_n56321_ = ~new_n56319_ & ~new_n56320_;
  assign ys__n43187 = new_n56211_ | ~new_n56321_;
  assign new_n56323_ = ~new_n56210_ & new_n56319_;
  assign new_n56324_ = new_n56210_ & ~new_n56318_;
  assign new_n56325_ = new_n56200_ & new_n56324_;
  assign new_n56326_ = ~new_n56210_ & new_n56318_;
  assign new_n56327_ = new_n56200_ & new_n56326_;
  assign new_n56328_ = new_n56210_ & new_n56318_;
  assign new_n56329_ = ~new_n56200_ & new_n56328_;
  assign new_n56330_ = ~new_n56327_ & ~new_n56329_;
  assign new_n56331_ = ~new_n56325_ & new_n56330_;
  assign ys__n43192 = new_n56323_ | ~new_n56331_;
  assign new_n56333_ = ~new_n56271_ & new_n56315_;
  assign new_n56334_ = new_n56271_ & ~new_n56314_;
  assign new_n56335_ = new_n56221_ & new_n56334_;
  assign new_n56336_ = ~new_n56271_ & new_n56314_;
  assign new_n56337_ = new_n56221_ & new_n56336_;
  assign new_n56338_ = new_n56271_ & new_n56314_;
  assign new_n56339_ = ~new_n56221_ & new_n56338_;
  assign new_n56340_ = ~new_n56337_ & ~new_n56339_;
  assign new_n56341_ = ~new_n56335_ & new_n56340_;
  assign new_n56342_ = ~new_n56333_ & new_n56341_;
  assign new_n56343_ = ~new_n56109_ & new_n56126_;
  assign new_n56344_ = new_n56094_ & new_n56125_;
  assign new_n56345_ = ~new_n56109_ & new_n56344_;
  assign new_n56346_ = ~new_n56343_ & ~new_n56345_;
  assign new_n56347_ = ~new_n56094_ & new_n56125_;
  assign new_n56348_ = new_n56109_ & new_n56347_;
  assign new_n56349_ = new_n56094_ & ~new_n56125_;
  assign new_n56350_ = new_n56109_ & new_n56349_;
  assign new_n56351_ = ~new_n56348_ & ~new_n56350_;
  assign new_n56352_ = new_n56346_ & new_n56351_;
  assign new_n56353_ = ~new_n56342_ & ~new_n56352_;
  assign new_n56354_ = ~new_n56302_ & new_n56311_;
  assign new_n56355_ = new_n56287_ & new_n56310_;
  assign new_n56356_ = ~new_n56302_ & new_n56355_;
  assign new_n56357_ = ~new_n56354_ & ~new_n56356_;
  assign new_n56358_ = ~new_n56287_ & new_n56310_;
  assign new_n56359_ = new_n56302_ & new_n56358_;
  assign new_n56360_ = new_n56287_ & ~new_n56310_;
  assign new_n56361_ = new_n56302_ & new_n56360_;
  assign new_n56362_ = ~new_n56359_ & ~new_n56361_;
  assign new_n56363_ = new_n56357_ & new_n56362_;
  assign new_n56364_ = ys__n39758 & new_n53834_;
  assign new_n56365_ = ys__n39756 & new_n53833_;
  assign new_n56366_ = ~new_n56364_ & ~new_n56365_;
  assign new_n56367_ = ys__n33723 & new_n53847_;
  assign new_n56368_ = ~ys__n33723 & new_n53850_;
  assign new_n56369_ = ~new_n56367_ & ~new_n56368_;
  assign new_n56370_ = new_n56366_ & new_n56369_;
  assign new_n56371_ = ys__n24807 & new_n53839_;
  assign new_n56372_ = ys__n24804 & new_n53842_;
  assign new_n56373_ = ~new_n56371_ & ~new_n56372_;
  assign new_n56374_ = ys__n24801 & new_n53841_;
  assign new_n56375_ = ys__n39760 & new_n53831_;
  assign new_n56376_ = ~new_n56374_ & ~new_n56375_;
  assign new_n56377_ = new_n56373_ & new_n56376_;
  assign new_n56378_ = new_n56370_ & new_n56377_;
  assign new_n56379_ = ys__n39764 & new_n53723_;
  assign new_n56380_ = ys__n39762 & new_n53726_;
  assign new_n56381_ = ~new_n56379_ & ~new_n56380_;
  assign new_n56382_ = ys__n33729 & new_n53730_;
  assign new_n56383_ = ~ys__n33729 & new_n53733_;
  assign new_n56384_ = ~new_n56382_ & ~new_n56383_;
  assign new_n56385_ = new_n56381_ & new_n56384_;
  assign new_n56386_ = ys__n24816 & new_n53738_;
  assign new_n56387_ = ys__n24813 & new_n53740_;
  assign new_n56388_ = ~new_n56386_ & ~new_n56387_;
  assign new_n56389_ = ys__n24810 & new_n53744_;
  assign new_n56390_ = ys__n39766 & new_n53746_;
  assign new_n56391_ = ~new_n56389_ & ~new_n56390_;
  assign new_n56392_ = new_n56388_ & new_n56391_;
  assign new_n56393_ = new_n56385_ & new_n56392_;
  assign new_n56394_ = ~new_n56378_ & ~new_n56393_;
  assign new_n56395_ = ys__n39752 & new_n53871_;
  assign new_n56396_ = ys__n39750 & new_n53870_;
  assign new_n56397_ = ~new_n56395_ & ~new_n56396_;
  assign new_n56398_ = ys__n33717 & new_n53884_;
  assign new_n56399_ = ~ys__n33717 & new_n53887_;
  assign new_n56400_ = ~new_n56398_ & ~new_n56399_;
  assign new_n56401_ = new_n56397_ & new_n56400_;
  assign new_n56402_ = ys__n24798 & new_n53876_;
  assign new_n56403_ = ys__n24795 & new_n53879_;
  assign new_n56404_ = ~new_n56402_ & ~new_n56403_;
  assign new_n56405_ = ys__n24792 & new_n53878_;
  assign new_n56406_ = ys__n39754 & new_n53868_;
  assign new_n56407_ = ~new_n56405_ & ~new_n56406_;
  assign new_n56408_ = new_n56404_ & new_n56407_;
  assign new_n56409_ = new_n56401_ & new_n56408_;
  assign new_n56410_ = ~new_n56378_ & ~new_n56409_;
  assign new_n56411_ = ~new_n56393_ & ~new_n56409_;
  assign new_n56412_ = ~new_n56410_ & ~new_n56411_;
  assign new_n56413_ = ~new_n56394_ & new_n56412_;
  assign new_n56414_ = ~new_n56363_ & ~new_n56413_;
  assign new_n56415_ = ys__n39740 & new_n53781_;
  assign new_n56416_ = ys__n39738 & new_n53780_;
  assign new_n56417_ = ~new_n56415_ & ~new_n56416_;
  assign new_n56418_ = ys__n33705 & new_n53794_;
  assign new_n56419_ = ~ys__n33705 & new_n53797_;
  assign new_n56420_ = ~new_n56418_ & ~new_n56419_;
  assign new_n56421_ = new_n56417_ & new_n56420_;
  assign new_n56422_ = ys__n24780 & new_n53786_;
  assign new_n56423_ = ys__n24777 & new_n53789_;
  assign new_n56424_ = ~new_n56422_ & ~new_n56423_;
  assign new_n56425_ = ys__n24774 & new_n53788_;
  assign new_n56426_ = ys__n39742 & new_n53778_;
  assign new_n56427_ = ~new_n56425_ & ~new_n56426_;
  assign new_n56428_ = new_n56424_ & new_n56427_;
  assign new_n56429_ = new_n56421_ & new_n56428_;
  assign new_n56430_ = ys__n39746 & new_n53756_;
  assign new_n56431_ = ys__n39744 & new_n53755_;
  assign new_n56432_ = ~new_n56430_ & ~new_n56431_;
  assign new_n56433_ = ys__n33711 & new_n53769_;
  assign new_n56434_ = ~ys__n33711 & new_n53772_;
  assign new_n56435_ = ~new_n56433_ & ~new_n56434_;
  assign new_n56436_ = new_n56432_ & new_n56435_;
  assign new_n56437_ = ys__n24789 & new_n53761_;
  assign new_n56438_ = ys__n24786 & new_n53764_;
  assign new_n56439_ = ~new_n56437_ & ~new_n56438_;
  assign new_n56440_ = ys__n24783 & new_n53763_;
  assign new_n56441_ = ys__n39748 & new_n53753_;
  assign new_n56442_ = ~new_n56440_ & ~new_n56441_;
  assign new_n56443_ = new_n56439_ & new_n56442_;
  assign new_n56444_ = new_n56436_ & new_n56443_;
  assign new_n56445_ = ~new_n56429_ & ~new_n56444_;
  assign new_n56446_ = ys__n24771 & new_n53805_;
  assign new_n56447_ = ys__n24768 & new_n53806_;
  assign new_n56448_ = ~new_n56446_ & ~new_n56447_;
  assign new_n56449_ = ys__n39736 & new_n53813_;
  assign new_n56450_ = ys__n39734 & new_n53814_;
  assign new_n56451_ = ~new_n56449_ & ~new_n56450_;
  assign new_n56452_ = new_n56448_ & new_n56451_;
  assign new_n56453_ = ~new_n56429_ & ~new_n56452_;
  assign new_n56454_ = ~new_n56444_ & ~new_n56452_;
  assign new_n56455_ = ~new_n56453_ & ~new_n56454_;
  assign new_n56456_ = ~new_n56445_ & new_n56455_;
  assign new_n56457_ = ~new_n56363_ & ~new_n56456_;
  assign new_n56458_ = ~new_n56413_ & ~new_n56456_;
  assign new_n56459_ = ~new_n56457_ & ~new_n56458_;
  assign new_n56460_ = ~new_n56414_ & new_n56459_;
  assign new_n56461_ = ~new_n56342_ & ~new_n56460_;
  assign new_n56462_ = ~new_n56352_ & ~new_n56460_;
  assign new_n56463_ = ~new_n56461_ & ~new_n56462_;
  assign ys__n43241 = new_n56353_ | ~new_n56463_;
  assign new_n56465_ = ~new_n56352_ & new_n56461_;
  assign new_n56466_ = new_n56352_ & ~new_n56460_;
  assign new_n56467_ = new_n56342_ & new_n56466_;
  assign new_n56468_ = ~new_n56352_ & new_n56460_;
  assign new_n56469_ = new_n56342_ & new_n56468_;
  assign new_n56470_ = new_n56352_ & new_n56460_;
  assign new_n56471_ = ~new_n56342_ & new_n56470_;
  assign new_n56472_ = ~new_n56469_ & ~new_n56471_;
  assign new_n56473_ = ~new_n56467_ & new_n56472_;
  assign ys__n43246 = new_n56465_ | ~new_n56473_;
  assign new_n56475_ = ~new_n56413_ & new_n56457_;
  assign new_n56476_ = new_n56413_ & ~new_n56456_;
  assign new_n56477_ = new_n56363_ & new_n56476_;
  assign new_n56478_ = ~new_n56413_ & new_n56456_;
  assign new_n56479_ = new_n56363_ & new_n56478_;
  assign new_n56480_ = new_n56413_ & new_n56456_;
  assign new_n56481_ = ~new_n56363_ & new_n56480_;
  assign new_n56482_ = ~new_n56479_ & ~new_n56481_;
  assign new_n56483_ = ~new_n56477_ & new_n56482_;
  assign new_n56484_ = ~new_n56475_ & new_n56483_;
  assign new_n56485_ = ~new_n56251_ & new_n56268_;
  assign new_n56486_ = new_n56236_ & new_n56267_;
  assign new_n56487_ = ~new_n56251_ & new_n56486_;
  assign new_n56488_ = ~new_n56485_ & ~new_n56487_;
  assign new_n56489_ = ~new_n56236_ & new_n56267_;
  assign new_n56490_ = new_n56251_ & new_n56489_;
  assign new_n56491_ = new_n56236_ & ~new_n56267_;
  assign new_n56492_ = new_n56251_ & new_n56491_;
  assign new_n56493_ = ~new_n56490_ & ~new_n56492_;
  assign new_n56494_ = new_n56488_ & new_n56493_;
  assign new_n56495_ = ~new_n56484_ & ~new_n56494_;
  assign new_n56496_ = ~new_n56444_ & new_n56453_;
  assign new_n56497_ = new_n56429_ & new_n56452_;
  assign new_n56498_ = ~new_n56444_ & new_n56497_;
  assign new_n56499_ = ~new_n56496_ & ~new_n56498_;
  assign new_n56500_ = ~new_n56429_ & new_n56452_;
  assign new_n56501_ = new_n56444_ & new_n56500_;
  assign new_n56502_ = new_n56429_ & ~new_n56452_;
  assign new_n56503_ = new_n56444_ & new_n56502_;
  assign new_n56504_ = ~new_n56501_ & ~new_n56503_;
  assign new_n56505_ = new_n56499_ & new_n56504_;
  assign new_n56506_ = ys__n39756 & new_n53834_;
  assign new_n56507_ = ys__n39754 & new_n53833_;
  assign new_n56508_ = ~new_n56506_ & ~new_n56507_;
  assign new_n56509_ = ys__n33721 & new_n53847_;
  assign new_n56510_ = ~ys__n33721 & new_n53850_;
  assign new_n56511_ = ~new_n56509_ & ~new_n56510_;
  assign new_n56512_ = new_n56508_ & new_n56511_;
  assign new_n56513_ = ys__n24804 & new_n53839_;
  assign new_n56514_ = ys__n24801 & new_n53842_;
  assign new_n56515_ = ~new_n56513_ & ~new_n56514_;
  assign new_n56516_ = ys__n24798 & new_n53841_;
  assign new_n56517_ = ys__n39758 & new_n53831_;
  assign new_n56518_ = ~new_n56516_ & ~new_n56517_;
  assign new_n56519_ = new_n56515_ & new_n56518_;
  assign new_n56520_ = new_n56512_ & new_n56519_;
  assign new_n56521_ = ys__n39762 & new_n53723_;
  assign new_n56522_ = ys__n39760 & new_n53726_;
  assign new_n56523_ = ~new_n56521_ & ~new_n56522_;
  assign new_n56524_ = ys__n33727 & new_n53730_;
  assign new_n56525_ = ~ys__n33727 & new_n53733_;
  assign new_n56526_ = ~new_n56524_ & ~new_n56525_;
  assign new_n56527_ = new_n56523_ & new_n56526_;
  assign new_n56528_ = ys__n24813 & new_n53738_;
  assign new_n56529_ = ys__n24810 & new_n53740_;
  assign new_n56530_ = ~new_n56528_ & ~new_n56529_;
  assign new_n56531_ = ys__n24807 & new_n53744_;
  assign new_n56532_ = ys__n39764 & new_n53746_;
  assign new_n56533_ = ~new_n56531_ & ~new_n56532_;
  assign new_n56534_ = new_n56530_ & new_n56533_;
  assign new_n56535_ = new_n56527_ & new_n56534_;
  assign new_n56536_ = ~new_n56520_ & ~new_n56535_;
  assign new_n56537_ = ys__n39750 & new_n53871_;
  assign new_n56538_ = ys__n39748 & new_n53870_;
  assign new_n56539_ = ~new_n56537_ & ~new_n56538_;
  assign new_n56540_ = ys__n33715 & new_n53884_;
  assign new_n56541_ = ~ys__n33715 & new_n53887_;
  assign new_n56542_ = ~new_n56540_ & ~new_n56541_;
  assign new_n56543_ = new_n56539_ & new_n56542_;
  assign new_n56544_ = ys__n24795 & new_n53876_;
  assign new_n56545_ = ys__n24792 & new_n53879_;
  assign new_n56546_ = ~new_n56544_ & ~new_n56545_;
  assign new_n56547_ = ys__n24789 & new_n53878_;
  assign new_n56548_ = ys__n39752 & new_n53868_;
  assign new_n56549_ = ~new_n56547_ & ~new_n56548_;
  assign new_n56550_ = new_n56546_ & new_n56549_;
  assign new_n56551_ = new_n56543_ & new_n56550_;
  assign new_n56552_ = ~new_n56520_ & ~new_n56551_;
  assign new_n56553_ = ~new_n56535_ & ~new_n56551_;
  assign new_n56554_ = ~new_n56552_ & ~new_n56553_;
  assign new_n56555_ = ~new_n56536_ & new_n56554_;
  assign new_n56556_ = ~new_n56505_ & ~new_n56555_;
  assign new_n56557_ = ys__n39738 & new_n53781_;
  assign new_n56558_ = ys__n39736 & new_n53780_;
  assign new_n56559_ = ~new_n56557_ & ~new_n56558_;
  assign new_n56560_ = ys__n33703 & new_n53794_;
  assign new_n56561_ = ~ys__n33703 & new_n53797_;
  assign new_n56562_ = ~new_n56560_ & ~new_n56561_;
  assign new_n56563_ = new_n56559_ & new_n56562_;
  assign new_n56564_ = ys__n24777 & new_n53786_;
  assign new_n56565_ = ys__n24774 & new_n53789_;
  assign new_n56566_ = ~new_n56564_ & ~new_n56565_;
  assign new_n56567_ = ys__n24771 & new_n53788_;
  assign new_n56568_ = ys__n39740 & new_n53778_;
  assign new_n56569_ = ~new_n56567_ & ~new_n56568_;
  assign new_n56570_ = new_n56566_ & new_n56569_;
  assign new_n56571_ = new_n56563_ & new_n56570_;
  assign new_n56572_ = ys__n39744 & new_n53756_;
  assign new_n56573_ = ys__n39742 & new_n53755_;
  assign new_n56574_ = ~new_n56572_ & ~new_n56573_;
  assign new_n56575_ = ys__n33709 & new_n53769_;
  assign new_n56576_ = ~ys__n33709 & new_n53772_;
  assign new_n56577_ = ~new_n56575_ & ~new_n56576_;
  assign new_n56578_ = new_n56574_ & new_n56577_;
  assign new_n56579_ = ys__n24786 & new_n53761_;
  assign new_n56580_ = ys__n24783 & new_n53764_;
  assign new_n56581_ = ~new_n56579_ & ~new_n56580_;
  assign new_n56582_ = ys__n24780 & new_n53763_;
  assign new_n56583_ = ys__n39746 & new_n53753_;
  assign new_n56584_ = ~new_n56582_ & ~new_n56583_;
  assign new_n56585_ = new_n56581_ & new_n56584_;
  assign new_n56586_ = new_n56578_ & new_n56585_;
  assign new_n56587_ = ~new_n56571_ & ~new_n56586_;
  assign new_n56588_ = ys__n24768 & new_n53805_;
  assign new_n56589_ = ys__n24765 & new_n53806_;
  assign new_n56590_ = ~new_n56588_ & ~new_n56589_;
  assign new_n56591_ = ys__n39734 & new_n53813_;
  assign new_n56592_ = ys__n39732 & new_n53814_;
  assign new_n56593_ = ~new_n56591_ & ~new_n56592_;
  assign new_n56594_ = new_n56590_ & new_n56593_;
  assign new_n56595_ = ~new_n56571_ & ~new_n56594_;
  assign new_n56596_ = ~new_n56586_ & ~new_n56594_;
  assign new_n56597_ = ~new_n56595_ & ~new_n56596_;
  assign new_n56598_ = ~new_n56587_ & new_n56597_;
  assign new_n56599_ = ~new_n56505_ & ~new_n56598_;
  assign new_n56600_ = ~new_n56555_ & ~new_n56598_;
  assign new_n56601_ = ~new_n56599_ & ~new_n56600_;
  assign new_n56602_ = ~new_n56556_ & new_n56601_;
  assign new_n56603_ = ~new_n56484_ & ~new_n56602_;
  assign new_n56604_ = ~new_n56494_ & ~new_n56602_;
  assign new_n56605_ = ~new_n56603_ & ~new_n56604_;
  assign ys__n43295 = new_n56495_ | ~new_n56605_;
  assign new_n56607_ = ~new_n56494_ & new_n56603_;
  assign new_n56608_ = new_n56494_ & ~new_n56602_;
  assign new_n56609_ = new_n56484_ & new_n56608_;
  assign new_n56610_ = ~new_n56494_ & new_n56602_;
  assign new_n56611_ = new_n56484_ & new_n56610_;
  assign new_n56612_ = new_n56494_ & new_n56602_;
  assign new_n56613_ = ~new_n56484_ & new_n56612_;
  assign new_n56614_ = ~new_n56611_ & ~new_n56613_;
  assign new_n56615_ = ~new_n56609_ & new_n56614_;
  assign ys__n43300 = new_n56607_ | ~new_n56615_;
  assign new_n56617_ = ~new_n56555_ & new_n56599_;
  assign new_n56618_ = new_n56555_ & ~new_n56598_;
  assign new_n56619_ = new_n56505_ & new_n56618_;
  assign new_n56620_ = ~new_n56555_ & new_n56598_;
  assign new_n56621_ = new_n56505_ & new_n56620_;
  assign new_n56622_ = new_n56555_ & new_n56598_;
  assign new_n56623_ = ~new_n56505_ & new_n56622_;
  assign new_n56624_ = ~new_n56621_ & ~new_n56623_;
  assign new_n56625_ = ~new_n56619_ & new_n56624_;
  assign new_n56626_ = ~new_n56617_ & new_n56625_;
  assign new_n56627_ = ~new_n56393_ & new_n56410_;
  assign new_n56628_ = new_n56378_ & new_n56409_;
  assign new_n56629_ = ~new_n56393_ & new_n56628_;
  assign new_n56630_ = ~new_n56627_ & ~new_n56629_;
  assign new_n56631_ = ~new_n56378_ & new_n56409_;
  assign new_n56632_ = new_n56393_ & new_n56631_;
  assign new_n56633_ = new_n56378_ & ~new_n56409_;
  assign new_n56634_ = new_n56393_ & new_n56633_;
  assign new_n56635_ = ~new_n56632_ & ~new_n56634_;
  assign new_n56636_ = new_n56630_ & new_n56635_;
  assign new_n56637_ = ~new_n56626_ & ~new_n56636_;
  assign new_n56638_ = ~new_n56586_ & new_n56595_;
  assign new_n56639_ = new_n56571_ & new_n56594_;
  assign new_n56640_ = ~new_n56586_ & new_n56639_;
  assign new_n56641_ = ~new_n56638_ & ~new_n56640_;
  assign new_n56642_ = ~new_n56571_ & new_n56594_;
  assign new_n56643_ = new_n56586_ & new_n56642_;
  assign new_n56644_ = new_n56571_ & ~new_n56594_;
  assign new_n56645_ = new_n56586_ & new_n56644_;
  assign new_n56646_ = ~new_n56643_ & ~new_n56645_;
  assign new_n56647_ = new_n56641_ & new_n56646_;
  assign new_n56648_ = ys__n39754 & new_n53834_;
  assign new_n56649_ = ys__n39752 & new_n53833_;
  assign new_n56650_ = ~new_n56648_ & ~new_n56649_;
  assign new_n56651_ = ys__n33719 & new_n53847_;
  assign new_n56652_ = ~ys__n33719 & new_n53850_;
  assign new_n56653_ = ~new_n56651_ & ~new_n56652_;
  assign new_n56654_ = new_n56650_ & new_n56653_;
  assign new_n56655_ = ys__n24801 & new_n53839_;
  assign new_n56656_ = ys__n24798 & new_n53842_;
  assign new_n56657_ = ~new_n56655_ & ~new_n56656_;
  assign new_n56658_ = ys__n24795 & new_n53841_;
  assign new_n56659_ = ys__n39756 & new_n53831_;
  assign new_n56660_ = ~new_n56658_ & ~new_n56659_;
  assign new_n56661_ = new_n56657_ & new_n56660_;
  assign new_n56662_ = new_n56654_ & new_n56661_;
  assign new_n56663_ = ys__n39760 & new_n53723_;
  assign new_n56664_ = ys__n39758 & new_n53726_;
  assign new_n56665_ = ~new_n56663_ & ~new_n56664_;
  assign new_n56666_ = ys__n33725 & new_n53730_;
  assign new_n56667_ = ~ys__n33725 & new_n53733_;
  assign new_n56668_ = ~new_n56666_ & ~new_n56667_;
  assign new_n56669_ = new_n56665_ & new_n56668_;
  assign new_n56670_ = ys__n24810 & new_n53738_;
  assign new_n56671_ = ys__n24807 & new_n53740_;
  assign new_n56672_ = ~new_n56670_ & ~new_n56671_;
  assign new_n56673_ = ys__n24804 & new_n53744_;
  assign new_n56674_ = ys__n39762 & new_n53746_;
  assign new_n56675_ = ~new_n56673_ & ~new_n56674_;
  assign new_n56676_ = new_n56672_ & new_n56675_;
  assign new_n56677_ = new_n56669_ & new_n56676_;
  assign new_n56678_ = ~new_n56662_ & ~new_n56677_;
  assign new_n56679_ = ys__n39748 & new_n53871_;
  assign new_n56680_ = ys__n39746 & new_n53870_;
  assign new_n56681_ = ~new_n56679_ & ~new_n56680_;
  assign new_n56682_ = ys__n33713 & new_n53884_;
  assign new_n56683_ = ~ys__n33713 & new_n53887_;
  assign new_n56684_ = ~new_n56682_ & ~new_n56683_;
  assign new_n56685_ = new_n56681_ & new_n56684_;
  assign new_n56686_ = ys__n24792 & new_n53876_;
  assign new_n56687_ = ys__n24789 & new_n53879_;
  assign new_n56688_ = ~new_n56686_ & ~new_n56687_;
  assign new_n56689_ = ys__n24786 & new_n53878_;
  assign new_n56690_ = ys__n39750 & new_n53868_;
  assign new_n56691_ = ~new_n56689_ & ~new_n56690_;
  assign new_n56692_ = new_n56688_ & new_n56691_;
  assign new_n56693_ = new_n56685_ & new_n56692_;
  assign new_n56694_ = ~new_n56662_ & ~new_n56693_;
  assign new_n56695_ = ~new_n56677_ & ~new_n56693_;
  assign new_n56696_ = ~new_n56694_ & ~new_n56695_;
  assign new_n56697_ = ~new_n56678_ & new_n56696_;
  assign new_n56698_ = ~new_n56647_ & ~new_n56697_;
  assign new_n56699_ = ys__n39736 & new_n53781_;
  assign new_n56700_ = ys__n39734 & new_n53780_;
  assign new_n56701_ = ~new_n56699_ & ~new_n56700_;
  assign new_n56702_ = ys__n33701 & new_n53794_;
  assign new_n56703_ = ~ys__n33701 & new_n53797_;
  assign new_n56704_ = ~new_n56702_ & ~new_n56703_;
  assign new_n56705_ = new_n56701_ & new_n56704_;
  assign new_n56706_ = ys__n24774 & new_n53786_;
  assign new_n56707_ = ys__n24771 & new_n53789_;
  assign new_n56708_ = ~new_n56706_ & ~new_n56707_;
  assign new_n56709_ = ys__n24768 & new_n53788_;
  assign new_n56710_ = ys__n39738 & new_n53778_;
  assign new_n56711_ = ~new_n56709_ & ~new_n56710_;
  assign new_n56712_ = new_n56708_ & new_n56711_;
  assign new_n56713_ = new_n56705_ & new_n56712_;
  assign new_n56714_ = ys__n39742 & new_n53756_;
  assign new_n56715_ = ys__n39740 & new_n53755_;
  assign new_n56716_ = ~new_n56714_ & ~new_n56715_;
  assign new_n56717_ = ys__n33707 & new_n53769_;
  assign new_n56718_ = ~ys__n33707 & new_n53772_;
  assign new_n56719_ = ~new_n56717_ & ~new_n56718_;
  assign new_n56720_ = new_n56716_ & new_n56719_;
  assign new_n56721_ = ys__n24783 & new_n53761_;
  assign new_n56722_ = ys__n24780 & new_n53764_;
  assign new_n56723_ = ~new_n56721_ & ~new_n56722_;
  assign new_n56724_ = ys__n24777 & new_n53763_;
  assign new_n56725_ = ys__n39744 & new_n53753_;
  assign new_n56726_ = ~new_n56724_ & ~new_n56725_;
  assign new_n56727_ = new_n56723_ & new_n56726_;
  assign new_n56728_ = new_n56720_ & new_n56727_;
  assign new_n56729_ = ~new_n56713_ & ~new_n56728_;
  assign new_n56730_ = ys__n24765 & new_n53805_;
  assign new_n56731_ = ys__n24762 & new_n53806_;
  assign new_n56732_ = ~new_n56730_ & ~new_n56731_;
  assign new_n56733_ = ys__n39732 & new_n53813_;
  assign new_n56734_ = ys__n39730 & new_n53814_;
  assign new_n56735_ = ~new_n56733_ & ~new_n56734_;
  assign new_n56736_ = new_n56732_ & new_n56735_;
  assign new_n56737_ = ~new_n56713_ & ~new_n56736_;
  assign new_n56738_ = ~new_n56728_ & ~new_n56736_;
  assign new_n56739_ = ~new_n56737_ & ~new_n56738_;
  assign new_n56740_ = ~new_n56729_ & new_n56739_;
  assign new_n56741_ = ~new_n56647_ & ~new_n56740_;
  assign new_n56742_ = ~new_n56697_ & ~new_n56740_;
  assign new_n56743_ = ~new_n56741_ & ~new_n56742_;
  assign new_n56744_ = ~new_n56698_ & new_n56743_;
  assign new_n56745_ = ~new_n56626_ & ~new_n56744_;
  assign new_n56746_ = ~new_n56636_ & ~new_n56744_;
  assign new_n56747_ = ~new_n56745_ & ~new_n56746_;
  assign ys__n43349 = new_n56637_ | ~new_n56747_;
  assign new_n56749_ = ~new_n56636_ & new_n56745_;
  assign new_n56750_ = new_n56636_ & ~new_n56744_;
  assign new_n56751_ = new_n56626_ & new_n56750_;
  assign new_n56752_ = ~new_n56636_ & new_n56744_;
  assign new_n56753_ = new_n56626_ & new_n56752_;
  assign new_n56754_ = new_n56636_ & new_n56744_;
  assign new_n56755_ = ~new_n56626_ & new_n56754_;
  assign new_n56756_ = ~new_n56753_ & ~new_n56755_;
  assign new_n56757_ = ~new_n56751_ & new_n56756_;
  assign ys__n43354 = new_n56749_ | ~new_n56757_;
  assign new_n56759_ = ~new_n56697_ & new_n56741_;
  assign new_n56760_ = new_n56697_ & ~new_n56740_;
  assign new_n56761_ = new_n56647_ & new_n56760_;
  assign new_n56762_ = ~new_n56697_ & new_n56740_;
  assign new_n56763_ = new_n56647_ & new_n56762_;
  assign new_n56764_ = new_n56697_ & new_n56740_;
  assign new_n56765_ = ~new_n56647_ & new_n56764_;
  assign new_n56766_ = ~new_n56763_ & ~new_n56765_;
  assign new_n56767_ = ~new_n56761_ & new_n56766_;
  assign new_n56768_ = ~new_n56759_ & new_n56767_;
  assign new_n56769_ = ~new_n56535_ & new_n56552_;
  assign new_n56770_ = new_n56520_ & new_n56551_;
  assign new_n56771_ = ~new_n56535_ & new_n56770_;
  assign new_n56772_ = ~new_n56769_ & ~new_n56771_;
  assign new_n56773_ = ~new_n56520_ & new_n56551_;
  assign new_n56774_ = new_n56535_ & new_n56773_;
  assign new_n56775_ = new_n56520_ & ~new_n56551_;
  assign new_n56776_ = new_n56535_ & new_n56775_;
  assign new_n56777_ = ~new_n56774_ & ~new_n56776_;
  assign new_n56778_ = new_n56772_ & new_n56777_;
  assign new_n56779_ = ~new_n56768_ & ~new_n56778_;
  assign new_n56780_ = ~new_n56728_ & new_n56737_;
  assign new_n56781_ = new_n56713_ & new_n56736_;
  assign new_n56782_ = ~new_n56728_ & new_n56781_;
  assign new_n56783_ = ~new_n56780_ & ~new_n56782_;
  assign new_n56784_ = ~new_n56713_ & new_n56736_;
  assign new_n56785_ = new_n56728_ & new_n56784_;
  assign new_n56786_ = new_n56713_ & ~new_n56736_;
  assign new_n56787_ = new_n56728_ & new_n56786_;
  assign new_n56788_ = ~new_n56785_ & ~new_n56787_;
  assign new_n56789_ = new_n56783_ & new_n56788_;
  assign new_n56790_ = ys__n39752 & new_n53834_;
  assign new_n56791_ = ys__n39750 & new_n53833_;
  assign new_n56792_ = ~new_n56790_ & ~new_n56791_;
  assign new_n56793_ = ys__n33717 & new_n53847_;
  assign new_n56794_ = ~ys__n33717 & new_n53850_;
  assign new_n56795_ = ~new_n56793_ & ~new_n56794_;
  assign new_n56796_ = new_n56792_ & new_n56795_;
  assign new_n56797_ = ys__n24798 & new_n53839_;
  assign new_n56798_ = ys__n24795 & new_n53842_;
  assign new_n56799_ = ~new_n56797_ & ~new_n56798_;
  assign new_n56800_ = ys__n24792 & new_n53841_;
  assign new_n56801_ = ys__n39754 & new_n53831_;
  assign new_n56802_ = ~new_n56800_ & ~new_n56801_;
  assign new_n56803_ = new_n56799_ & new_n56802_;
  assign new_n56804_ = new_n56796_ & new_n56803_;
  assign new_n56805_ = ys__n39758 & new_n53723_;
  assign new_n56806_ = ys__n39756 & new_n53726_;
  assign new_n56807_ = ~new_n56805_ & ~new_n56806_;
  assign new_n56808_ = ys__n33723 & new_n53730_;
  assign new_n56809_ = ~ys__n33723 & new_n53733_;
  assign new_n56810_ = ~new_n56808_ & ~new_n56809_;
  assign new_n56811_ = new_n56807_ & new_n56810_;
  assign new_n56812_ = ys__n24807 & new_n53738_;
  assign new_n56813_ = ys__n24804 & new_n53740_;
  assign new_n56814_ = ~new_n56812_ & ~new_n56813_;
  assign new_n56815_ = ys__n24801 & new_n53744_;
  assign new_n56816_ = ys__n39760 & new_n53746_;
  assign new_n56817_ = ~new_n56815_ & ~new_n56816_;
  assign new_n56818_ = new_n56814_ & new_n56817_;
  assign new_n56819_ = new_n56811_ & new_n56818_;
  assign new_n56820_ = ~new_n56804_ & ~new_n56819_;
  assign new_n56821_ = ys__n39746 & new_n53871_;
  assign new_n56822_ = ys__n39744 & new_n53870_;
  assign new_n56823_ = ~new_n56821_ & ~new_n56822_;
  assign new_n56824_ = ys__n33711 & new_n53884_;
  assign new_n56825_ = ~ys__n33711 & new_n53887_;
  assign new_n56826_ = ~new_n56824_ & ~new_n56825_;
  assign new_n56827_ = new_n56823_ & new_n56826_;
  assign new_n56828_ = ys__n24789 & new_n53876_;
  assign new_n56829_ = ys__n24786 & new_n53879_;
  assign new_n56830_ = ~new_n56828_ & ~new_n56829_;
  assign new_n56831_ = ys__n24783 & new_n53878_;
  assign new_n56832_ = ys__n39748 & new_n53868_;
  assign new_n56833_ = ~new_n56831_ & ~new_n56832_;
  assign new_n56834_ = new_n56830_ & new_n56833_;
  assign new_n56835_ = new_n56827_ & new_n56834_;
  assign new_n56836_ = ~new_n56804_ & ~new_n56835_;
  assign new_n56837_ = ~new_n56819_ & ~new_n56835_;
  assign new_n56838_ = ~new_n56836_ & ~new_n56837_;
  assign new_n56839_ = ~new_n56820_ & new_n56838_;
  assign new_n56840_ = ~new_n56789_ & ~new_n56839_;
  assign new_n56841_ = ys__n39734 & new_n53781_;
  assign new_n56842_ = ys__n39732 & new_n53780_;
  assign new_n56843_ = ~new_n56841_ & ~new_n56842_;
  assign new_n56844_ = ys__n33699 & new_n53794_;
  assign new_n56845_ = ~ys__n33699 & new_n53797_;
  assign new_n56846_ = ~new_n56844_ & ~new_n56845_;
  assign new_n56847_ = new_n56843_ & new_n56846_;
  assign new_n56848_ = ys__n24771 & new_n53786_;
  assign new_n56849_ = ys__n24768 & new_n53789_;
  assign new_n56850_ = ~new_n56848_ & ~new_n56849_;
  assign new_n56851_ = ys__n24765 & new_n53788_;
  assign new_n56852_ = ys__n39736 & new_n53778_;
  assign new_n56853_ = ~new_n56851_ & ~new_n56852_;
  assign new_n56854_ = new_n56850_ & new_n56853_;
  assign new_n56855_ = new_n56847_ & new_n56854_;
  assign new_n56856_ = ys__n39740 & new_n53756_;
  assign new_n56857_ = ys__n39738 & new_n53755_;
  assign new_n56858_ = ~new_n56856_ & ~new_n56857_;
  assign new_n56859_ = ys__n33705 & new_n53769_;
  assign new_n56860_ = ~ys__n33705 & new_n53772_;
  assign new_n56861_ = ~new_n56859_ & ~new_n56860_;
  assign new_n56862_ = new_n56858_ & new_n56861_;
  assign new_n56863_ = ys__n24780 & new_n53761_;
  assign new_n56864_ = ys__n24777 & new_n53764_;
  assign new_n56865_ = ~new_n56863_ & ~new_n56864_;
  assign new_n56866_ = ys__n24774 & new_n53763_;
  assign new_n56867_ = ys__n39742 & new_n53753_;
  assign new_n56868_ = ~new_n56866_ & ~new_n56867_;
  assign new_n56869_ = new_n56865_ & new_n56868_;
  assign new_n56870_ = new_n56862_ & new_n56869_;
  assign new_n56871_ = ~new_n56855_ & ~new_n56870_;
  assign new_n56872_ = ys__n24762 & new_n53805_;
  assign new_n56873_ = ys__n24759 & new_n53806_;
  assign new_n56874_ = ~new_n56872_ & ~new_n56873_;
  assign new_n56875_ = ys__n39730 & new_n53813_;
  assign new_n56876_ = ys__n39728 & new_n53814_;
  assign new_n56877_ = ~new_n56875_ & ~new_n56876_;
  assign new_n56878_ = new_n56874_ & new_n56877_;
  assign new_n56879_ = ~new_n56855_ & ~new_n56878_;
  assign new_n56880_ = ~new_n56870_ & ~new_n56878_;
  assign new_n56881_ = ~new_n56879_ & ~new_n56880_;
  assign new_n56882_ = ~new_n56871_ & new_n56881_;
  assign new_n56883_ = ~new_n56789_ & ~new_n56882_;
  assign new_n56884_ = ~new_n56839_ & ~new_n56882_;
  assign new_n56885_ = ~new_n56883_ & ~new_n56884_;
  assign new_n56886_ = ~new_n56840_ & new_n56885_;
  assign new_n56887_ = ~new_n56768_ & ~new_n56886_;
  assign new_n56888_ = ~new_n56778_ & ~new_n56886_;
  assign new_n56889_ = ~new_n56887_ & ~new_n56888_;
  assign ys__n43403 = new_n56779_ | ~new_n56889_;
  assign new_n56891_ = ~new_n56778_ & new_n56887_;
  assign new_n56892_ = new_n56778_ & ~new_n56886_;
  assign new_n56893_ = new_n56768_ & new_n56892_;
  assign new_n56894_ = ~new_n56778_ & new_n56886_;
  assign new_n56895_ = new_n56768_ & new_n56894_;
  assign new_n56896_ = new_n56778_ & new_n56886_;
  assign new_n56897_ = ~new_n56768_ & new_n56896_;
  assign new_n56898_ = ~new_n56895_ & ~new_n56897_;
  assign new_n56899_ = ~new_n56893_ & new_n56898_;
  assign ys__n43408 = new_n56891_ | ~new_n56899_;
  assign new_n56901_ = ~new_n56839_ & new_n56883_;
  assign new_n56902_ = new_n56839_ & ~new_n56882_;
  assign new_n56903_ = new_n56789_ & new_n56902_;
  assign new_n56904_ = ~new_n56839_ & new_n56882_;
  assign new_n56905_ = new_n56789_ & new_n56904_;
  assign new_n56906_ = new_n56839_ & new_n56882_;
  assign new_n56907_ = ~new_n56789_ & new_n56906_;
  assign new_n56908_ = ~new_n56905_ & ~new_n56907_;
  assign new_n56909_ = ~new_n56903_ & new_n56908_;
  assign new_n56910_ = ~new_n56901_ & new_n56909_;
  assign new_n56911_ = ~new_n56677_ & new_n56694_;
  assign new_n56912_ = new_n56662_ & new_n56693_;
  assign new_n56913_ = ~new_n56677_ & new_n56912_;
  assign new_n56914_ = ~new_n56911_ & ~new_n56913_;
  assign new_n56915_ = ~new_n56662_ & new_n56693_;
  assign new_n56916_ = new_n56677_ & new_n56915_;
  assign new_n56917_ = new_n56662_ & ~new_n56693_;
  assign new_n56918_ = new_n56677_ & new_n56917_;
  assign new_n56919_ = ~new_n56916_ & ~new_n56918_;
  assign new_n56920_ = new_n56914_ & new_n56919_;
  assign new_n56921_ = ~new_n56910_ & ~new_n56920_;
  assign new_n56922_ = ~new_n56870_ & new_n56879_;
  assign new_n56923_ = new_n56855_ & new_n56878_;
  assign new_n56924_ = ~new_n56870_ & new_n56923_;
  assign new_n56925_ = ~new_n56922_ & ~new_n56924_;
  assign new_n56926_ = ~new_n56855_ & new_n56878_;
  assign new_n56927_ = new_n56870_ & new_n56926_;
  assign new_n56928_ = new_n56855_ & ~new_n56878_;
  assign new_n56929_ = new_n56870_ & new_n56928_;
  assign new_n56930_ = ~new_n56927_ & ~new_n56929_;
  assign new_n56931_ = new_n56925_ & new_n56930_;
  assign new_n56932_ = ys__n39750 & new_n53834_;
  assign new_n56933_ = ys__n39748 & new_n53833_;
  assign new_n56934_ = ~new_n56932_ & ~new_n56933_;
  assign new_n56935_ = ys__n33715 & new_n53847_;
  assign new_n56936_ = ~ys__n33715 & new_n53850_;
  assign new_n56937_ = ~new_n56935_ & ~new_n56936_;
  assign new_n56938_ = new_n56934_ & new_n56937_;
  assign new_n56939_ = ys__n24795 & new_n53839_;
  assign new_n56940_ = ys__n24792 & new_n53842_;
  assign new_n56941_ = ~new_n56939_ & ~new_n56940_;
  assign new_n56942_ = ys__n24789 & new_n53841_;
  assign new_n56943_ = ys__n39752 & new_n53831_;
  assign new_n56944_ = ~new_n56942_ & ~new_n56943_;
  assign new_n56945_ = new_n56941_ & new_n56944_;
  assign new_n56946_ = new_n56938_ & new_n56945_;
  assign new_n56947_ = ys__n39756 & new_n53723_;
  assign new_n56948_ = ys__n39754 & new_n53726_;
  assign new_n56949_ = ~new_n56947_ & ~new_n56948_;
  assign new_n56950_ = ys__n33721 & new_n53730_;
  assign new_n56951_ = ~ys__n33721 & new_n53733_;
  assign new_n56952_ = ~new_n56950_ & ~new_n56951_;
  assign new_n56953_ = new_n56949_ & new_n56952_;
  assign new_n56954_ = ys__n24804 & new_n53738_;
  assign new_n56955_ = ys__n24801 & new_n53740_;
  assign new_n56956_ = ~new_n56954_ & ~new_n56955_;
  assign new_n56957_ = ys__n24798 & new_n53744_;
  assign new_n56958_ = ys__n39758 & new_n53746_;
  assign new_n56959_ = ~new_n56957_ & ~new_n56958_;
  assign new_n56960_ = new_n56956_ & new_n56959_;
  assign new_n56961_ = new_n56953_ & new_n56960_;
  assign new_n56962_ = ~new_n56946_ & ~new_n56961_;
  assign new_n56963_ = ys__n39744 & new_n53871_;
  assign new_n56964_ = ys__n39742 & new_n53870_;
  assign new_n56965_ = ~new_n56963_ & ~new_n56964_;
  assign new_n56966_ = ys__n33709 & new_n53884_;
  assign new_n56967_ = ~ys__n33709 & new_n53887_;
  assign new_n56968_ = ~new_n56966_ & ~new_n56967_;
  assign new_n56969_ = new_n56965_ & new_n56968_;
  assign new_n56970_ = ys__n24786 & new_n53876_;
  assign new_n56971_ = ys__n24783 & new_n53879_;
  assign new_n56972_ = ~new_n56970_ & ~new_n56971_;
  assign new_n56973_ = ys__n24780 & new_n53878_;
  assign new_n56974_ = ys__n39746 & new_n53868_;
  assign new_n56975_ = ~new_n56973_ & ~new_n56974_;
  assign new_n56976_ = new_n56972_ & new_n56975_;
  assign new_n56977_ = new_n56969_ & new_n56976_;
  assign new_n56978_ = ~new_n56946_ & ~new_n56977_;
  assign new_n56979_ = ~new_n56961_ & ~new_n56977_;
  assign new_n56980_ = ~new_n56978_ & ~new_n56979_;
  assign new_n56981_ = ~new_n56962_ & new_n56980_;
  assign new_n56982_ = ~new_n56931_ & ~new_n56981_;
  assign new_n56983_ = ys__n39732 & new_n53781_;
  assign new_n56984_ = ys__n39730 & new_n53780_;
  assign new_n56985_ = ~new_n56983_ & ~new_n56984_;
  assign new_n56986_ = ys__n33697 & new_n53794_;
  assign new_n56987_ = ~ys__n33697 & new_n53797_;
  assign new_n56988_ = ~new_n56986_ & ~new_n56987_;
  assign new_n56989_ = new_n56985_ & new_n56988_;
  assign new_n56990_ = ys__n24768 & new_n53786_;
  assign new_n56991_ = ys__n24765 & new_n53789_;
  assign new_n56992_ = ~new_n56990_ & ~new_n56991_;
  assign new_n56993_ = ys__n24762 & new_n53788_;
  assign new_n56994_ = ys__n39734 & new_n53778_;
  assign new_n56995_ = ~new_n56993_ & ~new_n56994_;
  assign new_n56996_ = new_n56992_ & new_n56995_;
  assign new_n56997_ = new_n56989_ & new_n56996_;
  assign new_n56998_ = ys__n39738 & new_n53756_;
  assign new_n56999_ = ys__n39736 & new_n53755_;
  assign new_n57000_ = ~new_n56998_ & ~new_n56999_;
  assign new_n57001_ = ys__n33703 & new_n53769_;
  assign new_n57002_ = ~ys__n33703 & new_n53772_;
  assign new_n57003_ = ~new_n57001_ & ~new_n57002_;
  assign new_n57004_ = new_n57000_ & new_n57003_;
  assign new_n57005_ = ys__n24777 & new_n53761_;
  assign new_n57006_ = ys__n24774 & new_n53764_;
  assign new_n57007_ = ~new_n57005_ & ~new_n57006_;
  assign new_n57008_ = ys__n24771 & new_n53763_;
  assign new_n57009_ = ys__n39740 & new_n53753_;
  assign new_n57010_ = ~new_n57008_ & ~new_n57009_;
  assign new_n57011_ = new_n57007_ & new_n57010_;
  assign new_n57012_ = new_n57004_ & new_n57011_;
  assign new_n57013_ = ~new_n56997_ & ~new_n57012_;
  assign new_n57014_ = ys__n24759 & new_n53805_;
  assign new_n57015_ = ys__n24756 & new_n53806_;
  assign new_n57016_ = ~new_n57014_ & ~new_n57015_;
  assign new_n57017_ = ys__n39728 & new_n53813_;
  assign new_n57018_ = ys__n39726 & new_n53814_;
  assign new_n57019_ = ~new_n57017_ & ~new_n57018_;
  assign new_n57020_ = new_n57016_ & new_n57019_;
  assign new_n57021_ = ~new_n56997_ & ~new_n57020_;
  assign new_n57022_ = ~new_n57012_ & ~new_n57020_;
  assign new_n57023_ = ~new_n57021_ & ~new_n57022_;
  assign new_n57024_ = ~new_n57013_ & new_n57023_;
  assign new_n57025_ = ~new_n56931_ & ~new_n57024_;
  assign new_n57026_ = ~new_n56981_ & ~new_n57024_;
  assign new_n57027_ = ~new_n57025_ & ~new_n57026_;
  assign new_n57028_ = ~new_n56982_ & new_n57027_;
  assign new_n57029_ = ~new_n56910_ & ~new_n57028_;
  assign new_n57030_ = ~new_n56920_ & ~new_n57028_;
  assign new_n57031_ = ~new_n57029_ & ~new_n57030_;
  assign ys__n43457 = new_n56921_ | ~new_n57031_;
  assign new_n57033_ = ~new_n56920_ & new_n57029_;
  assign new_n57034_ = new_n56920_ & ~new_n57028_;
  assign new_n57035_ = new_n56910_ & new_n57034_;
  assign new_n57036_ = ~new_n56920_ & new_n57028_;
  assign new_n57037_ = new_n56910_ & new_n57036_;
  assign new_n57038_ = new_n56920_ & new_n57028_;
  assign new_n57039_ = ~new_n56910_ & new_n57038_;
  assign new_n57040_ = ~new_n57037_ & ~new_n57039_;
  assign new_n57041_ = ~new_n57035_ & new_n57040_;
  assign ys__n43462 = new_n57033_ | ~new_n57041_;
  assign new_n57043_ = ~new_n56981_ & new_n57025_;
  assign new_n57044_ = new_n56981_ & ~new_n57024_;
  assign new_n57045_ = new_n56931_ & new_n57044_;
  assign new_n57046_ = ~new_n56981_ & new_n57024_;
  assign new_n57047_ = new_n56931_ & new_n57046_;
  assign new_n57048_ = new_n56981_ & new_n57024_;
  assign new_n57049_ = ~new_n56931_ & new_n57048_;
  assign new_n57050_ = ~new_n57047_ & ~new_n57049_;
  assign new_n57051_ = ~new_n57045_ & new_n57050_;
  assign new_n57052_ = ~new_n57043_ & new_n57051_;
  assign new_n57053_ = ~new_n56819_ & new_n56836_;
  assign new_n57054_ = new_n56804_ & new_n56835_;
  assign new_n57055_ = ~new_n56819_ & new_n57054_;
  assign new_n57056_ = ~new_n57053_ & ~new_n57055_;
  assign new_n57057_ = ~new_n56804_ & new_n56835_;
  assign new_n57058_ = new_n56819_ & new_n57057_;
  assign new_n57059_ = new_n56804_ & ~new_n56835_;
  assign new_n57060_ = new_n56819_ & new_n57059_;
  assign new_n57061_ = ~new_n57058_ & ~new_n57060_;
  assign new_n57062_ = new_n57056_ & new_n57061_;
  assign new_n57063_ = ~new_n57052_ & ~new_n57062_;
  assign new_n57064_ = ~new_n57012_ & new_n57021_;
  assign new_n57065_ = new_n56997_ & new_n57020_;
  assign new_n57066_ = ~new_n57012_ & new_n57065_;
  assign new_n57067_ = ~new_n57064_ & ~new_n57066_;
  assign new_n57068_ = ~new_n56997_ & new_n57020_;
  assign new_n57069_ = new_n57012_ & new_n57068_;
  assign new_n57070_ = new_n56997_ & ~new_n57020_;
  assign new_n57071_ = new_n57012_ & new_n57070_;
  assign new_n57072_ = ~new_n57069_ & ~new_n57071_;
  assign new_n57073_ = new_n57067_ & new_n57072_;
  assign new_n57074_ = ys__n39748 & new_n53834_;
  assign new_n57075_ = ys__n39746 & new_n53833_;
  assign new_n57076_ = ~new_n57074_ & ~new_n57075_;
  assign new_n57077_ = ys__n33713 & new_n53847_;
  assign new_n57078_ = ~ys__n33713 & new_n53850_;
  assign new_n57079_ = ~new_n57077_ & ~new_n57078_;
  assign new_n57080_ = new_n57076_ & new_n57079_;
  assign new_n57081_ = ys__n24792 & new_n53839_;
  assign new_n57082_ = ys__n24789 & new_n53842_;
  assign new_n57083_ = ~new_n57081_ & ~new_n57082_;
  assign new_n57084_ = ys__n24786 & new_n53841_;
  assign new_n57085_ = ys__n39750 & new_n53831_;
  assign new_n57086_ = ~new_n57084_ & ~new_n57085_;
  assign new_n57087_ = new_n57083_ & new_n57086_;
  assign new_n57088_ = new_n57080_ & new_n57087_;
  assign new_n57089_ = ys__n39754 & new_n53723_;
  assign new_n57090_ = ys__n39752 & new_n53726_;
  assign new_n57091_ = ~new_n57089_ & ~new_n57090_;
  assign new_n57092_ = ys__n33719 & new_n53730_;
  assign new_n57093_ = ~ys__n33719 & new_n53733_;
  assign new_n57094_ = ~new_n57092_ & ~new_n57093_;
  assign new_n57095_ = new_n57091_ & new_n57094_;
  assign new_n57096_ = ys__n24801 & new_n53738_;
  assign new_n57097_ = ys__n24798 & new_n53740_;
  assign new_n57098_ = ~new_n57096_ & ~new_n57097_;
  assign new_n57099_ = ys__n24795 & new_n53744_;
  assign new_n57100_ = ys__n39756 & new_n53746_;
  assign new_n57101_ = ~new_n57099_ & ~new_n57100_;
  assign new_n57102_ = new_n57098_ & new_n57101_;
  assign new_n57103_ = new_n57095_ & new_n57102_;
  assign new_n57104_ = ~new_n57088_ & ~new_n57103_;
  assign new_n57105_ = ys__n39742 & new_n53871_;
  assign new_n57106_ = ys__n39740 & new_n53870_;
  assign new_n57107_ = ~new_n57105_ & ~new_n57106_;
  assign new_n57108_ = ys__n33707 & new_n53884_;
  assign new_n57109_ = ~ys__n33707 & new_n53887_;
  assign new_n57110_ = ~new_n57108_ & ~new_n57109_;
  assign new_n57111_ = new_n57107_ & new_n57110_;
  assign new_n57112_ = ys__n24783 & new_n53876_;
  assign new_n57113_ = ys__n24780 & new_n53879_;
  assign new_n57114_ = ~new_n57112_ & ~new_n57113_;
  assign new_n57115_ = ys__n24777 & new_n53878_;
  assign new_n57116_ = ys__n39744 & new_n53868_;
  assign new_n57117_ = ~new_n57115_ & ~new_n57116_;
  assign new_n57118_ = new_n57114_ & new_n57117_;
  assign new_n57119_ = new_n57111_ & new_n57118_;
  assign new_n57120_ = ~new_n57088_ & ~new_n57119_;
  assign new_n57121_ = ~new_n57103_ & ~new_n57119_;
  assign new_n57122_ = ~new_n57120_ & ~new_n57121_;
  assign new_n57123_ = ~new_n57104_ & new_n57122_;
  assign new_n57124_ = ~new_n57073_ & ~new_n57123_;
  assign new_n57125_ = ys__n39730 & new_n53781_;
  assign new_n57126_ = ys__n39728 & new_n53780_;
  assign new_n57127_ = ~new_n57125_ & ~new_n57126_;
  assign new_n57128_ = ys__n33695 & new_n53794_;
  assign new_n57129_ = ~ys__n33695 & new_n53797_;
  assign new_n57130_ = ~new_n57128_ & ~new_n57129_;
  assign new_n57131_ = new_n57127_ & new_n57130_;
  assign new_n57132_ = ys__n24765 & new_n53786_;
  assign new_n57133_ = ys__n24762 & new_n53789_;
  assign new_n57134_ = ~new_n57132_ & ~new_n57133_;
  assign new_n57135_ = ys__n24759 & new_n53788_;
  assign new_n57136_ = ys__n39732 & new_n53778_;
  assign new_n57137_ = ~new_n57135_ & ~new_n57136_;
  assign new_n57138_ = new_n57134_ & new_n57137_;
  assign new_n57139_ = new_n57131_ & new_n57138_;
  assign new_n57140_ = ys__n39736 & new_n53756_;
  assign new_n57141_ = ys__n39734 & new_n53755_;
  assign new_n57142_ = ~new_n57140_ & ~new_n57141_;
  assign new_n57143_ = ys__n33701 & new_n53769_;
  assign new_n57144_ = ~ys__n33701 & new_n53772_;
  assign new_n57145_ = ~new_n57143_ & ~new_n57144_;
  assign new_n57146_ = new_n57142_ & new_n57145_;
  assign new_n57147_ = ys__n24774 & new_n53761_;
  assign new_n57148_ = ys__n24771 & new_n53764_;
  assign new_n57149_ = ~new_n57147_ & ~new_n57148_;
  assign new_n57150_ = ys__n24768 & new_n53763_;
  assign new_n57151_ = ys__n39738 & new_n53753_;
  assign new_n57152_ = ~new_n57150_ & ~new_n57151_;
  assign new_n57153_ = new_n57149_ & new_n57152_;
  assign new_n57154_ = new_n57146_ & new_n57153_;
  assign new_n57155_ = ~new_n57139_ & ~new_n57154_;
  assign new_n57156_ = ys__n24756 & new_n53805_;
  assign new_n57157_ = ys__n24753 & new_n53806_;
  assign new_n57158_ = ~new_n57156_ & ~new_n57157_;
  assign new_n57159_ = ys__n39726 & new_n53813_;
  assign new_n57160_ = ys__n39724 & new_n53814_;
  assign new_n57161_ = ~new_n57159_ & ~new_n57160_;
  assign new_n57162_ = new_n57158_ & new_n57161_;
  assign new_n57163_ = ~new_n57139_ & ~new_n57162_;
  assign new_n57164_ = ~new_n57154_ & ~new_n57162_;
  assign new_n57165_ = ~new_n57163_ & ~new_n57164_;
  assign new_n57166_ = ~new_n57155_ & new_n57165_;
  assign new_n57167_ = ~new_n57073_ & ~new_n57166_;
  assign new_n57168_ = ~new_n57123_ & ~new_n57166_;
  assign new_n57169_ = ~new_n57167_ & ~new_n57168_;
  assign new_n57170_ = ~new_n57124_ & new_n57169_;
  assign new_n57171_ = ~new_n57052_ & ~new_n57170_;
  assign new_n57172_ = ~new_n57062_ & ~new_n57170_;
  assign new_n57173_ = ~new_n57171_ & ~new_n57172_;
  assign ys__n43511 = new_n57063_ | ~new_n57173_;
  assign new_n57175_ = ~new_n57062_ & new_n57171_;
  assign new_n57176_ = new_n57062_ & ~new_n57170_;
  assign new_n57177_ = new_n57052_ & new_n57176_;
  assign new_n57178_ = ~new_n57062_ & new_n57170_;
  assign new_n57179_ = new_n57052_ & new_n57178_;
  assign new_n57180_ = new_n57062_ & new_n57170_;
  assign new_n57181_ = ~new_n57052_ & new_n57180_;
  assign new_n57182_ = ~new_n57179_ & ~new_n57181_;
  assign new_n57183_ = ~new_n57177_ & new_n57182_;
  assign ys__n43516 = new_n57175_ | ~new_n57183_;
  assign new_n57185_ = ~new_n57123_ & new_n57167_;
  assign new_n57186_ = new_n57123_ & ~new_n57166_;
  assign new_n57187_ = new_n57073_ & new_n57186_;
  assign new_n57188_ = ~new_n57123_ & new_n57166_;
  assign new_n57189_ = new_n57073_ & new_n57188_;
  assign new_n57190_ = new_n57123_ & new_n57166_;
  assign new_n57191_ = ~new_n57073_ & new_n57190_;
  assign new_n57192_ = ~new_n57189_ & ~new_n57191_;
  assign new_n57193_ = ~new_n57187_ & new_n57192_;
  assign new_n57194_ = ~new_n57185_ & new_n57193_;
  assign new_n57195_ = ~new_n56961_ & new_n56978_;
  assign new_n57196_ = new_n56946_ & new_n56977_;
  assign new_n57197_ = ~new_n56961_ & new_n57196_;
  assign new_n57198_ = ~new_n57195_ & ~new_n57197_;
  assign new_n57199_ = ~new_n56946_ & new_n56977_;
  assign new_n57200_ = new_n56961_ & new_n57199_;
  assign new_n57201_ = new_n56946_ & ~new_n56977_;
  assign new_n57202_ = new_n56961_ & new_n57201_;
  assign new_n57203_ = ~new_n57200_ & ~new_n57202_;
  assign new_n57204_ = new_n57198_ & new_n57203_;
  assign new_n57205_ = ~new_n57194_ & ~new_n57204_;
  assign new_n57206_ = ~new_n57154_ & new_n57163_;
  assign new_n57207_ = new_n57139_ & new_n57162_;
  assign new_n57208_ = ~new_n57154_ & new_n57207_;
  assign new_n57209_ = ~new_n57206_ & ~new_n57208_;
  assign new_n57210_ = ~new_n57139_ & new_n57162_;
  assign new_n57211_ = new_n57154_ & new_n57210_;
  assign new_n57212_ = new_n57139_ & ~new_n57162_;
  assign new_n57213_ = new_n57154_ & new_n57212_;
  assign new_n57214_ = ~new_n57211_ & ~new_n57213_;
  assign new_n57215_ = new_n57209_ & new_n57214_;
  assign new_n57216_ = ys__n39746 & new_n53834_;
  assign new_n57217_ = ys__n39744 & new_n53833_;
  assign new_n57218_ = ~new_n57216_ & ~new_n57217_;
  assign new_n57219_ = ys__n33711 & new_n53847_;
  assign new_n57220_ = ~ys__n33711 & new_n53850_;
  assign new_n57221_ = ~new_n57219_ & ~new_n57220_;
  assign new_n57222_ = new_n57218_ & new_n57221_;
  assign new_n57223_ = ys__n24789 & new_n53839_;
  assign new_n57224_ = ys__n24786 & new_n53842_;
  assign new_n57225_ = ~new_n57223_ & ~new_n57224_;
  assign new_n57226_ = ys__n24783 & new_n53841_;
  assign new_n57227_ = ys__n39748 & new_n53831_;
  assign new_n57228_ = ~new_n57226_ & ~new_n57227_;
  assign new_n57229_ = new_n57225_ & new_n57228_;
  assign new_n57230_ = new_n57222_ & new_n57229_;
  assign new_n57231_ = ys__n39752 & new_n53723_;
  assign new_n57232_ = ys__n39750 & new_n53726_;
  assign new_n57233_ = ~new_n57231_ & ~new_n57232_;
  assign new_n57234_ = ys__n33717 & new_n53730_;
  assign new_n57235_ = ~ys__n33717 & new_n53733_;
  assign new_n57236_ = ~new_n57234_ & ~new_n57235_;
  assign new_n57237_ = new_n57233_ & new_n57236_;
  assign new_n57238_ = ys__n24798 & new_n53738_;
  assign new_n57239_ = ys__n24795 & new_n53740_;
  assign new_n57240_ = ~new_n57238_ & ~new_n57239_;
  assign new_n57241_ = ys__n24792 & new_n53744_;
  assign new_n57242_ = ys__n39754 & new_n53746_;
  assign new_n57243_ = ~new_n57241_ & ~new_n57242_;
  assign new_n57244_ = new_n57240_ & new_n57243_;
  assign new_n57245_ = new_n57237_ & new_n57244_;
  assign new_n57246_ = ~new_n57230_ & ~new_n57245_;
  assign new_n57247_ = ys__n39740 & new_n53871_;
  assign new_n57248_ = ys__n39738 & new_n53870_;
  assign new_n57249_ = ~new_n57247_ & ~new_n57248_;
  assign new_n57250_ = ys__n33705 & new_n53884_;
  assign new_n57251_ = ~ys__n33705 & new_n53887_;
  assign new_n57252_ = ~new_n57250_ & ~new_n57251_;
  assign new_n57253_ = new_n57249_ & new_n57252_;
  assign new_n57254_ = ys__n24780 & new_n53876_;
  assign new_n57255_ = ys__n24777 & new_n53879_;
  assign new_n57256_ = ~new_n57254_ & ~new_n57255_;
  assign new_n57257_ = ys__n24774 & new_n53878_;
  assign new_n57258_ = ys__n39742 & new_n53868_;
  assign new_n57259_ = ~new_n57257_ & ~new_n57258_;
  assign new_n57260_ = new_n57256_ & new_n57259_;
  assign new_n57261_ = new_n57253_ & new_n57260_;
  assign new_n57262_ = ~new_n57230_ & ~new_n57261_;
  assign new_n57263_ = ~new_n57245_ & ~new_n57261_;
  assign new_n57264_ = ~new_n57262_ & ~new_n57263_;
  assign new_n57265_ = ~new_n57246_ & new_n57264_;
  assign new_n57266_ = ~new_n57215_ & ~new_n57265_;
  assign new_n57267_ = ys__n39728 & new_n53781_;
  assign new_n57268_ = ys__n39726 & new_n53780_;
  assign new_n57269_ = ~new_n57267_ & ~new_n57268_;
  assign new_n57270_ = ys__n33693 & new_n53794_;
  assign new_n57271_ = ~ys__n33693 & new_n53797_;
  assign new_n57272_ = ~new_n57270_ & ~new_n57271_;
  assign new_n57273_ = new_n57269_ & new_n57272_;
  assign new_n57274_ = ys__n24762 & new_n53786_;
  assign new_n57275_ = ys__n24759 & new_n53789_;
  assign new_n57276_ = ~new_n57274_ & ~new_n57275_;
  assign new_n57277_ = ys__n24756 & new_n53788_;
  assign new_n57278_ = ys__n39730 & new_n53778_;
  assign new_n57279_ = ~new_n57277_ & ~new_n57278_;
  assign new_n57280_ = new_n57276_ & new_n57279_;
  assign new_n57281_ = new_n57273_ & new_n57280_;
  assign new_n57282_ = ys__n39734 & new_n53756_;
  assign new_n57283_ = ys__n39732 & new_n53755_;
  assign new_n57284_ = ~new_n57282_ & ~new_n57283_;
  assign new_n57285_ = ys__n33699 & new_n53769_;
  assign new_n57286_ = ~ys__n33699 & new_n53772_;
  assign new_n57287_ = ~new_n57285_ & ~new_n57286_;
  assign new_n57288_ = new_n57284_ & new_n57287_;
  assign new_n57289_ = ys__n24771 & new_n53761_;
  assign new_n57290_ = ys__n24768 & new_n53764_;
  assign new_n57291_ = ~new_n57289_ & ~new_n57290_;
  assign new_n57292_ = ys__n24765 & new_n53763_;
  assign new_n57293_ = ys__n39736 & new_n53753_;
  assign new_n57294_ = ~new_n57292_ & ~new_n57293_;
  assign new_n57295_ = new_n57291_ & new_n57294_;
  assign new_n57296_ = new_n57288_ & new_n57295_;
  assign new_n57297_ = ~new_n57281_ & ~new_n57296_;
  assign new_n57298_ = ys__n24753 & new_n53805_;
  assign new_n57299_ = ys__n24750 & new_n53806_;
  assign new_n57300_ = ~new_n57298_ & ~new_n57299_;
  assign new_n57301_ = ys__n39724 & new_n53813_;
  assign new_n57302_ = ys__n39722 & new_n53814_;
  assign new_n57303_ = ~new_n57301_ & ~new_n57302_;
  assign new_n57304_ = new_n57300_ & new_n57303_;
  assign new_n57305_ = ~new_n57281_ & ~new_n57304_;
  assign new_n57306_ = ~new_n57296_ & ~new_n57304_;
  assign new_n57307_ = ~new_n57305_ & ~new_n57306_;
  assign new_n57308_ = ~new_n57297_ & new_n57307_;
  assign new_n57309_ = ~new_n57215_ & ~new_n57308_;
  assign new_n57310_ = ~new_n57265_ & ~new_n57308_;
  assign new_n57311_ = ~new_n57309_ & ~new_n57310_;
  assign new_n57312_ = ~new_n57266_ & new_n57311_;
  assign new_n57313_ = ~new_n57194_ & ~new_n57312_;
  assign new_n57314_ = ~new_n57204_ & ~new_n57312_;
  assign new_n57315_ = ~new_n57313_ & ~new_n57314_;
  assign ys__n43565 = new_n57205_ | ~new_n57315_;
  assign new_n57317_ = ~new_n57204_ & new_n57313_;
  assign new_n57318_ = new_n57204_ & ~new_n57312_;
  assign new_n57319_ = new_n57194_ & new_n57318_;
  assign new_n57320_ = ~new_n57204_ & new_n57312_;
  assign new_n57321_ = new_n57194_ & new_n57320_;
  assign new_n57322_ = new_n57204_ & new_n57312_;
  assign new_n57323_ = ~new_n57194_ & new_n57322_;
  assign new_n57324_ = ~new_n57321_ & ~new_n57323_;
  assign new_n57325_ = ~new_n57319_ & new_n57324_;
  assign ys__n43570 = new_n57317_ | ~new_n57325_;
  assign new_n57327_ = ~new_n57265_ & new_n57309_;
  assign new_n57328_ = new_n57265_ & ~new_n57308_;
  assign new_n57329_ = new_n57215_ & new_n57328_;
  assign new_n57330_ = ~new_n57265_ & new_n57308_;
  assign new_n57331_ = new_n57215_ & new_n57330_;
  assign new_n57332_ = new_n57265_ & new_n57308_;
  assign new_n57333_ = ~new_n57215_ & new_n57332_;
  assign new_n57334_ = ~new_n57331_ & ~new_n57333_;
  assign new_n57335_ = ~new_n57329_ & new_n57334_;
  assign new_n57336_ = ~new_n57327_ & new_n57335_;
  assign new_n57337_ = ~new_n57103_ & new_n57120_;
  assign new_n57338_ = new_n57088_ & new_n57119_;
  assign new_n57339_ = ~new_n57103_ & new_n57338_;
  assign new_n57340_ = ~new_n57337_ & ~new_n57339_;
  assign new_n57341_ = ~new_n57088_ & new_n57119_;
  assign new_n57342_ = new_n57103_ & new_n57341_;
  assign new_n57343_ = new_n57088_ & ~new_n57119_;
  assign new_n57344_ = new_n57103_ & new_n57343_;
  assign new_n57345_ = ~new_n57342_ & ~new_n57344_;
  assign new_n57346_ = new_n57340_ & new_n57345_;
  assign new_n57347_ = ~new_n57336_ & ~new_n57346_;
  assign new_n57348_ = ~new_n57296_ & new_n57305_;
  assign new_n57349_ = new_n57281_ & new_n57304_;
  assign new_n57350_ = ~new_n57296_ & new_n57349_;
  assign new_n57351_ = ~new_n57348_ & ~new_n57350_;
  assign new_n57352_ = ~new_n57281_ & new_n57304_;
  assign new_n57353_ = new_n57296_ & new_n57352_;
  assign new_n57354_ = new_n57281_ & ~new_n57304_;
  assign new_n57355_ = new_n57296_ & new_n57354_;
  assign new_n57356_ = ~new_n57353_ & ~new_n57355_;
  assign new_n57357_ = new_n57351_ & new_n57356_;
  assign new_n57358_ = ys__n39744 & new_n53834_;
  assign new_n57359_ = ys__n39742 & new_n53833_;
  assign new_n57360_ = ~new_n57358_ & ~new_n57359_;
  assign new_n57361_ = ys__n33709 & new_n53847_;
  assign new_n57362_ = ~ys__n33709 & new_n53850_;
  assign new_n57363_ = ~new_n57361_ & ~new_n57362_;
  assign new_n57364_ = new_n57360_ & new_n57363_;
  assign new_n57365_ = ys__n24786 & new_n53839_;
  assign new_n57366_ = ys__n24783 & new_n53842_;
  assign new_n57367_ = ~new_n57365_ & ~new_n57366_;
  assign new_n57368_ = ys__n24780 & new_n53841_;
  assign new_n57369_ = ys__n39746 & new_n53831_;
  assign new_n57370_ = ~new_n57368_ & ~new_n57369_;
  assign new_n57371_ = new_n57367_ & new_n57370_;
  assign new_n57372_ = new_n57364_ & new_n57371_;
  assign new_n57373_ = ys__n39750 & new_n53723_;
  assign new_n57374_ = ys__n39748 & new_n53726_;
  assign new_n57375_ = ~new_n57373_ & ~new_n57374_;
  assign new_n57376_ = ys__n33715 & new_n53730_;
  assign new_n57377_ = ~ys__n33715 & new_n53733_;
  assign new_n57378_ = ~new_n57376_ & ~new_n57377_;
  assign new_n57379_ = new_n57375_ & new_n57378_;
  assign new_n57380_ = ys__n24795 & new_n53738_;
  assign new_n57381_ = ys__n24792 & new_n53740_;
  assign new_n57382_ = ~new_n57380_ & ~new_n57381_;
  assign new_n57383_ = ys__n24789 & new_n53744_;
  assign new_n57384_ = ys__n39752 & new_n53746_;
  assign new_n57385_ = ~new_n57383_ & ~new_n57384_;
  assign new_n57386_ = new_n57382_ & new_n57385_;
  assign new_n57387_ = new_n57379_ & new_n57386_;
  assign new_n57388_ = ~new_n57372_ & ~new_n57387_;
  assign new_n57389_ = ys__n39738 & new_n53871_;
  assign new_n57390_ = ys__n39736 & new_n53870_;
  assign new_n57391_ = ~new_n57389_ & ~new_n57390_;
  assign new_n57392_ = ys__n33703 & new_n53884_;
  assign new_n57393_ = ~ys__n33703 & new_n53887_;
  assign new_n57394_ = ~new_n57392_ & ~new_n57393_;
  assign new_n57395_ = new_n57391_ & new_n57394_;
  assign new_n57396_ = ys__n24777 & new_n53876_;
  assign new_n57397_ = ys__n24774 & new_n53879_;
  assign new_n57398_ = ~new_n57396_ & ~new_n57397_;
  assign new_n57399_ = ys__n24771 & new_n53878_;
  assign new_n57400_ = ys__n39740 & new_n53868_;
  assign new_n57401_ = ~new_n57399_ & ~new_n57400_;
  assign new_n57402_ = new_n57398_ & new_n57401_;
  assign new_n57403_ = new_n57395_ & new_n57402_;
  assign new_n57404_ = ~new_n57372_ & ~new_n57403_;
  assign new_n57405_ = ~new_n57387_ & ~new_n57403_;
  assign new_n57406_ = ~new_n57404_ & ~new_n57405_;
  assign new_n57407_ = ~new_n57388_ & new_n57406_;
  assign new_n57408_ = ~new_n57357_ & ~new_n57407_;
  assign new_n57409_ = ys__n39726 & new_n53781_;
  assign new_n57410_ = ys__n39724 & new_n53780_;
  assign new_n57411_ = ~new_n57409_ & ~new_n57410_;
  assign new_n57412_ = ys__n33691 & new_n53794_;
  assign new_n57413_ = ~ys__n33691 & new_n53797_;
  assign new_n57414_ = ~new_n57412_ & ~new_n57413_;
  assign new_n57415_ = new_n57411_ & new_n57414_;
  assign new_n57416_ = ys__n24759 & new_n53786_;
  assign new_n57417_ = ys__n24756 & new_n53789_;
  assign new_n57418_ = ~new_n57416_ & ~new_n57417_;
  assign new_n57419_ = ys__n24753 & new_n53788_;
  assign new_n57420_ = ys__n39728 & new_n53778_;
  assign new_n57421_ = ~new_n57419_ & ~new_n57420_;
  assign new_n57422_ = new_n57418_ & new_n57421_;
  assign new_n57423_ = new_n57415_ & new_n57422_;
  assign new_n57424_ = ys__n39732 & new_n53756_;
  assign new_n57425_ = ys__n39730 & new_n53755_;
  assign new_n57426_ = ~new_n57424_ & ~new_n57425_;
  assign new_n57427_ = ys__n33697 & new_n53769_;
  assign new_n57428_ = ~ys__n33697 & new_n53772_;
  assign new_n57429_ = ~new_n57427_ & ~new_n57428_;
  assign new_n57430_ = new_n57426_ & new_n57429_;
  assign new_n57431_ = ys__n24768 & new_n53761_;
  assign new_n57432_ = ys__n24765 & new_n53764_;
  assign new_n57433_ = ~new_n57431_ & ~new_n57432_;
  assign new_n57434_ = ys__n24762 & new_n53763_;
  assign new_n57435_ = ys__n39734 & new_n53753_;
  assign new_n57436_ = ~new_n57434_ & ~new_n57435_;
  assign new_n57437_ = new_n57433_ & new_n57436_;
  assign new_n57438_ = new_n57430_ & new_n57437_;
  assign new_n57439_ = ~new_n57423_ & ~new_n57438_;
  assign new_n57440_ = ys__n24750 & new_n53805_;
  assign new_n57441_ = ys__n24747 & new_n53806_;
  assign new_n57442_ = ~new_n57440_ & ~new_n57441_;
  assign new_n57443_ = ys__n39722 & new_n53813_;
  assign new_n57444_ = ys__n39720 & new_n53814_;
  assign new_n57445_ = ~new_n57443_ & ~new_n57444_;
  assign new_n57446_ = new_n57442_ & new_n57445_;
  assign new_n57447_ = ~new_n57423_ & ~new_n57446_;
  assign new_n57448_ = ~new_n57438_ & ~new_n57446_;
  assign new_n57449_ = ~new_n57447_ & ~new_n57448_;
  assign new_n57450_ = ~new_n57439_ & new_n57449_;
  assign new_n57451_ = ~new_n57357_ & ~new_n57450_;
  assign new_n57452_ = ~new_n57407_ & ~new_n57450_;
  assign new_n57453_ = ~new_n57451_ & ~new_n57452_;
  assign new_n57454_ = ~new_n57408_ & new_n57453_;
  assign new_n57455_ = ~new_n57336_ & ~new_n57454_;
  assign new_n57456_ = ~new_n57346_ & ~new_n57454_;
  assign new_n57457_ = ~new_n57455_ & ~new_n57456_;
  assign ys__n43619 = new_n57347_ | ~new_n57457_;
  assign new_n57459_ = ~new_n57346_ & new_n57455_;
  assign new_n57460_ = new_n57346_ & ~new_n57454_;
  assign new_n57461_ = new_n57336_ & new_n57460_;
  assign new_n57462_ = ~new_n57346_ & new_n57454_;
  assign new_n57463_ = new_n57336_ & new_n57462_;
  assign new_n57464_ = new_n57346_ & new_n57454_;
  assign new_n57465_ = ~new_n57336_ & new_n57464_;
  assign new_n57466_ = ~new_n57463_ & ~new_n57465_;
  assign new_n57467_ = ~new_n57461_ & new_n57466_;
  assign ys__n43624 = new_n57459_ | ~new_n57467_;
  assign new_n57469_ = ~new_n57407_ & new_n57451_;
  assign new_n57470_ = new_n57407_ & ~new_n57450_;
  assign new_n57471_ = new_n57357_ & new_n57470_;
  assign new_n57472_ = ~new_n57407_ & new_n57450_;
  assign new_n57473_ = new_n57357_ & new_n57472_;
  assign new_n57474_ = new_n57407_ & new_n57450_;
  assign new_n57475_ = ~new_n57357_ & new_n57474_;
  assign new_n57476_ = ~new_n57473_ & ~new_n57475_;
  assign new_n57477_ = ~new_n57471_ & new_n57476_;
  assign new_n57478_ = ~new_n57469_ & new_n57477_;
  assign new_n57479_ = ~new_n57245_ & new_n57262_;
  assign new_n57480_ = new_n57230_ & new_n57261_;
  assign new_n57481_ = ~new_n57245_ & new_n57480_;
  assign new_n57482_ = ~new_n57479_ & ~new_n57481_;
  assign new_n57483_ = ~new_n57230_ & new_n57261_;
  assign new_n57484_ = new_n57245_ & new_n57483_;
  assign new_n57485_ = new_n57230_ & ~new_n57261_;
  assign new_n57486_ = new_n57245_ & new_n57485_;
  assign new_n57487_ = ~new_n57484_ & ~new_n57486_;
  assign new_n57488_ = new_n57482_ & new_n57487_;
  assign new_n57489_ = ~new_n57478_ & ~new_n57488_;
  assign new_n57490_ = ~new_n57438_ & new_n57447_;
  assign new_n57491_ = new_n57423_ & new_n57446_;
  assign new_n57492_ = ~new_n57438_ & new_n57491_;
  assign new_n57493_ = ~new_n57490_ & ~new_n57492_;
  assign new_n57494_ = ~new_n57423_ & new_n57446_;
  assign new_n57495_ = new_n57438_ & new_n57494_;
  assign new_n57496_ = new_n57423_ & ~new_n57446_;
  assign new_n57497_ = new_n57438_ & new_n57496_;
  assign new_n57498_ = ~new_n57495_ & ~new_n57497_;
  assign new_n57499_ = new_n57493_ & new_n57498_;
  assign new_n57500_ = ys__n39742 & new_n53834_;
  assign new_n57501_ = ys__n39740 & new_n53833_;
  assign new_n57502_ = ~new_n57500_ & ~new_n57501_;
  assign new_n57503_ = ys__n33707 & new_n53847_;
  assign new_n57504_ = ~ys__n33707 & new_n53850_;
  assign new_n57505_ = ~new_n57503_ & ~new_n57504_;
  assign new_n57506_ = new_n57502_ & new_n57505_;
  assign new_n57507_ = ys__n24783 & new_n53839_;
  assign new_n57508_ = ys__n24780 & new_n53842_;
  assign new_n57509_ = ~new_n57507_ & ~new_n57508_;
  assign new_n57510_ = ys__n24777 & new_n53841_;
  assign new_n57511_ = ys__n39744 & new_n53831_;
  assign new_n57512_ = ~new_n57510_ & ~new_n57511_;
  assign new_n57513_ = new_n57509_ & new_n57512_;
  assign new_n57514_ = new_n57506_ & new_n57513_;
  assign new_n57515_ = ys__n39748 & new_n53723_;
  assign new_n57516_ = ys__n39746 & new_n53726_;
  assign new_n57517_ = ~new_n57515_ & ~new_n57516_;
  assign new_n57518_ = ys__n33713 & new_n53730_;
  assign new_n57519_ = ~ys__n33713 & new_n53733_;
  assign new_n57520_ = ~new_n57518_ & ~new_n57519_;
  assign new_n57521_ = new_n57517_ & new_n57520_;
  assign new_n57522_ = ys__n24792 & new_n53738_;
  assign new_n57523_ = ys__n24789 & new_n53740_;
  assign new_n57524_ = ~new_n57522_ & ~new_n57523_;
  assign new_n57525_ = ys__n24786 & new_n53744_;
  assign new_n57526_ = ys__n39750 & new_n53746_;
  assign new_n57527_ = ~new_n57525_ & ~new_n57526_;
  assign new_n57528_ = new_n57524_ & new_n57527_;
  assign new_n57529_ = new_n57521_ & new_n57528_;
  assign new_n57530_ = ~new_n57514_ & ~new_n57529_;
  assign new_n57531_ = ys__n39736 & new_n53871_;
  assign new_n57532_ = ys__n39734 & new_n53870_;
  assign new_n57533_ = ~new_n57531_ & ~new_n57532_;
  assign new_n57534_ = ys__n33701 & new_n53884_;
  assign new_n57535_ = ~ys__n33701 & new_n53887_;
  assign new_n57536_ = ~new_n57534_ & ~new_n57535_;
  assign new_n57537_ = new_n57533_ & new_n57536_;
  assign new_n57538_ = ys__n24774 & new_n53876_;
  assign new_n57539_ = ys__n24771 & new_n53879_;
  assign new_n57540_ = ~new_n57538_ & ~new_n57539_;
  assign new_n57541_ = ys__n24768 & new_n53878_;
  assign new_n57542_ = ys__n39738 & new_n53868_;
  assign new_n57543_ = ~new_n57541_ & ~new_n57542_;
  assign new_n57544_ = new_n57540_ & new_n57543_;
  assign new_n57545_ = new_n57537_ & new_n57544_;
  assign new_n57546_ = ~new_n57514_ & ~new_n57545_;
  assign new_n57547_ = ~new_n57529_ & ~new_n57545_;
  assign new_n57548_ = ~new_n57546_ & ~new_n57547_;
  assign new_n57549_ = ~new_n57530_ & new_n57548_;
  assign new_n57550_ = ~new_n57499_ & ~new_n57549_;
  assign new_n57551_ = ys__n39724 & new_n53781_;
  assign new_n57552_ = ys__n39722 & new_n53780_;
  assign new_n57553_ = ~new_n57551_ & ~new_n57552_;
  assign new_n57554_ = ys__n33689 & new_n53794_;
  assign new_n57555_ = ~ys__n33689 & new_n53797_;
  assign new_n57556_ = ~new_n57554_ & ~new_n57555_;
  assign new_n57557_ = new_n57553_ & new_n57556_;
  assign new_n57558_ = ys__n24756 & new_n53786_;
  assign new_n57559_ = ys__n24753 & new_n53789_;
  assign new_n57560_ = ~new_n57558_ & ~new_n57559_;
  assign new_n57561_ = ys__n24750 & new_n53788_;
  assign new_n57562_ = ys__n39726 & new_n53778_;
  assign new_n57563_ = ~new_n57561_ & ~new_n57562_;
  assign new_n57564_ = new_n57560_ & new_n57563_;
  assign new_n57565_ = new_n57557_ & new_n57564_;
  assign new_n57566_ = ys__n39730 & new_n53756_;
  assign new_n57567_ = ys__n39728 & new_n53755_;
  assign new_n57568_ = ~new_n57566_ & ~new_n57567_;
  assign new_n57569_ = ys__n33695 & new_n53769_;
  assign new_n57570_ = ~ys__n33695 & new_n53772_;
  assign new_n57571_ = ~new_n57569_ & ~new_n57570_;
  assign new_n57572_ = new_n57568_ & new_n57571_;
  assign new_n57573_ = ys__n24765 & new_n53761_;
  assign new_n57574_ = ys__n24762 & new_n53764_;
  assign new_n57575_ = ~new_n57573_ & ~new_n57574_;
  assign new_n57576_ = ys__n24759 & new_n53763_;
  assign new_n57577_ = ys__n39732 & new_n53753_;
  assign new_n57578_ = ~new_n57576_ & ~new_n57577_;
  assign new_n57579_ = new_n57575_ & new_n57578_;
  assign new_n57580_ = new_n57572_ & new_n57579_;
  assign new_n57581_ = ~new_n57565_ & ~new_n57580_;
  assign new_n57582_ = ys__n24747 & new_n53805_;
  assign new_n57583_ = ys__n24744 & new_n53806_;
  assign new_n57584_ = ~new_n57582_ & ~new_n57583_;
  assign new_n57585_ = ys__n39720 & new_n53813_;
  assign new_n57586_ = ys__n39718 & new_n53814_;
  assign new_n57587_ = ~new_n57585_ & ~new_n57586_;
  assign new_n57588_ = new_n57584_ & new_n57587_;
  assign new_n57589_ = ~new_n57565_ & ~new_n57588_;
  assign new_n57590_ = ~new_n57580_ & ~new_n57588_;
  assign new_n57591_ = ~new_n57589_ & ~new_n57590_;
  assign new_n57592_ = ~new_n57581_ & new_n57591_;
  assign new_n57593_ = ~new_n57499_ & ~new_n57592_;
  assign new_n57594_ = ~new_n57549_ & ~new_n57592_;
  assign new_n57595_ = ~new_n57593_ & ~new_n57594_;
  assign new_n57596_ = ~new_n57550_ & new_n57595_;
  assign new_n57597_ = ~new_n57478_ & ~new_n57596_;
  assign new_n57598_ = ~new_n57488_ & ~new_n57596_;
  assign new_n57599_ = ~new_n57597_ & ~new_n57598_;
  assign ys__n43673 = new_n57489_ | ~new_n57599_;
  assign new_n57601_ = ~new_n57488_ & new_n57597_;
  assign new_n57602_ = new_n57488_ & ~new_n57596_;
  assign new_n57603_ = new_n57478_ & new_n57602_;
  assign new_n57604_ = ~new_n57488_ & new_n57596_;
  assign new_n57605_ = new_n57478_ & new_n57604_;
  assign new_n57606_ = new_n57488_ & new_n57596_;
  assign new_n57607_ = ~new_n57478_ & new_n57606_;
  assign new_n57608_ = ~new_n57605_ & ~new_n57607_;
  assign new_n57609_ = ~new_n57603_ & new_n57608_;
  assign ys__n43678 = new_n57601_ | ~new_n57609_;
  assign new_n57611_ = ~new_n57549_ & new_n57593_;
  assign new_n57612_ = new_n57549_ & ~new_n57592_;
  assign new_n57613_ = new_n57499_ & new_n57612_;
  assign new_n57614_ = ~new_n57549_ & new_n57592_;
  assign new_n57615_ = new_n57499_ & new_n57614_;
  assign new_n57616_ = new_n57549_ & new_n57592_;
  assign new_n57617_ = ~new_n57499_ & new_n57616_;
  assign new_n57618_ = ~new_n57615_ & ~new_n57617_;
  assign new_n57619_ = ~new_n57613_ & new_n57618_;
  assign new_n57620_ = ~new_n57611_ & new_n57619_;
  assign new_n57621_ = ~new_n57387_ & new_n57404_;
  assign new_n57622_ = new_n57372_ & new_n57403_;
  assign new_n57623_ = ~new_n57387_ & new_n57622_;
  assign new_n57624_ = ~new_n57621_ & ~new_n57623_;
  assign new_n57625_ = ~new_n57372_ & new_n57403_;
  assign new_n57626_ = new_n57387_ & new_n57625_;
  assign new_n57627_ = new_n57372_ & ~new_n57403_;
  assign new_n57628_ = new_n57387_ & new_n57627_;
  assign new_n57629_ = ~new_n57626_ & ~new_n57628_;
  assign new_n57630_ = new_n57624_ & new_n57629_;
  assign new_n57631_ = ~new_n57620_ & ~new_n57630_;
  assign new_n57632_ = ~new_n57580_ & new_n57589_;
  assign new_n57633_ = new_n57565_ & new_n57588_;
  assign new_n57634_ = ~new_n57580_ & new_n57633_;
  assign new_n57635_ = ~new_n57632_ & ~new_n57634_;
  assign new_n57636_ = ~new_n57565_ & new_n57588_;
  assign new_n57637_ = new_n57580_ & new_n57636_;
  assign new_n57638_ = new_n57565_ & ~new_n57588_;
  assign new_n57639_ = new_n57580_ & new_n57638_;
  assign new_n57640_ = ~new_n57637_ & ~new_n57639_;
  assign new_n57641_ = new_n57635_ & new_n57640_;
  assign new_n57642_ = ys__n39740 & new_n53834_;
  assign new_n57643_ = ys__n39738 & new_n53833_;
  assign new_n57644_ = ~new_n57642_ & ~new_n57643_;
  assign new_n57645_ = ys__n33705 & new_n53847_;
  assign new_n57646_ = ~ys__n33705 & new_n53850_;
  assign new_n57647_ = ~new_n57645_ & ~new_n57646_;
  assign new_n57648_ = new_n57644_ & new_n57647_;
  assign new_n57649_ = ys__n24780 & new_n53839_;
  assign new_n57650_ = ys__n24777 & new_n53842_;
  assign new_n57651_ = ~new_n57649_ & ~new_n57650_;
  assign new_n57652_ = ys__n24774 & new_n53841_;
  assign new_n57653_ = ys__n39742 & new_n53831_;
  assign new_n57654_ = ~new_n57652_ & ~new_n57653_;
  assign new_n57655_ = new_n57651_ & new_n57654_;
  assign new_n57656_ = new_n57648_ & new_n57655_;
  assign new_n57657_ = ys__n39746 & new_n53723_;
  assign new_n57658_ = ys__n39744 & new_n53726_;
  assign new_n57659_ = ~new_n57657_ & ~new_n57658_;
  assign new_n57660_ = ys__n33711 & new_n53730_;
  assign new_n57661_ = ~ys__n33711 & new_n53733_;
  assign new_n57662_ = ~new_n57660_ & ~new_n57661_;
  assign new_n57663_ = new_n57659_ & new_n57662_;
  assign new_n57664_ = ys__n24789 & new_n53738_;
  assign new_n57665_ = ys__n24786 & new_n53740_;
  assign new_n57666_ = ~new_n57664_ & ~new_n57665_;
  assign new_n57667_ = ys__n24783 & new_n53744_;
  assign new_n57668_ = ys__n39748 & new_n53746_;
  assign new_n57669_ = ~new_n57667_ & ~new_n57668_;
  assign new_n57670_ = new_n57666_ & new_n57669_;
  assign new_n57671_ = new_n57663_ & new_n57670_;
  assign new_n57672_ = ~new_n57656_ & ~new_n57671_;
  assign new_n57673_ = ys__n39734 & new_n53871_;
  assign new_n57674_ = ys__n39732 & new_n53870_;
  assign new_n57675_ = ~new_n57673_ & ~new_n57674_;
  assign new_n57676_ = ys__n33699 & new_n53884_;
  assign new_n57677_ = ~ys__n33699 & new_n53887_;
  assign new_n57678_ = ~new_n57676_ & ~new_n57677_;
  assign new_n57679_ = new_n57675_ & new_n57678_;
  assign new_n57680_ = ys__n24771 & new_n53876_;
  assign new_n57681_ = ys__n24768 & new_n53879_;
  assign new_n57682_ = ~new_n57680_ & ~new_n57681_;
  assign new_n57683_ = ys__n24765 & new_n53878_;
  assign new_n57684_ = ys__n39736 & new_n53868_;
  assign new_n57685_ = ~new_n57683_ & ~new_n57684_;
  assign new_n57686_ = new_n57682_ & new_n57685_;
  assign new_n57687_ = new_n57679_ & new_n57686_;
  assign new_n57688_ = ~new_n57656_ & ~new_n57687_;
  assign new_n57689_ = ~new_n57671_ & ~new_n57687_;
  assign new_n57690_ = ~new_n57688_ & ~new_n57689_;
  assign new_n57691_ = ~new_n57672_ & new_n57690_;
  assign new_n57692_ = ~new_n57641_ & ~new_n57691_;
  assign new_n57693_ = ys__n39722 & new_n53781_;
  assign new_n57694_ = ys__n39720 & new_n53780_;
  assign new_n57695_ = ~new_n57693_ & ~new_n57694_;
  assign new_n57696_ = ys__n33687 & new_n53794_;
  assign new_n57697_ = ~ys__n33687 & new_n53797_;
  assign new_n57698_ = ~new_n57696_ & ~new_n57697_;
  assign new_n57699_ = new_n57695_ & new_n57698_;
  assign new_n57700_ = ys__n24753 & new_n53786_;
  assign new_n57701_ = ys__n24750 & new_n53789_;
  assign new_n57702_ = ~new_n57700_ & ~new_n57701_;
  assign new_n57703_ = ys__n24747 & new_n53788_;
  assign new_n57704_ = ys__n39724 & new_n53778_;
  assign new_n57705_ = ~new_n57703_ & ~new_n57704_;
  assign new_n57706_ = new_n57702_ & new_n57705_;
  assign new_n57707_ = new_n57699_ & new_n57706_;
  assign new_n57708_ = ys__n39728 & new_n53756_;
  assign new_n57709_ = ys__n39726 & new_n53755_;
  assign new_n57710_ = ~new_n57708_ & ~new_n57709_;
  assign new_n57711_ = ys__n33693 & new_n53769_;
  assign new_n57712_ = ~ys__n33693 & new_n53772_;
  assign new_n57713_ = ~new_n57711_ & ~new_n57712_;
  assign new_n57714_ = new_n57710_ & new_n57713_;
  assign new_n57715_ = ys__n24762 & new_n53761_;
  assign new_n57716_ = ys__n24759 & new_n53764_;
  assign new_n57717_ = ~new_n57715_ & ~new_n57716_;
  assign new_n57718_ = ys__n24756 & new_n53763_;
  assign new_n57719_ = ys__n39730 & new_n53753_;
  assign new_n57720_ = ~new_n57718_ & ~new_n57719_;
  assign new_n57721_ = new_n57717_ & new_n57720_;
  assign new_n57722_ = new_n57714_ & new_n57721_;
  assign new_n57723_ = ~new_n57707_ & ~new_n57722_;
  assign new_n57724_ = ys__n24744 & new_n53805_;
  assign new_n57725_ = ys__n24741 & new_n53806_;
  assign new_n57726_ = ~new_n57724_ & ~new_n57725_;
  assign new_n57727_ = ys__n39718 & new_n53813_;
  assign new_n57728_ = ys__n24741 & new_n53814_;
  assign new_n57729_ = ~new_n57727_ & ~new_n57728_;
  assign new_n57730_ = new_n57726_ & new_n57729_;
  assign new_n57731_ = ~new_n57707_ & ~new_n57730_;
  assign new_n57732_ = ~new_n57722_ & ~new_n57730_;
  assign new_n57733_ = ~new_n57731_ & ~new_n57732_;
  assign new_n57734_ = ~new_n57723_ & new_n57733_;
  assign new_n57735_ = ~new_n57641_ & ~new_n57734_;
  assign new_n57736_ = ~new_n57691_ & ~new_n57734_;
  assign new_n57737_ = ~new_n57735_ & ~new_n57736_;
  assign new_n57738_ = ~new_n57692_ & new_n57737_;
  assign new_n57739_ = ~new_n57620_ & ~new_n57738_;
  assign new_n57740_ = ~new_n57630_ & ~new_n57738_;
  assign new_n57741_ = ~new_n57739_ & ~new_n57740_;
  assign ys__n43727 = new_n57631_ | ~new_n57741_;
  assign new_n57743_ = ~new_n57630_ & new_n57739_;
  assign new_n57744_ = new_n57630_ & ~new_n57738_;
  assign new_n57745_ = new_n57620_ & new_n57744_;
  assign new_n57746_ = ~new_n57630_ & new_n57738_;
  assign new_n57747_ = new_n57620_ & new_n57746_;
  assign new_n57748_ = new_n57630_ & new_n57738_;
  assign new_n57749_ = ~new_n57620_ & new_n57748_;
  assign new_n57750_ = ~new_n57747_ & ~new_n57749_;
  assign new_n57751_ = ~new_n57745_ & new_n57750_;
  assign ys__n43732 = new_n57743_ | ~new_n57751_;
  assign new_n57753_ = ~new_n57691_ & new_n57735_;
  assign new_n57754_ = new_n57691_ & ~new_n57734_;
  assign new_n57755_ = new_n57641_ & new_n57754_;
  assign new_n57756_ = ~new_n57691_ & new_n57734_;
  assign new_n57757_ = new_n57641_ & new_n57756_;
  assign new_n57758_ = new_n57691_ & new_n57734_;
  assign new_n57759_ = ~new_n57641_ & new_n57758_;
  assign new_n57760_ = ~new_n57757_ & ~new_n57759_;
  assign new_n57761_ = ~new_n57755_ & new_n57760_;
  assign new_n57762_ = ~new_n57753_ & new_n57761_;
  assign new_n57763_ = ~new_n57529_ & new_n57546_;
  assign new_n57764_ = new_n57514_ & new_n57545_;
  assign new_n57765_ = ~new_n57529_ & new_n57764_;
  assign new_n57766_ = ~new_n57763_ & ~new_n57765_;
  assign new_n57767_ = ~new_n57514_ & new_n57545_;
  assign new_n57768_ = new_n57529_ & new_n57767_;
  assign new_n57769_ = new_n57514_ & ~new_n57545_;
  assign new_n57770_ = new_n57529_ & new_n57769_;
  assign new_n57771_ = ~new_n57768_ & ~new_n57770_;
  assign new_n57772_ = new_n57766_ & new_n57771_;
  assign new_n57773_ = ~new_n57762_ & ~new_n57772_;
  assign new_n57774_ = ~new_n57722_ & new_n57731_;
  assign new_n57775_ = new_n57707_ & new_n57730_;
  assign new_n57776_ = ~new_n57722_ & new_n57775_;
  assign new_n57777_ = ~new_n57774_ & ~new_n57776_;
  assign new_n57778_ = ~new_n57707_ & new_n57730_;
  assign new_n57779_ = new_n57722_ & new_n57778_;
  assign new_n57780_ = new_n57707_ & ~new_n57730_;
  assign new_n57781_ = new_n57722_ & new_n57780_;
  assign new_n57782_ = ~new_n57779_ & ~new_n57781_;
  assign new_n57783_ = new_n57777_ & new_n57782_;
  assign new_n57784_ = ys__n39738 & new_n53834_;
  assign new_n57785_ = ys__n39736 & new_n53833_;
  assign new_n57786_ = ~new_n57784_ & ~new_n57785_;
  assign new_n57787_ = ys__n33703 & new_n53847_;
  assign new_n57788_ = ~ys__n33703 & new_n53850_;
  assign new_n57789_ = ~new_n57787_ & ~new_n57788_;
  assign new_n57790_ = new_n57786_ & new_n57789_;
  assign new_n57791_ = ys__n24777 & new_n53839_;
  assign new_n57792_ = ys__n24774 & new_n53842_;
  assign new_n57793_ = ~new_n57791_ & ~new_n57792_;
  assign new_n57794_ = ys__n24771 & new_n53841_;
  assign new_n57795_ = ys__n39740 & new_n53831_;
  assign new_n57796_ = ~new_n57794_ & ~new_n57795_;
  assign new_n57797_ = new_n57793_ & new_n57796_;
  assign new_n57798_ = new_n57790_ & new_n57797_;
  assign new_n57799_ = ys__n39744 & new_n53723_;
  assign new_n57800_ = ys__n39742 & new_n53726_;
  assign new_n57801_ = ~new_n57799_ & ~new_n57800_;
  assign new_n57802_ = ys__n33709 & new_n53730_;
  assign new_n57803_ = ~ys__n33709 & new_n53733_;
  assign new_n57804_ = ~new_n57802_ & ~new_n57803_;
  assign new_n57805_ = new_n57801_ & new_n57804_;
  assign new_n57806_ = ys__n24786 & new_n53738_;
  assign new_n57807_ = ys__n24783 & new_n53740_;
  assign new_n57808_ = ~new_n57806_ & ~new_n57807_;
  assign new_n57809_ = ys__n24780 & new_n53744_;
  assign new_n57810_ = ys__n39746 & new_n53746_;
  assign new_n57811_ = ~new_n57809_ & ~new_n57810_;
  assign new_n57812_ = new_n57808_ & new_n57811_;
  assign new_n57813_ = new_n57805_ & new_n57812_;
  assign new_n57814_ = ~new_n57798_ & ~new_n57813_;
  assign new_n57815_ = ys__n39732 & new_n53871_;
  assign new_n57816_ = ys__n39730 & new_n53870_;
  assign new_n57817_ = ~new_n57815_ & ~new_n57816_;
  assign new_n57818_ = ys__n33697 & new_n53884_;
  assign new_n57819_ = ~ys__n33697 & new_n53887_;
  assign new_n57820_ = ~new_n57818_ & ~new_n57819_;
  assign new_n57821_ = new_n57817_ & new_n57820_;
  assign new_n57822_ = ys__n24768 & new_n53876_;
  assign new_n57823_ = ys__n24765 & new_n53879_;
  assign new_n57824_ = ~new_n57822_ & ~new_n57823_;
  assign new_n57825_ = ys__n24762 & new_n53878_;
  assign new_n57826_ = ys__n39734 & new_n53868_;
  assign new_n57827_ = ~new_n57825_ & ~new_n57826_;
  assign new_n57828_ = new_n57824_ & new_n57827_;
  assign new_n57829_ = new_n57821_ & new_n57828_;
  assign new_n57830_ = ~new_n57798_ & ~new_n57829_;
  assign new_n57831_ = ~new_n57813_ & ~new_n57829_;
  assign new_n57832_ = ~new_n57830_ & ~new_n57831_;
  assign new_n57833_ = ~new_n57814_ & new_n57832_;
  assign new_n57834_ = ~new_n57783_ & ~new_n57833_;
  assign new_n57835_ = ys__n39720 & new_n53781_;
  assign new_n57836_ = ys__n39718 & new_n53780_;
  assign new_n57837_ = ~new_n57835_ & ~new_n57836_;
  assign new_n57838_ = ys__n33685 & new_n53794_;
  assign new_n57839_ = ~ys__n33685 & new_n53797_;
  assign new_n57840_ = ~new_n57838_ & ~new_n57839_;
  assign new_n57841_ = new_n57837_ & new_n57840_;
  assign new_n57842_ = ys__n24750 & new_n53786_;
  assign new_n57843_ = ys__n24747 & new_n53789_;
  assign new_n57844_ = ~new_n57842_ & ~new_n57843_;
  assign new_n57845_ = ys__n24744 & new_n53788_;
  assign new_n57846_ = ys__n39722 & new_n53778_;
  assign new_n57847_ = ~new_n57845_ & ~new_n57846_;
  assign new_n57848_ = new_n57844_ & new_n57847_;
  assign new_n57849_ = new_n57841_ & new_n57848_;
  assign new_n57850_ = ys__n39726 & new_n53756_;
  assign new_n57851_ = ys__n39724 & new_n53755_;
  assign new_n57852_ = ~new_n57850_ & ~new_n57851_;
  assign new_n57853_ = ys__n33691 & new_n53769_;
  assign new_n57854_ = ~ys__n33691 & new_n53772_;
  assign new_n57855_ = ~new_n57853_ & ~new_n57854_;
  assign new_n57856_ = new_n57852_ & new_n57855_;
  assign new_n57857_ = ys__n24759 & new_n53761_;
  assign new_n57858_ = ys__n24756 & new_n53764_;
  assign new_n57859_ = ~new_n57857_ & ~new_n57858_;
  assign new_n57860_ = ys__n24753 & new_n53763_;
  assign new_n57861_ = ys__n39728 & new_n53753_;
  assign new_n57862_ = ~new_n57860_ & ~new_n57861_;
  assign new_n57863_ = new_n57859_ & new_n57862_;
  assign new_n57864_ = new_n57856_ & new_n57863_;
  assign new_n57865_ = ~new_n57849_ & ~new_n57864_;
  assign new_n57866_ = ys__n24741 & new_n53805_;
  assign new_n57867_ = ys__n24741 & new_n53813_;
  assign new_n57868_ = ~new_n57866_ & ~new_n57867_;
  assign new_n57869_ = ~new_n57849_ & ~new_n57868_;
  assign new_n57870_ = ~new_n57864_ & ~new_n57868_;
  assign new_n57871_ = ~new_n57869_ & ~new_n57870_;
  assign new_n57872_ = ~new_n57865_ & new_n57871_;
  assign new_n57873_ = ~new_n57783_ & ~new_n57872_;
  assign new_n57874_ = ~new_n57833_ & ~new_n57872_;
  assign new_n57875_ = ~new_n57873_ & ~new_n57874_;
  assign new_n57876_ = ~new_n57834_ & new_n57875_;
  assign new_n57877_ = ~new_n57762_ & ~new_n57876_;
  assign new_n57878_ = ~new_n57772_ & ~new_n57876_;
  assign new_n57879_ = ~new_n57877_ & ~new_n57878_;
  assign ys__n43781 = new_n57773_ | ~new_n57879_;
  assign new_n57881_ = ~new_n57772_ & new_n57877_;
  assign new_n57882_ = new_n57772_ & ~new_n57876_;
  assign new_n57883_ = new_n57762_ & new_n57882_;
  assign new_n57884_ = ~new_n57772_ & new_n57876_;
  assign new_n57885_ = new_n57762_ & new_n57884_;
  assign new_n57886_ = new_n57772_ & new_n57876_;
  assign new_n57887_ = ~new_n57762_ & new_n57886_;
  assign new_n57888_ = ~new_n57885_ & ~new_n57887_;
  assign new_n57889_ = ~new_n57883_ & new_n57888_;
  assign ys__n43786 = new_n57881_ | ~new_n57889_;
  assign new_n57891_ = ~new_n57833_ & new_n57873_;
  assign new_n57892_ = new_n57833_ & ~new_n57872_;
  assign new_n57893_ = new_n57783_ & new_n57892_;
  assign new_n57894_ = ~new_n57833_ & new_n57872_;
  assign new_n57895_ = new_n57783_ & new_n57894_;
  assign new_n57896_ = new_n57833_ & new_n57872_;
  assign new_n57897_ = ~new_n57783_ & new_n57896_;
  assign new_n57898_ = ~new_n57895_ & ~new_n57897_;
  assign new_n57899_ = ~new_n57893_ & new_n57898_;
  assign new_n57900_ = ~new_n57891_ & new_n57899_;
  assign new_n57901_ = ~new_n57671_ & new_n57688_;
  assign new_n57902_ = new_n57656_ & new_n57687_;
  assign new_n57903_ = ~new_n57671_ & new_n57902_;
  assign new_n57904_ = ~new_n57901_ & ~new_n57903_;
  assign new_n57905_ = ~new_n57656_ & new_n57687_;
  assign new_n57906_ = new_n57671_ & new_n57905_;
  assign new_n57907_ = new_n57656_ & ~new_n57687_;
  assign new_n57908_ = new_n57671_ & new_n57907_;
  assign new_n57909_ = ~new_n57906_ & ~new_n57908_;
  assign new_n57910_ = new_n57904_ & new_n57909_;
  assign new_n57911_ = ~new_n57900_ & ~new_n57910_;
  assign new_n57912_ = ~new_n57864_ & new_n57869_;
  assign new_n57913_ = new_n57849_ & new_n57868_;
  assign new_n57914_ = ~new_n57864_ & new_n57913_;
  assign new_n57915_ = ~new_n57912_ & ~new_n57914_;
  assign new_n57916_ = ~new_n57849_ & new_n57868_;
  assign new_n57917_ = new_n57864_ & new_n57916_;
  assign new_n57918_ = new_n57849_ & ~new_n57868_;
  assign new_n57919_ = new_n57864_ & new_n57918_;
  assign new_n57920_ = ~new_n57917_ & ~new_n57919_;
  assign new_n57921_ = new_n57915_ & new_n57920_;
  assign new_n57922_ = ys__n39736 & new_n53834_;
  assign new_n57923_ = ys__n39734 & new_n53833_;
  assign new_n57924_ = ~new_n57922_ & ~new_n57923_;
  assign new_n57925_ = ys__n33701 & new_n53847_;
  assign new_n57926_ = ~ys__n33701 & new_n53850_;
  assign new_n57927_ = ~new_n57925_ & ~new_n57926_;
  assign new_n57928_ = new_n57924_ & new_n57927_;
  assign new_n57929_ = ys__n24774 & new_n53839_;
  assign new_n57930_ = ys__n24771 & new_n53842_;
  assign new_n57931_ = ~new_n57929_ & ~new_n57930_;
  assign new_n57932_ = ys__n24768 & new_n53841_;
  assign new_n57933_ = ys__n39738 & new_n53831_;
  assign new_n57934_ = ~new_n57932_ & ~new_n57933_;
  assign new_n57935_ = new_n57931_ & new_n57934_;
  assign new_n57936_ = new_n57928_ & new_n57935_;
  assign new_n57937_ = ys__n39742 & new_n53723_;
  assign new_n57938_ = ys__n39740 & new_n53726_;
  assign new_n57939_ = ~new_n57937_ & ~new_n57938_;
  assign new_n57940_ = ys__n33707 & new_n53730_;
  assign new_n57941_ = ~ys__n33707 & new_n53733_;
  assign new_n57942_ = ~new_n57940_ & ~new_n57941_;
  assign new_n57943_ = new_n57939_ & new_n57942_;
  assign new_n57944_ = ys__n24783 & new_n53738_;
  assign new_n57945_ = ys__n24780 & new_n53740_;
  assign new_n57946_ = ~new_n57944_ & ~new_n57945_;
  assign new_n57947_ = ys__n24777 & new_n53744_;
  assign new_n57948_ = ys__n39744 & new_n53746_;
  assign new_n57949_ = ~new_n57947_ & ~new_n57948_;
  assign new_n57950_ = new_n57946_ & new_n57949_;
  assign new_n57951_ = new_n57943_ & new_n57950_;
  assign new_n57952_ = ~new_n57936_ & ~new_n57951_;
  assign new_n57953_ = ys__n39730 & new_n53871_;
  assign new_n57954_ = ys__n39728 & new_n53870_;
  assign new_n57955_ = ~new_n57953_ & ~new_n57954_;
  assign new_n57956_ = ys__n33695 & new_n53884_;
  assign new_n57957_ = ~ys__n33695 & new_n53887_;
  assign new_n57958_ = ~new_n57956_ & ~new_n57957_;
  assign new_n57959_ = new_n57955_ & new_n57958_;
  assign new_n57960_ = ys__n24765 & new_n53876_;
  assign new_n57961_ = ys__n24762 & new_n53879_;
  assign new_n57962_ = ~new_n57960_ & ~new_n57961_;
  assign new_n57963_ = ys__n24759 & new_n53878_;
  assign new_n57964_ = ys__n39732 & new_n53868_;
  assign new_n57965_ = ~new_n57963_ & ~new_n57964_;
  assign new_n57966_ = new_n57962_ & new_n57965_;
  assign new_n57967_ = new_n57959_ & new_n57966_;
  assign new_n57968_ = ~new_n57936_ & ~new_n57967_;
  assign new_n57969_ = ~new_n57951_ & ~new_n57967_;
  assign new_n57970_ = ~new_n57968_ & ~new_n57969_;
  assign new_n57971_ = ~new_n57952_ & new_n57970_;
  assign new_n57972_ = ~new_n57921_ & ~new_n57971_;
  assign new_n57973_ = ys__n39718 & new_n53781_;
  assign new_n57974_ = ys__n24741 & new_n53780_;
  assign new_n57975_ = ~new_n57973_ & ~new_n57974_;
  assign new_n57976_ = ys__n33683 & new_n53794_;
  assign new_n57977_ = ~ys__n33683 & new_n53797_;
  assign new_n57978_ = ~new_n57976_ & ~new_n57977_;
  assign new_n57979_ = new_n57975_ & new_n57978_;
  assign new_n57980_ = ys__n24747 & new_n53786_;
  assign new_n57981_ = ys__n24744 & new_n53789_;
  assign new_n57982_ = ~new_n57980_ & ~new_n57981_;
  assign new_n57983_ = ys__n24741 & new_n53788_;
  assign new_n57984_ = ys__n39720 & new_n53778_;
  assign new_n57985_ = ~new_n57983_ & ~new_n57984_;
  assign new_n57986_ = new_n57982_ & new_n57985_;
  assign new_n57987_ = new_n57979_ & new_n57986_;
  assign new_n57988_ = ys__n39724 & new_n53756_;
  assign new_n57989_ = ys__n39722 & new_n53755_;
  assign new_n57990_ = ~new_n57988_ & ~new_n57989_;
  assign new_n57991_ = ys__n33689 & new_n53769_;
  assign new_n57992_ = ~ys__n33689 & new_n53772_;
  assign new_n57993_ = ~new_n57991_ & ~new_n57992_;
  assign new_n57994_ = new_n57990_ & new_n57993_;
  assign new_n57995_ = ys__n24756 & new_n53761_;
  assign new_n57996_ = ys__n24753 & new_n53764_;
  assign new_n57997_ = ~new_n57995_ & ~new_n57996_;
  assign new_n57998_ = ys__n24750 & new_n53763_;
  assign new_n57999_ = ys__n39726 & new_n53753_;
  assign new_n58000_ = ~new_n57998_ & ~new_n57999_;
  assign new_n58001_ = new_n57997_ & new_n58000_;
  assign new_n58002_ = new_n57994_ & new_n58001_;
  assign new_n58003_ = ~new_n57987_ & ~new_n58002_;
  assign new_n58004_ = ~new_n57921_ & new_n58003_;
  assign new_n58005_ = ~new_n57971_ & new_n58003_;
  assign new_n58006_ = ~new_n58004_ & ~new_n58005_;
  assign new_n58007_ = ~new_n57972_ & new_n58006_;
  assign new_n58008_ = ~new_n57900_ & ~new_n58007_;
  assign new_n58009_ = ~new_n57910_ & ~new_n58007_;
  assign new_n58010_ = ~new_n58008_ & ~new_n58009_;
  assign ys__n43835 = new_n57911_ | ~new_n58010_;
  assign new_n58012_ = ~new_n57910_ & new_n58008_;
  assign new_n58013_ = new_n57910_ & ~new_n58007_;
  assign new_n58014_ = new_n57900_ & new_n58013_;
  assign new_n58015_ = ~new_n57910_ & new_n58007_;
  assign new_n58016_ = new_n57900_ & new_n58015_;
  assign new_n58017_ = new_n57910_ & new_n58007_;
  assign new_n58018_ = ~new_n57900_ & new_n58017_;
  assign new_n58019_ = ~new_n58016_ & ~new_n58018_;
  assign new_n58020_ = ~new_n58014_ & new_n58019_;
  assign ys__n43840 = new_n58012_ | ~new_n58020_;
  assign new_n58022_ = ~new_n57971_ & new_n58004_;
  assign new_n58023_ = new_n57971_ & new_n58003_;
  assign new_n58024_ = new_n57921_ & new_n58023_;
  assign new_n58025_ = ~new_n57971_ & ~new_n58003_;
  assign new_n58026_ = new_n57921_ & new_n58025_;
  assign new_n58027_ = new_n57971_ & ~new_n58003_;
  assign new_n58028_ = ~new_n57921_ & new_n58027_;
  assign new_n58029_ = ~new_n58026_ & ~new_n58028_;
  assign new_n58030_ = ~new_n58024_ & new_n58029_;
  assign new_n58031_ = ~new_n58022_ & new_n58030_;
  assign new_n58032_ = ~new_n57813_ & new_n57830_;
  assign new_n58033_ = new_n57798_ & new_n57829_;
  assign new_n58034_ = ~new_n57813_ & new_n58033_;
  assign new_n58035_ = ~new_n58032_ & ~new_n58034_;
  assign new_n58036_ = ~new_n57798_ & new_n57829_;
  assign new_n58037_ = new_n57813_ & new_n58036_;
  assign new_n58038_ = new_n57798_ & ~new_n57829_;
  assign new_n58039_ = new_n57813_ & new_n58038_;
  assign new_n58040_ = ~new_n58037_ & ~new_n58039_;
  assign new_n58041_ = new_n58035_ & new_n58040_;
  assign new_n58042_ = ~new_n58031_ & ~new_n58041_;
  assign new_n58043_ = new_n57987_ & ~new_n58002_;
  assign new_n58044_ = ~new_n57987_ & new_n58002_;
  assign new_n58045_ = ~new_n58043_ & ~new_n58044_;
  assign new_n58046_ = ys__n39734 & new_n53834_;
  assign new_n58047_ = ys__n39732 & new_n53833_;
  assign new_n58048_ = ~new_n58046_ & ~new_n58047_;
  assign new_n58049_ = ys__n33699 & new_n53847_;
  assign new_n58050_ = ~ys__n33699 & new_n53850_;
  assign new_n58051_ = ~new_n58049_ & ~new_n58050_;
  assign new_n58052_ = new_n58048_ & new_n58051_;
  assign new_n58053_ = ys__n24771 & new_n53839_;
  assign new_n58054_ = ys__n24768 & new_n53842_;
  assign new_n58055_ = ~new_n58053_ & ~new_n58054_;
  assign new_n58056_ = ys__n24765 & new_n53841_;
  assign new_n58057_ = ys__n39736 & new_n53831_;
  assign new_n58058_ = ~new_n58056_ & ~new_n58057_;
  assign new_n58059_ = new_n58055_ & new_n58058_;
  assign new_n58060_ = new_n58052_ & new_n58059_;
  assign new_n58061_ = ys__n39740 & new_n53723_;
  assign new_n58062_ = ys__n39738 & new_n53726_;
  assign new_n58063_ = ~new_n58061_ & ~new_n58062_;
  assign new_n58064_ = ys__n33705 & new_n53730_;
  assign new_n58065_ = ~ys__n33705 & new_n53733_;
  assign new_n58066_ = ~new_n58064_ & ~new_n58065_;
  assign new_n58067_ = new_n58063_ & new_n58066_;
  assign new_n58068_ = ys__n24780 & new_n53738_;
  assign new_n58069_ = ys__n24777 & new_n53740_;
  assign new_n58070_ = ~new_n58068_ & ~new_n58069_;
  assign new_n58071_ = ys__n24774 & new_n53744_;
  assign new_n58072_ = ys__n39742 & new_n53746_;
  assign new_n58073_ = ~new_n58071_ & ~new_n58072_;
  assign new_n58074_ = new_n58070_ & new_n58073_;
  assign new_n58075_ = new_n58067_ & new_n58074_;
  assign new_n58076_ = ~new_n58060_ & ~new_n58075_;
  assign new_n58077_ = ys__n39728 & new_n53871_;
  assign new_n58078_ = ys__n39726 & new_n53870_;
  assign new_n58079_ = ~new_n58077_ & ~new_n58078_;
  assign new_n58080_ = ys__n33693 & new_n53884_;
  assign new_n58081_ = ~ys__n33693 & new_n53887_;
  assign new_n58082_ = ~new_n58080_ & ~new_n58081_;
  assign new_n58083_ = new_n58079_ & new_n58082_;
  assign new_n58084_ = ys__n24762 & new_n53876_;
  assign new_n58085_ = ys__n24759 & new_n53879_;
  assign new_n58086_ = ~new_n58084_ & ~new_n58085_;
  assign new_n58087_ = ys__n24756 & new_n53878_;
  assign new_n58088_ = ys__n39730 & new_n53868_;
  assign new_n58089_ = ~new_n58087_ & ~new_n58088_;
  assign new_n58090_ = new_n58086_ & new_n58089_;
  assign new_n58091_ = new_n58083_ & new_n58090_;
  assign new_n58092_ = ~new_n58060_ & ~new_n58091_;
  assign new_n58093_ = ~new_n58075_ & ~new_n58091_;
  assign new_n58094_ = ~new_n58092_ & ~new_n58093_;
  assign new_n58095_ = ~new_n58076_ & new_n58094_;
  assign new_n58096_ = ~new_n58045_ & ~new_n58095_;
  assign new_n58097_ = ys__n24744 & new_n53786_;
  assign new_n58098_ = ys__n24741 & new_n53789_;
  assign new_n58099_ = ~new_n58097_ & ~new_n58098_;
  assign new_n58100_ = ys__n39718 & new_n53778_;
  assign new_n58101_ = ys__n24741 & new_n53781_;
  assign new_n58102_ = ~new_n58100_ & ~new_n58101_;
  assign new_n58103_ = ys__n33681 & new_n53794_;
  assign new_n58104_ = ~ys__n33681 & new_n53797_;
  assign new_n58105_ = ~new_n58103_ & ~new_n58104_;
  assign new_n58106_ = new_n58102_ & new_n58105_;
  assign new_n58107_ = new_n58099_ & new_n58106_;
  assign new_n58108_ = ys__n39722 & new_n53756_;
  assign new_n58109_ = ys__n39720 & new_n53755_;
  assign new_n58110_ = ~new_n58108_ & ~new_n58109_;
  assign new_n58111_ = ys__n33687 & new_n53769_;
  assign new_n58112_ = ~ys__n33687 & new_n53772_;
  assign new_n58113_ = ~new_n58111_ & ~new_n58112_;
  assign new_n58114_ = new_n58110_ & new_n58113_;
  assign new_n58115_ = ys__n24753 & new_n53761_;
  assign new_n58116_ = ys__n24750 & new_n53764_;
  assign new_n58117_ = ~new_n58115_ & ~new_n58116_;
  assign new_n58118_ = ys__n24747 & new_n53763_;
  assign new_n58119_ = ys__n39724 & new_n53753_;
  assign new_n58120_ = ~new_n58118_ & ~new_n58119_;
  assign new_n58121_ = new_n58117_ & new_n58120_;
  assign new_n58122_ = new_n58114_ & new_n58121_;
  assign new_n58123_ = ~new_n58107_ & ~new_n58122_;
  assign new_n58124_ = ~new_n58045_ & new_n58123_;
  assign new_n58125_ = ~new_n58095_ & new_n58123_;
  assign new_n58126_ = ~new_n58124_ & ~new_n58125_;
  assign new_n58127_ = ~new_n58096_ & new_n58126_;
  assign new_n58128_ = ~new_n58031_ & ~new_n58127_;
  assign new_n58129_ = ~new_n58041_ & ~new_n58127_;
  assign new_n58130_ = ~new_n58128_ & ~new_n58129_;
  assign ys__n43889 = new_n58042_ | ~new_n58130_;
  assign new_n58132_ = ~new_n58041_ & new_n58128_;
  assign new_n58133_ = new_n58041_ & ~new_n58127_;
  assign new_n58134_ = new_n58031_ & new_n58133_;
  assign new_n58135_ = ~new_n58041_ & new_n58127_;
  assign new_n58136_ = new_n58031_ & new_n58135_;
  assign new_n58137_ = new_n58041_ & new_n58127_;
  assign new_n58138_ = ~new_n58031_ & new_n58137_;
  assign new_n58139_ = ~new_n58136_ & ~new_n58138_;
  assign new_n58140_ = ~new_n58134_ & new_n58139_;
  assign ys__n43894 = new_n58132_ | ~new_n58140_;
  assign new_n58142_ = ~new_n58095_ & new_n58124_;
  assign new_n58143_ = new_n58045_ & ~new_n58123_;
  assign new_n58144_ = ~new_n58095_ & new_n58143_;
  assign new_n58145_ = ~new_n58142_ & ~new_n58144_;
  assign new_n58146_ = ~new_n58045_ & ~new_n58123_;
  assign new_n58147_ = new_n58095_ & new_n58146_;
  assign new_n58148_ = new_n58045_ & new_n58123_;
  assign new_n58149_ = new_n58095_ & new_n58148_;
  assign new_n58150_ = ~new_n58147_ & ~new_n58149_;
  assign new_n58151_ = new_n58145_ & new_n58150_;
  assign new_n58152_ = ~new_n57951_ & new_n57968_;
  assign new_n58153_ = new_n57936_ & new_n57967_;
  assign new_n58154_ = ~new_n57951_ & new_n58153_;
  assign new_n58155_ = ~new_n58152_ & ~new_n58154_;
  assign new_n58156_ = ~new_n57936_ & new_n57967_;
  assign new_n58157_ = new_n57951_ & new_n58156_;
  assign new_n58158_ = new_n57936_ & ~new_n57967_;
  assign new_n58159_ = new_n57951_ & new_n58158_;
  assign new_n58160_ = ~new_n58157_ & ~new_n58159_;
  assign new_n58161_ = new_n58155_ & new_n58160_;
  assign new_n58162_ = ~new_n58151_ & ~new_n58161_;
  assign new_n58163_ = new_n58107_ & ~new_n58122_;
  assign new_n58164_ = ~new_n58107_ & new_n58122_;
  assign new_n58165_ = ~new_n58163_ & ~new_n58164_;
  assign new_n58166_ = ys__n39732 & new_n53834_;
  assign new_n58167_ = ys__n39730 & new_n53833_;
  assign new_n58168_ = ~new_n58166_ & ~new_n58167_;
  assign new_n58169_ = ys__n33697 & new_n53847_;
  assign new_n58170_ = ~ys__n33697 & new_n53850_;
  assign new_n58171_ = ~new_n58169_ & ~new_n58170_;
  assign new_n58172_ = new_n58168_ & new_n58171_;
  assign new_n58173_ = ys__n24768 & new_n53839_;
  assign new_n58174_ = ys__n24765 & new_n53842_;
  assign new_n58175_ = ~new_n58173_ & ~new_n58174_;
  assign new_n58176_ = ys__n24762 & new_n53841_;
  assign new_n58177_ = ys__n39734 & new_n53831_;
  assign new_n58178_ = ~new_n58176_ & ~new_n58177_;
  assign new_n58179_ = new_n58175_ & new_n58178_;
  assign new_n58180_ = new_n58172_ & new_n58179_;
  assign new_n58181_ = ys__n39738 & new_n53723_;
  assign new_n58182_ = ys__n39736 & new_n53726_;
  assign new_n58183_ = ~new_n58181_ & ~new_n58182_;
  assign new_n58184_ = ys__n33703 & new_n53730_;
  assign new_n58185_ = ~ys__n33703 & new_n53733_;
  assign new_n58186_ = ~new_n58184_ & ~new_n58185_;
  assign new_n58187_ = new_n58183_ & new_n58186_;
  assign new_n58188_ = ys__n24777 & new_n53738_;
  assign new_n58189_ = ys__n24774 & new_n53740_;
  assign new_n58190_ = ~new_n58188_ & ~new_n58189_;
  assign new_n58191_ = ys__n24771 & new_n53744_;
  assign new_n58192_ = ys__n39740 & new_n53746_;
  assign new_n58193_ = ~new_n58191_ & ~new_n58192_;
  assign new_n58194_ = new_n58190_ & new_n58193_;
  assign new_n58195_ = new_n58187_ & new_n58194_;
  assign new_n58196_ = ~new_n58180_ & ~new_n58195_;
  assign new_n58197_ = ys__n39726 & new_n53871_;
  assign new_n58198_ = ys__n39724 & new_n53870_;
  assign new_n58199_ = ~new_n58197_ & ~new_n58198_;
  assign new_n58200_ = ys__n33691 & new_n53884_;
  assign new_n58201_ = ~ys__n33691 & new_n53887_;
  assign new_n58202_ = ~new_n58200_ & ~new_n58201_;
  assign new_n58203_ = new_n58199_ & new_n58202_;
  assign new_n58204_ = ys__n24759 & new_n53876_;
  assign new_n58205_ = ys__n24756 & new_n53879_;
  assign new_n58206_ = ~new_n58204_ & ~new_n58205_;
  assign new_n58207_ = ys__n24753 & new_n53878_;
  assign new_n58208_ = ys__n39728 & new_n53868_;
  assign new_n58209_ = ~new_n58207_ & ~new_n58208_;
  assign new_n58210_ = new_n58206_ & new_n58209_;
  assign new_n58211_ = new_n58203_ & new_n58210_;
  assign new_n58212_ = ~new_n58180_ & ~new_n58211_;
  assign new_n58213_ = ~new_n58195_ & ~new_n58211_;
  assign new_n58214_ = ~new_n58212_ & ~new_n58213_;
  assign new_n58215_ = ~new_n58196_ & new_n58214_;
  assign new_n58216_ = ~new_n58165_ & ~new_n58215_;
  assign new_n58217_ = ys__n24741 & new_n53786_;
  assign new_n58218_ = ys__n24741 & new_n53778_;
  assign new_n58219_ = ~new_n58217_ & ~new_n58218_;
  assign new_n58220_ = ys__n24741 & new_n53794_;
  assign new_n58221_ = ~ys__n24741 & new_n53797_;
  assign new_n58222_ = ~new_n58220_ & ~new_n58221_;
  assign new_n58223_ = new_n58219_ & new_n58222_;
  assign new_n58224_ = ys__n39720 & new_n53756_;
  assign new_n58225_ = ys__n39718 & new_n53755_;
  assign new_n58226_ = ~new_n58224_ & ~new_n58225_;
  assign new_n58227_ = ys__n33685 & new_n53769_;
  assign new_n58228_ = ~ys__n33685 & new_n53772_;
  assign new_n58229_ = ~new_n58227_ & ~new_n58228_;
  assign new_n58230_ = new_n58226_ & new_n58229_;
  assign new_n58231_ = ys__n24750 & new_n53761_;
  assign new_n58232_ = ys__n24747 & new_n53764_;
  assign new_n58233_ = ~new_n58231_ & ~new_n58232_;
  assign new_n58234_ = ys__n24744 & new_n53763_;
  assign new_n58235_ = ys__n39722 & new_n53753_;
  assign new_n58236_ = ~new_n58234_ & ~new_n58235_;
  assign new_n58237_ = new_n58233_ & new_n58236_;
  assign new_n58238_ = new_n58230_ & new_n58237_;
  assign new_n58239_ = ~new_n58223_ & ~new_n58238_;
  assign new_n58240_ = new_n53797_ & ~new_n58223_;
  assign new_n58241_ = new_n53797_ & ~new_n58238_;
  assign new_n58242_ = ~new_n58240_ & ~new_n58241_;
  assign new_n58243_ = ~new_n58239_ & new_n58242_;
  assign new_n58244_ = ~new_n58165_ & ~new_n58243_;
  assign new_n58245_ = ~new_n58215_ & ~new_n58243_;
  assign new_n58246_ = ~new_n58244_ & ~new_n58245_;
  assign new_n58247_ = ~new_n58216_ & new_n58246_;
  assign new_n58248_ = ~new_n58151_ & ~new_n58247_;
  assign new_n58249_ = ~new_n58161_ & ~new_n58247_;
  assign new_n58250_ = ~new_n58248_ & ~new_n58249_;
  assign ys__n43932 = new_n58162_ | ~new_n58250_;
  assign new_n58252_ = ~new_n58161_ & new_n58248_;
  assign new_n58253_ = ~new_n58161_ & new_n58247_;
  assign new_n58254_ = new_n58151_ & new_n58253_;
  assign new_n58255_ = ~new_n58252_ & ~new_n58254_;
  assign new_n58256_ = new_n58161_ & new_n58247_;
  assign new_n58257_ = ~new_n58151_ & new_n58256_;
  assign new_n58258_ = new_n58161_ & ~new_n58247_;
  assign new_n58259_ = new_n58151_ & new_n58258_;
  assign new_n58260_ = ~new_n58257_ & ~new_n58259_;
  assign ys__n43937 = ~new_n58255_ | ~new_n58260_;
  assign new_n58262_ = ~new_n58215_ & new_n58244_;
  assign new_n58263_ = new_n58165_ & new_n58243_;
  assign new_n58264_ = ~new_n58215_ & new_n58263_;
  assign new_n58265_ = ~new_n58262_ & ~new_n58264_;
  assign new_n58266_ = ~new_n58165_ & new_n58243_;
  assign new_n58267_ = new_n58215_ & new_n58266_;
  assign new_n58268_ = new_n58165_ & ~new_n58243_;
  assign new_n58269_ = new_n58215_ & new_n58268_;
  assign new_n58270_ = ~new_n58267_ & ~new_n58269_;
  assign new_n58271_ = new_n58265_ & new_n58270_;
  assign new_n58272_ = ~new_n58075_ & new_n58092_;
  assign new_n58273_ = new_n58060_ & new_n58091_;
  assign new_n58274_ = ~new_n58075_ & new_n58273_;
  assign new_n58275_ = ~new_n58272_ & ~new_n58274_;
  assign new_n58276_ = ~new_n58060_ & new_n58091_;
  assign new_n58277_ = new_n58075_ & new_n58276_;
  assign new_n58278_ = new_n58060_ & ~new_n58091_;
  assign new_n58279_ = new_n58075_ & new_n58278_;
  assign new_n58280_ = ~new_n58277_ & ~new_n58279_;
  assign new_n58281_ = new_n58275_ & new_n58280_;
  assign new_n58282_ = ~new_n58271_ & ~new_n58281_;
  assign new_n58283_ = ~new_n58238_ & new_n58240_;
  assign new_n58284_ = ~new_n53797_ & new_n58223_;
  assign new_n58285_ = ~new_n58238_ & new_n58284_;
  assign new_n58286_ = ~new_n58283_ & ~new_n58285_;
  assign new_n58287_ = ~new_n53797_ & ~new_n58223_;
  assign new_n58288_ = new_n58238_ & new_n58287_;
  assign new_n58289_ = new_n53797_ & new_n58223_;
  assign new_n58290_ = new_n58238_ & new_n58289_;
  assign new_n58291_ = ~new_n58288_ & ~new_n58290_;
  assign new_n58292_ = new_n58286_ & new_n58291_;
  assign new_n58293_ = ys__n39730 & new_n53834_;
  assign new_n58294_ = ys__n39728 & new_n53833_;
  assign new_n58295_ = ~new_n58293_ & ~new_n58294_;
  assign new_n58296_ = ys__n33695 & new_n53847_;
  assign new_n58297_ = ~ys__n33695 & new_n53850_;
  assign new_n58298_ = ~new_n58296_ & ~new_n58297_;
  assign new_n58299_ = new_n58295_ & new_n58298_;
  assign new_n58300_ = ys__n24765 & new_n53839_;
  assign new_n58301_ = ys__n24762 & new_n53842_;
  assign new_n58302_ = ~new_n58300_ & ~new_n58301_;
  assign new_n58303_ = ys__n24759 & new_n53841_;
  assign new_n58304_ = ys__n39732 & new_n53831_;
  assign new_n58305_ = ~new_n58303_ & ~new_n58304_;
  assign new_n58306_ = new_n58302_ & new_n58305_;
  assign new_n58307_ = new_n58299_ & new_n58306_;
  assign new_n58308_ = ys__n39736 & new_n53723_;
  assign new_n58309_ = ys__n39734 & new_n53726_;
  assign new_n58310_ = ~new_n58308_ & ~new_n58309_;
  assign new_n58311_ = ys__n33701 & new_n53730_;
  assign new_n58312_ = ~ys__n33701 & new_n53733_;
  assign new_n58313_ = ~new_n58311_ & ~new_n58312_;
  assign new_n58314_ = new_n58310_ & new_n58313_;
  assign new_n58315_ = ys__n24774 & new_n53738_;
  assign new_n58316_ = ys__n24771 & new_n53740_;
  assign new_n58317_ = ~new_n58315_ & ~new_n58316_;
  assign new_n58318_ = ys__n24768 & new_n53744_;
  assign new_n58319_ = ys__n39738 & new_n53746_;
  assign new_n58320_ = ~new_n58318_ & ~new_n58319_;
  assign new_n58321_ = new_n58317_ & new_n58320_;
  assign new_n58322_ = new_n58314_ & new_n58321_;
  assign new_n58323_ = ~new_n58307_ & ~new_n58322_;
  assign new_n58324_ = ys__n39724 & new_n53871_;
  assign new_n58325_ = ys__n39722 & new_n53870_;
  assign new_n58326_ = ~new_n58324_ & ~new_n58325_;
  assign new_n58327_ = ys__n33689 & new_n53884_;
  assign new_n58328_ = ~ys__n33689 & new_n53887_;
  assign new_n58329_ = ~new_n58327_ & ~new_n58328_;
  assign new_n58330_ = new_n58326_ & new_n58329_;
  assign new_n58331_ = ys__n24756 & new_n53876_;
  assign new_n58332_ = ys__n24753 & new_n53879_;
  assign new_n58333_ = ~new_n58331_ & ~new_n58332_;
  assign new_n58334_ = ys__n24750 & new_n53878_;
  assign new_n58335_ = ys__n39726 & new_n53868_;
  assign new_n58336_ = ~new_n58334_ & ~new_n58335_;
  assign new_n58337_ = new_n58333_ & new_n58336_;
  assign new_n58338_ = new_n58330_ & new_n58337_;
  assign new_n58339_ = ~new_n58307_ & ~new_n58338_;
  assign new_n58340_ = ~new_n58322_ & ~new_n58338_;
  assign new_n58341_ = ~new_n58339_ & ~new_n58340_;
  assign new_n58342_ = ~new_n58323_ & new_n58341_;
  assign new_n58343_ = ~new_n58292_ & ~new_n58342_;
  assign new_n58344_ = ~new_n58271_ & new_n58343_;
  assign new_n58345_ = ~new_n58281_ & new_n58343_;
  assign new_n58346_ = ~new_n58344_ & ~new_n58345_;
  assign ys__n43975 = new_n58282_ | ~new_n58346_;
  assign new_n58348_ = ~new_n58281_ & new_n58344_;
  assign new_n58349_ = new_n58281_ & new_n58343_;
  assign new_n58350_ = new_n58271_ & new_n58349_;
  assign new_n58351_ = ~new_n58281_ & ~new_n58343_;
  assign new_n58352_ = new_n58271_ & new_n58351_;
  assign new_n58353_ = new_n58281_ & ~new_n58343_;
  assign new_n58354_ = ~new_n58271_ & new_n58353_;
  assign new_n58355_ = ~new_n58352_ & ~new_n58354_;
  assign new_n58356_ = ~new_n58350_ & new_n58355_;
  assign ys__n43980 = new_n58348_ | ~new_n58356_;
  assign new_n58358_ = new_n58292_ & ~new_n58342_;
  assign new_n58359_ = ~new_n58292_ & new_n58342_;
  assign new_n58360_ = ~new_n58358_ & ~new_n58359_;
  assign new_n58361_ = ~new_n58195_ & new_n58212_;
  assign new_n58362_ = new_n58180_ & new_n58211_;
  assign new_n58363_ = ~new_n58195_ & new_n58362_;
  assign new_n58364_ = ~new_n58361_ & ~new_n58363_;
  assign new_n58365_ = ~new_n58180_ & new_n58211_;
  assign new_n58366_ = new_n58195_ & new_n58365_;
  assign new_n58367_ = new_n58180_ & ~new_n58211_;
  assign new_n58368_ = new_n58195_ & new_n58367_;
  assign new_n58369_ = ~new_n58366_ & ~new_n58368_;
  assign new_n58370_ = new_n58364_ & new_n58369_;
  assign new_n58371_ = ~new_n58360_ & ~new_n58370_;
  assign new_n58372_ = ys__n39718 & new_n53756_;
  assign new_n58373_ = ys__n24741 & new_n53755_;
  assign new_n58374_ = ~new_n58372_ & ~new_n58373_;
  assign new_n58375_ = ys__n33683 & new_n53769_;
  assign new_n58376_ = ~ys__n33683 & new_n53772_;
  assign new_n58377_ = ~new_n58375_ & ~new_n58376_;
  assign new_n58378_ = new_n58374_ & new_n58377_;
  assign new_n58379_ = ys__n24747 & new_n53761_;
  assign new_n58380_ = ys__n24744 & new_n53764_;
  assign new_n58381_ = ~new_n58379_ & ~new_n58380_;
  assign new_n58382_ = ys__n24741 & new_n53763_;
  assign new_n58383_ = ys__n39720 & new_n53753_;
  assign new_n58384_ = ~new_n58382_ & ~new_n58383_;
  assign new_n58385_ = new_n58381_ & new_n58384_;
  assign new_n58386_ = new_n58378_ & new_n58385_;
  assign new_n58387_ = ys__n39728 & new_n53834_;
  assign new_n58388_ = ys__n39726 & new_n53833_;
  assign new_n58389_ = ~new_n58387_ & ~new_n58388_;
  assign new_n58390_ = ys__n33693 & new_n53847_;
  assign new_n58391_ = ~ys__n33693 & new_n53850_;
  assign new_n58392_ = ~new_n58390_ & ~new_n58391_;
  assign new_n58393_ = new_n58389_ & new_n58392_;
  assign new_n58394_ = ys__n24762 & new_n53839_;
  assign new_n58395_ = ys__n24759 & new_n53842_;
  assign new_n58396_ = ~new_n58394_ & ~new_n58395_;
  assign new_n58397_ = ys__n24756 & new_n53841_;
  assign new_n58398_ = ys__n39730 & new_n53831_;
  assign new_n58399_ = ~new_n58397_ & ~new_n58398_;
  assign new_n58400_ = new_n58396_ & new_n58399_;
  assign new_n58401_ = new_n58393_ & new_n58400_;
  assign new_n58402_ = ys__n39734 & new_n53723_;
  assign new_n58403_ = ys__n39732 & new_n53726_;
  assign new_n58404_ = ~new_n58402_ & ~new_n58403_;
  assign new_n58405_ = ys__n33699 & new_n53730_;
  assign new_n58406_ = ~ys__n33699 & new_n53733_;
  assign new_n58407_ = ~new_n58405_ & ~new_n58406_;
  assign new_n58408_ = new_n58404_ & new_n58407_;
  assign new_n58409_ = ys__n24771 & new_n53738_;
  assign new_n58410_ = ys__n24768 & new_n53740_;
  assign new_n58411_ = ~new_n58409_ & ~new_n58410_;
  assign new_n58412_ = ys__n24765 & new_n53744_;
  assign new_n58413_ = ys__n39736 & new_n53746_;
  assign new_n58414_ = ~new_n58412_ & ~new_n58413_;
  assign new_n58415_ = new_n58411_ & new_n58414_;
  assign new_n58416_ = new_n58408_ & new_n58415_;
  assign new_n58417_ = ~new_n58401_ & ~new_n58416_;
  assign new_n58418_ = ys__n39722 & new_n53871_;
  assign new_n58419_ = ys__n39720 & new_n53870_;
  assign new_n58420_ = ~new_n58418_ & ~new_n58419_;
  assign new_n58421_ = ys__n33687 & new_n53884_;
  assign new_n58422_ = ~ys__n33687 & new_n53887_;
  assign new_n58423_ = ~new_n58421_ & ~new_n58422_;
  assign new_n58424_ = new_n58420_ & new_n58423_;
  assign new_n58425_ = ys__n24753 & new_n53876_;
  assign new_n58426_ = ys__n24750 & new_n53879_;
  assign new_n58427_ = ~new_n58425_ & ~new_n58426_;
  assign new_n58428_ = ys__n24747 & new_n53878_;
  assign new_n58429_ = ys__n39724 & new_n53868_;
  assign new_n58430_ = ~new_n58428_ & ~new_n58429_;
  assign new_n58431_ = new_n58427_ & new_n58430_;
  assign new_n58432_ = new_n58424_ & new_n58431_;
  assign new_n58433_ = ~new_n58401_ & ~new_n58432_;
  assign new_n58434_ = ~new_n58416_ & ~new_n58432_;
  assign new_n58435_ = ~new_n58433_ & ~new_n58434_;
  assign new_n58436_ = ~new_n58417_ & new_n58435_;
  assign new_n58437_ = ~new_n58386_ & ~new_n58436_;
  assign new_n58438_ = ~new_n58360_ & new_n58437_;
  assign new_n58439_ = ~new_n58370_ & new_n58437_;
  assign new_n58440_ = ~new_n58438_ & ~new_n58439_;
  assign ys__n44018 = new_n58371_ | ~new_n58440_;
  assign new_n58442_ = ~new_n58370_ & new_n58438_;
  assign new_n58443_ = new_n58370_ & new_n58437_;
  assign new_n58444_ = new_n58360_ & new_n58443_;
  assign new_n58445_ = ~new_n58370_ & ~new_n58437_;
  assign new_n58446_ = new_n58360_ & new_n58445_;
  assign new_n58447_ = new_n58370_ & ~new_n58437_;
  assign new_n58448_ = ~new_n58360_ & new_n58447_;
  assign new_n58449_ = ~new_n58446_ & ~new_n58448_;
  assign new_n58450_ = ~new_n58444_ & new_n58449_;
  assign ys__n44023 = new_n58442_ | ~new_n58450_;
  assign new_n58452_ = ys__n24744 & new_n53761_;
  assign new_n58453_ = ys__n24741 & new_n53764_;
  assign new_n58454_ = ~new_n58452_ & ~new_n58453_;
  assign new_n58455_ = ys__n39718 & new_n53753_;
  assign new_n58456_ = ys__n24741 & new_n53756_;
  assign new_n58457_ = ~new_n58455_ & ~new_n58456_;
  assign new_n58458_ = ys__n33681 & new_n53769_;
  assign new_n58459_ = ~ys__n33681 & new_n53772_;
  assign new_n58460_ = ~new_n58458_ & ~new_n58459_;
  assign new_n58461_ = new_n58457_ & new_n58460_;
  assign new_n58462_ = new_n58454_ & new_n58461_;
  assign new_n58463_ = ys__n39726 & new_n53834_;
  assign new_n58464_ = ys__n39724 & new_n53833_;
  assign new_n58465_ = ~new_n58463_ & ~new_n58464_;
  assign new_n58466_ = ys__n33691 & new_n53847_;
  assign new_n58467_ = ~ys__n33691 & new_n53850_;
  assign new_n58468_ = ~new_n58466_ & ~new_n58467_;
  assign new_n58469_ = new_n58465_ & new_n58468_;
  assign new_n58470_ = ys__n24759 & new_n53839_;
  assign new_n58471_ = ys__n24756 & new_n53842_;
  assign new_n58472_ = ~new_n58470_ & ~new_n58471_;
  assign new_n58473_ = ys__n24753 & new_n53841_;
  assign new_n58474_ = ys__n39728 & new_n53831_;
  assign new_n58475_ = ~new_n58473_ & ~new_n58474_;
  assign new_n58476_ = new_n58472_ & new_n58475_;
  assign new_n58477_ = new_n58469_ & new_n58476_;
  assign new_n58478_ = ys__n39732 & new_n53723_;
  assign new_n58479_ = ys__n39730 & new_n53726_;
  assign new_n58480_ = ~new_n58478_ & ~new_n58479_;
  assign new_n58481_ = ys__n33697 & new_n53730_;
  assign new_n58482_ = ~ys__n33697 & new_n53733_;
  assign new_n58483_ = ~new_n58481_ & ~new_n58482_;
  assign new_n58484_ = new_n58480_ & new_n58483_;
  assign new_n58485_ = ys__n24768 & new_n53738_;
  assign new_n58486_ = ys__n24765 & new_n53740_;
  assign new_n58487_ = ~new_n58485_ & ~new_n58486_;
  assign new_n58488_ = ys__n24762 & new_n53744_;
  assign new_n58489_ = ys__n39734 & new_n53746_;
  assign new_n58490_ = ~new_n58488_ & ~new_n58489_;
  assign new_n58491_ = new_n58487_ & new_n58490_;
  assign new_n58492_ = new_n58484_ & new_n58491_;
  assign new_n58493_ = ~new_n58477_ & ~new_n58492_;
  assign new_n58494_ = ys__n39720 & new_n53871_;
  assign new_n58495_ = ys__n39718 & new_n53870_;
  assign new_n58496_ = ~new_n58494_ & ~new_n58495_;
  assign new_n58497_ = ys__n33685 & new_n53884_;
  assign new_n58498_ = ~ys__n33685 & new_n53887_;
  assign new_n58499_ = ~new_n58497_ & ~new_n58498_;
  assign new_n58500_ = new_n58496_ & new_n58499_;
  assign new_n58501_ = ys__n24750 & new_n53876_;
  assign new_n58502_ = ys__n24747 & new_n53879_;
  assign new_n58503_ = ~new_n58501_ & ~new_n58502_;
  assign new_n58504_ = ys__n24744 & new_n53878_;
  assign new_n58505_ = ys__n39722 & new_n53868_;
  assign new_n58506_ = ~new_n58504_ & ~new_n58505_;
  assign new_n58507_ = new_n58503_ & new_n58506_;
  assign new_n58508_ = new_n58500_ & new_n58507_;
  assign new_n58509_ = ~new_n58477_ & ~new_n58508_;
  assign new_n58510_ = ~new_n58492_ & ~new_n58508_;
  assign new_n58511_ = ~new_n58509_ & ~new_n58510_;
  assign new_n58512_ = ~new_n58493_ & new_n58511_;
  assign new_n58513_ = ~new_n58462_ & ~new_n58512_;
  assign new_n58514_ = ys__n24741 & new_n53761_;
  assign new_n58515_ = ys__n24741 & new_n53753_;
  assign new_n58516_ = ~new_n58514_ & ~new_n58515_;
  assign new_n58517_ = ys__n24741 & new_n53769_;
  assign new_n58518_ = ~ys__n24741 & new_n53772_;
  assign new_n58519_ = ~new_n58517_ & ~new_n58518_;
  assign new_n58520_ = new_n58516_ & new_n58519_;
  assign new_n58521_ = new_n53772_ & ~new_n58520_;
  assign new_n58522_ = ~new_n58462_ & new_n58521_;
  assign new_n58523_ = ~new_n58512_ & new_n58521_;
  assign new_n58524_ = ~new_n58522_ & ~new_n58523_;
  assign new_n58525_ = ~new_n58513_ & new_n58524_;
  assign new_n58526_ = ~new_n58322_ & new_n58339_;
  assign new_n58527_ = new_n58307_ & new_n58338_;
  assign new_n58528_ = ~new_n58322_ & new_n58527_;
  assign new_n58529_ = ~new_n58526_ & ~new_n58528_;
  assign new_n58530_ = ~new_n58307_ & new_n58338_;
  assign new_n58531_ = new_n58322_ & new_n58530_;
  assign new_n58532_ = new_n58307_ & ~new_n58338_;
  assign new_n58533_ = new_n58322_ & new_n58532_;
  assign new_n58534_ = ~new_n58531_ & ~new_n58533_;
  assign new_n58535_ = new_n58529_ & new_n58534_;
  assign new_n58536_ = ~new_n58525_ & ~new_n58535_;
  assign new_n58537_ = new_n58386_ & ~new_n58436_;
  assign new_n58538_ = ~new_n58386_ & new_n58436_;
  assign new_n58539_ = ~new_n58537_ & ~new_n58538_;
  assign new_n58540_ = ~new_n58525_ & ~new_n58539_;
  assign new_n58541_ = ~new_n58535_ & ~new_n58539_;
  assign new_n58542_ = ~new_n58540_ & ~new_n58541_;
  assign ys__n44048 = new_n58536_ | ~new_n58542_;
  assign new_n58544_ = ~new_n58535_ & new_n58540_;
  assign new_n58545_ = new_n58535_ & new_n58539_;
  assign new_n58546_ = ~new_n58525_ & new_n58545_;
  assign new_n58547_ = ~new_n58535_ & new_n58539_;
  assign new_n58548_ = new_n58525_ & new_n58547_;
  assign new_n58549_ = new_n58535_ & ~new_n58539_;
  assign new_n58550_ = new_n58525_ & new_n58549_;
  assign new_n58551_ = ~new_n58548_ & ~new_n58550_;
  assign new_n58552_ = ~new_n58546_ & new_n58551_;
  assign ys__n44053 = new_n58544_ | ~new_n58552_;
  assign new_n58554_ = ~new_n58512_ & new_n58522_;
  assign new_n58555_ = new_n58462_ & ~new_n58521_;
  assign new_n58556_ = ~new_n58512_ & new_n58555_;
  assign new_n58557_ = ~new_n58554_ & ~new_n58556_;
  assign new_n58558_ = ~new_n58462_ & ~new_n58521_;
  assign new_n58559_ = new_n58512_ & new_n58558_;
  assign new_n58560_ = new_n58462_ & new_n58521_;
  assign new_n58561_ = new_n58512_ & new_n58560_;
  assign new_n58562_ = ~new_n58559_ & ~new_n58561_;
  assign new_n58563_ = new_n58557_ & new_n58562_;
  assign new_n58564_ = ~new_n58416_ & new_n58433_;
  assign new_n58565_ = new_n58401_ & new_n58432_;
  assign new_n58566_ = ~new_n58416_ & new_n58565_;
  assign new_n58567_ = ~new_n58564_ & ~new_n58566_;
  assign new_n58568_ = ~new_n58401_ & new_n58432_;
  assign new_n58569_ = new_n58416_ & new_n58568_;
  assign new_n58570_ = new_n58401_ & ~new_n58432_;
  assign new_n58571_ = new_n58416_ & new_n58570_;
  assign new_n58572_ = ~new_n58569_ & ~new_n58571_;
  assign new_n58573_ = new_n58567_ & new_n58572_;
  assign new_n58574_ = ~new_n58563_ & ~new_n58573_;
  assign new_n58575_ = ~new_n53772_ & ~new_n58520_;
  assign new_n58576_ = new_n53772_ & new_n58520_;
  assign new_n58577_ = ~new_n58575_ & ~new_n58576_;
  assign new_n58578_ = ys__n39724 & new_n53834_;
  assign new_n58579_ = ys__n39722 & new_n53833_;
  assign new_n58580_ = ~new_n58578_ & ~new_n58579_;
  assign new_n58581_ = ys__n33689 & new_n53847_;
  assign new_n58582_ = ~ys__n33689 & new_n53850_;
  assign new_n58583_ = ~new_n58581_ & ~new_n58582_;
  assign new_n58584_ = new_n58580_ & new_n58583_;
  assign new_n58585_ = ys__n24756 & new_n53839_;
  assign new_n58586_ = ys__n24753 & new_n53842_;
  assign new_n58587_ = ~new_n58585_ & ~new_n58586_;
  assign new_n58588_ = ys__n24750 & new_n53841_;
  assign new_n58589_ = ys__n39726 & new_n53831_;
  assign new_n58590_ = ~new_n58588_ & ~new_n58589_;
  assign new_n58591_ = new_n58587_ & new_n58590_;
  assign new_n58592_ = new_n58584_ & new_n58591_;
  assign new_n58593_ = ys__n39730 & new_n53723_;
  assign new_n58594_ = ys__n39728 & new_n53726_;
  assign new_n58595_ = ~new_n58593_ & ~new_n58594_;
  assign new_n58596_ = ys__n33695 & new_n53730_;
  assign new_n58597_ = ~ys__n33695 & new_n53733_;
  assign new_n58598_ = ~new_n58596_ & ~new_n58597_;
  assign new_n58599_ = new_n58595_ & new_n58598_;
  assign new_n58600_ = ys__n24765 & new_n53738_;
  assign new_n58601_ = ys__n24762 & new_n53740_;
  assign new_n58602_ = ~new_n58600_ & ~new_n58601_;
  assign new_n58603_ = ys__n24759 & new_n53744_;
  assign new_n58604_ = ys__n39732 & new_n53746_;
  assign new_n58605_ = ~new_n58603_ & ~new_n58604_;
  assign new_n58606_ = new_n58602_ & new_n58605_;
  assign new_n58607_ = new_n58599_ & new_n58606_;
  assign new_n58608_ = ~new_n58592_ & ~new_n58607_;
  assign new_n58609_ = ys__n39718 & new_n53871_;
  assign new_n58610_ = ys__n24741 & new_n53870_;
  assign new_n58611_ = ~new_n58609_ & ~new_n58610_;
  assign new_n58612_ = ys__n33683 & new_n53884_;
  assign new_n58613_ = ~ys__n33683 & new_n53887_;
  assign new_n58614_ = ~new_n58612_ & ~new_n58613_;
  assign new_n58615_ = new_n58611_ & new_n58614_;
  assign new_n58616_ = ys__n24747 & new_n53876_;
  assign new_n58617_ = ys__n24744 & new_n53879_;
  assign new_n58618_ = ~new_n58616_ & ~new_n58617_;
  assign new_n58619_ = ys__n24741 & new_n53878_;
  assign new_n58620_ = ys__n39720 & new_n53868_;
  assign new_n58621_ = ~new_n58619_ & ~new_n58620_;
  assign new_n58622_ = new_n58618_ & new_n58621_;
  assign new_n58623_ = new_n58615_ & new_n58622_;
  assign new_n58624_ = ~new_n58592_ & ~new_n58623_;
  assign new_n58625_ = ~new_n58607_ & ~new_n58623_;
  assign new_n58626_ = ~new_n58624_ & ~new_n58625_;
  assign new_n58627_ = ~new_n58608_ & new_n58626_;
  assign new_n58628_ = ~new_n58577_ & ~new_n58627_;
  assign new_n58629_ = ~new_n58563_ & new_n58628_;
  assign new_n58630_ = ~new_n58573_ & new_n58628_;
  assign new_n58631_ = ~new_n58629_ & ~new_n58630_;
  assign ys__n44089 = new_n58574_ | ~new_n58631_;
  assign new_n58633_ = ~new_n58573_ & new_n58629_;
  assign new_n58634_ = new_n58573_ & new_n58628_;
  assign new_n58635_ = new_n58563_ & new_n58634_;
  assign new_n58636_ = ~new_n58573_ & ~new_n58628_;
  assign new_n58637_ = new_n58563_ & new_n58636_;
  assign new_n58638_ = new_n58573_ & ~new_n58628_;
  assign new_n58639_ = ~new_n58563_ & new_n58638_;
  assign new_n58640_ = ~new_n58637_ & ~new_n58639_;
  assign new_n58641_ = ~new_n58635_ & new_n58640_;
  assign ys__n44094 = new_n58633_ | ~new_n58641_;
  assign new_n58643_ = new_n58577_ & ~new_n58627_;
  assign new_n58644_ = ~new_n58577_ & new_n58627_;
  assign new_n58645_ = ~new_n58643_ & ~new_n58644_;
  assign new_n58646_ = ~new_n58492_ & new_n58509_;
  assign new_n58647_ = new_n58477_ & new_n58508_;
  assign new_n58648_ = ~new_n58492_ & new_n58647_;
  assign new_n58649_ = ~new_n58646_ & ~new_n58648_;
  assign new_n58650_ = ~new_n58477_ & new_n58508_;
  assign new_n58651_ = new_n58492_ & new_n58650_;
  assign new_n58652_ = new_n58477_ & ~new_n58508_;
  assign new_n58653_ = new_n58492_ & new_n58652_;
  assign new_n58654_ = ~new_n58651_ & ~new_n58653_;
  assign new_n58655_ = new_n58649_ & new_n58654_;
  assign ys__n44119 = ~new_n58645_ & ~new_n58655_;
  assign new_n58657_ = new_n58645_ & ~new_n58655_;
  assign new_n58658_ = ~new_n58645_ & new_n58655_;
  assign ys__n44122 = new_n58657_ | new_n58658_;
  assign new_n58660_ = ys__n39722 & new_n53834_;
  assign new_n58661_ = ys__n39720 & new_n53833_;
  assign new_n58662_ = ~new_n58660_ & ~new_n58661_;
  assign new_n58663_ = ys__n33687 & new_n53847_;
  assign new_n58664_ = ~ys__n33687 & new_n53850_;
  assign new_n58665_ = ~new_n58663_ & ~new_n58664_;
  assign new_n58666_ = new_n58662_ & new_n58665_;
  assign new_n58667_ = ys__n24753 & new_n53839_;
  assign new_n58668_ = ys__n24750 & new_n53842_;
  assign new_n58669_ = ~new_n58667_ & ~new_n58668_;
  assign new_n58670_ = ys__n24747 & new_n53841_;
  assign new_n58671_ = ys__n39724 & new_n53831_;
  assign new_n58672_ = ~new_n58670_ & ~new_n58671_;
  assign new_n58673_ = new_n58669_ & new_n58672_;
  assign new_n58674_ = new_n58666_ & new_n58673_;
  assign new_n58675_ = ys__n39728 & new_n53723_;
  assign new_n58676_ = ys__n39726 & new_n53726_;
  assign new_n58677_ = ~new_n58675_ & ~new_n58676_;
  assign new_n58678_ = ys__n33693 & new_n53730_;
  assign new_n58679_ = ~ys__n33693 & new_n53733_;
  assign new_n58680_ = ~new_n58678_ & ~new_n58679_;
  assign new_n58681_ = new_n58677_ & new_n58680_;
  assign new_n58682_ = ys__n24762 & new_n53738_;
  assign new_n58683_ = ys__n24759 & new_n53740_;
  assign new_n58684_ = ~new_n58682_ & ~new_n58683_;
  assign new_n58685_ = ys__n24756 & new_n53744_;
  assign new_n58686_ = ys__n39730 & new_n53746_;
  assign new_n58687_ = ~new_n58685_ & ~new_n58686_;
  assign new_n58688_ = new_n58684_ & new_n58687_;
  assign new_n58689_ = new_n58681_ & new_n58688_;
  assign new_n58690_ = ~new_n58674_ & ~new_n58689_;
  assign new_n58691_ = ys__n24744 & new_n53876_;
  assign new_n58692_ = ys__n24741 & new_n53879_;
  assign new_n58693_ = ~new_n58691_ & ~new_n58692_;
  assign new_n58694_ = ys__n39718 & new_n53868_;
  assign new_n58695_ = ys__n24741 & new_n53871_;
  assign new_n58696_ = ~new_n58694_ & ~new_n58695_;
  assign new_n58697_ = ys__n33681 & new_n53884_;
  assign new_n58698_ = ~ys__n33681 & new_n53887_;
  assign new_n58699_ = ~new_n58697_ & ~new_n58698_;
  assign new_n58700_ = new_n58696_ & new_n58699_;
  assign new_n58701_ = new_n58693_ & new_n58700_;
  assign new_n58702_ = ~new_n58674_ & ~new_n58701_;
  assign new_n58703_ = ~new_n58689_ & ~new_n58701_;
  assign new_n58704_ = ~new_n58702_ & ~new_n58703_;
  assign new_n58705_ = ~new_n58690_ & new_n58704_;
  assign new_n58706_ = ~new_n58607_ & new_n58624_;
  assign new_n58707_ = new_n58592_ & new_n58623_;
  assign new_n58708_ = ~new_n58607_ & new_n58707_;
  assign new_n58709_ = ~new_n58706_ & ~new_n58708_;
  assign new_n58710_ = ~new_n58592_ & new_n58623_;
  assign new_n58711_ = new_n58607_ & new_n58710_;
  assign new_n58712_ = new_n58592_ & ~new_n58623_;
  assign new_n58713_ = new_n58607_ & new_n58712_;
  assign new_n58714_ = ~new_n58711_ & ~new_n58713_;
  assign new_n58715_ = new_n58709_ & new_n58714_;
  assign ys__n44136 = ~new_n58705_ & ~new_n58715_;
  assign new_n58717_ = new_n58705_ & ~new_n58715_;
  assign new_n58718_ = ~new_n58705_ & new_n58715_;
  assign ys__n44139 = new_n58717_ | new_n58718_;
  assign new_n58720_ = ys__n39720 & new_n53834_;
  assign new_n58721_ = ys__n39718 & new_n53833_;
  assign new_n58722_ = ~new_n58720_ & ~new_n58721_;
  assign new_n58723_ = ys__n33685 & new_n53847_;
  assign new_n58724_ = ~ys__n33685 & new_n53850_;
  assign new_n58725_ = ~new_n58723_ & ~new_n58724_;
  assign new_n58726_ = new_n58722_ & new_n58725_;
  assign new_n58727_ = ys__n24750 & new_n53839_;
  assign new_n58728_ = ys__n24747 & new_n53842_;
  assign new_n58729_ = ~new_n58727_ & ~new_n58728_;
  assign new_n58730_ = ys__n24744 & new_n53841_;
  assign new_n58731_ = ys__n39722 & new_n53831_;
  assign new_n58732_ = ~new_n58730_ & ~new_n58731_;
  assign new_n58733_ = new_n58729_ & new_n58732_;
  assign new_n58734_ = new_n58726_ & new_n58733_;
  assign new_n58735_ = ys__n39726 & new_n53723_;
  assign new_n58736_ = ys__n39724 & new_n53726_;
  assign new_n58737_ = ~new_n58735_ & ~new_n58736_;
  assign new_n58738_ = ys__n33691 & new_n53730_;
  assign new_n58739_ = ~ys__n33691 & new_n53733_;
  assign new_n58740_ = ~new_n58738_ & ~new_n58739_;
  assign new_n58741_ = new_n58737_ & new_n58740_;
  assign new_n58742_ = ys__n24759 & new_n53738_;
  assign new_n58743_ = ys__n24756 & new_n53740_;
  assign new_n58744_ = ~new_n58742_ & ~new_n58743_;
  assign new_n58745_ = ys__n24753 & new_n53744_;
  assign new_n58746_ = ys__n39728 & new_n53746_;
  assign new_n58747_ = ~new_n58745_ & ~new_n58746_;
  assign new_n58748_ = new_n58744_ & new_n58747_;
  assign new_n58749_ = new_n58741_ & new_n58748_;
  assign new_n58750_ = ~new_n58734_ & ~new_n58749_;
  assign new_n58751_ = ys__n24741 & new_n53876_;
  assign new_n58752_ = ys__n24741 & new_n53868_;
  assign new_n58753_ = ~new_n58751_ & ~new_n58752_;
  assign new_n58754_ = ys__n24741 & new_n53884_;
  assign new_n58755_ = ~ys__n24741 & new_n53887_;
  assign new_n58756_ = ~new_n58754_ & ~new_n58755_;
  assign new_n58757_ = new_n58753_ & new_n58756_;
  assign new_n58758_ = ~new_n58734_ & ~new_n58757_;
  assign new_n58759_ = ~new_n58749_ & ~new_n58757_;
  assign new_n58760_ = ~new_n58758_ & ~new_n58759_;
  assign new_n58761_ = ~new_n58750_ & new_n58760_;
  assign new_n58762_ = ~new_n58689_ & new_n58702_;
  assign new_n58763_ = new_n58674_ & new_n58701_;
  assign new_n58764_ = ~new_n58689_ & new_n58763_;
  assign new_n58765_ = ~new_n58762_ & ~new_n58764_;
  assign new_n58766_ = ~new_n58674_ & new_n58701_;
  assign new_n58767_ = new_n58689_ & new_n58766_;
  assign new_n58768_ = new_n58674_ & ~new_n58701_;
  assign new_n58769_ = new_n58689_ & new_n58768_;
  assign new_n58770_ = ~new_n58767_ & ~new_n58769_;
  assign new_n58771_ = new_n58765_ & new_n58770_;
  assign new_n58772_ = ~new_n58761_ & ~new_n58771_;
  assign new_n58773_ = ys__n39718 & new_n53834_;
  assign new_n58774_ = ys__n24741 & new_n53833_;
  assign new_n58775_ = ~new_n58773_ & ~new_n58774_;
  assign new_n58776_ = ys__n33683 & new_n53847_;
  assign new_n58777_ = ~ys__n33683 & new_n53850_;
  assign new_n58778_ = ~new_n58776_ & ~new_n58777_;
  assign new_n58779_ = new_n58775_ & new_n58778_;
  assign new_n58780_ = ys__n24747 & new_n53839_;
  assign new_n58781_ = ys__n24744 & new_n53842_;
  assign new_n58782_ = ~new_n58780_ & ~new_n58781_;
  assign new_n58783_ = ys__n24741 & new_n53841_;
  assign new_n58784_ = ys__n39720 & new_n53831_;
  assign new_n58785_ = ~new_n58783_ & ~new_n58784_;
  assign new_n58786_ = new_n58782_ & new_n58785_;
  assign new_n58787_ = new_n58779_ & new_n58786_;
  assign new_n58788_ = ys__n39724 & new_n53723_;
  assign new_n58789_ = ys__n39722 & new_n53726_;
  assign new_n58790_ = ~new_n58788_ & ~new_n58789_;
  assign new_n58791_ = ys__n33689 & new_n53730_;
  assign new_n58792_ = ~ys__n33689 & new_n53733_;
  assign new_n58793_ = ~new_n58791_ & ~new_n58792_;
  assign new_n58794_ = new_n58790_ & new_n58793_;
  assign new_n58795_ = ys__n24756 & new_n53738_;
  assign new_n58796_ = ys__n24753 & new_n53740_;
  assign new_n58797_ = ~new_n58795_ & ~new_n58796_;
  assign new_n58798_ = ys__n24750 & new_n53744_;
  assign new_n58799_ = ys__n39726 & new_n53746_;
  assign new_n58800_ = ~new_n58798_ & ~new_n58799_;
  assign new_n58801_ = new_n58797_ & new_n58800_;
  assign new_n58802_ = new_n58794_ & new_n58801_;
  assign new_n58803_ = ~new_n58787_ & ~new_n58802_;
  assign new_n58804_ = new_n53887_ & new_n58803_;
  assign new_n58805_ = ~new_n58761_ & new_n58804_;
  assign new_n58806_ = ~new_n58771_ & new_n58804_;
  assign new_n58807_ = ~new_n58805_ & ~new_n58806_;
  assign ys__n44155 = new_n58772_ | ~new_n58807_;
  assign new_n58809_ = ~new_n58771_ & new_n58805_;
  assign new_n58810_ = new_n58761_ & ~new_n58804_;
  assign new_n58811_ = ~new_n58771_ & new_n58810_;
  assign new_n58812_ = ~new_n58809_ & ~new_n58811_;
  assign new_n58813_ = ~new_n58761_ & ~new_n58804_;
  assign new_n58814_ = new_n58771_ & new_n58813_;
  assign new_n58815_ = new_n58761_ & new_n58804_;
  assign new_n58816_ = new_n58771_ & new_n58815_;
  assign new_n58817_ = ~new_n58814_ & ~new_n58816_;
  assign ys__n44160 = ~new_n58812_ | ~new_n58817_;
  assign new_n58819_ = ~new_n53887_ & new_n58803_;
  assign new_n58820_ = new_n53887_ & ~new_n58803_;
  assign new_n58821_ = ~new_n58819_ & ~new_n58820_;
  assign new_n58822_ = ~new_n58749_ & new_n58758_;
  assign new_n58823_ = new_n58734_ & new_n58757_;
  assign new_n58824_ = ~new_n58749_ & new_n58823_;
  assign new_n58825_ = ~new_n58822_ & ~new_n58824_;
  assign new_n58826_ = ~new_n58734_ & new_n58757_;
  assign new_n58827_ = new_n58749_ & new_n58826_;
  assign new_n58828_ = new_n58734_ & ~new_n58757_;
  assign new_n58829_ = new_n58749_ & new_n58828_;
  assign new_n58830_ = ~new_n58827_ & ~new_n58829_;
  assign new_n58831_ = new_n58825_ & new_n58830_;
  assign ys__n44183 = ~new_n58821_ & ~new_n58831_;
  assign new_n58833_ = new_n58821_ & ~new_n58831_;
  assign new_n58834_ = ~new_n58821_ & new_n58831_;
  assign ys__n44186 = new_n58833_ | new_n58834_;
  assign new_n58836_ = ys__n24744 & new_n53839_;
  assign new_n58837_ = ys__n24741 & new_n53842_;
  assign new_n58838_ = ~new_n58836_ & ~new_n58837_;
  assign new_n58839_ = ys__n39718 & new_n53831_;
  assign new_n58840_ = ys__n24741 & new_n53834_;
  assign new_n58841_ = ~new_n58839_ & ~new_n58840_;
  assign new_n58842_ = ys__n33681 & new_n53847_;
  assign new_n58843_ = ~ys__n33681 & new_n53850_;
  assign new_n58844_ = ~new_n58842_ & ~new_n58843_;
  assign new_n58845_ = new_n58841_ & new_n58844_;
  assign new_n58846_ = new_n58838_ & new_n58845_;
  assign new_n58847_ = ys__n39722 & new_n53723_;
  assign new_n58848_ = ys__n39720 & new_n53726_;
  assign new_n58849_ = ~new_n58847_ & ~new_n58848_;
  assign new_n58850_ = ys__n33687 & new_n53730_;
  assign new_n58851_ = ~ys__n33687 & new_n53733_;
  assign new_n58852_ = ~new_n58850_ & ~new_n58851_;
  assign new_n58853_ = new_n58849_ & new_n58852_;
  assign new_n58854_ = ys__n24753 & new_n53738_;
  assign new_n58855_ = ys__n24750 & new_n53740_;
  assign new_n58856_ = ~new_n58854_ & ~new_n58855_;
  assign new_n58857_ = ys__n24747 & new_n53744_;
  assign new_n58858_ = ys__n39724 & new_n53746_;
  assign new_n58859_ = ~new_n58857_ & ~new_n58858_;
  assign new_n58860_ = new_n58856_ & new_n58859_;
  assign new_n58861_ = new_n58853_ & new_n58860_;
  assign new_n58862_ = ~new_n58846_ & ~new_n58861_;
  assign new_n58863_ = new_n58787_ & ~new_n58802_;
  assign new_n58864_ = ~new_n58787_ & new_n58802_;
  assign new_n58865_ = ~new_n58863_ & ~new_n58864_;
  assign ys__n44189 = new_n58862_ & ~new_n58865_;
  assign new_n58867_ = ~new_n58862_ & ~new_n58865_;
  assign new_n58868_ = new_n58862_ & new_n58865_;
  assign ys__n44192 = new_n58867_ | new_n58868_;
  assign new_n58870_ = ys__n24741 & new_n53839_;
  assign new_n58871_ = ys__n24741 & new_n53831_;
  assign new_n58872_ = ~new_n58870_ & ~new_n58871_;
  assign new_n58873_ = ys__n24741 & new_n53847_;
  assign new_n58874_ = ~ys__n24741 & new_n53850_;
  assign new_n58875_ = ~new_n58873_ & ~new_n58874_;
  assign new_n58876_ = new_n58872_ & new_n58875_;
  assign new_n58877_ = ys__n39720 & new_n53723_;
  assign new_n58878_ = ys__n39718 & new_n53726_;
  assign new_n58879_ = ~new_n58877_ & ~new_n58878_;
  assign new_n58880_ = ys__n33685 & new_n53730_;
  assign new_n58881_ = ~ys__n33685 & new_n53733_;
  assign new_n58882_ = ~new_n58880_ & ~new_n58881_;
  assign new_n58883_ = new_n58879_ & new_n58882_;
  assign new_n58884_ = ys__n24750 & new_n53738_;
  assign new_n58885_ = ys__n24747 & new_n53740_;
  assign new_n58886_ = ~new_n58884_ & ~new_n58885_;
  assign new_n58887_ = ys__n24744 & new_n53744_;
  assign new_n58888_ = ys__n39722 & new_n53746_;
  assign new_n58889_ = ~new_n58887_ & ~new_n58888_;
  assign new_n58890_ = new_n58886_ & new_n58889_;
  assign new_n58891_ = new_n58883_ & new_n58890_;
  assign new_n58892_ = ~new_n58876_ & ~new_n58891_;
  assign new_n58893_ = new_n53850_ & ~new_n58876_;
  assign new_n58894_ = new_n53850_ & ~new_n58891_;
  assign new_n58895_ = ~new_n58893_ & ~new_n58894_;
  assign new_n58896_ = ~new_n58892_ & new_n58895_;
  assign new_n58897_ = new_n58846_ & ~new_n58861_;
  assign new_n58898_ = ~new_n58846_ & new_n58861_;
  assign new_n58899_ = ~new_n58897_ & ~new_n58898_;
  assign ys__n44195 = ~new_n58896_ & ~new_n58899_;
  assign new_n58901_ = new_n58896_ & ~new_n58899_;
  assign new_n58902_ = ~new_n58896_ & new_n58899_;
  assign ys__n44198 = new_n58901_ | new_n58902_;
  assign new_n58904_ = ~new_n58891_ & new_n58893_;
  assign new_n58905_ = ~new_n53850_ & new_n58876_;
  assign new_n58906_ = ~new_n58891_ & new_n58905_;
  assign new_n58907_ = ~new_n58904_ & ~new_n58906_;
  assign new_n58908_ = ~new_n53850_ & ~new_n58876_;
  assign new_n58909_ = new_n58891_ & new_n58908_;
  assign new_n58910_ = new_n53850_ & new_n58876_;
  assign new_n58911_ = new_n58891_ & new_n58910_;
  assign new_n58912_ = ~new_n58909_ & ~new_n58911_;
  assign ys__n44205 = ~new_n58907_ | ~new_n58912_;
  assign new_n58914_ = ys__n24741 & new_n53738_;
  assign new_n58915_ = ys__n24741 & new_n53746_;
  assign new_n58916_ = ~new_n58914_ & ~new_n58915_;
  assign new_n58917_ = ys__n24741 & new_n53730_;
  assign new_n58918_ = ~ys__n24741 & new_n53733_;
  assign new_n58919_ = ~new_n58917_ & ~new_n58918_;
  assign new_n58920_ = new_n58916_ & new_n58919_;
  assign new_n58921_ = new_n53733_ & ~new_n58920_;
  assign new_n58922_ = ys__n24744 & new_n53738_;
  assign new_n58923_ = ys__n24741 & new_n53740_;
  assign new_n58924_ = ~new_n58922_ & ~new_n58923_;
  assign new_n58925_ = ys__n39718 & new_n53746_;
  assign new_n58926_ = ys__n24741 & new_n53723_;
  assign new_n58927_ = ~new_n58925_ & ~new_n58926_;
  assign new_n58928_ = ys__n33681 & new_n53730_;
  assign new_n58929_ = ~ys__n33681 & new_n53733_;
  assign new_n58930_ = ~new_n58928_ & ~new_n58929_;
  assign new_n58931_ = new_n58927_ & new_n58930_;
  assign new_n58932_ = new_n58924_ & new_n58931_;
  assign ys__n44213 = new_n58921_ & ~new_n58932_;
  assign new_n58934_ = ~new_n58921_ & ~new_n58932_;
  assign new_n58935_ = new_n58921_ & new_n58932_;
  assign ys__n44216 = new_n58934_ | new_n58935_;
  assign new_n58937_ = ~new_n53733_ & ~new_n58920_;
  assign new_n58938_ = new_n53733_ & new_n58920_;
  assign ys__n44219 = new_n58937_ | new_n58938_;
  assign new_n58940_ = new_n13472_ & new_n13741_;
  assign new_n58941_ = ys__n948 & new_n58940_;
  assign ys__n44838 = ys__n44836 | new_n58941_;
  assign ys__n44841 = ys__n44840 & ~ys__n4566;
  assign ys__n44843 = ys__n44842 & ~ys__n4566;
  assign new_n58945_ = ys__n160 & ys__n344;
  assign new_n58946_ = ys__n352 & new_n58945_;
  assign new_n58947_ = new_n13734_ & new_n58946_;
  assign new_n58948_ = new_n13483_ & new_n58947_;
  assign new_n58949_ = new_n42818_ & ~new_n58948_;
  assign ys__n44844 = ys__n948 & ~new_n58949_;
  assign ys__n44845 = ys__n948 & ~new_n53251_;
  assign new_n58952_ = new_n13726_ & new_n53239_;
  assign new_n58953_ = new_n53241_ & new_n58952_;
  assign new_n58954_ = new_n53243_ & new_n58952_;
  assign new_n58955_ = ~new_n58953_ & ~new_n58954_;
  assign new_n58956_ = new_n13732_ & new_n58952_;
  assign new_n58957_ = ys__n352 & new_n53247_;
  assign new_n58958_ = new_n58952_ & new_n58957_;
  assign new_n58959_ = ~new_n58956_ & ~new_n58958_;
  assign new_n58960_ = new_n58955_ & new_n58959_;
  assign ys__n44846 = ys__n948 & ~new_n58960_;
  assign ys__n44848 = ys__n44847 & ~ys__n4566;
  assign ys__n44850 = ys__n44849 & ~ys__n4566;
  assign new_n58964_ = new_n13738_ & new_n53252_;
  assign new_n58965_ = ~new_n42817_ & ~new_n53244_;
  assign new_n58966_ = ~new_n53249_ & ~new_n58954_;
  assign new_n58967_ = ~new_n58958_ & new_n58966_;
  assign new_n58968_ = new_n58965_ & new_n58967_;
  assign new_n58969_ = new_n58964_ & new_n58968_;
  assign new_n58970_ = ~new_n42816_ & ~new_n53242_;
  assign new_n58971_ = ~new_n53246_ & ~new_n58953_;
  assign new_n58972_ = ~new_n58956_ & new_n58971_;
  assign new_n58973_ = new_n58970_ & new_n58972_;
  assign new_n58974_ = new_n58969_ & new_n58973_;
  assign new_n58975_ = ~new_n58969_ & ~new_n58974_;
  assign ys__n44851 = ys__n948 & new_n58975_;
  assign new_n58977_ = new_n58964_ & new_n58973_;
  assign new_n58978_ = ~new_n58974_ & ~new_n58977_;
  assign ys__n44852 = ys__n948 & new_n58978_;
  assign ys__n44853 = ys__n948 & ~new_n42812_;
  assign new_n58981_ = ~new_n53244_ & ~new_n58954_;
  assign new_n58982_ = ~new_n53242_ & ~new_n58953_;
  assign new_n58983_ = new_n42812_ & new_n58982_;
  assign new_n58984_ = new_n58981_ & new_n58983_;
  assign new_n58985_ = ys__n948 & ~new_n58981_;
  assign ys__n44854 = ~new_n58984_ & new_n58985_;
  assign new_n58987_ = ys__n948 & ~new_n58983_;
  assign ys__n44855 = ~new_n58984_ & new_n58987_;
  assign new_n58989_ = ys__n152 & ~ys__n158;
  assign new_n58990_ = ys__n148 & new_n42796_;
  assign new_n58991_ = new_n58989_ & new_n58990_;
  assign new_n58992_ = new_n42792_ & new_n58990_;
  assign new_n58993_ = ~new_n58991_ & ~new_n58992_;
  assign new_n58994_ = new_n42802_ & new_n58993_;
  assign new_n58995_ = new_n42795_ & new_n58994_;
  assign new_n58996_ = ~new_n42791_ & new_n58994_;
  assign new_n58997_ = ~ys__n30837 & ~new_n58996_;
  assign new_n58998_ = ~new_n58995_ & new_n58997_;
  assign new_n58999_ = ~new_n42794_ & new_n58994_;
  assign new_n59000_ = ~ys__n30837 & ~new_n58995_;
  assign new_n59001_ = ~new_n58999_ & new_n59000_;
  assign new_n59002_ = ~new_n58998_ & ~new_n59001_;
  assign new_n59003_ = ~ys__n4839 & ~ys__n4840;
  assign new_n59004_ = ~ys__n402 & ~new_n17381_;
  assign new_n59005_ = new_n17402_ & new_n59004_;
  assign new_n59006_ = new_n59003_ & ~new_n59005_;
  assign new_n59007_ = ~new_n59002_ & new_n59006_;
  assign new_n59008_ = new_n58978_ & new_n58998_;
  assign new_n59009_ = new_n58975_ & new_n59001_;
  assign new_n59010_ = ~new_n59008_ & ~new_n59009_;
  assign new_n59011_ = new_n53254_ & ~new_n58940_;
  assign new_n59012_ = ~new_n59010_ & ~new_n59011_;
  assign new_n59013_ = ~new_n59007_ & ~new_n59012_;
  assign new_n59014_ = ys__n948 & ~new_n59013_;
  assign new_n59015_ = new_n42789_ & new_n42797_;
  assign new_n59016_ = ys__n148 & new_n59015_;
  assign new_n59017_ = new_n42789_ & new_n58989_;
  assign new_n59018_ = ys__n148 & new_n59017_;
  assign new_n59019_ = ~new_n59016_ & ~new_n59018_;
  assign new_n59020_ = ~ys__n30837 & new_n59018_;
  assign new_n59021_ = ~new_n59019_ & new_n59020_;
  assign new_n59022_ = new_n58975_ & new_n59021_;
  assign new_n59023_ = ~ys__n30837 & new_n59016_;
  assign new_n59024_ = ~new_n59019_ & new_n59023_;
  assign new_n59025_ = new_n58978_ & new_n59024_;
  assign new_n59026_ = ~new_n59021_ & ~new_n59024_;
  assign new_n59027_ = ~new_n59005_ & ~new_n59026_;
  assign new_n59028_ = new_n59003_ & new_n59027_;
  assign new_n59029_ = ys__n30820 & new_n59024_;
  assign new_n59030_ = ys__n30819 & new_n59021_;
  assign new_n59031_ = ~new_n59029_ & ~new_n59030_;
  assign new_n59032_ = ys__n2779 & ~new_n59031_;
  assign new_n59033_ = ys__n44849 & new_n59024_;
  assign new_n59034_ = ys__n44847 & new_n59021_;
  assign new_n59035_ = ~new_n59033_ & ~new_n59034_;
  assign new_n59036_ = ~new_n59032_ & new_n59035_;
  assign new_n59037_ = ~new_n59028_ & new_n59036_;
  assign new_n59038_ = ~new_n59025_ & new_n59037_;
  assign new_n59039_ = ~new_n59022_ & new_n59038_;
  assign new_n59040_ = ys__n948 & ~new_n59039_;
  assign new_n59041_ = new_n17401_ & new_n42824_;
  assign new_n59042_ = new_n42812_ & new_n59041_;
  assign new_n59043_ = new_n58973_ & new_n59042_;
  assign new_n59044_ = new_n58968_ & new_n58973_;
  assign new_n59045_ = new_n59042_ & new_n59044_;
  assign new_n59046_ = ~new_n59043_ & ~new_n59045_;
  assign new_n59047_ = new_n58968_ & new_n59042_;
  assign new_n59048_ = ~new_n59045_ & ~new_n59047_;
  assign new_n59049_ = ~new_n59046_ & ~new_n59048_;
  assign new_n59050_ = ~ys__n4836 & ~ys__n4837;
  assign new_n59051_ = ~new_n59004_ & new_n59050_;
  assign new_n59052_ = ~ys__n4566 & ys__n30832;
  assign new_n59053_ = new_n59051_ & new_n59052_;
  assign new_n59054_ = ~new_n59049_ & new_n59053_;
  assign new_n59055_ = new_n13476_ & new_n42813_;
  assign new_n59056_ = new_n13476_ & new_n42806_;
  assign new_n59057_ = ~new_n59055_ & ~new_n59056_;
  assign new_n59058_ = new_n59055_ & ~new_n59057_;
  assign new_n59059_ = ys__n30819 & new_n59058_;
  assign new_n59060_ = new_n59056_ & ~new_n59057_;
  assign new_n59061_ = ys__n30820 & new_n59060_;
  assign new_n59062_ = ~new_n59059_ & ~new_n59061_;
  assign new_n59063_ = ys__n2779 & ~new_n59062_;
  assign new_n59064_ = ~new_n59058_ & ~new_n59060_;
  assign new_n59065_ = new_n59051_ & ~new_n59064_;
  assign new_n59066_ = ys__n44847 & new_n59058_;
  assign new_n59067_ = ys__n44849 & new_n59060_;
  assign new_n59068_ = ~new_n59066_ & ~new_n59067_;
  assign new_n59069_ = ~new_n59065_ & new_n59068_;
  assign new_n59070_ = ~new_n59063_ & new_n59069_;
  assign new_n59071_ = new_n59052_ & ~new_n59070_;
  assign new_n59072_ = ~new_n59004_ & new_n59052_;
  assign new_n59073_ = ~new_n17402_ & new_n59072_;
  assign new_n59074_ = ~ys__n30837 & ~new_n58993_;
  assign new_n59075_ = ~ys__n4566 & new_n59074_;
  assign new_n59076_ = ~ys__n30832 & new_n59075_;
  assign new_n59077_ = ~new_n59005_ & new_n59076_;
  assign new_n59078_ = new_n42805_ & ~new_n53254_;
  assign new_n59079_ = ~new_n59077_ & ~new_n59078_;
  assign new_n59080_ = ~new_n59073_ & new_n59079_;
  assign new_n59081_ = ~new_n59071_ & new_n59080_;
  assign new_n59082_ = ~new_n59054_ & new_n59081_;
  assign new_n59083_ = ~new_n59040_ & new_n59082_;
  assign ys__n44858 = new_n59014_ | ~new_n59083_;
  assign ys__n44948 = ~ys__n4566 & new_n59021_;
  assign ys__n44949 = ~ys__n4566 & new_n59024_;
  assign new_n59087_ = new_n42795_ & new_n59019_;
  assign new_n59088_ = new_n58994_ & new_n59087_;
  assign new_n59089_ = ~ys__n30837 & ~ys__n30832;
  assign new_n59090_ = ~new_n59088_ & new_n59089_;
  assign new_n59091_ = ys__n352 & ys__n30832;
  assign new_n59092_ = ~new_n59090_ & ~new_n59091_;
  assign ys__n44950 = ~ys__n4566 & ~new_n59092_;
  assign new_n59094_ = ~ys__n22792 & ys__n38927;
  assign ys__n44985 = ys__n46954 & new_n59094_;
  assign new_n59096_ = ~ys__n38236 & ~ys__n38237;
  assign new_n59097_ = ~ys__n33364 & ~new_n59096_;
  assign ys__n44987 = new_n15018_ & new_n59097_;
  assign new_n59099_ = ~new_n52541_ & new_n52549_;
  assign ys__n46131 = ys__n46130 | new_n59099_;
  assign new_n59101_ = ~new_n52541_ & new_n52548_;
  assign ys__n46133 = ys__n46132 | new_n59101_;
  assign new_n59103_ = ~new_n52541_ & new_n52546_;
  assign ys__n46135 = ys__n46134 | new_n59103_;
  assign new_n59105_ = ~new_n52541_ & new_n52545_;
  assign ys__n46137 = ys__n46136 | new_n59105_;
  assign new_n59107_ = ~ys__n35028 & ys__n26573;
  assign new_n59108_ = ~ys__n30863 & ~new_n59107_;
  assign new_n59109_ = ~ys__n46141 & ys__n46142;
  assign new_n59110_ = ys__n46141 & ~ys__n46142;
  assign new_n59111_ = ~new_n59109_ & ~new_n59110_;
  assign ys__n46143 = ~new_n59108_ & new_n59111_;
  assign new_n59113_ = ~ys__n34988 & ys__n26555;
  assign new_n59114_ = ~ys__n34966 & new_n59113_;
  assign new_n59115_ = ys__n34966 & ~new_n59113_;
  assign ys__n46146 = new_n59114_ | new_n59115_;
  assign new_n59117_ = ys__n18317 & ~new_n33481_;
  assign ys__n46159 = ~ys__n34962 & new_n59117_;
  assign new_n59119_ = ~ys__n35033 & ys__n46159;
  assign new_n59120_ = ~ys__n35047 & ~new_n59119_;
  assign new_n59121_ = ~ys__n46152 & ys__n46153;
  assign new_n59122_ = ys__n46152 & ~ys__n46153;
  assign new_n59123_ = ~new_n59121_ & ~new_n59122_;
  assign ys__n46154 = ~new_n59120_ & new_n59123_;
  assign new_n59125_ = ys__n46150 & ~ys__n46151;
  assign new_n59126_ = ~ys__n46150 & ys__n46151;
  assign new_n59127_ = ~ys__n26565 & ~new_n59126_;
  assign new_n59128_ = ~new_n59125_ & new_n59127_;
  assign new_n59129_ = ~ys__n30941 & ~ys__n35031;
  assign ys__n46163 = ~ys__n26291 & new_n59129_;
  assign new_n59131_ = ~ys__n34976 & ys__n46163;
  assign ys__n46155 = ~new_n59128_ & ~new_n59131_;
  assign new_n59133_ = ~ys__n34972 & new_n59119_;
  assign new_n59134_ = ys__n34972 & ~new_n59119_;
  assign ys__n46158 = new_n59133_ | new_n59134_;
  assign new_n59136_ = ~ys__n34978 & new_n59131_;
  assign new_n59137_ = ys__n34978 & ~new_n59131_;
  assign ys__n46162 = new_n59136_ | new_n59137_;
  assign new_n59139_ = ~ys__n35035 & ys__n26288;
  assign new_n59140_ = ~ys__n26561 & ~new_n59139_;
  assign new_n59141_ = ~ys__n46170 & ys__n46171;
  assign new_n59142_ = ys__n46170 & ~ys__n46171;
  assign new_n59143_ = ~new_n59141_ & ~new_n59142_;
  assign ys__n46172 = ~new_n59140_ & new_n59143_;
  assign new_n59145_ = ys__n46168 & ~ys__n46169;
  assign new_n59146_ = ~ys__n46168 & ys__n46169;
  assign new_n59147_ = ~ys__n46166 & ~new_n59146_;
  assign new_n59148_ = ~new_n59145_ & new_n59147_;
  assign ys__n46173 = ~new_n59113_ & ~new_n59148_;
  assign new_n59150_ = ~ys__n34984 & new_n59139_;
  assign new_n59151_ = ys__n34984 & ~new_n59139_;
  assign ys__n46176 = new_n59150_ | new_n59151_;
  assign new_n59153_ = ~ys__n34990 & new_n59113_;
  assign new_n59154_ = ys__n34990 & ~new_n59113_;
  assign ys__n46179 = new_n59153_ | new_n59154_;
  assign new_n59156_ = ~ys__n35037 & ys__n26294;
  assign new_n59157_ = ~ys__n46180 & ~new_n59156_;
  assign new_n59158_ = ~ys__n46186 & ys__n46187;
  assign new_n59159_ = ys__n46186 & ~ys__n46187;
  assign new_n59160_ = ~new_n59158_ & ~new_n59159_;
  assign ys__n46188 = ~new_n59157_ & new_n59160_;
  assign new_n59162_ = ys__n46184 & ~ys__n46185;
  assign new_n59163_ = ~ys__n46184 & ys__n46185;
  assign new_n59164_ = ~ys__n26553 & ~new_n59163_;
  assign new_n59165_ = ~new_n59162_ & new_n59164_;
  assign new_n59166_ = ~ys__n35000 & ys__n26282;
  assign ys__n46189 = ~new_n59165_ & ~new_n59166_;
  assign new_n59168_ = ~ys__n34996 & new_n59156_;
  assign new_n59169_ = ys__n34996 & ~new_n59156_;
  assign ys__n46192 = new_n59168_ | new_n59169_;
  assign new_n59171_ = ~ys__n35002 & new_n59166_;
  assign new_n59172_ = ys__n35002 & ~new_n59166_;
  assign ys__n46195 = new_n59171_ | new_n59172_;
  assign new_n59174_ = ~ys__n35039 & ys__n26284;
  assign new_n59175_ = ~ys__n26554 & ~new_n59174_;
  assign new_n59176_ = ~ys__n46202 & ys__n46203;
  assign new_n59177_ = ys__n46202 & ~ys__n46203;
  assign new_n59178_ = ~new_n59176_ & ~new_n59177_;
  assign ys__n46204 = ~new_n59175_ & new_n59178_;
  assign new_n59180_ = ys__n46200 & ~ys__n46201;
  assign new_n59181_ = ~ys__n46200 & ys__n46201;
  assign new_n59182_ = ~ys__n46198 & ~new_n59181_;
  assign new_n59183_ = ~new_n59180_ & new_n59182_;
  assign new_n59184_ = ~ys__n35012 & ys__n26293;
  assign ys__n46205 = ~new_n59183_ & ~new_n59184_;
  assign new_n59186_ = ~ys__n35008 & new_n59174_;
  assign new_n59187_ = ys__n35008 & ~new_n59174_;
  assign ys__n46208 = new_n59186_ | new_n59187_;
  assign new_n59189_ = ~ys__n35014 & new_n59184_;
  assign new_n59190_ = ys__n35014 & ~new_n59184_;
  assign ys__n46211 = new_n59189_ | new_n59190_;
  assign new_n59192_ = ~ys__n35041 & ys__n26286;
  assign new_n59193_ = ~ys__n26560 & ~new_n59192_;
  assign new_n59194_ = ~ys__n46218 & ys__n46219;
  assign new_n59195_ = ys__n46218 & ~ys__n46219;
  assign new_n59196_ = ~new_n59194_ & ~new_n59195_;
  assign ys__n46220 = ~new_n59193_ & new_n59196_;
  assign new_n59198_ = ys__n46216 & ~ys__n46217;
  assign new_n59199_ = ~ys__n46216 & ys__n46217;
  assign new_n59200_ = ~ys__n46214 & ~new_n59199_;
  assign new_n59201_ = ~new_n59198_ & new_n59200_;
  assign new_n59202_ = ~ys__n35024 & ys__n37738;
  assign ys__n46221 = ~new_n59201_ & ~new_n59202_;
  assign new_n59204_ = ~ys__n35020 & new_n59192_;
  assign new_n59205_ = ys__n35020 & ~new_n59192_;
  assign ys__n46224 = new_n59204_ | new_n59205_;
  assign new_n59207_ = ~ys__n35026 & new_n59202_;
  assign new_n59208_ = ys__n35026 & ~new_n59202_;
  assign ys__n46227 = new_n59207_ | new_n59208_;
  assign ys__n46233 = ~ys__n26562 & ys__n26563;
  assign new_n59211_ = ~ys__n25470 & ys__n30863;
  assign ys__n46234 = ys__n46166 | new_n59211_;
  assign new_n59213_ = ys__n312 & ~ys__n622;
  assign new_n59214_ = ~ys__n312 & ys__n622;
  assign ys__n48339 = new_n59213_ | new_n59214_;
  assign new_n59216_ = ~ys__n620 & new_n17624_;
  assign new_n59217_ = ys__n620 & ~new_n17624_;
  assign ys__n48340 = new_n59216_ | new_n59217_;
  assign new_n59219_ = ys__n620 & new_n17624_;
  assign new_n59220_ = ~ys__n618 & new_n59219_;
  assign new_n59221_ = ys__n618 & ~new_n59219_;
  assign ys__n48341 = new_n59220_ | new_n59221_;
  assign new_n59223_ = ~ys__n614 & new_n17626_;
  assign new_n59224_ = ys__n614 & ~new_n17626_;
  assign ys__n48342 = new_n59223_ | new_n59224_;
  assign new_n59226_ = ys__n614 & new_n17626_;
  assign new_n59227_ = ~ys__n612 & new_n59226_;
  assign new_n59228_ = ys__n612 & ~new_n59226_;
  assign ys__n48343 = new_n59227_ | new_n59228_;
  assign new_n59230_ = new_n17626_ & new_n17627_;
  assign new_n59231_ = ~ys__n616 & new_n59230_;
  assign new_n59232_ = ys__n616 & ~new_n59230_;
  assign ys__n48344 = new_n59231_ | new_n59232_;
  assign new_n59234_ = new_n42095_ & new_n42111_;
  assign new_n59235_ = ~new_n42095_ & ~new_n42111_;
  assign ys__n48349 = new_n59234_ | new_n59235_;
  assign new_n59237_ = ~new_n42095_ & new_n42111_;
  assign new_n59238_ = ~new_n42115_ & ~new_n59237_;
  assign new_n59239_ = new_n42104_ & ~new_n59238_;
  assign new_n59240_ = ~new_n42104_ & new_n59238_;
  assign ys__n48350 = new_n59239_ | new_n59240_;
  assign new_n59242_ = ~new_n42118_ & new_n42155_;
  assign new_n59243_ = new_n42118_ & ~new_n42155_;
  assign ys__n48351 = new_n59242_ | new_n59243_;
  assign new_n59245_ = ~new_n42118_ & ~new_n42155_;
  assign new_n59246_ = ~new_n42160_ & ~new_n59245_;
  assign new_n59247_ = new_n42152_ & ~new_n59246_;
  assign new_n59248_ = ~new_n42152_ & new_n59246_;
  assign ys__n48352 = new_n59247_ | new_n59248_;
  assign new_n59250_ = ~new_n42118_ & new_n42156_;
  assign new_n59251_ = new_n42162_ & ~new_n59250_;
  assign new_n59252_ = new_n42142_ & ~new_n59251_;
  assign new_n59253_ = ~new_n42142_ & new_n59251_;
  assign ys__n48353 = new_n59252_ | new_n59253_;
  assign new_n59255_ = ~new_n42142_ & ~new_n59251_;
  assign new_n59256_ = ~new_n42165_ & ~new_n59255_;
  assign new_n59257_ = new_n42133_ & ~new_n59256_;
  assign new_n59258_ = ~new_n42133_ & new_n59256_;
  assign ys__n48354 = new_n59257_ | new_n59258_;
  assign new_n59260_ = ~new_n42169_ & new_n42239_;
  assign new_n59261_ = new_n42169_ & ~new_n42239_;
  assign ys__n48355 = new_n59260_ | new_n59261_;
  assign new_n59263_ = ~new_n42169_ & ~new_n42239_;
  assign new_n59264_ = ~new_n42245_ & ~new_n59263_;
  assign new_n59265_ = new_n42236_ & ~new_n59264_;
  assign new_n59266_ = ~new_n42236_ & new_n59264_;
  assign ys__n48356 = new_n59265_ | new_n59266_;
  assign new_n59268_ = ~new_n42169_ & new_n42240_;
  assign new_n59269_ = new_n42247_ & ~new_n59268_;
  assign new_n59270_ = new_n42226_ & ~new_n59269_;
  assign new_n59271_ = ~new_n42226_ & new_n59269_;
  assign ys__n48357 = new_n59270_ | new_n59271_;
  assign new_n59273_ = ~new_n42226_ & ~new_n59269_;
  assign new_n59274_ = ~new_n42250_ & ~new_n59273_;
  assign new_n59275_ = new_n42217_ & ~new_n59274_;
  assign new_n59276_ = ~new_n42217_ & new_n59274_;
  assign ys__n48358 = new_n59275_ | new_n59276_;
  assign new_n59278_ = ~new_n42169_ & new_n42241_;
  assign new_n59279_ = new_n42253_ & ~new_n59278_;
  assign new_n59280_ = new_n42206_ & ~new_n59279_;
  assign new_n59281_ = ~new_n42206_ & new_n59279_;
  assign ys__n48359 = new_n59280_ | new_n59281_;
  assign new_n59283_ = ~new_n42206_ & ~new_n59279_;
  assign new_n59284_ = ~new_n42256_ & ~new_n59283_;
  assign new_n59285_ = new_n42197_ & ~new_n59284_;
  assign new_n59286_ = ~new_n42197_ & new_n59284_;
  assign ys__n48360 = new_n59285_ | new_n59286_;
  assign new_n59288_ = new_n42207_ & ~new_n59279_;
  assign new_n59289_ = new_n42258_ & ~new_n59288_;
  assign new_n59290_ = new_n42187_ & ~new_n59289_;
  assign new_n59291_ = ~new_n42187_ & new_n59289_;
  assign ys__n48361 = new_n59290_ | new_n59291_;
  assign new_n59293_ = ~new_n42187_ & ~new_n59289_;
  assign new_n59294_ = ~new_n42261_ & ~new_n59293_;
  assign new_n59295_ = new_n42178_ & ~new_n59294_;
  assign new_n59296_ = ~new_n42178_ & new_n59294_;
  assign ys__n48362 = new_n59295_ | new_n59296_;
  assign ys__n264 = 1'b0;
  assign ys__n28247 = 1'b0;
  assign ys__n28249 = 1'b1;
  assign ys__n28250 = 1'b0;
  assign ys__n28251 = 1'b0;
  assign ys__n28252 = 1'b0;
  assign ys__n28254 = 1'b0;
  assign ys__n28256 = 1'b1;
  assign ys__n28259 = 1'b0;
  assign ys__n28261 = 1'b0;
  assign ys__n28263 = 1'b0;
  assign ys__n28265 = 1'b0;
  assign ys__n28266 = 1'b0;
  assign ys__n28268 = 1'b0;
  assign ys__n28270 = 1'b0;
  assign ys__n28271 = 1'b0;
  assign ys__n28272 = 1'b0;
  assign ys__n28274 = 1'b0;
  assign ys__n28858 = 1'b0;
  assign ys__n30836 = 1'b0;
  assign ys__n30856 = 1'b0;
  assign ys__n30858 = 1'b0;
  assign ys__n30860 = 1'b0;
  assign ys__n38185 = 1'b0;
  assign ys__n38186 = 1'b0;
  assign ys__n38188 = 1'b0;
  assign ys__n38191 = 1'b0;
  assign ys__n280 = ~ys__n20273;
  assign ys__n313 = ~ys__n312;
  assign ys__n319 = ~ys__n318;
  assign ys__n415 = ~ys__n414;
  assign ys__n417 = ~ys__n416;
  assign ys__n455 = ~ys__n454;
  assign ys__n457 = ~ys__n456;
  assign ys__n565 = ~ys__n564;
  assign ys__n890 = ~ys__n874;
  assign ys__n18131 = ~ys__n33515;
  assign ys__n18386 = ~ys__n33324;
  assign ys__n18391 = ~ys__n33317;
  assign ys__n23340 = ~ys__n28243;
  assign ys__n33329 = ~ys__n33328;
  assign ys__n33331 = ~ys__n33330;
  assign ys__n33333 = ~ys__n33332;
  assign ys__n33335 = ~ys__n33334;
  assign ys__n33337 = ~ys__n33336;
  assign ys__n33339 = ~ys__n33338;
  assign ys__n33420 = ~ys__n18121;
  assign ys__n33437 = ~ys__n33438;
  assign ys__n33439 = ~ys__n24177;
  assign ys__n33453 = ~ys__n33454;
  assign ys__n33456 = ~ys__n33455;
  assign ys__n33513 = ~ys__n33514;
  assign ys__n33535 = ~ys__n24590;
  assign ys__n4175 = ys__n738;
  assign ys__n28269 = ys__n23340;
  assign ys__n28334 = ys__n28276;
  assign ys__n38338 = ys__n38334;
  assign ys__n48348 = ys__n35144;
endmodule


